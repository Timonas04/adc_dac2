VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 112.465 219.150 113.275 219.290 ;
        RECT 112.275 218.980 113.275 219.150 ;
        RECT 112.465 217.920 113.275 218.980 ;
        RECT 112.465 217.770 113.275 217.910 ;
        RECT 112.275 217.600 113.275 217.770 ;
        RECT 112.465 212.400 113.275 217.600 ;
        RECT 112.465 212.250 113.275 212.390 ;
        RECT 112.275 212.080 113.275 212.250 ;
        RECT 112.465 208.720 113.275 212.080 ;
        RECT 112.305 208.455 112.415 208.575 ;
        RECT 112.465 208.110 113.145 208.250 ;
        RECT 112.275 207.940 113.145 208.110 ;
        RECT 112.465 207.765 113.145 207.940 ;
        RECT 112.465 206.420 113.375 207.765 ;
        RECT 112.550 205.970 113.335 206.400 ;
        RECT 112.305 205.695 112.415 205.815 ;
        RECT 112.465 204.145 113.375 205.490 ;
        RECT 112.465 203.970 113.145 204.145 ;
        RECT 112.275 203.800 113.145 203.970 ;
        RECT 112.465 203.660 113.145 203.800 ;
        RECT 112.465 203.510 113.145 203.650 ;
        RECT 112.275 203.340 113.145 203.510 ;
      LAYER nwell ;
        RECT 11.760 200.455 90.800 202.060 ;
      LAYER pwell ;
        RECT 11.955 199.255 13.325 200.065 ;
        RECT 13.335 199.255 18.845 200.065 ;
        RECT 18.855 199.255 24.365 200.065 ;
        RECT 24.845 199.340 25.275 200.125 ;
        RECT 25.295 199.255 30.805 200.065 ;
        RECT 30.815 199.255 36.325 200.065 ;
        RECT 36.335 199.255 37.705 200.065 ;
        RECT 37.725 199.340 38.155 200.125 ;
        RECT 38.175 199.255 43.685 200.065 ;
        RECT 43.695 199.255 49.205 200.065 ;
        RECT 49.215 199.255 50.585 200.065 ;
        RECT 50.605 199.340 51.035 200.125 ;
        RECT 51.055 199.255 56.565 200.065 ;
        RECT 56.575 199.935 57.495 200.165 ;
        RECT 112.465 200.135 113.145 203.340 ;
        RECT 56.575 199.255 58.865 199.935 ;
        RECT 58.875 199.255 61.625 200.065 ;
        RECT 61.635 199.255 63.005 200.035 ;
        RECT 63.485 199.340 63.915 200.125 ;
        RECT 63.935 199.255 69.445 200.065 ;
        RECT 69.455 199.255 71.285 200.065 ;
        RECT 71.295 199.255 72.665 200.035 ;
        RECT 72.675 199.255 76.345 200.065 ;
        RECT 76.365 199.340 76.795 200.125 ;
        RECT 76.815 199.255 82.325 200.065 ;
        RECT 82.335 199.255 87.845 200.065 ;
        RECT 87.855 199.255 89.225 200.065 ;
        RECT 89.235 199.255 90.605 200.065 ;
        RECT 12.095 199.045 12.265 199.255 ;
        RECT 13.475 199.045 13.645 199.255 ;
        RECT 18.995 199.045 19.165 199.255 ;
        RECT 24.515 199.205 24.685 199.235 ;
        RECT 24.510 199.095 24.685 199.205 ;
        RECT 24.515 199.045 24.685 199.095 ;
        RECT 25.435 199.065 25.605 199.255 ;
        RECT 30.035 199.045 30.205 199.235 ;
        RECT 30.955 199.065 31.125 199.255 ;
        RECT 35.555 199.045 35.725 199.235 ;
        RECT 36.475 199.065 36.645 199.255 ;
        RECT 37.390 199.095 37.510 199.205 ;
        RECT 38.315 199.045 38.485 199.255 ;
        RECT 41.990 199.045 42.160 199.235 ;
        RECT 42.455 199.045 42.625 199.235 ;
        RECT 43.835 199.065 44.005 199.255 ;
        RECT 44.755 199.045 44.925 199.235 ;
        RECT 49.355 199.065 49.525 199.255 ;
        RECT 51.195 199.065 51.365 199.255 ;
        RECT 52.115 199.045 52.285 199.235 ;
        RECT 55.795 199.045 55.965 199.235 ;
        RECT 58.555 199.065 58.725 199.255 ;
        RECT 59.015 199.065 59.185 199.255 ;
        RECT 61.775 199.065 61.945 199.255 ;
        RECT 63.150 199.095 63.270 199.205 ;
        RECT 64.075 199.045 64.245 199.255 ;
        RECT 65.910 199.095 66.030 199.205 ;
        RECT 69.595 199.065 69.765 199.255 ;
        RECT 72.355 199.065 72.525 199.255 ;
        RECT 72.815 199.065 72.985 199.255 ;
        RECT 73.275 199.045 73.445 199.235 ;
        RECT 73.735 199.045 73.905 199.235 ;
        RECT 76.955 199.065 77.125 199.255 ;
        RECT 79.255 199.045 79.425 199.235 ;
        RECT 82.475 199.065 82.645 199.255 ;
        RECT 84.775 199.045 84.945 199.235 ;
        RECT 87.995 199.065 88.165 199.255 ;
        RECT 88.465 199.090 88.625 199.200 ;
        RECT 90.295 199.045 90.465 199.255 ;
        RECT 112.465 199.225 113.365 200.135 ;
        RECT 11.955 198.235 13.325 199.045 ;
        RECT 13.335 198.235 18.845 199.045 ;
        RECT 18.855 198.235 24.365 199.045 ;
        RECT 24.375 198.235 29.885 199.045 ;
        RECT 29.895 198.235 35.405 199.045 ;
        RECT 35.415 198.235 37.245 199.045 ;
        RECT 37.725 198.175 38.155 198.960 ;
        RECT 38.175 198.235 40.925 199.045 ;
        RECT 40.955 198.135 42.305 199.045 ;
        RECT 42.315 198.365 44.605 199.045 ;
        RECT 44.615 198.365 51.925 199.045 ;
        RECT 43.685 198.135 44.605 198.365 ;
        RECT 48.130 198.145 49.040 198.365 ;
        RECT 50.575 198.135 51.925 198.365 ;
        RECT 51.975 198.235 55.645 199.045 ;
        RECT 55.655 198.365 62.965 199.045 ;
        RECT 59.170 198.145 60.080 198.365 ;
        RECT 61.615 198.135 62.965 198.365 ;
        RECT 63.485 198.175 63.915 198.960 ;
        RECT 63.935 198.235 65.765 199.045 ;
        RECT 66.275 198.365 73.585 199.045 ;
        RECT 66.275 198.135 67.625 198.365 ;
        RECT 69.160 198.145 70.070 198.365 ;
        RECT 73.595 198.235 79.105 199.045 ;
        RECT 79.115 198.235 84.625 199.045 ;
        RECT 84.635 198.235 88.305 199.045 ;
        RECT 89.235 198.235 90.605 199.045 ;
      LAYER nwell ;
        RECT 11.760 195.015 90.800 197.845 ;
      LAYER pwell ;
        RECT 112.465 197.690 113.145 199.225 ;
        RECT 112.465 196.340 113.375 197.690 ;
        RECT 112.465 194.945 113.375 196.290 ;
        RECT 112.465 194.770 113.145 194.945 ;
        RECT 11.955 193.815 13.325 194.625 ;
        RECT 13.335 193.815 18.845 194.625 ;
        RECT 18.855 193.815 24.365 194.625 ;
        RECT 24.845 193.900 25.275 194.685 ;
        RECT 25.295 193.815 30.805 194.625 ;
        RECT 30.815 193.815 36.325 194.625 ;
        RECT 40.310 194.495 41.220 194.715 ;
        RECT 42.755 194.495 44.105 194.725 ;
        RECT 36.795 193.815 44.105 194.495 ;
        RECT 44.615 194.495 45.535 194.725 ;
        RECT 44.615 193.815 46.905 194.495 ;
        RECT 46.915 193.815 48.265 194.725 ;
        RECT 49.665 194.495 50.585 194.725 ;
        RECT 48.295 193.815 50.585 194.495 ;
        RECT 50.605 193.900 51.035 194.685 ;
        RECT 54.570 194.495 55.480 194.715 ;
        RECT 57.015 194.495 58.365 194.725 ;
        RECT 51.055 193.815 58.365 194.495 ;
        RECT 59.355 193.815 60.705 194.725 ;
        RECT 61.655 193.815 63.005 194.725 ;
        RECT 63.015 193.815 64.385 194.625 ;
        RECT 64.415 193.815 65.765 194.725 ;
        RECT 67.145 194.495 68.065 194.725 ;
        RECT 65.775 193.815 68.065 194.495 ;
        RECT 69.035 194.495 70.385 194.725 ;
        RECT 71.920 194.495 72.830 194.715 ;
        RECT 69.035 193.815 76.345 194.495 ;
        RECT 76.365 193.900 76.795 194.685 ;
        RECT 76.815 193.815 82.325 194.625 ;
        RECT 82.335 193.815 87.845 194.625 ;
        RECT 87.855 193.815 89.225 194.625 ;
        RECT 89.235 193.815 90.605 194.625 ;
        RECT 112.275 194.600 113.145 194.770 ;
        RECT 112.465 194.460 113.145 194.600 ;
        RECT 112.310 194.140 112.420 194.300 ;
        RECT 12.095 193.605 12.265 193.815 ;
        RECT 13.475 193.605 13.645 193.815 ;
        RECT 18.995 193.605 19.165 193.815 ;
        RECT 24.515 193.765 24.685 193.795 ;
        RECT 24.510 193.655 24.685 193.765 ;
        RECT 24.515 193.605 24.685 193.655 ;
        RECT 25.435 193.625 25.605 193.815 ;
        RECT 30.035 193.605 30.205 193.795 ;
        RECT 30.955 193.625 31.125 193.815 ;
        RECT 35.555 193.605 35.725 193.795 ;
        RECT 36.470 193.655 36.590 193.765 ;
        RECT 36.935 193.625 37.105 193.815 ;
        RECT 37.390 193.655 37.510 193.765 ;
        RECT 38.315 193.605 38.485 193.795 ;
        RECT 41.535 193.605 41.705 193.795 ;
        RECT 42.000 193.605 42.170 193.795 ;
        RECT 43.375 193.605 43.545 193.795 ;
        RECT 44.290 193.655 44.410 193.765 ;
        RECT 46.595 193.605 46.765 193.815 ;
        RECT 47.060 193.625 47.230 193.815 ;
        RECT 48.435 193.625 48.605 193.815 ;
        RECT 51.195 193.605 51.365 193.815 ;
        RECT 51.655 193.605 51.825 193.795 ;
        RECT 57.175 193.605 57.345 193.795 ;
        RECT 58.565 193.660 58.725 193.770 ;
        RECT 60.390 193.625 60.560 193.815 ;
        RECT 60.865 193.660 61.025 193.770 ;
        RECT 62.690 193.625 62.860 193.815 ;
        RECT 63.155 193.605 63.325 193.815 ;
        RECT 64.075 193.605 64.245 193.795 ;
        RECT 65.450 193.625 65.620 193.815 ;
        RECT 65.915 193.625 66.085 193.815 ;
        RECT 67.295 193.605 67.465 193.795 ;
        RECT 68.225 193.660 68.385 193.770 ;
        RECT 69.135 193.605 69.305 193.795 ;
        RECT 72.355 193.625 72.525 193.795 ;
        RECT 72.360 193.605 72.525 193.625 ;
        RECT 74.655 193.605 74.825 193.795 ;
        RECT 76.035 193.625 76.205 193.815 ;
        RECT 76.955 193.625 77.125 193.815 ;
        RECT 80.175 193.605 80.345 193.795 ;
        RECT 82.475 193.625 82.645 193.815 ;
        RECT 85.695 193.605 85.865 193.795 ;
        RECT 87.995 193.625 88.165 193.815 ;
        RECT 90.295 193.605 90.465 193.815 ;
        RECT 11.955 192.795 13.325 193.605 ;
        RECT 13.335 192.795 18.845 193.605 ;
        RECT 18.855 192.795 24.365 193.605 ;
        RECT 24.375 192.795 29.885 193.605 ;
        RECT 29.895 192.795 35.405 193.605 ;
        RECT 35.415 192.795 37.245 193.605 ;
        RECT 37.725 192.735 38.155 193.520 ;
        RECT 38.175 192.795 39.545 193.605 ;
        RECT 39.555 192.925 41.845 193.605 ;
        RECT 39.555 192.695 40.475 192.925 ;
        RECT 41.855 192.695 43.205 193.605 ;
        RECT 43.235 192.925 46.445 193.605 ;
        RECT 45.310 192.695 46.445 192.925 ;
        RECT 46.470 192.695 48.285 193.605 ;
        RECT 48.295 192.695 51.465 193.605 ;
        RECT 51.515 192.795 57.025 193.605 ;
        RECT 57.035 192.795 60.705 193.605 ;
        RECT 60.725 192.925 63.465 193.605 ;
        RECT 63.485 192.735 63.915 193.520 ;
        RECT 63.935 192.925 67.145 193.605 ;
        RECT 66.010 192.695 67.145 192.925 ;
        RECT 67.170 192.695 68.985 193.605 ;
        RECT 68.995 192.925 72.205 193.605 ;
        RECT 72.360 192.925 74.195 193.605 ;
        RECT 71.070 192.695 72.205 192.925 ;
        RECT 73.265 192.695 74.195 192.925 ;
        RECT 74.515 192.795 80.025 193.605 ;
        RECT 80.035 192.795 85.545 193.605 ;
        RECT 85.555 192.795 89.225 193.605 ;
        RECT 89.235 192.795 90.605 193.605 ;
        RECT 112.550 193.090 113.335 193.520 ;
        RECT 112.310 192.760 112.420 192.920 ;
      LAYER nwell ;
        RECT 11.760 189.575 90.800 192.405 ;
      LAYER pwell ;
        RECT 112.465 192.010 113.145 192.150 ;
        RECT 112.275 191.840 113.145 192.010 ;
        RECT 112.465 191.665 113.145 191.840 ;
        RECT 112.465 190.320 113.375 191.665 ;
        RECT 11.955 188.375 13.325 189.185 ;
        RECT 13.335 188.375 18.845 189.185 ;
        RECT 18.855 188.375 24.365 189.185 ;
        RECT 24.845 188.460 25.275 189.245 ;
        RECT 25.295 188.375 30.805 189.185 ;
        RECT 30.815 188.375 36.325 189.185 ;
        RECT 36.335 188.375 40.005 189.185 ;
        RECT 40.015 189.055 40.935 189.285 ;
        RECT 40.015 188.375 42.305 189.055 ;
        RECT 42.315 188.375 47.825 189.185 ;
        RECT 47.835 188.375 50.585 189.185 ;
        RECT 50.605 188.460 51.035 189.245 ;
        RECT 51.055 188.375 54.725 189.185 ;
        RECT 55.655 188.375 57.470 189.285 ;
        RECT 57.495 188.375 60.705 189.285 ;
        RECT 60.715 188.375 63.465 189.285 ;
        RECT 63.935 189.055 64.855 189.285 ;
        RECT 63.935 188.375 66.225 189.055 ;
        RECT 66.235 188.375 68.985 189.185 ;
        RECT 69.475 188.375 70.825 189.285 ;
        RECT 112.465 189.260 113.245 190.310 ;
        RECT 70.835 188.375 76.345 189.185 ;
        RECT 76.365 188.460 76.795 189.245 ;
        RECT 76.815 188.375 82.325 189.185 ;
        RECT 82.335 188.375 87.845 189.185 ;
        RECT 87.855 188.375 89.225 189.185 ;
        RECT 89.235 188.375 90.605 189.185 ;
        RECT 112.275 189.090 113.245 189.260 ;
        RECT 112.465 188.940 113.245 189.090 ;
        RECT 112.310 188.620 112.420 188.780 ;
        RECT 12.095 188.165 12.265 188.375 ;
        RECT 13.475 188.165 13.645 188.375 ;
        RECT 18.995 188.165 19.165 188.375 ;
        RECT 22.215 188.165 22.385 188.355 ;
        RECT 22.675 188.165 22.845 188.355 ;
        RECT 24.510 188.215 24.630 188.325 ;
        RECT 25.435 188.185 25.605 188.375 ;
        RECT 26.355 188.165 26.525 188.355 ;
        RECT 30.955 188.185 31.125 188.375 ;
        RECT 33.715 188.165 33.885 188.355 ;
        RECT 36.475 188.185 36.645 188.375 ;
        RECT 37.390 188.215 37.510 188.325 ;
        RECT 38.315 188.165 38.485 188.355 ;
        RECT 41.995 188.185 42.165 188.375 ;
        RECT 42.455 188.185 42.625 188.375 ;
        RECT 45.675 188.165 45.845 188.355 ;
        RECT 47.975 188.185 48.145 188.375 ;
        RECT 51.195 188.165 51.365 188.375 ;
        RECT 54.885 188.325 55.045 188.330 ;
        RECT 54.870 188.220 55.045 188.325 ;
        RECT 54.870 188.215 54.990 188.220 ;
        RECT 56.715 188.165 56.885 188.355 ;
        RECT 57.175 188.165 57.345 188.375 ;
        RECT 57.635 188.185 57.805 188.375 ;
        RECT 59.010 188.215 59.130 188.325 ;
        RECT 59.480 188.165 59.650 188.355 ;
        RECT 60.855 188.185 61.025 188.375 ;
        RECT 61.315 188.165 61.485 188.355 ;
        RECT 63.150 188.215 63.270 188.325 ;
        RECT 63.610 188.215 63.730 188.325 ;
        RECT 64.075 188.165 64.245 188.355 ;
        RECT 65.915 188.185 66.085 188.375 ;
        RECT 66.375 188.185 66.545 188.375 ;
        RECT 69.590 188.355 69.760 188.375 ;
        RECT 69.130 188.215 69.250 188.325 ;
        RECT 69.590 188.185 69.765 188.355 ;
        RECT 70.975 188.185 71.145 188.375 ;
        RECT 69.595 188.165 69.765 188.185 ;
        RECT 75.115 188.165 75.285 188.355 ;
        RECT 76.955 188.185 77.125 188.375 ;
        RECT 80.635 188.165 80.805 188.355 ;
        RECT 82.475 188.185 82.645 188.375 ;
        RECT 86.155 188.165 86.325 188.355 ;
        RECT 87.995 188.185 88.165 188.375 ;
        RECT 88.910 188.215 89.030 188.325 ;
        RECT 90.295 188.165 90.465 188.375 ;
        RECT 11.955 187.355 13.325 188.165 ;
        RECT 13.335 187.355 18.845 188.165 ;
        RECT 18.855 187.355 20.225 188.165 ;
        RECT 20.235 187.485 22.525 188.165 ;
        RECT 20.235 187.255 21.155 187.485 ;
        RECT 22.535 187.355 26.205 188.165 ;
        RECT 26.215 187.485 33.525 188.165 ;
        RECT 29.730 187.265 30.640 187.485 ;
        RECT 32.175 187.255 33.525 187.485 ;
        RECT 33.575 187.355 37.245 188.165 ;
        RECT 37.725 187.295 38.155 188.080 ;
        RECT 38.175 187.485 45.485 188.165 ;
        RECT 41.690 187.265 42.600 187.485 ;
        RECT 44.135 187.255 45.485 187.485 ;
        RECT 45.535 187.355 51.045 188.165 ;
        RECT 51.055 187.355 54.725 188.165 ;
        RECT 55.195 187.255 57.010 188.165 ;
        RECT 57.035 187.355 58.865 188.165 ;
        RECT 59.335 187.255 61.165 188.165 ;
        RECT 61.175 187.355 63.005 188.165 ;
        RECT 63.485 187.295 63.915 188.080 ;
        RECT 63.935 187.355 69.445 188.165 ;
        RECT 69.455 187.355 74.965 188.165 ;
        RECT 74.975 187.355 80.485 188.165 ;
        RECT 80.495 187.355 86.005 188.165 ;
        RECT 86.015 187.355 88.765 188.165 ;
        RECT 89.235 187.355 90.605 188.165 ;
        RECT 112.465 187.870 113.145 188.010 ;
        RECT 112.275 187.700 113.145 187.870 ;
      LAYER nwell ;
        RECT 11.760 184.135 90.800 186.965 ;
      LAYER pwell ;
        RECT 112.465 186.190 113.145 187.700 ;
        RECT 112.465 185.260 113.375 186.190 ;
        RECT 112.305 184.995 112.415 185.115 ;
        RECT 11.955 182.935 13.325 183.745 ;
        RECT 13.335 182.935 16.085 183.745 ;
        RECT 16.115 182.935 17.465 183.845 ;
        RECT 17.515 183.615 18.865 183.845 ;
        RECT 20.400 183.615 21.310 183.835 ;
        RECT 17.515 182.935 24.825 183.615 ;
        RECT 24.845 183.020 25.275 183.805 ;
        RECT 26.215 183.615 27.135 183.845 ;
        RECT 26.215 182.935 28.505 183.615 ;
        RECT 28.515 182.935 31.435 183.845 ;
        RECT 31.745 182.935 34.475 183.845 ;
        RECT 34.695 183.755 35.645 183.845 ;
        RECT 34.695 182.935 36.625 183.755 ;
        RECT 36.795 182.935 38.625 183.845 ;
        RECT 38.675 182.935 41.845 183.845 ;
        RECT 41.855 182.935 45.525 183.745 ;
        RECT 45.535 182.935 47.365 183.615 ;
        RECT 47.375 182.935 50.125 183.745 ;
        RECT 50.605 183.020 51.035 183.805 ;
        RECT 51.065 182.935 53.795 183.845 ;
        RECT 53.815 182.935 57.485 183.745 ;
        RECT 57.955 182.935 61.615 183.845 ;
        RECT 61.835 183.755 62.785 183.845 ;
        RECT 61.835 182.935 63.765 183.755 ;
        RECT 63.945 182.935 65.295 183.845 ;
        RECT 65.775 183.645 66.705 183.845 ;
        RECT 68.035 183.645 68.985 183.845 ;
        RECT 65.775 183.165 68.985 183.645 ;
        RECT 65.920 182.965 68.985 183.165 ;
        RECT 12.095 182.725 12.265 182.935 ;
        RECT 13.475 182.725 13.645 182.935 ;
        RECT 16.230 182.745 16.400 182.935 ;
        RECT 18.995 182.725 19.165 182.915 ;
        RECT 22.675 182.745 22.845 182.915 ;
        RECT 22.675 182.725 22.840 182.745 ;
        RECT 23.135 182.725 23.305 182.915 ;
        RECT 24.515 182.745 24.685 182.935 ;
        RECT 25.445 182.780 25.605 182.890 ;
        RECT 28.195 182.745 28.365 182.935 ;
        RECT 28.660 182.885 28.830 182.935 ;
        RECT 28.650 182.775 28.830 182.885 ;
        RECT 28.660 182.745 28.830 182.775 ;
        RECT 31.875 182.725 32.045 182.935 ;
        RECT 36.475 182.915 36.625 182.935 ;
        RECT 32.330 182.775 32.450 182.885 ;
        RECT 32.795 182.725 32.965 182.915 ;
        RECT 36.015 182.725 36.185 182.915 ;
        RECT 36.475 182.745 36.645 182.915 ;
        RECT 38.310 182.880 38.480 182.935 ;
        RECT 38.310 182.770 38.485 182.880 ;
        RECT 38.310 182.745 38.480 182.770 ;
        RECT 38.775 182.745 38.945 182.935 ;
        RECT 39.235 182.725 39.405 182.915 ;
        RECT 41.995 182.745 42.165 182.935 ;
        RECT 43.380 182.725 43.550 182.915 ;
        RECT 43.835 182.745 44.005 182.915 ;
        RECT 43.840 182.725 44.005 182.745 ;
        RECT 46.135 182.725 46.305 182.915 ;
        RECT 47.055 182.745 47.225 182.935 ;
        RECT 47.515 182.745 47.685 182.935 ;
        RECT 49.820 182.725 49.990 182.915 ;
        RECT 50.270 182.775 50.390 182.885 ;
        RECT 51.195 182.745 51.365 182.935 ;
        RECT 53.955 182.745 54.125 182.935 ;
        RECT 55.790 182.725 55.960 182.915 ;
        RECT 56.255 182.725 56.425 182.915 ;
        RECT 57.630 182.775 57.750 182.885 ;
        RECT 59.930 182.775 60.050 182.885 ;
        RECT 11.955 181.915 13.325 182.725 ;
        RECT 13.335 181.915 18.845 182.725 ;
        RECT 18.855 181.915 20.685 182.725 ;
        RECT 21.005 182.045 22.840 182.725 ;
        RECT 21.005 181.815 21.935 182.045 ;
        RECT 22.995 181.915 28.505 182.725 ;
        RECT 28.975 182.045 32.185 182.725 ;
        RECT 28.975 181.815 30.110 182.045 ;
        RECT 32.735 181.815 35.735 182.725 ;
        RECT 35.875 181.915 37.705 182.725 ;
        RECT 37.725 181.855 38.155 182.640 ;
        RECT 39.195 181.815 42.305 182.725 ;
        RECT 42.315 181.815 43.665 182.725 ;
        RECT 43.840 182.045 45.675 182.725 ;
        RECT 45.995 182.045 49.665 182.725 ;
        RECT 44.745 181.815 45.675 182.045 ;
        RECT 48.735 181.815 49.665 182.045 ;
        RECT 49.675 181.815 51.505 182.725 ;
        RECT 51.715 181.815 56.105 182.725 ;
        RECT 56.115 181.815 59.785 182.725 ;
        RECT 60.395 182.695 60.565 182.915 ;
        RECT 61.320 182.745 61.490 182.935 ;
        RECT 63.615 182.915 63.765 182.935 ;
        RECT 63.615 182.745 63.785 182.915 ;
        RECT 64.075 182.745 64.245 182.935 ;
        RECT 65.450 182.775 65.570 182.885 ;
        RECT 65.920 182.745 66.090 182.965 ;
        RECT 68.050 182.935 68.985 182.965 ;
        RECT 69.035 183.615 70.385 183.845 ;
        RECT 71.920 183.615 72.830 183.835 ;
        RECT 69.035 182.935 76.345 183.615 ;
        RECT 76.365 183.020 76.795 183.805 ;
        RECT 76.815 182.935 82.325 183.745 ;
        RECT 82.335 182.935 87.845 183.745 ;
        RECT 87.855 182.935 89.225 183.745 ;
        RECT 89.235 182.935 90.605 183.745 ;
        RECT 112.465 183.730 113.275 184.790 ;
        RECT 112.275 183.560 113.275 183.730 ;
        RECT 112.465 183.420 113.275 183.560 ;
      LAYER nwell ;
        RECT 113.665 183.225 116.495 219.485 ;
      LAYER pwell ;
        RECT 116.885 219.150 117.695 219.290 ;
        RECT 117.905 219.150 118.715 219.290 ;
        RECT 116.885 218.980 118.715 219.150 ;
        RECT 116.885 217.920 117.695 218.980 ;
        RECT 117.905 217.920 118.715 218.980 ;
        RECT 116.785 216.565 117.695 217.910 ;
        RECT 117.015 216.390 117.695 216.565 ;
        RECT 117.905 216.520 118.815 217.870 ;
        RECT 117.015 216.220 117.885 216.390 ;
        RECT 117.015 216.080 117.695 216.220 ;
        RECT 117.740 215.760 117.850 215.920 ;
        RECT 116.785 214.735 117.695 215.150 ;
        RECT 117.905 214.985 118.585 216.520 ;
        RECT 116.785 214.565 117.885 214.735 ;
        RECT 116.785 214.220 117.695 214.565 ;
        RECT 117.015 211.250 117.695 214.220 ;
        RECT 117.905 214.075 118.805 214.985 ;
        RECT 116.885 210.870 117.695 211.010 ;
        RECT 117.905 210.870 118.585 214.075 ;
        RECT 116.885 210.700 118.585 210.870 ;
        RECT 116.885 207.340 117.695 210.700 ;
        RECT 117.905 210.560 118.585 210.700 ;
        RECT 117.905 210.410 118.715 210.550 ;
        RECT 117.715 210.240 118.715 210.410 ;
        RECT 116.885 207.190 117.695 207.330 ;
        RECT 116.885 207.020 117.885 207.190 ;
        RECT 116.885 205.960 117.695 207.020 ;
        RECT 117.905 206.880 118.715 210.240 ;
        RECT 117.745 206.615 117.855 206.735 ;
        RECT 117.990 205.970 118.775 206.400 ;
        RECT 116.785 204.560 117.695 205.910 ;
        RECT 117.905 205.810 118.585 205.950 ;
        RECT 117.715 205.640 118.585 205.810 ;
        RECT 117.015 203.025 117.695 204.560 ;
        RECT 116.795 202.115 117.695 203.025 ;
        RECT 117.015 198.910 117.695 202.115 ;
        RECT 117.015 198.740 117.885 198.910 ;
        RECT 117.015 198.600 117.695 198.740 ;
        RECT 116.785 198.175 117.695 198.590 ;
        RECT 116.785 198.005 117.885 198.175 ;
        RECT 116.785 197.660 117.695 198.005 ;
        RECT 117.015 194.690 117.695 197.660 ;
        RECT 117.905 196.845 118.585 205.640 ;
        RECT 117.905 196.610 118.715 196.750 ;
        RECT 117.715 196.440 118.715 196.610 ;
        RECT 117.905 195.380 118.715 196.440 ;
        RECT 117.905 195.230 118.685 195.370 ;
        RECT 117.715 195.060 118.685 195.230 ;
        RECT 117.740 194.140 117.850 194.300 ;
        RECT 117.905 194.000 118.685 195.060 ;
        RECT 117.905 193.850 118.685 193.990 ;
        RECT 117.715 193.680 118.685 193.850 ;
        RECT 116.825 193.090 117.610 193.520 ;
        RECT 116.785 192.055 117.695 192.975 ;
        RECT 117.905 192.620 118.685 193.680 ;
        RECT 117.905 192.470 118.685 192.610 ;
        RECT 117.715 192.300 118.685 192.470 ;
        RECT 117.015 189.710 117.695 192.055 ;
        RECT 117.905 191.240 118.685 192.300 ;
        RECT 117.905 191.090 118.685 191.230 ;
        RECT 117.715 190.920 118.685 191.090 ;
        RECT 117.905 189.860 118.685 190.920 ;
        RECT 117.015 189.540 117.885 189.710 ;
        RECT 117.015 189.510 117.695 189.540 ;
        RECT 117.740 189.080 117.850 189.240 ;
        RECT 117.905 188.795 118.815 189.830 ;
        RECT 117.715 188.625 118.815 188.795 ;
        RECT 117.905 188.480 118.815 188.625 ;
        RECT 116.785 186.030 117.695 188.470 ;
        RECT 117.905 188.330 118.815 188.390 ;
        RECT 117.715 188.160 118.815 188.330 ;
        RECT 116.785 185.860 117.885 186.030 ;
        RECT 116.785 185.720 117.695 185.860 ;
        RECT 117.740 185.400 117.850 185.560 ;
        RECT 117.905 184.940 118.815 188.160 ;
        RECT 116.885 183.730 117.695 184.790 ;
        RECT 117.905 183.730 118.715 184.790 ;
        RECT 116.885 183.560 118.715 183.730 ;
        RECT 116.885 183.420 117.695 183.560 ;
        RECT 117.905 183.420 118.715 183.560 ;
      LAYER nwell ;
        RECT 119.105 183.225 121.935 219.485 ;
      LAYER pwell ;
        RECT 122.325 219.150 123.135 219.290 ;
        RECT 123.345 219.150 124.155 219.290 ;
        RECT 122.325 218.980 124.155 219.150 ;
        RECT 122.325 217.920 123.135 218.980 ;
        RECT 123.345 217.920 124.155 218.980 ;
        RECT 122.225 216.565 123.135 217.910 ;
        RECT 123.345 217.770 124.025 217.910 ;
        RECT 123.155 217.600 124.025 217.770 ;
        RECT 122.455 216.390 123.135 216.565 ;
        RECT 122.455 216.220 123.325 216.390 ;
        RECT 122.455 216.080 123.135 216.220 ;
        RECT 123.180 215.760 123.290 215.920 ;
        RECT 122.455 215.010 123.135 215.040 ;
        RECT 122.455 214.840 123.325 215.010 ;
        RECT 122.455 212.495 123.135 214.840 ;
        RECT 122.225 211.575 123.135 212.495 ;
        RECT 123.345 214.395 124.025 217.600 ;
        RECT 123.345 213.485 124.245 214.395 ;
        RECT 123.345 211.950 124.025 213.485 ;
        RECT 123.180 211.160 123.290 211.320 ;
        RECT 123.345 210.600 124.255 211.950 ;
        RECT 122.455 210.410 123.135 210.440 ;
        RECT 123.345 210.410 124.155 210.550 ;
        RECT 122.455 210.240 124.155 210.410 ;
        RECT 122.455 207.895 123.135 210.240 ;
        RECT 122.225 206.975 123.135 207.895 ;
        RECT 123.345 206.880 124.155 210.240 ;
        RECT 122.455 203.670 123.135 206.640 ;
        RECT 123.185 206.615 123.295 206.735 ;
        RECT 123.430 205.970 124.215 206.400 ;
        RECT 123.345 205.810 124.025 205.950 ;
        RECT 123.155 205.640 124.025 205.810 ;
        RECT 122.225 203.325 123.135 203.670 ;
        RECT 122.225 203.155 123.325 203.325 ;
        RECT 122.225 202.740 123.135 203.155 ;
        RECT 122.325 202.590 123.135 202.730 ;
        RECT 122.325 202.420 123.325 202.590 ;
        RECT 123.345 202.435 124.025 205.640 ;
        RECT 122.325 200.900 123.135 202.420 ;
        RECT 123.345 201.525 124.245 202.435 ;
        RECT 122.455 200.750 123.135 200.890 ;
        RECT 122.455 200.580 123.325 200.750 ;
        RECT 122.455 197.375 123.135 200.580 ;
        RECT 123.345 199.990 124.025 201.525 ;
        RECT 123.345 198.640 124.255 199.990 ;
        RECT 123.345 198.445 124.025 198.590 ;
        RECT 123.155 198.275 124.025 198.445 ;
        RECT 122.235 196.465 123.135 197.375 ;
        RECT 122.455 194.930 123.135 196.465 ;
        RECT 123.345 196.745 124.025 198.275 ;
        RECT 123.345 195.380 124.255 196.745 ;
        RECT 123.345 195.230 124.155 195.370 ;
        RECT 123.155 195.060 124.155 195.230 ;
        RECT 122.225 193.580 123.135 194.930 ;
        RECT 122.265 193.090 123.050 193.520 ;
        RECT 122.225 192.655 123.135 193.070 ;
        RECT 122.225 192.485 123.325 192.655 ;
        RECT 123.345 192.620 124.155 195.060 ;
        RECT 122.225 192.140 123.135 192.485 ;
        RECT 123.185 192.355 123.295 192.475 ;
        RECT 122.455 189.170 123.135 192.140 ;
        RECT 123.345 192.010 124.025 192.040 ;
        RECT 123.155 191.840 124.025 192.010 ;
        RECT 123.345 189.495 124.025 191.840 ;
        RECT 122.355 188.790 123.135 188.930 ;
        RECT 122.355 188.620 123.325 188.790 ;
        RECT 122.355 187.560 123.135 188.620 ;
        RECT 123.345 188.575 124.255 189.495 ;
        RECT 123.345 188.330 124.255 188.390 ;
        RECT 123.155 188.160 124.255 188.330 ;
        RECT 122.225 186.605 123.135 187.550 ;
        RECT 122.425 185.115 123.105 186.605 ;
        RECT 123.345 185.390 124.255 188.160 ;
        RECT 122.425 184.945 123.325 185.115 ;
        RECT 122.425 184.800 123.105 184.945 ;
        RECT 122.325 183.730 123.135 184.790 ;
        RECT 123.345 183.730 124.155 184.790 ;
        RECT 122.325 183.560 124.155 183.730 ;
        RECT 122.325 183.420 123.135 183.560 ;
        RECT 123.345 183.420 124.155 183.560 ;
      LAYER nwell ;
        RECT 124.545 183.225 127.375 219.485 ;
      LAYER pwell ;
        RECT 127.765 219.150 128.575 219.290 ;
        RECT 128.785 219.150 129.595 219.290 ;
        RECT 127.765 218.980 129.595 219.150 ;
        RECT 127.765 217.920 128.575 218.980 ;
        RECT 128.785 217.920 129.595 218.980 ;
        RECT 127.665 216.565 128.575 217.910 ;
        RECT 128.785 217.770 129.595 217.910 ;
        RECT 128.595 217.600 129.595 217.770 ;
        RECT 127.895 216.390 128.575 216.565 ;
        RECT 128.785 216.540 129.595 217.600 ;
        RECT 128.785 216.390 129.465 216.420 ;
        RECT 127.895 216.220 129.465 216.390 ;
        RECT 127.895 216.080 128.575 216.220 ;
        RECT 128.625 215.815 128.735 215.935 ;
        RECT 127.665 215.195 128.575 215.610 ;
        RECT 127.665 215.025 128.765 215.195 ;
        RECT 127.665 214.680 128.575 215.025 ;
        RECT 127.895 211.710 128.575 214.680 ;
        RECT 128.785 213.875 129.465 216.220 ;
        RECT 128.785 212.955 129.695 213.875 ;
        RECT 128.785 211.835 129.695 212.755 ;
        RECT 127.895 211.330 128.575 211.470 ;
        RECT 127.895 211.160 128.765 211.330 ;
        RECT 127.895 207.955 128.575 211.160 ;
        RECT 128.785 209.490 129.465 211.835 ;
        RECT 128.595 209.320 129.465 209.490 ;
        RECT 128.785 209.290 129.465 209.320 ;
        RECT 128.785 209.030 129.595 209.170 ;
        RECT 128.595 208.860 129.595 209.030 ;
        RECT 127.675 207.045 128.575 207.955 ;
        RECT 127.895 205.510 128.575 207.045 ;
        RECT 128.785 206.420 129.595 208.860 ;
        RECT 128.870 205.970 129.655 206.400 ;
        RECT 127.665 204.160 128.575 205.510 ;
        RECT 128.785 204.895 129.695 205.930 ;
        RECT 128.595 204.725 129.695 204.895 ;
        RECT 128.785 204.580 129.695 204.725 ;
        RECT 127.665 203.695 128.575 204.110 ;
        RECT 127.665 203.525 128.765 203.695 ;
        RECT 127.665 203.180 128.575 203.525 ;
        RECT 127.895 200.210 128.575 203.180 ;
        RECT 128.785 200.750 129.695 204.500 ;
        RECT 128.595 200.580 129.695 200.750 ;
        RECT 128.785 200.440 129.695 200.580 ;
        RECT 127.665 198.955 128.575 199.875 ;
        RECT 127.895 196.610 128.575 198.955 ;
        RECT 128.785 199.415 129.695 200.335 ;
        RECT 128.785 197.070 129.465 199.415 ;
        RECT 128.595 196.900 129.465 197.070 ;
        RECT 128.785 196.870 129.465 196.900 ;
        RECT 128.785 196.610 129.595 196.750 ;
        RECT 127.895 196.440 129.595 196.610 ;
        RECT 127.895 196.410 128.575 196.440 ;
        RECT 127.765 196.150 128.575 196.290 ;
        RECT 127.765 195.980 128.765 196.150 ;
        RECT 127.765 193.540 128.575 195.980 ;
        RECT 128.785 195.380 129.595 196.440 ;
        RECT 128.785 194.420 129.695 195.370 ;
        RECT 127.705 193.090 128.490 193.520 ;
        RECT 127.665 190.175 128.575 192.780 ;
        RECT 128.815 192.015 129.495 194.420 ;
        RECT 128.595 191.845 129.495 192.015 ;
        RECT 128.815 191.700 129.495 191.845 ;
        RECT 128.785 191.545 129.695 191.690 ;
        RECT 128.595 191.375 129.695 191.545 ;
        RECT 128.785 190.340 129.695 191.375 ;
        RECT 127.665 190.160 128.765 190.175 ;
        RECT 128.785 190.160 129.565 190.310 ;
        RECT 127.665 190.005 129.565 190.160 ;
        RECT 127.665 189.860 128.575 190.005 ;
        RECT 128.595 189.990 129.565 190.005 ;
        RECT 128.620 189.540 128.730 189.700 ;
        RECT 128.785 188.940 129.565 189.990 ;
        RECT 127.665 185.570 128.575 188.790 ;
        RECT 128.785 185.570 129.695 188.790 ;
        RECT 127.665 185.400 129.695 185.570 ;
        RECT 127.665 185.340 128.575 185.400 ;
        RECT 128.785 185.340 129.695 185.400 ;
        RECT 128.625 184.995 128.735 185.115 ;
        RECT 127.765 183.730 128.575 184.790 ;
        RECT 128.785 183.730 129.595 184.790 ;
        RECT 127.765 183.560 129.595 183.730 ;
        RECT 127.765 183.420 128.575 183.560 ;
        RECT 128.785 183.420 129.595 183.560 ;
      LAYER nwell ;
        RECT 129.985 183.225 132.815 219.485 ;
      LAYER pwell ;
        RECT 133.205 219.150 134.015 219.290 ;
        RECT 134.225 219.150 135.035 219.290 ;
        RECT 133.205 218.980 135.035 219.150 ;
        RECT 133.205 217.920 134.015 218.980 ;
        RECT 134.225 217.920 135.035 218.980 ;
        RECT 133.105 216.520 134.015 217.870 ;
        RECT 134.225 217.495 135.135 217.910 ;
        RECT 134.035 217.325 135.135 217.495 ;
        RECT 133.335 214.985 134.015 216.520 ;
        RECT 133.115 214.075 134.015 214.985 ;
        RECT 133.335 210.870 134.015 214.075 ;
        RECT 134.225 216.980 135.135 217.325 ;
        RECT 134.225 214.010 134.905 216.980 ;
        RECT 134.225 213.630 134.905 213.770 ;
        RECT 134.035 213.460 134.905 213.630 ;
        RECT 133.335 210.700 134.205 210.870 ;
        RECT 133.335 210.560 134.015 210.700 ;
        RECT 133.205 210.410 134.015 210.550 ;
        RECT 133.205 210.240 134.205 210.410 ;
        RECT 134.225 210.255 134.905 213.460 ;
        RECT 133.205 207.800 134.015 210.240 ;
        RECT 134.225 209.345 135.125 210.255 ;
        RECT 134.225 207.810 134.905 209.345 ;
        RECT 134.065 207.535 134.175 207.655 ;
        RECT 133.335 207.190 134.015 207.330 ;
        RECT 133.335 207.020 134.205 207.190 ;
        RECT 133.335 198.225 134.015 207.020 ;
        RECT 134.225 206.460 135.135 207.810 ;
        RECT 134.310 205.970 135.095 206.400 ;
        RECT 134.225 205.810 134.905 205.950 ;
        RECT 134.035 205.640 134.905 205.810 ;
        RECT 134.225 202.435 134.905 205.640 ;
        RECT 134.225 201.525 135.125 202.435 ;
        RECT 134.225 199.990 134.905 201.525 ;
        RECT 134.225 198.640 135.135 199.990 ;
        RECT 134.065 198.335 134.175 198.455 ;
        RECT 133.105 197.115 134.015 198.035 ;
        RECT 133.335 194.770 134.015 197.115 ;
        RECT 134.225 196.765 135.135 198.130 ;
        RECT 134.225 195.235 134.905 196.765 ;
        RECT 134.035 195.065 134.905 195.235 ;
        RECT 134.225 194.920 134.905 195.065 ;
        RECT 133.335 194.600 134.205 194.770 ;
        RECT 133.335 194.570 134.015 194.600 ;
        RECT 134.060 194.140 134.170 194.300 ;
        RECT 134.225 193.850 135.135 193.910 ;
        RECT 134.035 193.680 135.135 193.850 ;
        RECT 133.145 193.090 133.930 193.520 ;
        RECT 133.305 192.935 133.985 193.060 ;
        RECT 133.305 192.765 134.205 192.935 ;
        RECT 133.305 191.735 133.985 192.765 ;
        RECT 133.105 190.780 134.015 191.735 ;
        RECT 134.225 190.910 135.135 193.680 ;
        RECT 133.205 190.630 134.015 190.770 ;
        RECT 133.205 190.625 134.205 190.630 ;
        RECT 134.225 190.625 135.135 190.770 ;
        RECT 133.205 190.460 135.135 190.625 ;
        RECT 133.205 188.020 134.015 190.460 ;
        RECT 134.035 190.455 135.135 190.460 ;
        RECT 134.225 189.420 135.135 190.455 ;
        RECT 134.065 189.135 134.175 189.255 ;
        RECT 134.225 188.790 135.135 188.850 ;
        RECT 134.035 188.620 135.135 188.790 ;
        RECT 134.065 187.755 134.175 187.875 ;
        RECT 133.105 186.495 134.015 187.530 ;
        RECT 133.105 186.325 134.205 186.495 ;
        RECT 133.105 186.180 134.015 186.325 ;
        RECT 133.235 185.110 134.015 186.170 ;
        RECT 134.225 185.400 135.135 188.620 ;
        RECT 134.065 185.110 134.175 185.115 ;
        RECT 133.235 184.940 134.205 185.110 ;
        RECT 133.235 184.800 134.015 184.940 ;
        RECT 133.205 183.730 134.015 184.790 ;
        RECT 134.225 183.730 135.035 184.790 ;
        RECT 133.205 183.560 135.035 183.730 ;
        RECT 133.205 183.420 134.015 183.560 ;
        RECT 134.225 183.420 135.035 183.560 ;
      LAYER nwell ;
        RECT 135.425 183.225 138.255 219.485 ;
      LAYER pwell ;
        RECT 138.645 219.150 139.455 219.290 ;
        RECT 139.665 219.150 140.475 219.290 ;
        RECT 138.645 218.980 140.475 219.150 ;
        RECT 138.645 217.920 139.455 218.980 ;
        RECT 139.665 217.920 140.475 218.980 ;
        RECT 138.545 216.565 139.455 217.910 ;
        RECT 139.665 217.770 140.345 217.910 ;
        RECT 139.475 217.600 140.345 217.770 ;
        RECT 138.775 216.390 139.455 216.565 ;
        RECT 138.775 216.220 139.645 216.390 ;
        RECT 138.775 216.080 139.455 216.220 ;
        RECT 138.545 215.655 139.455 216.070 ;
        RECT 138.545 215.485 139.645 215.655 ;
        RECT 138.545 215.140 139.455 215.485 ;
        RECT 138.775 212.170 139.455 215.140 ;
        RECT 139.665 214.395 140.345 217.600 ;
        RECT 139.665 213.485 140.565 214.395 ;
        RECT 139.665 211.950 140.345 213.485 ;
        RECT 138.645 211.790 139.455 211.930 ;
        RECT 138.645 211.620 139.645 211.790 ;
        RECT 138.645 210.560 139.455 211.620 ;
        RECT 139.665 210.600 140.575 211.950 ;
        RECT 138.775 201.670 139.455 210.465 ;
        RECT 139.665 209.535 140.575 210.455 ;
        RECT 139.665 207.190 140.345 209.535 ;
        RECT 139.475 207.020 140.345 207.190 ;
        RECT 139.665 206.990 140.345 207.020 ;
        RECT 139.505 206.615 139.615 206.735 ;
        RECT 139.750 205.970 140.535 206.400 ;
        RECT 139.665 205.535 140.575 205.950 ;
        RECT 139.475 205.365 140.575 205.535 ;
        RECT 139.665 205.020 140.575 205.365 ;
        RECT 139.665 202.050 140.345 205.020 ;
        RECT 139.505 201.670 139.615 201.675 ;
        RECT 138.775 201.500 139.645 201.670 ;
        RECT 138.775 201.360 139.455 201.500 ;
        RECT 138.545 200.335 139.455 201.255 ;
        RECT 139.475 201.205 139.645 201.210 ;
        RECT 139.475 201.040 140.345 201.205 ;
        RECT 138.775 197.990 139.455 200.335 ;
        RECT 139.665 200.300 140.345 201.040 ;
        RECT 139.665 199.370 140.575 200.300 ;
        RECT 139.665 197.990 140.575 199.040 ;
        RECT 138.775 197.820 140.575 197.990 ;
        RECT 138.775 197.790 139.455 197.820 ;
        RECT 139.665 197.690 140.575 197.820 ;
        RECT 138.645 197.530 139.455 197.670 ;
        RECT 139.665 197.530 140.345 197.670 ;
        RECT 138.645 197.360 140.345 197.530 ;
        RECT 138.645 196.300 139.455 197.360 ;
        RECT 138.745 196.145 139.425 196.290 ;
        RECT 138.745 195.975 139.645 196.145 ;
        RECT 138.745 194.485 139.425 195.975 ;
        RECT 138.545 193.540 139.455 194.485 ;
        RECT 139.665 194.155 140.345 197.360 ;
        RECT 138.585 193.090 139.370 193.520 ;
        RECT 139.665 193.245 140.565 194.155 ;
        RECT 138.545 192.930 139.455 192.990 ;
        RECT 138.545 192.760 139.645 192.930 ;
        RECT 138.545 189.540 139.455 192.760 ;
        RECT 139.665 191.710 140.345 193.245 ;
        RECT 139.665 190.360 140.575 191.710 ;
        RECT 139.505 190.055 139.615 190.175 ;
        RECT 139.475 189.705 139.645 189.710 ;
        RECT 139.475 189.540 140.345 189.705 ;
        RECT 138.545 189.250 139.455 189.310 ;
        RECT 138.545 189.080 139.645 189.250 ;
        RECT 138.545 185.860 139.455 189.080 ;
        RECT 139.665 188.800 140.345 189.540 ;
        RECT 139.665 187.870 140.575 188.800 ;
        RECT 139.665 187.410 140.445 187.550 ;
        RECT 139.475 187.240 140.445 187.410 ;
        RECT 139.665 186.180 140.445 187.240 ;
        RECT 139.500 185.400 139.610 185.560 ;
        RECT 139.665 185.120 140.445 186.170 ;
        RECT 139.475 184.950 140.445 185.120 ;
        RECT 139.665 184.800 140.445 184.950 ;
        RECT 138.645 183.730 139.455 184.790 ;
        RECT 139.665 183.730 140.475 184.790 ;
        RECT 138.645 183.560 140.475 183.730 ;
        RECT 138.645 183.420 139.455 183.560 ;
        RECT 139.665 183.420 140.475 183.560 ;
      LAYER nwell ;
        RECT 140.865 183.225 143.695 219.485 ;
      LAYER pwell ;
        RECT 144.085 219.150 144.895 219.290 ;
        RECT 145.105 219.150 145.915 219.290 ;
        RECT 144.085 218.980 145.915 219.150 ;
        RECT 144.085 217.920 144.895 218.980 ;
        RECT 145.105 217.920 145.915 218.980 ;
        RECT 144.085 217.770 144.895 217.910 ;
        RECT 145.105 217.770 145.915 217.910 ;
        RECT 144.085 217.600 145.915 217.770 ;
        RECT 144.085 214.240 144.895 217.600 ;
        RECT 144.945 213.975 145.055 214.095 ;
        RECT 143.985 212.380 144.895 213.730 ;
        RECT 145.105 212.400 145.915 217.600 ;
        RECT 144.215 210.845 144.895 212.380 ;
        RECT 144.950 212.080 145.060 212.240 ;
        RECT 145.105 211.330 145.785 211.470 ;
        RECT 144.915 211.160 145.785 211.330 ;
        RECT 143.995 209.935 144.895 210.845 ;
        RECT 144.215 206.730 144.895 209.935 ;
        RECT 145.105 210.985 145.785 211.160 ;
        RECT 145.105 209.640 146.015 210.985 ;
        RECT 145.105 206.730 146.015 209.500 ;
        RECT 144.215 206.560 146.015 206.730 ;
        RECT 144.215 206.420 144.895 206.560 ;
        RECT 145.105 206.500 146.015 206.560 ;
        RECT 144.215 206.270 144.895 206.410 ;
        RECT 144.215 206.100 145.085 206.270 ;
        RECT 144.215 202.895 144.895 206.100 ;
        RECT 145.190 205.970 145.975 206.400 ;
        RECT 144.950 205.640 145.060 205.800 ;
        RECT 145.105 204.890 145.785 204.920 ;
        RECT 144.915 204.720 145.785 204.890 ;
        RECT 143.995 201.985 144.895 202.895 ;
        RECT 144.215 200.450 144.895 201.985 ;
        RECT 145.105 202.375 145.785 204.720 ;
        RECT 145.105 201.455 146.015 202.375 ;
        RECT 144.950 201.040 145.060 201.200 ;
        RECT 143.985 199.100 144.895 200.450 ;
        RECT 145.105 199.085 146.015 200.430 ;
        RECT 145.105 198.910 145.785 199.085 ;
        RECT 144.915 198.740 145.785 198.910 ;
        RECT 143.985 197.810 144.895 198.740 ;
        RECT 145.105 198.600 145.785 198.740 ;
        RECT 145.105 198.450 145.785 198.480 ;
        RECT 144.915 198.280 145.785 198.450 ;
        RECT 144.215 197.070 144.895 197.810 ;
        RECT 144.215 196.905 145.085 197.070 ;
        RECT 144.915 196.900 145.085 196.905 ;
        RECT 144.215 196.610 144.895 196.750 ;
        RECT 144.215 196.440 145.085 196.610 ;
        RECT 144.215 196.265 144.895 196.440 ;
        RECT 143.985 194.920 144.895 196.265 ;
        RECT 145.105 195.935 145.785 198.280 ;
        RECT 145.105 195.015 146.015 195.935 ;
        RECT 143.985 194.770 144.895 194.900 ;
        RECT 143.985 194.760 145.085 194.770 ;
        RECT 145.105 194.760 145.885 194.910 ;
        RECT 143.985 194.600 145.885 194.760 ;
        RECT 143.985 193.550 144.895 194.600 ;
        RECT 144.915 194.590 145.885 194.600 ;
        RECT 145.105 193.540 145.885 194.590 ;
        RECT 144.025 193.090 144.810 193.520 ;
        RECT 145.190 193.090 145.975 193.520 ;
        RECT 143.985 192.930 144.895 192.990 ;
        RECT 143.985 192.760 145.085 192.930 ;
        RECT 143.985 189.990 144.895 192.760 ;
        RECT 145.105 190.805 146.015 192.150 ;
        RECT 145.105 190.630 145.785 190.805 ;
        RECT 144.915 190.460 145.785 190.630 ;
        RECT 145.105 190.320 145.785 190.460 ;
        RECT 145.105 190.170 145.915 190.310 ;
        RECT 144.915 190.000 145.915 190.170 ;
        RECT 144.215 189.710 144.895 189.740 ;
        RECT 144.215 189.540 145.085 189.710 ;
        RECT 144.215 187.195 144.895 189.540 ;
        RECT 145.105 188.940 145.915 190.000 ;
        RECT 145.105 187.870 145.885 188.930 ;
        RECT 144.915 187.700 145.885 187.870 ;
        RECT 145.105 187.560 145.885 187.700 ;
        RECT 143.985 186.275 144.895 187.195 ;
        RECT 145.105 186.490 145.885 187.550 ;
        RECT 144.915 186.320 145.885 186.490 ;
        RECT 145.105 186.180 145.885 186.320 ;
        RECT 144.115 185.120 144.895 186.170 ;
        RECT 145.105 185.120 145.885 186.170 ;
        RECT 144.115 184.950 145.885 185.120 ;
        RECT 144.115 184.800 144.895 184.950 ;
        RECT 145.105 184.800 145.885 184.950 ;
        RECT 144.085 183.730 144.895 184.790 ;
        RECT 145.105 183.730 145.915 184.790 ;
        RECT 144.085 183.560 145.915 183.730 ;
        RECT 144.085 183.420 144.895 183.560 ;
        RECT 145.105 183.420 145.915 183.560 ;
      LAYER nwell ;
        RECT 146.305 183.225 147.910 219.485 ;
      LAYER pwell ;
        RECT 62.520 182.695 63.465 182.725 ;
        RECT 60.395 182.495 63.465 182.695 ;
        RECT 63.935 182.695 64.870 182.725 ;
        RECT 66.830 182.695 67.000 182.915 ;
        RECT 67.295 182.725 67.465 182.915 ;
        RECT 69.595 182.725 69.765 182.915 ;
        RECT 76.035 182.745 76.205 182.935 ;
        RECT 76.955 182.725 77.125 182.935 ;
        RECT 82.475 182.725 82.645 182.935 ;
        RECT 87.995 182.725 88.165 182.935 ;
        RECT 90.295 182.725 90.465 182.935 ;
        RECT 60.255 182.015 63.465 182.495 ;
        RECT 60.255 181.815 61.185 182.015 ;
        RECT 62.520 181.815 63.465 182.015 ;
        RECT 63.485 181.855 63.915 182.640 ;
        RECT 63.935 182.495 67.000 182.695 ;
        RECT 63.935 182.015 67.145 182.495 ;
        RECT 67.155 182.045 69.445 182.725 ;
        RECT 69.455 182.045 76.765 182.725 ;
        RECT 63.935 181.815 64.885 182.015 ;
        RECT 66.215 181.815 67.145 182.015 ;
        RECT 68.525 181.815 69.445 182.045 ;
        RECT 72.970 181.825 73.880 182.045 ;
        RECT 75.415 181.815 76.765 182.045 ;
        RECT 76.815 181.915 82.325 182.725 ;
        RECT 82.335 181.915 87.845 182.725 ;
        RECT 87.855 181.915 89.225 182.725 ;
        RECT 89.235 181.915 90.605 182.725 ;
      LAYER nwell ;
        RECT 11.760 178.695 90.800 181.525 ;
      LAYER pwell ;
        RECT 11.955 177.495 13.325 178.305 ;
        RECT 13.335 177.495 17.005 178.305 ;
        RECT 17.515 178.175 18.865 178.405 ;
        RECT 20.400 178.175 21.310 178.395 ;
        RECT 17.515 177.495 24.825 178.175 ;
        RECT 24.845 177.580 25.275 178.365 ;
        RECT 25.295 178.205 26.225 178.405 ;
        RECT 27.555 178.205 28.505 178.405 ;
        RECT 25.295 177.725 28.505 178.205 ;
        RECT 32.030 178.175 32.940 178.395 ;
        RECT 34.475 178.175 35.825 178.405 ;
        RECT 25.440 177.525 28.505 177.725 ;
        RECT 12.095 177.285 12.265 177.495 ;
        RECT 13.475 177.285 13.645 177.495 ;
        RECT 17.150 177.335 17.270 177.445 ;
        RECT 18.990 177.335 19.110 177.445 ;
        RECT 19.455 177.285 19.625 177.475 ;
        RECT 22.215 177.285 22.385 177.475 ;
        RECT 24.515 177.305 24.685 177.495 ;
        RECT 25.440 177.305 25.610 177.525 ;
        RECT 27.570 177.495 28.505 177.525 ;
        RECT 28.515 177.495 35.825 178.175 ;
        RECT 36.335 178.175 37.265 178.405 ;
        RECT 36.335 177.495 39.085 178.175 ;
        RECT 39.095 177.495 44.605 178.305 ;
        RECT 45.665 178.175 46.595 178.405 ;
        RECT 49.180 178.205 50.125 178.405 ;
        RECT 44.760 177.495 46.595 178.175 ;
        RECT 47.375 177.525 50.125 178.205 ;
        RECT 50.605 177.580 51.035 178.365 ;
        RECT 27.735 177.285 27.905 177.475 ;
        RECT 28.655 177.305 28.825 177.495 ;
        RECT 33.255 177.285 33.425 177.475 ;
        RECT 36.010 177.335 36.130 177.445 ;
        RECT 36.945 177.330 37.105 177.440 ;
        RECT 38.315 177.285 38.485 177.475 ;
        RECT 38.775 177.305 38.945 177.495 ;
        RECT 39.235 177.305 39.405 177.495 ;
        RECT 44.760 177.475 44.925 177.495 ;
        RECT 41.995 177.285 42.165 177.475 ;
        RECT 43.380 177.285 43.550 177.475 ;
        RECT 44.755 177.285 44.925 177.475 ;
        RECT 47.050 177.335 47.170 177.445 ;
        RECT 47.520 177.305 47.690 177.525 ;
        RECT 49.180 177.495 50.125 177.525 ;
        RECT 51.055 177.495 54.265 178.405 ;
        RECT 54.735 177.495 56.085 178.405 ;
        RECT 56.115 178.175 57.035 178.405 ;
        RECT 56.115 177.495 58.405 178.175 ;
        RECT 58.475 177.495 60.245 178.405 ;
        RECT 61.175 177.495 64.650 178.405 ;
        RECT 64.855 177.495 68.525 178.305 ;
        RECT 68.555 177.495 69.905 178.405 ;
        RECT 69.915 177.495 71.265 178.405 ;
        RECT 71.295 177.495 74.965 178.305 ;
        RECT 74.975 177.495 76.345 178.305 ;
        RECT 76.365 177.580 76.795 178.365 ;
        RECT 76.815 177.495 82.325 178.305 ;
        RECT 82.335 177.495 87.845 178.305 ;
        RECT 87.855 177.495 89.225 178.305 ;
        RECT 89.235 177.495 90.605 178.305 ;
        RECT 50.275 177.445 50.445 177.475 ;
        RECT 50.270 177.335 50.445 177.445 ;
        RECT 50.275 177.285 50.445 177.335 ;
        RECT 51.195 177.305 51.365 177.495 ;
        RECT 55.800 177.475 55.970 177.495 ;
        RECT 54.410 177.335 54.530 177.445 ;
        RECT 55.795 177.305 55.970 177.475 ;
        RECT 58.095 177.305 58.265 177.495 ;
        RECT 59.930 177.305 60.100 177.495 ;
        RECT 61.320 177.475 61.490 177.495 ;
        RECT 60.405 177.340 60.565 177.450 ;
        RECT 61.315 177.305 61.490 177.475 ;
        RECT 63.150 177.335 63.270 177.445 ;
        RECT 55.795 177.285 55.965 177.305 ;
        RECT 61.315 177.285 61.485 177.305 ;
        RECT 64.075 177.285 64.245 177.475 ;
        RECT 64.995 177.305 65.165 177.495 ;
        RECT 67.755 177.285 67.925 177.475 ;
        RECT 68.225 177.330 68.385 177.440 ;
        RECT 69.140 177.285 69.310 177.475 ;
        RECT 69.590 177.305 69.760 177.495 ;
        RECT 70.060 177.305 70.230 177.495 ;
        RECT 71.435 177.475 71.605 177.495 ;
        RECT 71.430 177.305 71.605 177.475 ;
        RECT 71.430 177.285 71.600 177.305 ;
        RECT 72.820 177.285 72.990 177.475 ;
        RECT 73.275 177.285 73.445 177.475 ;
        RECT 75.115 177.305 75.285 177.495 ;
        RECT 76.955 177.305 77.125 177.495 ;
        RECT 78.795 177.285 78.965 177.475 ;
        RECT 82.475 177.305 82.645 177.495 ;
        RECT 84.315 177.285 84.485 177.475 ;
        RECT 87.995 177.285 88.165 177.495 ;
        RECT 90.295 177.285 90.465 177.495 ;
        RECT 11.955 176.475 13.325 177.285 ;
        RECT 13.335 176.475 18.845 177.285 ;
        RECT 19.315 176.605 22.065 177.285 ;
        RECT 21.135 176.375 22.065 176.605 ;
        RECT 22.075 176.475 27.585 177.285 ;
        RECT 27.595 176.475 33.105 177.285 ;
        RECT 33.115 176.475 36.785 177.285 ;
        RECT 37.725 176.415 38.155 177.200 ;
        RECT 38.175 176.475 41.845 177.285 ;
        RECT 41.855 176.475 43.225 177.285 ;
        RECT 43.235 176.375 44.585 177.285 ;
        RECT 44.615 176.475 50.125 177.285 ;
        RECT 50.135 176.475 55.645 177.285 ;
        RECT 55.655 176.475 61.165 177.285 ;
        RECT 61.175 176.475 63.005 177.285 ;
        RECT 63.485 176.415 63.915 177.200 ;
        RECT 63.935 176.475 66.685 177.285 ;
        RECT 66.705 176.375 68.055 177.285 ;
        RECT 68.995 176.375 70.345 177.285 ;
        RECT 70.395 176.375 71.745 177.285 ;
        RECT 71.755 176.375 73.105 177.285 ;
        RECT 73.135 176.475 78.645 177.285 ;
        RECT 78.655 176.475 84.165 177.285 ;
        RECT 84.175 176.475 87.845 177.285 ;
        RECT 87.855 176.475 89.225 177.285 ;
        RECT 89.235 176.475 90.605 177.285 ;
      LAYER nwell ;
        RECT 11.760 173.255 90.800 176.085 ;
      LAYER pwell ;
        RECT 11.955 172.055 13.325 172.865 ;
        RECT 13.335 172.055 18.845 172.865 ;
        RECT 18.855 172.055 24.365 172.865 ;
        RECT 24.845 172.140 25.275 172.925 ;
        RECT 25.295 172.055 28.045 172.865 ;
        RECT 29.885 172.735 30.805 172.965 ;
        RECT 28.515 172.055 30.805 172.735 ;
        RECT 30.815 172.735 31.735 172.965 ;
        RECT 30.815 172.055 33.105 172.735 ;
        RECT 33.115 172.055 35.865 172.865 ;
        RECT 41.395 172.735 42.315 172.965 ;
        RECT 43.695 172.735 44.615 172.965 ;
        RECT 36.570 172.055 41.385 172.735 ;
        RECT 41.395 172.055 43.685 172.735 ;
        RECT 43.695 172.055 45.985 172.735 ;
        RECT 45.995 172.055 47.810 172.965 ;
        RECT 47.835 172.055 50.585 172.865 ;
        RECT 50.605 172.140 51.035 172.925 ;
        RECT 51.055 172.055 52.885 172.735 ;
        RECT 52.895 172.055 54.725 172.735 ;
        RECT 54.735 172.055 56.105 172.865 ;
        RECT 56.135 172.055 57.485 172.965 ;
        RECT 57.495 172.055 60.705 172.965 ;
        RECT 61.170 172.285 63.005 172.965 ;
        RECT 61.170 172.055 62.860 172.285 ;
        RECT 63.015 172.055 64.845 172.865 ;
        RECT 65.315 172.735 66.450 172.965 ;
        RECT 68.735 172.875 69.685 172.965 ;
        RECT 65.315 172.055 68.525 172.735 ;
        RECT 68.735 172.055 70.665 172.875 ;
        RECT 72.910 172.735 74.045 172.965 ;
        RECT 70.835 172.055 74.045 172.735 ;
        RECT 74.365 172.735 75.295 172.965 ;
        RECT 74.365 172.055 76.200 172.735 ;
        RECT 76.365 172.140 76.795 172.925 ;
        RECT 80.330 172.735 81.240 172.955 ;
        RECT 82.775 172.735 84.125 172.965 ;
        RECT 76.815 172.055 84.125 172.735 ;
        RECT 84.175 172.055 87.845 172.865 ;
        RECT 87.855 172.055 89.225 172.865 ;
        RECT 89.235 172.055 90.605 172.865 ;
        RECT 12.095 171.845 12.265 172.055 ;
        RECT 13.475 171.845 13.645 172.055 ;
        RECT 18.995 171.845 19.165 172.055 ;
        RECT 20.835 171.845 21.005 172.035 ;
        RECT 24.510 171.895 24.630 172.005 ;
        RECT 25.435 171.865 25.605 172.055 ;
        RECT 28.190 171.845 28.360 172.035 ;
        RECT 28.655 171.865 28.825 172.055 ;
        RECT 29.575 171.845 29.745 172.035 ;
        RECT 32.795 171.865 32.965 172.055 ;
        RECT 33.255 171.865 33.425 172.055 ;
        RECT 36.010 171.895 36.130 172.005 ;
        RECT 36.945 171.890 37.105 172.000 ;
        RECT 38.315 171.845 38.485 172.035 ;
        RECT 41.075 171.865 41.245 172.055 ;
        RECT 43.375 171.865 43.545 172.055 ;
        RECT 45.675 171.865 45.845 172.055 ;
        RECT 47.515 171.865 47.685 172.055 ;
        RECT 47.975 171.865 48.145 172.055 ;
        RECT 48.435 171.845 48.605 172.035 ;
        RECT 51.195 171.865 51.365 172.055 ;
        RECT 54.415 171.865 54.585 172.055 ;
        RECT 54.875 171.865 55.045 172.055 ;
        RECT 57.170 171.865 57.340 172.055 ;
        RECT 57.635 171.845 57.805 172.035 ;
        RECT 58.105 171.890 58.265 172.000 ;
        RECT 60.395 171.845 60.565 172.055 ;
        RECT 60.855 171.845 61.025 172.035 ;
        RECT 62.690 171.865 62.860 172.055 ;
        RECT 63.155 171.865 63.325 172.055 ;
        RECT 64.080 171.845 64.250 172.035 ;
        RECT 64.990 171.895 65.110 172.005 ;
        RECT 67.755 171.845 67.925 172.035 ;
        RECT 68.215 171.865 68.385 172.055 ;
        RECT 70.515 172.035 70.665 172.055 ;
        RECT 70.515 171.865 70.685 172.035 ;
        RECT 70.975 171.865 71.145 172.055 ;
        RECT 76.035 172.035 76.200 172.055 ;
        RECT 76.035 171.865 76.205 172.035 ;
        RECT 76.495 171.845 76.665 172.035 ;
        RECT 76.955 171.845 77.125 172.055 ;
        RECT 82.475 171.845 82.645 172.035 ;
        RECT 84.315 171.865 84.485 172.055 ;
        RECT 87.995 171.845 88.165 172.055 ;
        RECT 90.295 171.845 90.465 172.055 ;
        RECT 11.955 171.035 13.325 171.845 ;
        RECT 13.335 171.035 18.845 171.845 ;
        RECT 18.855 171.035 20.685 171.845 ;
        RECT 20.695 171.165 28.005 171.845 ;
        RECT 24.210 170.945 25.120 171.165 ;
        RECT 26.655 170.935 28.005 171.165 ;
        RECT 28.075 170.935 29.425 171.845 ;
        RECT 29.435 171.165 36.745 171.845 ;
        RECT 32.950 170.945 33.860 171.165 ;
        RECT 35.395 170.935 36.745 171.165 ;
        RECT 37.725 170.975 38.155 171.760 ;
        RECT 38.230 170.935 48.250 171.845 ;
        RECT 48.295 171.165 55.605 171.845 ;
        RECT 51.810 170.945 52.720 171.165 ;
        RECT 54.255 170.935 55.605 171.165 ;
        RECT 55.655 170.935 57.945 171.845 ;
        RECT 58.875 171.165 60.705 171.845 ;
        RECT 58.875 170.935 60.220 171.165 ;
        RECT 60.715 171.035 63.465 171.845 ;
        RECT 63.485 170.975 63.915 171.760 ;
        RECT 63.935 171.165 67.605 171.845 ;
        RECT 63.935 170.935 64.860 171.165 ;
        RECT 67.615 171.035 69.445 171.845 ;
        RECT 69.495 171.165 76.805 171.845 ;
        RECT 69.495 170.935 70.845 171.165 ;
        RECT 72.380 170.945 73.290 171.165 ;
        RECT 76.815 171.035 82.325 171.845 ;
        RECT 82.335 171.035 87.845 171.845 ;
        RECT 87.855 171.035 89.225 171.845 ;
        RECT 89.235 171.035 90.605 171.845 ;
      LAYER nwell ;
        RECT 11.760 167.815 90.800 170.645 ;
      LAYER pwell ;
        RECT 11.955 166.615 13.325 167.425 ;
        RECT 13.335 166.615 18.845 167.425 ;
        RECT 18.855 166.615 20.685 167.425 ;
        RECT 21.155 167.325 22.105 167.525 ;
        RECT 23.435 167.325 24.365 167.525 ;
        RECT 21.155 166.845 24.365 167.325 ;
        RECT 21.155 166.645 24.220 166.845 ;
        RECT 24.845 166.700 25.275 167.485 ;
        RECT 21.155 166.615 22.090 166.645 ;
        RECT 12.095 166.405 12.265 166.615 ;
        RECT 13.475 166.405 13.645 166.615 ;
        RECT 18.995 166.405 19.165 166.615 ;
        RECT 20.830 166.455 20.950 166.565 ;
        RECT 22.675 166.425 22.845 166.595 ;
        RECT 24.050 166.425 24.220 166.645 ;
        RECT 25.305 166.615 28.035 167.525 ;
        RECT 28.220 166.615 32.090 167.525 ;
        RECT 32.195 166.615 34.025 167.425 ;
        RECT 35.085 167.295 36.015 167.525 ;
        RECT 34.180 166.615 36.015 167.295 ;
        RECT 36.385 166.615 39.545 167.525 ;
        RECT 43.070 167.295 43.980 167.515 ;
        RECT 45.515 167.295 46.865 167.525 ;
        RECT 39.555 166.615 46.865 167.295 ;
        RECT 47.110 166.615 50.585 167.525 ;
        RECT 50.605 166.700 51.035 167.485 ;
        RECT 51.075 166.615 52.425 167.525 ;
        RECT 52.445 166.615 53.795 167.525 ;
        RECT 55.635 167.295 56.565 167.525 ;
        RECT 53.815 166.615 56.565 167.295 ;
        RECT 56.575 166.615 61.390 167.295 ;
        RECT 61.675 166.615 64.845 167.525 ;
        RECT 64.855 166.615 66.685 167.425 ;
        RECT 67.205 166.615 70.365 167.525 ;
        RECT 70.375 167.295 71.295 167.525 ;
        RECT 70.375 166.615 72.665 167.295 ;
        RECT 72.675 166.615 76.345 167.425 ;
        RECT 76.365 166.700 76.795 167.485 ;
        RECT 76.815 166.615 82.325 167.425 ;
        RECT 82.335 166.615 87.845 167.425 ;
        RECT 87.855 166.615 89.225 167.425 ;
        RECT 89.235 166.615 90.605 167.425 ;
        RECT 100.450 167.190 106.550 176.980 ;
        RECT 100.450 167.160 106.560 167.190 ;
        RECT 100.650 166.760 101.810 167.160 ;
        RECT 24.510 166.455 24.630 166.565 ;
        RECT 25.435 166.425 25.605 166.615 ;
        RECT 28.220 166.595 28.365 166.615 ;
        RECT 22.680 166.405 22.845 166.425 ;
        RECT 27.735 166.405 27.905 166.595 ;
        RECT 28.195 166.425 28.365 166.595 ;
        RECT 32.335 166.425 32.505 166.615 ;
        RECT 34.180 166.595 34.345 166.615 ;
        RECT 32.795 166.405 32.965 166.595 ;
        RECT 33.255 166.405 33.425 166.595 ;
        RECT 34.175 166.425 34.345 166.595 ;
        RECT 36.015 166.405 36.185 166.595 ;
        RECT 36.475 166.425 36.645 166.615 ;
        RECT 38.315 166.405 38.485 166.595 ;
        RECT 39.695 166.425 39.865 166.615 ;
        RECT 43.835 166.405 44.005 166.595 ;
        RECT 49.355 166.405 49.525 166.595 ;
        RECT 50.270 166.425 50.440 166.615 ;
        RECT 51.190 166.425 51.360 166.615 ;
        RECT 52.575 166.425 52.745 166.615 ;
        RECT 53.955 166.425 54.125 166.615 ;
        RECT 54.875 166.405 55.045 166.595 ;
        RECT 56.715 166.425 56.885 166.615 ;
        RECT 60.850 166.455 60.970 166.565 ;
        RECT 56.740 166.405 56.885 166.425 ;
        RECT 61.320 166.405 61.490 166.595 ;
        RECT 61.775 166.425 61.945 166.615 ;
        RECT 64.075 166.405 64.245 166.595 ;
        RECT 64.995 166.425 65.165 166.615 ;
        RECT 66.830 166.455 66.950 166.565 ;
        RECT 67.295 166.405 67.465 166.615 ;
        RECT 72.355 166.405 72.525 166.615 ;
        RECT 72.815 166.425 72.985 166.615 ;
        RECT 76.955 166.425 77.125 166.615 ;
        RECT 77.875 166.405 78.045 166.595 ;
        RECT 82.475 166.425 82.645 166.615 ;
        RECT 83.395 166.405 83.565 166.595 ;
        RECT 87.995 166.425 88.165 166.615 ;
        RECT 88.910 166.455 89.030 166.565 ;
        RECT 90.295 166.405 90.465 166.615 ;
        RECT 11.955 165.595 13.325 166.405 ;
        RECT 13.335 165.595 18.845 166.405 ;
        RECT 18.855 165.595 22.525 166.405 ;
        RECT 22.680 165.725 24.515 166.405 ;
        RECT 23.585 165.495 24.515 165.725 ;
        RECT 24.835 165.725 28.045 166.405 ;
        RECT 28.290 165.725 33.105 166.405 ;
        RECT 24.835 165.495 25.970 165.725 ;
        RECT 33.125 165.495 35.855 166.405 ;
        RECT 35.875 165.595 37.705 166.405 ;
        RECT 37.725 165.535 38.155 166.320 ;
        RECT 38.175 165.595 43.685 166.405 ;
        RECT 43.695 165.595 49.205 166.405 ;
        RECT 49.215 165.595 54.725 166.405 ;
        RECT 54.735 165.595 56.565 166.405 ;
        RECT 56.740 165.495 60.610 166.405 ;
        RECT 61.320 166.175 63.010 166.405 ;
        RECT 61.175 165.495 63.010 166.175 ;
        RECT 63.485 165.535 63.915 166.320 ;
        RECT 63.935 165.725 66.675 166.405 ;
        RECT 67.155 165.725 71.970 166.405 ;
        RECT 72.215 165.595 77.725 166.405 ;
        RECT 77.735 165.595 83.245 166.405 ;
        RECT 83.255 165.595 88.765 166.405 ;
        RECT 89.235 165.595 90.605 166.405 ;
      LAYER nwell ;
        RECT 11.760 162.375 90.800 165.205 ;
      LAYER pwell ;
        RECT 103.770 165.080 106.560 167.160 ;
      LAYER nwell ;
        RECT 101.660 162.970 106.500 165.080 ;
        RECT 107.780 164.740 117.970 176.990 ;
      LAYER pwell ;
        RECT 120.330 167.140 126.430 176.930 ;
        RECT 120.330 167.110 126.440 167.140 ;
        RECT 120.530 166.710 121.690 167.110 ;
        RECT 123.650 165.030 126.440 167.110 ;
      LAYER nwell ;
        RECT 121.540 162.920 126.380 165.030 ;
        RECT 127.660 164.690 137.850 176.940 ;
      LAYER pwell ;
        RECT 140.360 167.190 146.460 176.980 ;
        RECT 140.360 167.160 146.470 167.190 ;
        RECT 140.560 166.760 141.720 167.160 ;
        RECT 143.680 165.080 146.470 167.160 ;
      LAYER nwell ;
        RECT 141.570 162.970 146.410 165.080 ;
        RECT 147.690 164.740 157.880 176.990 ;
      LAYER pwell ;
        RECT 11.955 161.175 13.325 161.985 ;
        RECT 13.335 161.175 18.845 161.985 ;
        RECT 18.855 161.175 24.365 161.985 ;
        RECT 24.845 161.260 25.275 162.045 ;
        RECT 25.295 161.885 26.225 162.085 ;
        RECT 27.555 161.885 28.505 162.085 ;
        RECT 25.295 161.405 28.505 161.885 ;
        RECT 29.565 161.855 30.495 162.085 ;
        RECT 25.440 161.205 28.505 161.405 ;
        RECT 12.095 160.965 12.265 161.175 ;
        RECT 13.475 160.965 13.645 161.175 ;
        RECT 18.995 160.965 19.165 161.175 ;
        RECT 22.670 161.015 22.790 161.125 ;
        RECT 24.510 161.015 24.630 161.125 ;
        RECT 25.440 160.985 25.610 161.205 ;
        RECT 27.570 161.175 28.505 161.205 ;
        RECT 28.660 161.175 30.495 161.855 ;
        RECT 31.425 161.175 35.080 162.085 ;
        RECT 35.415 161.175 38.165 162.085 ;
        RECT 39.095 161.175 42.205 162.085 ;
        RECT 42.315 161.175 45.065 161.985 ;
        RECT 45.535 161.175 47.365 161.855 ;
        RECT 47.375 161.175 50.295 162.085 ;
        RECT 50.605 161.260 51.035 162.045 ;
        RECT 51.055 161.175 52.425 161.985 ;
        RECT 52.745 161.855 53.675 162.085 ;
        RECT 55.220 161.855 56.565 162.085 ;
        RECT 52.745 161.175 54.580 161.855 ;
        RECT 54.735 161.175 56.565 161.855 ;
        RECT 57.515 161.175 58.865 162.085 ;
        RECT 58.875 161.175 62.085 162.085 ;
        RECT 62.550 161.405 64.385 162.085 ;
        RECT 62.550 161.175 64.240 161.405 ;
        RECT 64.395 161.175 66.225 161.985 ;
        RECT 66.275 161.175 69.445 162.085 ;
        RECT 72.195 161.855 73.125 162.085 ;
        RECT 69.455 161.175 73.125 161.855 ;
        RECT 73.135 161.175 75.885 161.985 ;
        RECT 76.365 161.260 76.795 162.045 ;
        RECT 76.815 161.175 82.325 161.985 ;
        RECT 82.335 161.175 87.845 161.985 ;
        RECT 87.855 161.175 89.225 161.985 ;
        RECT 89.235 161.175 90.605 161.985 ;
        RECT 28.660 161.155 28.825 161.175 ;
        RECT 31.425 161.155 31.585 161.175 ;
        RECT 28.655 160.985 28.825 161.155 ;
        RECT 30.035 160.965 30.205 161.155 ;
        RECT 30.505 161.010 30.665 161.120 ;
        RECT 30.950 161.015 31.070 161.125 ;
        RECT 31.415 160.965 31.585 161.155 ;
        RECT 34.175 160.965 34.345 161.155 ;
        RECT 35.555 160.985 35.725 161.175 ;
        RECT 36.010 161.015 36.130 161.125 ;
        RECT 36.470 160.965 36.640 161.155 ;
        RECT 38.325 161.125 38.485 161.130 ;
        RECT 38.310 161.020 38.485 161.125 ;
        RECT 38.310 161.015 38.430 161.020 ;
        RECT 38.775 160.965 38.945 161.155 ;
        RECT 41.995 160.985 42.165 161.175 ;
        RECT 42.455 160.985 42.625 161.175 ;
        RECT 45.210 161.015 45.330 161.125 ;
        RECT 46.135 160.965 46.305 161.155 ;
        RECT 47.055 160.985 47.225 161.175 ;
        RECT 47.520 160.985 47.690 161.175 ;
        RECT 51.195 160.985 51.365 161.175 ;
        RECT 54.415 161.155 54.580 161.175 ;
        RECT 53.495 160.965 53.665 161.155 ;
        RECT 54.415 160.985 54.585 161.155 ;
        RECT 54.875 160.965 55.045 161.175 ;
        RECT 56.725 161.020 56.885 161.130 ;
        RECT 57.635 160.965 57.805 161.155 ;
        RECT 58.550 160.985 58.720 161.175 ;
        RECT 59.015 160.985 59.185 161.175 ;
        RECT 64.070 161.155 64.240 161.175 ;
        RECT 63.150 161.015 63.270 161.125 ;
        RECT 64.070 160.985 64.245 161.155 ;
        RECT 64.535 160.985 64.705 161.175 ;
        RECT 66.375 160.985 66.545 161.175 ;
        RECT 64.075 160.965 64.245 160.985 ;
        RECT 69.595 160.965 69.765 161.175 ;
        RECT 71.430 161.015 71.550 161.125 ;
        RECT 71.895 160.965 72.065 161.155 ;
        RECT 73.275 160.985 73.445 161.175 ;
        RECT 76.030 161.015 76.150 161.125 ;
        RECT 76.955 160.985 77.125 161.175 ;
        RECT 79.255 160.965 79.425 161.155 ;
        RECT 82.475 160.985 82.645 161.175 ;
        RECT 84.775 160.965 84.945 161.155 ;
        RECT 87.995 160.985 88.165 161.175 ;
        RECT 88.465 161.010 88.625 161.120 ;
        RECT 90.295 160.965 90.465 161.175 ;
        RECT 11.955 160.155 13.325 160.965 ;
        RECT 13.335 160.155 18.845 160.965 ;
        RECT 18.855 160.155 22.525 160.965 ;
        RECT 23.035 160.285 30.345 160.965 ;
        RECT 23.035 160.055 24.385 160.285 ;
        RECT 25.920 160.065 26.830 160.285 ;
        RECT 31.275 160.055 34.025 160.965 ;
        RECT 34.035 160.155 35.865 160.965 ;
        RECT 36.355 160.055 37.705 160.965 ;
        RECT 37.725 160.095 38.155 160.880 ;
        RECT 38.635 160.285 45.945 160.965 ;
        RECT 45.995 160.285 53.305 160.965 ;
        RECT 42.150 160.065 43.060 160.285 ;
        RECT 44.595 160.055 45.945 160.285 ;
        RECT 49.510 160.065 50.420 160.285 ;
        RECT 51.955 160.055 53.305 160.285 ;
        RECT 53.355 160.155 54.725 160.965 ;
        RECT 54.735 160.055 57.485 160.965 ;
        RECT 57.495 160.155 63.005 160.965 ;
        RECT 63.485 160.095 63.915 160.880 ;
        RECT 63.935 160.155 69.445 160.965 ;
        RECT 69.455 160.155 71.285 160.965 ;
        RECT 71.755 160.285 79.065 160.965 ;
        RECT 75.270 160.065 76.180 160.285 ;
        RECT 77.715 160.055 79.065 160.285 ;
        RECT 79.115 160.155 84.625 160.965 ;
        RECT 84.635 160.155 88.305 160.965 ;
        RECT 89.235 160.155 90.605 160.965 ;
      LAYER nwell ;
        RECT 11.760 156.935 90.800 159.765 ;
      LAYER pwell ;
        RECT 11.955 155.735 13.325 156.545 ;
        RECT 13.335 155.735 18.845 156.545 ;
        RECT 18.855 155.735 24.365 156.545 ;
        RECT 24.845 155.820 25.275 156.605 ;
        RECT 25.295 155.735 26.645 156.645 ;
        RECT 31.935 156.555 32.885 156.645 ;
        RECT 26.675 155.735 30.345 156.545 ;
        RECT 30.355 155.735 31.725 156.545 ;
        RECT 31.935 155.735 33.865 156.555 ;
        RECT 34.035 155.735 37.705 156.545 ;
        RECT 37.715 155.735 39.085 156.545 ;
        RECT 39.095 156.415 40.025 156.645 ;
        RECT 39.095 155.735 42.765 156.415 ;
        RECT 42.775 155.735 44.145 156.545 ;
        RECT 46.895 156.415 47.825 156.645 ;
        RECT 44.155 155.735 47.825 156.415 ;
        RECT 47.835 155.735 50.585 156.545 ;
        RECT 50.605 155.820 51.035 156.605 ;
        RECT 51.055 155.735 52.885 156.545 ;
        RECT 52.895 156.415 53.820 156.645 ;
        RECT 56.575 156.445 57.525 156.645 ;
        RECT 52.895 155.735 56.565 156.415 ;
        RECT 56.575 155.765 60.245 156.445 ;
        RECT 56.575 155.735 57.525 155.765 ;
        RECT 12.095 155.525 12.265 155.735 ;
        RECT 13.475 155.525 13.645 155.735 ;
        RECT 18.995 155.525 19.165 155.735 ;
        RECT 20.830 155.575 20.950 155.685 ;
        RECT 21.295 155.525 21.465 155.715 ;
        RECT 24.510 155.575 24.630 155.685 ;
        RECT 25.435 155.545 25.605 155.715 ;
        RECT 25.435 155.525 25.600 155.545 ;
        RECT 25.895 155.525 26.065 155.715 ;
        RECT 26.360 155.545 26.530 155.735 ;
        RECT 26.815 155.545 26.985 155.735 ;
        RECT 30.495 155.545 30.665 155.735 ;
        RECT 33.715 155.715 33.865 155.735 ;
        RECT 33.255 155.525 33.425 155.715 ;
        RECT 33.715 155.545 33.885 155.715 ;
        RECT 34.175 155.545 34.345 155.735 ;
        RECT 36.945 155.570 37.105 155.680 ;
        RECT 37.855 155.545 38.025 155.735 ;
        RECT 38.315 155.525 38.485 155.715 ;
        RECT 42.455 155.545 42.625 155.735 ;
        RECT 42.915 155.545 43.085 155.735 ;
        RECT 43.835 155.525 44.005 155.715 ;
        RECT 44.295 155.545 44.465 155.735 ;
        RECT 47.515 155.525 47.685 155.715 ;
        RECT 47.975 155.545 48.145 155.735 ;
        RECT 48.900 155.525 49.070 155.715 ;
        RECT 50.275 155.525 50.445 155.715 ;
        RECT 51.195 155.545 51.365 155.735 ;
        RECT 53.040 155.545 53.210 155.735 ;
        RECT 11.955 154.715 13.325 155.525 ;
        RECT 13.335 154.715 18.845 155.525 ;
        RECT 18.855 154.715 20.685 155.525 ;
        RECT 21.155 154.845 23.445 155.525 ;
        RECT 22.525 154.615 23.445 154.845 ;
        RECT 23.765 154.845 25.600 155.525 ;
        RECT 25.755 154.845 33.065 155.525 ;
        RECT 23.765 154.615 24.695 154.845 ;
        RECT 29.270 154.625 30.180 154.845 ;
        RECT 31.715 154.615 33.065 154.845 ;
        RECT 33.115 154.715 36.785 155.525 ;
        RECT 37.725 154.655 38.155 155.440 ;
        RECT 38.175 154.715 43.685 155.525 ;
        RECT 43.695 154.715 47.365 155.525 ;
        RECT 47.375 154.715 48.745 155.525 ;
        RECT 48.755 154.615 50.105 155.525 ;
        RECT 50.215 154.615 53.215 155.525 ;
        RECT 53.500 155.495 53.670 155.715 ;
        RECT 56.255 155.525 56.425 155.715 ;
        RECT 59.930 155.680 60.100 155.765 ;
        RECT 60.255 155.735 63.465 156.645 ;
        RECT 63.475 155.735 66.585 156.645 ;
        RECT 66.695 155.735 69.805 156.645 ;
        RECT 70.395 155.735 71.745 156.645 ;
        RECT 74.495 156.415 75.425 156.645 ;
        RECT 71.755 155.735 75.425 156.415 ;
        RECT 76.365 155.820 76.795 156.605 ;
        RECT 80.330 156.415 81.240 156.635 ;
        RECT 82.775 156.415 84.125 156.645 ;
        RECT 76.815 155.735 84.125 156.415 ;
        RECT 84.175 155.735 87.845 156.545 ;
        RECT 87.855 155.735 89.225 156.545 ;
        RECT 89.235 155.735 90.605 156.545 ;
        RECT 59.930 155.570 60.105 155.680 ;
        RECT 59.930 155.545 60.100 155.570 ;
        RECT 60.385 155.545 60.555 155.735 ;
        RECT 55.160 155.495 56.105 155.525 ;
        RECT 53.355 154.815 56.105 155.495 ;
        RECT 55.160 154.615 56.105 154.815 ;
        RECT 56.115 154.715 59.785 155.525 ;
        RECT 60.715 155.495 61.670 155.525 ;
        RECT 62.700 155.495 62.870 155.715 ;
        RECT 63.150 155.575 63.270 155.685 ;
        RECT 64.085 155.570 64.245 155.680 ;
        RECT 66.375 155.545 66.545 155.735 ;
        RECT 64.855 155.495 65.810 155.525 ;
        RECT 66.840 155.495 67.010 155.715 ;
        RECT 67.305 155.570 67.465 155.680 ;
        RECT 69.595 155.545 69.765 155.735 ;
        RECT 71.430 155.715 71.600 155.735 ;
        RECT 70.050 155.575 70.170 155.685 ;
        RECT 70.975 155.525 71.145 155.715 ;
        RECT 71.430 155.545 71.605 155.715 ;
        RECT 71.895 155.545 72.065 155.735 ;
        RECT 71.435 155.525 71.605 155.545 ;
        RECT 75.115 155.525 75.285 155.715 ;
        RECT 75.585 155.580 75.745 155.690 ;
        RECT 76.955 155.525 77.125 155.735 ;
        RECT 77.415 155.525 77.585 155.715 ;
        RECT 82.935 155.525 83.105 155.715 ;
        RECT 84.315 155.545 84.485 155.735 ;
        RECT 87.995 155.545 88.165 155.735 ;
        RECT 88.465 155.570 88.625 155.680 ;
        RECT 90.295 155.525 90.465 155.735 ;
        RECT 60.715 154.815 62.995 155.495 ;
        RECT 60.715 154.615 61.670 154.815 ;
        RECT 63.485 154.655 63.915 155.440 ;
        RECT 64.855 154.815 67.135 155.495 ;
        RECT 68.075 154.845 71.285 155.525 ;
        RECT 64.855 154.615 65.810 154.815 ;
        RECT 68.075 154.615 69.210 154.845 ;
        RECT 71.295 154.715 73.125 155.525 ;
        RECT 73.135 154.845 75.425 155.525 ;
        RECT 73.135 154.615 74.055 154.845 ;
        RECT 75.435 154.615 77.250 155.525 ;
        RECT 77.275 154.715 82.785 155.525 ;
        RECT 82.795 154.715 88.305 155.525 ;
        RECT 89.235 154.715 90.605 155.525 ;
      LAYER nwell ;
        RECT 11.760 151.495 90.800 154.325 ;
      LAYER pwell ;
        RECT 100.450 152.190 106.550 161.980 ;
        RECT 100.450 152.160 106.560 152.190 ;
        RECT 100.650 151.760 101.810 152.160 ;
        RECT 11.955 150.295 13.325 151.105 ;
        RECT 13.335 150.295 17.005 151.105 ;
        RECT 20.990 150.975 21.900 151.195 ;
        RECT 23.435 150.975 24.785 151.205 ;
        RECT 17.475 150.295 24.785 150.975 ;
        RECT 24.845 150.380 25.275 151.165 ;
        RECT 25.305 150.295 28.035 151.205 ;
        RECT 28.055 150.295 30.805 151.105 ;
        RECT 30.815 150.295 34.470 151.205 ;
        RECT 34.495 150.295 35.865 151.105 ;
        RECT 36.330 150.525 38.165 151.205 ;
        RECT 36.330 150.295 38.020 150.525 ;
        RECT 38.675 150.295 41.845 151.205 ;
        RECT 41.855 150.295 43.225 151.105 ;
        RECT 43.335 150.295 46.445 151.205 ;
        RECT 46.455 150.295 47.825 151.105 ;
        RECT 49.640 151.005 50.585 151.205 ;
        RECT 47.835 150.325 50.585 151.005 ;
        RECT 50.605 150.380 51.035 151.165 ;
        RECT 12.095 150.085 12.265 150.295 ;
        RECT 13.475 150.085 13.645 150.295 ;
        RECT 17.150 150.135 17.270 150.245 ;
        RECT 17.615 150.105 17.785 150.295 ;
        RECT 11.955 149.275 13.325 150.085 ;
        RECT 13.335 149.275 18.845 150.085 ;
        RECT 18.855 150.055 19.790 150.085 ;
        RECT 21.750 150.055 21.920 150.275 ;
        RECT 22.210 150.135 22.330 150.245 ;
        RECT 24.515 150.085 24.685 150.275 ;
        RECT 24.975 150.085 25.145 150.275 ;
        RECT 25.435 150.105 25.605 150.295 ;
        RECT 28.195 150.105 28.365 150.295 ;
        RECT 30.500 150.085 30.670 150.275 ;
        RECT 30.960 150.105 31.130 150.295 ;
        RECT 33.715 150.085 33.885 150.275 ;
        RECT 34.635 150.105 34.805 150.295 ;
        RECT 37.390 150.135 37.510 150.245 ;
        RECT 37.850 150.105 38.020 150.295 ;
        RECT 38.310 150.135 38.430 150.245 ;
        RECT 38.775 150.105 38.945 150.295 ;
        RECT 41.995 150.105 42.165 150.295 ;
        RECT 43.375 150.105 43.545 150.295 ;
        RECT 45.215 150.085 45.385 150.275 ;
        RECT 45.675 150.085 45.845 150.275 ;
        RECT 46.595 150.105 46.765 150.295 ;
        RECT 47.510 150.135 47.630 150.245 ;
        RECT 47.980 150.105 48.150 150.325 ;
        RECT 49.640 150.295 50.585 150.325 ;
        RECT 51.055 150.295 58.615 151.205 ;
        RECT 58.875 150.295 62.530 151.205 ;
        RECT 62.555 150.295 63.905 151.205 ;
        RECT 63.935 150.295 69.445 151.105 ;
        RECT 69.455 150.295 72.205 151.105 ;
        RECT 72.235 150.295 73.585 151.205 ;
        RECT 73.595 150.295 74.945 151.205 ;
        RECT 74.975 150.295 76.345 151.105 ;
        RECT 76.365 150.380 76.795 151.165 ;
        RECT 76.815 150.295 82.325 151.105 ;
        RECT 82.335 150.295 87.845 151.105 ;
        RECT 87.855 150.295 89.225 151.105 ;
        RECT 89.235 150.295 90.605 151.105 ;
        RECT 50.275 150.085 50.445 150.275 ;
        RECT 50.735 150.085 50.905 150.275 ;
        RECT 51.200 150.105 51.370 150.295 ;
        RECT 56.255 150.085 56.425 150.275 ;
        RECT 57.635 150.105 57.805 150.275 ;
        RECT 59.020 150.105 59.190 150.295 ;
        RECT 57.640 150.085 57.805 150.105 ;
        RECT 59.940 150.085 60.110 150.275 ;
        RECT 63.620 150.105 63.790 150.295 ;
        RECT 64.075 150.275 64.245 150.295 ;
        RECT 69.595 150.275 69.765 150.295 ;
        RECT 64.075 150.105 64.250 150.275 ;
        RECT 64.080 150.085 64.250 150.105 ;
        RECT 69.590 150.105 69.765 150.275 ;
        RECT 69.590 150.085 69.760 150.105 ;
        RECT 70.055 150.085 70.225 150.275 ;
        RECT 73.270 150.105 73.440 150.295 ;
        RECT 73.740 150.275 73.910 150.295 ;
        RECT 73.735 150.105 73.910 150.275 ;
        RECT 75.115 150.105 75.285 150.295 ;
        RECT 76.955 150.105 77.125 150.295 ;
        RECT 73.735 150.085 73.905 150.105 ;
        RECT 81.095 150.085 81.265 150.275 ;
        RECT 82.475 150.105 82.645 150.295 ;
        RECT 86.615 150.085 86.785 150.275 ;
        RECT 87.995 150.105 88.165 150.295 ;
        RECT 90.295 150.085 90.465 150.295 ;
        RECT 18.855 149.855 21.920 150.055 ;
        RECT 18.855 149.375 22.065 149.855 ;
        RECT 18.855 149.175 19.805 149.375 ;
        RECT 21.135 149.175 22.065 149.375 ;
        RECT 22.535 149.405 24.825 150.085 ;
        RECT 22.535 149.175 23.455 149.405 ;
        RECT 24.835 149.275 30.345 150.085 ;
        RECT 30.355 149.175 33.420 150.085 ;
        RECT 33.575 149.275 37.245 150.085 ;
        RECT 37.725 149.215 38.155 150.000 ;
        RECT 38.215 149.405 45.525 150.085 ;
        RECT 38.215 149.175 39.565 149.405 ;
        RECT 41.100 149.185 42.010 149.405 ;
        RECT 45.535 149.275 47.365 150.085 ;
        RECT 47.845 149.175 50.575 150.085 ;
        RECT 50.595 149.275 56.105 150.085 ;
        RECT 56.115 149.275 57.485 150.085 ;
        RECT 57.640 149.405 59.475 150.085 ;
        RECT 58.545 149.175 59.475 149.405 ;
        RECT 59.795 149.175 63.270 150.085 ;
        RECT 63.485 149.215 63.915 150.000 ;
        RECT 63.935 149.175 67.410 150.085 ;
        RECT 68.070 149.855 69.760 150.085 ;
        RECT 68.070 149.175 69.905 149.855 ;
        RECT 69.915 149.405 73.585 150.085 ;
        RECT 73.595 149.405 80.905 150.085 ;
        RECT 72.655 149.175 73.585 149.405 ;
        RECT 77.110 149.185 78.020 149.405 ;
        RECT 79.555 149.175 80.905 149.405 ;
        RECT 80.955 149.275 86.465 150.085 ;
        RECT 86.475 149.275 89.225 150.085 ;
        RECT 89.235 149.275 90.605 150.085 ;
        RECT 103.770 150.080 106.560 152.160 ;
      LAYER nwell ;
        RECT 11.760 146.055 90.800 148.885 ;
        RECT 101.660 147.970 106.500 150.080 ;
        RECT 107.780 149.740 117.970 161.990 ;
      LAYER pwell ;
        RECT 120.330 152.190 126.430 161.980 ;
        RECT 120.330 152.160 126.440 152.190 ;
        RECT 120.530 151.760 121.690 152.160 ;
        RECT 123.650 150.080 126.440 152.160 ;
      LAYER nwell ;
        RECT 121.540 147.970 126.380 150.080 ;
        RECT 127.660 149.740 137.850 161.990 ;
      LAYER pwell ;
        RECT 140.410 152.140 146.510 161.930 ;
        RECT 140.410 152.110 146.520 152.140 ;
        RECT 140.610 151.710 141.770 152.110 ;
        RECT 143.730 150.030 146.520 152.110 ;
      LAYER nwell ;
        RECT 141.620 147.920 146.460 150.030 ;
        RECT 147.740 149.690 157.930 161.940 ;
      LAYER pwell ;
        RECT 11.955 144.855 13.325 145.665 ;
        RECT 13.335 144.855 18.845 145.665 ;
        RECT 18.855 144.855 24.365 145.665 ;
        RECT 24.845 144.940 25.275 145.725 ;
        RECT 25.295 144.855 26.665 145.665 ;
        RECT 26.695 144.855 28.045 145.765 ;
        RECT 28.985 144.855 31.715 145.765 ;
        RECT 34.390 145.535 35.310 145.765 ;
        RECT 36.465 145.535 37.395 145.765 ;
        RECT 31.845 144.855 35.310 145.535 ;
        RECT 35.560 144.855 37.395 145.535 ;
        RECT 37.725 144.855 39.075 145.765 ;
        RECT 41.835 145.535 42.765 145.765 ;
        RECT 39.095 144.855 42.765 145.535 ;
        RECT 42.775 144.855 48.285 145.665 ;
        RECT 48.295 144.855 50.125 145.665 ;
        RECT 50.605 144.940 51.035 145.725 ;
        RECT 58.175 145.675 59.125 145.765 ;
        RECT 51.055 144.855 56.565 145.665 ;
        RECT 57.195 144.855 59.125 145.675 ;
        RECT 59.335 145.565 60.265 145.765 ;
        RECT 61.600 145.565 62.545 145.765 ;
        RECT 59.335 145.085 62.545 145.565 ;
        RECT 59.475 144.885 62.545 145.085 ;
        RECT 12.095 144.645 12.265 144.855 ;
        RECT 13.475 144.645 13.645 144.855 ;
        RECT 18.995 144.645 19.165 144.855 ;
        RECT 23.595 144.665 23.765 144.835 ;
        RECT 24.055 144.665 24.225 144.835 ;
        RECT 24.510 144.695 24.630 144.805 ;
        RECT 25.435 144.665 25.605 144.855 ;
        RECT 23.595 144.645 23.745 144.665 ;
        RECT 11.955 143.835 13.325 144.645 ;
        RECT 13.335 143.835 18.845 144.645 ;
        RECT 18.855 143.835 21.605 144.645 ;
        RECT 21.815 143.825 23.745 144.645 ;
        RECT 24.060 144.645 24.225 144.665 ;
        RECT 24.060 143.965 25.895 144.645 ;
        RECT 26.360 144.615 26.530 144.835 ;
        RECT 26.810 144.665 26.980 144.855 ;
        RECT 28.205 144.700 28.365 144.810 ;
        RECT 29.115 144.665 29.285 144.855 ;
        RECT 30.035 144.645 30.205 144.835 ;
        RECT 31.875 144.665 32.045 144.855 ;
        RECT 35.560 144.835 35.725 144.855 ;
        RECT 35.095 144.665 35.265 144.835 ;
        RECT 35.555 144.665 35.725 144.835 ;
        RECT 37.855 144.665 38.025 144.855 ;
        RECT 35.245 144.645 35.265 144.665 ;
        RECT 38.315 144.645 38.485 144.835 ;
        RECT 39.235 144.665 39.405 144.855 ;
        RECT 41.995 144.645 42.165 144.835 ;
        RECT 42.465 144.690 42.625 144.800 ;
        RECT 42.915 144.665 43.085 144.855 ;
        RECT 44.290 144.645 44.460 144.835 ;
        RECT 44.755 144.645 44.925 144.835 ;
        RECT 46.590 144.695 46.710 144.805 ;
        RECT 47.970 144.645 48.140 144.835 ;
        RECT 48.435 144.665 48.605 144.855 ;
        RECT 49.815 144.645 49.985 144.835 ;
        RECT 50.270 144.695 50.390 144.805 ;
        RECT 51.195 144.665 51.365 144.855 ;
        RECT 57.195 144.835 57.345 144.855 ;
        RECT 56.710 144.695 56.830 144.805 ;
        RECT 57.175 144.645 57.345 144.835 ;
        RECT 57.645 144.690 57.805 144.800 ;
        RECT 58.555 144.645 58.725 144.835 ;
        RECT 59.475 144.665 59.645 144.885 ;
        RECT 61.600 144.855 62.545 144.885 ;
        RECT 62.555 144.855 65.715 145.765 ;
        RECT 70.845 145.535 73.845 145.765 ;
        RECT 65.775 144.855 70.590 145.535 ;
        RECT 70.845 145.445 75.425 145.535 ;
        RECT 70.835 145.085 75.425 145.445 ;
        RECT 70.835 144.895 71.765 145.085 ;
        RECT 70.845 144.855 71.765 144.895 ;
        RECT 73.855 144.855 75.425 145.085 ;
        RECT 76.365 144.940 76.795 145.725 ;
        RECT 76.815 144.855 78.185 145.635 ;
        RECT 78.195 144.855 83.705 145.665 ;
        RECT 83.715 144.855 89.225 145.665 ;
        RECT 89.235 144.855 90.605 145.665 ;
        RECT 61.775 144.645 61.945 144.835 ;
        RECT 64.075 144.645 64.245 144.835 ;
        RECT 65.455 144.665 65.625 144.855 ;
        RECT 65.915 144.665 66.085 144.855 ;
        RECT 66.835 144.645 67.005 144.835 ;
        RECT 68.675 144.645 68.845 144.835 ;
        RECT 75.115 144.665 75.285 144.855 ;
        RECT 75.585 144.700 75.745 144.810 ;
        RECT 76.035 144.645 76.205 144.835 ;
        RECT 77.875 144.665 78.045 144.855 ;
        RECT 78.335 144.665 78.505 144.855 ;
        RECT 81.555 144.645 81.725 144.835 ;
        RECT 83.855 144.665 84.025 144.855 ;
        RECT 87.075 144.645 87.245 144.835 ;
        RECT 88.910 144.695 89.030 144.805 ;
        RECT 90.295 144.645 90.465 144.855 ;
        RECT 28.935 144.615 29.885 144.645 ;
        RECT 21.815 143.735 22.765 143.825 ;
        RECT 24.965 143.735 25.895 143.965 ;
        RECT 26.215 143.935 29.885 144.615 ;
        RECT 29.895 143.965 34.710 144.645 ;
        RECT 35.245 143.965 37.695 144.645 ;
        RECT 28.935 143.735 29.885 143.935 ;
        RECT 35.735 143.735 37.695 143.965 ;
        RECT 37.725 143.775 38.155 144.560 ;
        RECT 38.175 143.835 40.265 144.645 ;
        RECT 40.935 143.865 42.305 144.645 ;
        RECT 43.255 143.735 44.605 144.645 ;
        RECT 44.615 143.835 46.445 144.645 ;
        RECT 46.935 143.735 48.285 144.645 ;
        RECT 48.295 143.965 50.125 144.645 ;
        RECT 50.175 143.965 57.485 144.645 ;
        RECT 50.175 143.735 51.525 143.965 ;
        RECT 53.060 143.745 53.970 143.965 ;
        RECT 58.415 143.735 61.625 144.645 ;
        RECT 61.635 143.835 63.465 144.645 ;
        RECT 63.485 143.775 63.915 144.560 ;
        RECT 63.935 143.735 66.685 144.645 ;
        RECT 66.695 143.835 68.525 144.645 ;
        RECT 68.535 143.965 75.845 144.645 ;
        RECT 72.050 143.745 72.960 143.965 ;
        RECT 74.495 143.735 75.845 143.965 ;
        RECT 75.895 143.835 81.405 144.645 ;
        RECT 81.415 143.835 86.925 144.645 ;
        RECT 86.935 143.835 88.765 144.645 ;
        RECT 89.235 143.835 90.605 144.645 ;
      LAYER nwell ;
        RECT 11.760 140.615 90.800 143.445 ;
      LAYER pwell ;
        RECT 11.955 139.415 13.325 140.225 ;
        RECT 13.335 139.415 17.005 140.225 ;
        RECT 20.990 140.095 21.900 140.315 ;
        RECT 23.435 140.095 24.785 140.325 ;
        RECT 17.475 139.415 24.785 140.095 ;
        RECT 24.845 139.500 25.275 140.285 ;
        RECT 27.635 140.095 28.985 140.325 ;
        RECT 30.520 140.095 31.430 140.315 ;
        RECT 35.050 140.095 35.970 140.325 ;
        RECT 25.755 139.415 27.585 140.095 ;
        RECT 27.635 139.415 34.945 140.095 ;
        RECT 35.050 139.415 38.515 140.095 ;
        RECT 38.635 139.415 40.465 140.225 ;
        RECT 43.990 140.095 44.900 140.315 ;
        RECT 46.435 140.095 47.785 140.325 ;
        RECT 49.665 140.095 50.585 140.325 ;
        RECT 40.475 139.415 47.785 140.095 ;
        RECT 48.295 139.415 50.585 140.095 ;
        RECT 50.605 139.500 51.035 140.285 ;
        RECT 53.795 140.095 54.725 140.325 ;
        RECT 51.055 139.415 54.725 140.095 ;
        RECT 54.750 139.415 56.565 140.325 ;
        RECT 56.810 139.415 61.625 140.095 ;
        RECT 61.635 139.415 63.005 140.225 ;
        RECT 63.015 140.095 64.150 140.325 ;
        RECT 63.015 139.415 66.225 140.095 ;
        RECT 66.235 139.415 71.745 140.225 ;
        RECT 71.755 139.415 75.425 140.225 ;
        RECT 76.365 139.500 76.795 140.285 ;
        RECT 76.815 139.415 82.325 140.225 ;
        RECT 82.335 139.415 87.845 140.225 ;
        RECT 87.855 139.415 89.225 140.225 ;
        RECT 89.235 139.415 90.605 140.225 ;
        RECT 12.095 139.205 12.265 139.415 ;
        RECT 13.475 139.225 13.645 139.415 ;
        RECT 14.855 139.205 15.025 139.395 ;
        RECT 15.315 139.205 15.485 139.395 ;
        RECT 17.150 139.255 17.270 139.365 ;
        RECT 17.615 139.225 17.785 139.415 ;
        RECT 19.005 139.250 19.165 139.360 ;
        RECT 11.955 138.395 13.325 139.205 ;
        RECT 13.335 138.525 15.165 139.205 ;
        RECT 13.335 138.295 14.680 138.525 ;
        RECT 15.175 138.395 18.845 139.205 ;
        RECT 19.775 139.175 20.710 139.205 ;
        RECT 22.670 139.175 22.840 139.395 ;
        RECT 23.135 139.205 23.305 139.395 ;
        RECT 24.515 139.225 24.685 139.395 ;
        RECT 25.430 139.255 25.550 139.365 ;
        RECT 25.895 139.225 26.065 139.415 ;
        RECT 24.520 139.205 24.685 139.225 ;
        RECT 26.815 139.205 26.985 139.395 ;
        RECT 29.115 139.205 29.285 139.395 ;
        RECT 34.635 139.225 34.805 139.415 ;
        RECT 36.475 139.205 36.645 139.395 ;
        RECT 38.315 139.225 38.485 139.415 ;
        RECT 38.775 139.225 38.945 139.415 ;
        RECT 39.235 139.205 39.405 139.395 ;
        RECT 40.615 139.225 40.785 139.415 ;
        RECT 47.515 139.205 47.685 139.395 ;
        RECT 47.970 139.255 48.090 139.365 ;
        RECT 48.435 139.225 48.605 139.415 ;
        RECT 50.735 139.205 50.905 139.395 ;
        RECT 51.195 139.225 51.365 139.415 ;
        RECT 52.110 139.205 52.280 139.395 ;
        RECT 52.575 139.205 52.745 139.395 ;
        RECT 54.875 139.225 55.045 139.415 ;
        RECT 56.250 139.255 56.370 139.365 ;
        RECT 56.715 139.205 56.885 139.395 ;
        RECT 59.935 139.205 60.105 139.395 ;
        RECT 61.315 139.225 61.485 139.415 ;
        RECT 61.775 139.225 61.945 139.415 ;
        RECT 64.075 139.205 64.245 139.395 ;
        RECT 65.915 139.225 66.085 139.415 ;
        RECT 66.375 139.225 66.545 139.415 ;
        RECT 66.830 139.205 67.000 139.395 ;
        RECT 67.295 139.205 67.465 139.395 ;
        RECT 68.675 139.205 68.845 139.395 ;
        RECT 71.895 139.225 72.065 139.415 ;
        RECT 75.585 139.260 75.745 139.370 ;
        RECT 76.955 139.225 77.125 139.415 ;
        RECT 79.255 139.205 79.425 139.395 ;
        RECT 79.715 139.205 79.885 139.395 ;
        RECT 82.475 139.225 82.645 139.415 ;
        RECT 85.235 139.205 85.405 139.395 ;
        RECT 87.995 139.225 88.165 139.415 ;
        RECT 88.910 139.255 89.030 139.365 ;
        RECT 90.295 139.205 90.465 139.415 ;
        RECT 19.775 138.975 22.840 139.175 ;
        RECT 19.775 138.495 22.985 138.975 ;
        RECT 19.775 138.295 20.725 138.495 ;
        RECT 22.055 138.295 22.985 138.495 ;
        RECT 22.995 138.395 24.365 139.205 ;
        RECT 24.520 138.525 26.355 139.205 ;
        RECT 26.675 138.525 28.965 139.205 ;
        RECT 28.975 138.525 36.285 139.205 ;
        RECT 25.425 138.295 26.355 138.525 ;
        RECT 28.045 138.295 28.965 138.525 ;
        RECT 32.490 138.305 33.400 138.525 ;
        RECT 34.935 138.295 36.285 138.525 ;
        RECT 36.335 138.395 37.705 139.205 ;
        RECT 37.725 138.335 38.155 139.120 ;
        RECT 39.095 138.525 43.910 139.205 ;
        RECT 44.155 138.525 47.825 139.205 ;
        RECT 47.835 138.525 51.045 139.205 ;
        RECT 44.155 138.295 45.085 138.525 ;
        RECT 47.835 138.295 48.970 138.525 ;
        RECT 51.075 138.295 52.425 139.205 ;
        RECT 52.435 138.395 56.105 139.205 ;
        RECT 56.625 138.295 59.785 139.205 ;
        RECT 59.795 138.395 63.465 139.205 ;
        RECT 63.485 138.335 63.915 139.120 ;
        RECT 63.935 138.395 65.765 139.205 ;
        RECT 65.795 138.295 67.145 139.205 ;
        RECT 67.155 138.395 68.525 139.205 ;
        RECT 68.535 138.525 72.205 139.205 ;
        RECT 71.275 138.295 72.205 138.525 ;
        RECT 72.255 138.525 79.565 139.205 ;
        RECT 72.255 138.295 73.605 138.525 ;
        RECT 75.140 138.305 76.050 138.525 ;
        RECT 79.575 138.395 85.085 139.205 ;
        RECT 85.095 138.395 88.765 139.205 ;
        RECT 89.235 138.395 90.605 139.205 ;
      LAYER nwell ;
        RECT 11.760 135.175 90.800 138.005 ;
      LAYER pwell ;
        RECT 100.450 137.140 106.550 146.930 ;
        RECT 100.450 137.110 106.560 137.140 ;
        RECT 100.650 136.710 101.810 137.110 ;
        RECT 103.770 135.030 106.560 137.110 ;
        RECT 11.955 133.975 13.325 134.785 ;
        RECT 13.335 133.975 18.845 134.785 ;
        RECT 18.855 133.975 24.365 134.785 ;
        RECT 24.845 134.060 25.275 134.845 ;
        RECT 25.295 133.975 28.965 134.785 ;
        RECT 29.895 133.975 31.985 134.785 ;
        RECT 32.670 133.975 34.485 134.885 ;
        RECT 34.495 133.975 36.325 134.785 ;
        RECT 40.310 134.655 41.220 134.875 ;
        RECT 42.755 134.655 44.105 134.885 ;
        RECT 36.795 133.975 44.105 134.655 ;
        RECT 44.155 133.975 49.665 134.785 ;
        RECT 50.605 134.060 51.035 134.845 ;
        RECT 51.055 133.975 52.885 134.655 ;
        RECT 52.895 133.975 56.565 134.785 ;
        RECT 59.315 134.655 60.245 134.885 ;
        RECT 56.575 133.975 60.245 134.655 ;
        RECT 60.275 133.975 61.625 134.885 ;
        RECT 62.115 133.975 63.465 134.885 ;
        RECT 64.395 134.655 65.315 134.885 ;
        RECT 64.395 133.975 66.685 134.655 ;
        RECT 66.710 133.975 68.525 134.885 ;
        RECT 69.495 133.975 72.665 134.885 ;
        RECT 72.675 133.975 76.345 134.785 ;
        RECT 76.365 134.060 76.795 134.845 ;
        RECT 76.815 133.975 82.325 134.785 ;
        RECT 82.335 133.975 87.845 134.785 ;
        RECT 87.855 133.975 89.225 134.785 ;
        RECT 89.235 133.975 90.605 134.785 ;
        RECT 12.095 133.765 12.265 133.975 ;
        RECT 13.475 133.765 13.645 133.975 ;
        RECT 18.995 133.765 19.165 133.975 ;
        RECT 24.515 133.925 24.685 133.955 ;
        RECT 24.510 133.815 24.685 133.925 ;
        RECT 24.515 133.765 24.685 133.815 ;
        RECT 25.435 133.785 25.605 133.975 ;
        RECT 11.955 132.955 13.325 133.765 ;
        RECT 13.335 132.955 18.845 133.765 ;
        RECT 18.855 132.955 24.365 133.765 ;
        RECT 24.375 132.955 25.745 133.765 ;
        RECT 25.755 133.735 26.690 133.765 ;
        RECT 28.650 133.735 28.820 133.955 ;
        RECT 29.125 133.925 29.285 133.930 ;
        RECT 29.110 133.820 29.285 133.925 ;
        RECT 29.110 133.815 29.230 133.820 ;
        RECT 29.575 133.765 29.745 133.955 ;
        RECT 30.035 133.785 30.205 133.975 ;
        RECT 32.795 133.785 32.965 133.975 ;
        RECT 33.265 133.810 33.425 133.920 ;
        RECT 34.175 133.765 34.345 133.955 ;
        RECT 34.635 133.785 34.805 133.975 ;
        RECT 36.470 133.815 36.590 133.925 ;
        RECT 36.935 133.785 37.105 133.975 ;
        RECT 38.315 133.765 38.485 133.955 ;
        RECT 40.155 133.765 40.325 133.955 ;
        RECT 44.295 133.785 44.465 133.975 ;
        RECT 44.755 133.765 44.925 133.955 ;
        RECT 46.140 133.765 46.310 133.955 ;
        RECT 46.605 133.810 46.765 133.920 ;
        RECT 47.515 133.765 47.685 133.955 ;
        RECT 49.825 133.820 49.985 133.930 ;
        RECT 50.735 133.765 50.905 133.955 ;
        RECT 52.575 133.785 52.745 133.975 ;
        RECT 53.035 133.785 53.205 133.975 ;
        RECT 54.415 133.765 54.585 133.955 ;
        RECT 56.255 133.765 56.425 133.955 ;
        RECT 56.715 133.785 56.885 133.975 ;
        RECT 61.310 133.785 61.480 133.975 ;
        RECT 61.770 133.815 61.890 133.925 ;
        RECT 63.150 133.785 63.320 133.975 ;
        RECT 63.625 133.820 63.785 133.930 ;
        RECT 64.085 133.810 64.245 133.920 ;
        RECT 64.995 133.765 65.165 133.955 ;
        RECT 66.375 133.785 66.545 133.975 ;
        RECT 66.835 133.785 67.005 133.975 ;
        RECT 68.685 133.820 68.845 133.930 ;
        RECT 69.595 133.785 69.765 133.975 ;
        RECT 72.355 133.765 72.525 133.955 ;
        RECT 72.815 133.785 72.985 133.975 ;
        RECT 76.955 133.785 77.125 133.975 ;
        RECT 77.875 133.765 78.045 133.955 ;
        RECT 82.475 133.785 82.645 133.975 ;
        RECT 83.395 133.765 83.565 133.955 ;
        RECT 87.995 133.785 88.165 133.975 ;
        RECT 88.910 133.815 89.030 133.925 ;
        RECT 90.295 133.765 90.465 133.975 ;
        RECT 25.755 133.535 28.820 133.735 ;
        RECT 25.755 133.055 28.965 133.535 ;
        RECT 29.545 133.085 33.010 133.765 ;
        RECT 34.145 133.085 37.610 133.765 ;
        RECT 25.755 132.855 26.705 133.055 ;
        RECT 28.035 132.855 28.965 133.055 ;
        RECT 32.090 132.855 33.010 133.085 ;
        RECT 36.690 132.855 37.610 133.085 ;
        RECT 37.725 132.895 38.155 133.680 ;
        RECT 38.190 132.855 40.005 133.765 ;
        RECT 40.015 132.955 41.385 133.765 ;
        RECT 41.490 133.085 44.955 133.765 ;
        RECT 41.490 132.855 42.410 133.085 ;
        RECT 45.075 132.855 46.425 133.765 ;
        RECT 47.415 132.855 50.585 133.765 ;
        RECT 50.595 133.085 54.265 133.765 ;
        RECT 53.335 132.855 54.265 133.085 ;
        RECT 54.275 132.955 56.105 133.765 ;
        RECT 56.115 133.085 63.425 133.765 ;
        RECT 59.630 132.865 60.540 133.085 ;
        RECT 62.075 132.855 63.425 133.085 ;
        RECT 63.485 132.895 63.915 133.680 ;
        RECT 64.855 133.085 72.165 133.765 ;
        RECT 68.370 132.865 69.280 133.085 ;
        RECT 70.815 132.855 72.165 133.085 ;
        RECT 72.215 132.955 77.725 133.765 ;
        RECT 77.735 132.955 83.245 133.765 ;
        RECT 83.255 132.955 88.765 133.765 ;
        RECT 89.235 132.955 90.605 133.765 ;
      LAYER nwell ;
        RECT 101.660 132.920 106.500 135.030 ;
        RECT 107.780 134.690 117.970 146.940 ;
      LAYER pwell ;
        RECT 120.330 137.140 126.430 146.930 ;
        RECT 120.330 137.110 126.440 137.140 ;
        RECT 120.530 136.710 121.690 137.110 ;
        RECT 123.650 135.030 126.440 137.110 ;
      LAYER nwell ;
        RECT 121.540 132.920 126.380 135.030 ;
        RECT 127.660 134.690 137.850 146.940 ;
      LAYER pwell ;
        RECT 140.360 137.140 146.460 146.930 ;
        RECT 140.360 137.110 146.470 137.140 ;
        RECT 140.560 136.710 141.720 137.110 ;
        RECT 143.680 135.030 146.470 137.110 ;
      LAYER nwell ;
        RECT 141.570 132.920 146.410 135.030 ;
        RECT 147.690 134.690 157.880 146.940 ;
        RECT 11.760 129.735 90.800 132.565 ;
      LAYER pwell ;
        RECT 11.955 128.535 13.325 129.345 ;
        RECT 13.335 128.535 18.845 129.345 ;
        RECT 18.855 128.535 24.365 129.345 ;
        RECT 24.845 128.620 25.275 129.405 ;
        RECT 25.335 129.215 26.685 129.445 ;
        RECT 28.220 129.215 29.130 129.435 ;
        RECT 32.965 129.215 33.895 129.445 ;
        RECT 38.470 129.215 39.380 129.435 ;
        RECT 40.915 129.215 42.265 129.445 ;
        RECT 45.065 129.215 45.985 129.445 ;
        RECT 25.335 128.535 32.645 129.215 ;
        RECT 32.965 128.535 34.800 129.215 ;
        RECT 34.955 128.535 42.265 129.215 ;
        RECT 42.400 128.535 45.985 129.215 ;
        RECT 46.090 129.215 47.010 129.445 ;
        RECT 46.090 128.535 49.555 129.215 ;
        RECT 50.605 128.620 51.035 129.405 ;
        RECT 51.055 128.535 52.405 129.445 ;
        RECT 55.950 129.215 56.860 129.435 ;
        RECT 58.395 129.215 59.745 129.445 ;
        RECT 52.435 128.535 59.745 129.215 ;
        RECT 59.795 128.535 63.465 129.345 ;
        RECT 66.675 129.215 67.605 129.445 ;
        RECT 63.935 128.535 67.605 129.215 ;
        RECT 67.615 128.535 73.125 129.345 ;
        RECT 73.135 128.535 75.885 129.345 ;
        RECT 76.365 128.620 76.795 129.405 ;
        RECT 76.815 128.535 82.325 129.345 ;
        RECT 82.335 128.535 87.845 129.345 ;
        RECT 87.855 128.535 89.225 129.345 ;
        RECT 89.235 128.535 90.605 129.345 ;
        RECT 12.095 128.325 12.265 128.535 ;
        RECT 13.475 128.325 13.645 128.535 ;
        RECT 18.995 128.325 19.165 128.535 ;
        RECT 24.515 128.485 24.685 128.515 ;
        RECT 24.510 128.375 24.685 128.485 ;
        RECT 24.515 128.325 24.685 128.375 ;
        RECT 32.335 128.345 32.505 128.535 ;
        RECT 34.635 128.515 34.800 128.535 ;
        RECT 34.175 128.325 34.345 128.515 ;
        RECT 34.635 128.345 34.805 128.515 ;
        RECT 35.095 128.345 35.265 128.535 ;
        RECT 37.395 128.325 37.565 128.515 ;
        RECT 38.325 128.370 38.485 128.480 ;
        RECT 39.235 128.325 39.405 128.515 ;
        RECT 45.670 128.345 45.840 128.535 ;
        RECT 46.130 128.325 46.300 128.515 ;
        RECT 46.595 128.325 46.765 128.515 ;
        RECT 49.355 128.345 49.525 128.535 ;
        RECT 49.825 128.380 49.985 128.490 ;
        RECT 52.120 128.345 52.290 128.535 ;
        RECT 52.575 128.345 52.745 128.535 ;
        RECT 53.955 128.325 54.125 128.515 ;
        RECT 59.475 128.325 59.645 128.515 ;
        RECT 59.935 128.345 60.105 128.535 ;
        RECT 63.150 128.375 63.270 128.485 ;
        RECT 63.610 128.375 63.730 128.485 ;
        RECT 64.075 128.325 64.245 128.535 ;
        RECT 67.755 128.345 67.925 128.535 ;
        RECT 69.595 128.325 69.765 128.515 ;
        RECT 73.275 128.345 73.445 128.535 ;
        RECT 75.115 128.325 75.285 128.515 ;
        RECT 76.030 128.375 76.150 128.485 ;
        RECT 76.955 128.345 77.125 128.535 ;
        RECT 80.635 128.325 80.805 128.515 ;
        RECT 82.475 128.345 82.645 128.535 ;
        RECT 86.155 128.325 86.325 128.515 ;
        RECT 87.995 128.345 88.165 128.535 ;
        RECT 88.910 128.375 89.030 128.485 ;
        RECT 90.295 128.325 90.465 128.535 ;
        RECT 11.955 127.515 13.325 128.325 ;
        RECT 13.335 127.515 18.845 128.325 ;
        RECT 18.855 127.515 24.365 128.325 ;
        RECT 24.375 127.515 27.125 128.325 ;
        RECT 27.175 127.645 34.485 128.325 ;
        RECT 27.175 127.415 28.525 127.645 ;
        RECT 30.060 127.425 30.970 127.645 ;
        RECT 34.495 127.415 37.605 128.325 ;
        RECT 37.725 127.455 38.155 128.240 ;
        RECT 39.205 127.645 42.670 128.325 ;
        RECT 42.860 127.645 46.445 128.325 ;
        RECT 46.455 127.645 53.765 128.325 ;
        RECT 41.750 127.415 42.670 127.645 ;
        RECT 45.525 127.415 46.445 127.645 ;
        RECT 49.970 127.425 50.880 127.645 ;
        RECT 52.415 127.415 53.765 127.645 ;
        RECT 53.815 127.515 59.325 128.325 ;
        RECT 59.335 127.515 63.005 128.325 ;
        RECT 63.485 127.455 63.915 128.240 ;
        RECT 63.935 127.515 69.445 128.325 ;
        RECT 69.455 127.515 74.965 128.325 ;
        RECT 74.975 127.515 80.485 128.325 ;
        RECT 80.495 127.515 86.005 128.325 ;
        RECT 86.015 127.515 88.765 128.325 ;
        RECT 89.235 127.515 90.605 128.325 ;
      LAYER nwell ;
        RECT 11.760 124.295 90.800 127.125 ;
      LAYER pwell ;
        RECT 11.955 123.095 13.325 123.905 ;
        RECT 13.335 123.095 18.845 123.905 ;
        RECT 18.855 123.095 24.365 123.905 ;
        RECT 24.845 123.180 25.275 123.965 ;
        RECT 25.295 123.095 26.665 123.905 ;
        RECT 29.330 123.775 30.250 124.005 ;
        RECT 26.785 123.095 30.250 123.775 ;
        RECT 30.355 123.095 33.105 123.905 ;
        RECT 33.585 123.095 37.245 124.005 ;
        RECT 37.285 123.095 40.005 124.005 ;
        RECT 43.530 123.775 44.440 123.995 ;
        RECT 45.975 123.775 47.325 124.005 ;
        RECT 48.710 123.805 49.665 124.005 ;
        RECT 40.015 123.095 47.325 123.775 ;
        RECT 47.385 123.125 49.665 123.805 ;
        RECT 50.605 123.180 51.035 123.965 ;
        RECT 12.095 122.885 12.265 123.095 ;
        RECT 13.475 122.885 13.645 123.095 ;
        RECT 18.995 122.885 19.165 123.095 ;
        RECT 21.755 122.885 21.925 123.075 ;
        RECT 24.510 122.935 24.630 123.045 ;
        RECT 25.435 122.905 25.605 123.095 ;
        RECT 26.815 122.905 26.985 123.095 ;
        RECT 29.115 122.885 29.285 123.075 ;
        RECT 30.495 122.905 30.665 123.095 ;
        RECT 33.250 122.935 33.370 123.045 ;
        RECT 33.710 122.905 33.880 123.095 ;
        RECT 34.635 122.885 34.805 123.075 ;
        RECT 37.390 122.935 37.510 123.045 ;
        RECT 38.315 122.885 38.485 123.075 ;
        RECT 39.695 122.905 39.865 123.095 ;
        RECT 40.155 122.905 40.325 123.095 ;
        RECT 45.675 122.905 45.845 123.075 ;
        RECT 45.675 122.885 45.840 122.905 ;
        RECT 47.055 122.885 47.225 123.075 ;
        RECT 47.510 122.905 47.680 123.125 ;
        RECT 48.710 123.095 49.665 123.125 ;
        RECT 51.055 123.095 53.795 123.775 ;
        RECT 53.815 123.095 55.645 123.905 ;
        RECT 55.750 123.775 56.670 124.005 ;
        RECT 55.750 123.095 59.215 123.775 ;
        RECT 59.335 123.095 61.165 123.905 ;
        RECT 61.270 123.775 62.190 124.005 ;
        RECT 61.270 123.095 64.735 123.775 ;
        RECT 64.855 123.095 68.330 124.005 ;
        RECT 68.535 123.095 74.045 123.905 ;
        RECT 74.055 123.095 75.885 123.905 ;
        RECT 76.365 123.180 76.795 123.965 ;
        RECT 76.815 123.095 82.325 123.905 ;
        RECT 82.335 123.095 87.845 123.905 ;
        RECT 87.855 123.095 89.225 123.905 ;
        RECT 89.235 123.095 90.605 123.905 ;
        RECT 48.430 122.885 48.600 123.075 ;
        RECT 48.895 122.885 49.065 123.075 ;
        RECT 49.825 122.940 49.985 123.050 ;
        RECT 51.195 122.905 51.365 123.095 ;
        RECT 52.575 122.885 52.745 123.075 ;
        RECT 53.955 122.885 54.125 123.095 ;
        RECT 59.015 122.905 59.185 123.095 ;
        RECT 59.475 122.905 59.645 123.095 ;
        RECT 61.320 122.885 61.490 123.075 ;
        RECT 62.705 122.930 62.865 123.040 ;
        RECT 64.075 122.885 64.245 123.075 ;
        RECT 64.535 122.905 64.705 123.095 ;
        RECT 65.000 122.905 65.170 123.095 ;
        RECT 68.675 122.905 68.845 123.095 ;
        RECT 72.815 122.885 72.985 123.075 ;
        RECT 73.275 122.885 73.445 123.075 ;
        RECT 74.195 122.905 74.365 123.095 ;
        RECT 76.030 122.935 76.150 123.045 ;
        RECT 76.955 122.905 77.125 123.095 ;
        RECT 78.795 122.885 78.965 123.075 ;
        RECT 82.475 122.905 82.645 123.095 ;
        RECT 84.315 122.885 84.485 123.075 ;
        RECT 87.995 122.885 88.165 123.095 ;
        RECT 90.295 122.885 90.465 123.095 ;
        RECT 11.955 122.075 13.325 122.885 ;
        RECT 13.335 122.075 18.845 122.885 ;
        RECT 18.855 122.075 21.605 122.885 ;
        RECT 21.615 122.205 28.925 122.885 ;
        RECT 25.130 121.985 26.040 122.205 ;
        RECT 27.575 121.975 28.925 122.205 ;
        RECT 28.975 122.075 34.485 122.885 ;
        RECT 34.495 122.075 37.245 122.885 ;
        RECT 37.725 122.015 38.155 122.800 ;
        RECT 38.175 122.075 43.685 122.885 ;
        RECT 44.005 122.205 45.840 122.885 ;
        RECT 44.005 121.975 44.935 122.205 ;
        RECT 46.005 121.975 47.355 122.885 ;
        RECT 47.395 121.975 48.745 122.885 ;
        RECT 48.755 122.075 52.425 122.885 ;
        RECT 52.435 122.075 53.805 122.885 ;
        RECT 53.815 122.205 61.125 122.885 ;
        RECT 57.330 121.985 58.240 122.205 ;
        RECT 59.775 121.975 61.125 122.205 ;
        RECT 61.175 121.975 62.525 122.885 ;
        RECT 63.485 122.015 63.915 122.800 ;
        RECT 63.935 122.075 65.765 122.885 ;
        RECT 65.815 122.205 73.125 122.885 ;
        RECT 65.815 121.975 67.165 122.205 ;
        RECT 68.700 121.985 69.610 122.205 ;
        RECT 73.135 122.075 78.645 122.885 ;
        RECT 78.655 122.075 84.165 122.885 ;
        RECT 84.175 122.075 87.845 122.885 ;
        RECT 87.855 122.075 89.225 122.885 ;
        RECT 89.235 122.075 90.605 122.885 ;
        RECT 100.450 122.140 106.550 131.930 ;
        RECT 100.450 122.110 106.560 122.140 ;
        RECT 100.650 121.710 101.810 122.110 ;
      LAYER nwell ;
        RECT 11.760 118.855 90.800 121.685 ;
      LAYER pwell ;
        RECT 103.770 120.030 106.560 122.110 ;
        RECT 11.955 117.655 13.325 118.465 ;
        RECT 13.335 117.655 14.705 118.465 ;
        RECT 14.755 118.335 16.105 118.565 ;
        RECT 17.640 118.335 18.550 118.555 ;
        RECT 14.755 117.655 22.065 118.335 ;
        RECT 22.075 117.655 24.825 118.565 ;
        RECT 24.845 117.740 25.275 118.525 ;
        RECT 28.810 118.335 29.720 118.555 ;
        RECT 31.255 118.335 32.605 118.565 ;
        RECT 25.295 117.655 32.605 118.335 ;
        RECT 32.750 118.335 33.670 118.565 ;
        RECT 36.890 118.335 37.810 118.565 ;
        RECT 32.750 117.655 36.215 118.335 ;
        RECT 36.890 117.655 40.355 118.335 ;
        RECT 40.475 117.655 45.985 118.465 ;
        RECT 45.995 117.655 49.665 118.465 ;
        RECT 50.605 117.740 51.035 118.525 ;
        RECT 54.570 118.335 55.480 118.555 ;
        RECT 57.015 118.335 58.365 118.565 ;
        RECT 62.390 118.335 63.300 118.555 ;
        RECT 64.835 118.335 66.185 118.565 ;
        RECT 51.055 117.655 58.365 118.335 ;
        RECT 58.875 117.655 66.185 118.335 ;
        RECT 66.330 118.335 67.250 118.565 ;
        RECT 66.330 117.655 69.795 118.335 ;
        RECT 69.915 117.655 73.125 118.565 ;
        RECT 73.135 117.655 75.885 118.465 ;
        RECT 76.365 117.740 76.795 118.525 ;
        RECT 76.815 117.655 82.325 118.465 ;
        RECT 82.335 117.655 87.845 118.465 ;
        RECT 87.855 117.655 89.225 118.465 ;
        RECT 89.235 117.655 90.605 118.465 ;
      LAYER nwell ;
        RECT 101.660 117.920 106.500 120.030 ;
        RECT 107.780 119.690 117.970 131.940 ;
      LAYER pwell ;
        RECT 120.330 122.200 126.430 131.990 ;
        RECT 120.330 122.170 126.440 122.200 ;
        RECT 120.530 121.770 121.690 122.170 ;
        RECT 123.650 120.090 126.440 122.170 ;
      LAYER nwell ;
        RECT 121.540 117.980 126.380 120.090 ;
        RECT 127.660 119.750 137.850 132.000 ;
      LAYER pwell ;
        RECT 140.360 122.200 146.460 131.990 ;
        RECT 140.360 122.170 146.470 122.200 ;
        RECT 140.560 121.770 141.720 122.170 ;
        RECT 143.680 120.090 146.470 122.170 ;
      LAYER nwell ;
        RECT 141.570 117.980 146.410 120.090 ;
        RECT 147.690 119.750 157.880 132.000 ;
      LAYER pwell ;
        RECT 12.095 117.445 12.265 117.655 ;
        RECT 13.475 117.445 13.645 117.655 ;
        RECT 15.315 117.445 15.485 117.635 ;
        RECT 20.835 117.445 21.005 117.635 ;
        RECT 21.755 117.465 21.925 117.655 ;
        RECT 22.215 117.465 22.385 117.655 ;
        RECT 22.675 117.445 22.845 117.635 ;
        RECT 25.435 117.465 25.605 117.655 ;
        RECT 26.355 117.445 26.525 117.635 ;
        RECT 30.035 117.445 30.205 117.635 ;
        RECT 30.500 117.445 30.670 117.635 ;
        RECT 31.875 117.445 32.045 117.635 ;
        RECT 34.640 117.445 34.810 117.635 ;
        RECT 36.015 117.465 36.185 117.655 ;
        RECT 36.470 117.495 36.590 117.605 ;
        RECT 38.310 117.495 38.430 117.605 ;
        RECT 39.700 117.445 39.870 117.635 ;
        RECT 40.155 117.445 40.325 117.655 ;
        RECT 40.615 117.465 40.785 117.655 ;
        RECT 43.830 117.445 44.000 117.635 ;
        RECT 46.135 117.465 46.305 117.655 ;
        RECT 48.435 117.445 48.605 117.635 ;
        RECT 48.895 117.445 49.065 117.635 ;
        RECT 49.825 117.500 49.985 117.610 ;
        RECT 51.195 117.465 51.365 117.655 ;
        RECT 56.255 117.445 56.425 117.635 ;
        RECT 58.550 117.495 58.670 117.605 ;
        RECT 59.015 117.465 59.185 117.655 ;
        RECT 61.775 117.445 61.945 117.635 ;
        RECT 64.070 117.495 64.190 117.605 ;
        RECT 65.460 117.445 65.630 117.635 ;
        RECT 65.915 117.445 66.085 117.635 ;
        RECT 67.300 117.445 67.470 117.635 ;
        RECT 68.675 117.445 68.845 117.635 ;
        RECT 69.595 117.465 69.765 117.655 ;
        RECT 70.055 117.465 70.225 117.655 ;
        RECT 70.510 117.495 70.630 117.605 ;
        RECT 70.975 117.445 71.145 117.635 ;
        RECT 73.275 117.465 73.445 117.655 ;
        RECT 73.735 117.445 73.905 117.635 ;
        RECT 76.030 117.495 76.150 117.605 ;
        RECT 76.955 117.465 77.125 117.655 ;
        RECT 79.255 117.445 79.425 117.635 ;
        RECT 82.475 117.465 82.645 117.655 ;
        RECT 84.775 117.445 84.945 117.635 ;
        RECT 87.535 117.445 87.705 117.635 ;
        RECT 87.995 117.465 88.165 117.655 ;
        RECT 90.295 117.445 90.465 117.655 ;
        RECT 11.955 116.635 13.325 117.445 ;
        RECT 13.335 116.765 15.165 117.445 ;
        RECT 15.175 116.635 20.685 117.445 ;
        RECT 20.695 116.635 22.525 117.445 ;
        RECT 22.550 116.535 24.365 117.445 ;
        RECT 24.375 116.765 26.665 117.445 ;
        RECT 26.770 116.765 30.235 117.445 ;
        RECT 24.375 116.535 25.295 116.765 ;
        RECT 26.770 116.535 27.690 116.765 ;
        RECT 30.355 116.535 31.705 117.445 ;
        RECT 31.735 116.635 34.485 117.445 ;
        RECT 34.495 116.535 37.415 117.445 ;
        RECT 37.725 116.575 38.155 117.360 ;
        RECT 38.635 116.535 39.985 117.445 ;
        RECT 40.125 116.765 43.590 117.445 ;
        RECT 42.670 116.535 43.590 116.765 ;
        RECT 43.715 116.535 45.065 117.445 ;
        RECT 45.170 116.765 48.635 117.445 ;
        RECT 48.755 116.765 56.065 117.445 ;
        RECT 45.170 116.535 46.090 116.765 ;
        RECT 52.270 116.545 53.180 116.765 ;
        RECT 54.715 116.535 56.065 116.765 ;
        RECT 56.115 116.635 61.625 117.445 ;
        RECT 61.635 116.635 63.465 117.445 ;
        RECT 63.485 116.575 63.915 117.360 ;
        RECT 64.395 116.535 65.745 117.445 ;
        RECT 65.775 116.635 67.145 117.445 ;
        RECT 67.155 116.535 68.505 117.445 ;
        RECT 68.535 116.635 70.365 117.445 ;
        RECT 70.835 116.765 73.585 117.445 ;
        RECT 72.655 116.535 73.585 116.765 ;
        RECT 73.595 116.635 79.105 117.445 ;
        RECT 79.115 116.635 84.625 117.445 ;
        RECT 84.635 116.635 87.385 117.445 ;
        RECT 87.395 116.765 89.225 117.445 ;
        RECT 87.880 116.535 89.225 116.765 ;
        RECT 89.235 116.635 90.605 117.445 ;
      LAYER nwell ;
        RECT 11.760 113.415 90.800 116.245 ;
      LAYER pwell ;
        RECT 11.955 112.215 13.325 113.025 ;
        RECT 13.995 112.895 17.925 113.125 ;
        RECT 13.510 112.215 17.925 112.895 ;
        RECT 18.030 112.895 18.950 113.125 ;
        RECT 18.030 112.215 21.495 112.895 ;
        RECT 21.615 112.215 24.365 113.025 ;
        RECT 24.845 112.300 25.275 113.085 ;
        RECT 25.295 112.215 30.805 113.025 ;
        RECT 30.815 112.215 32.645 113.025 ;
        RECT 36.630 112.895 37.540 113.115 ;
        RECT 39.075 112.895 40.425 113.125 ;
        RECT 33.115 112.215 40.425 112.895 ;
        RECT 40.485 112.215 43.215 113.125 ;
        RECT 46.750 112.895 47.660 113.115 ;
        RECT 49.195 112.895 50.545 113.125 ;
        RECT 43.235 112.215 50.545 112.895 ;
        RECT 50.605 112.300 51.035 113.085 ;
        RECT 51.055 112.215 53.805 113.025 ;
        RECT 53.815 112.925 54.745 113.125 ;
        RECT 56.075 112.925 57.025 113.125 ;
        RECT 53.815 112.445 57.025 112.925 ;
        RECT 60.550 112.895 61.460 113.115 ;
        RECT 62.995 112.895 64.345 113.125 ;
        RECT 53.960 112.245 57.025 112.445 ;
        RECT 12.095 112.005 12.265 112.215 ;
        RECT 13.510 112.195 13.620 112.215 ;
        RECT 13.450 112.025 13.645 112.195 ;
        RECT 13.475 112.005 13.645 112.025 ;
        RECT 14.860 112.005 15.030 112.195 ;
        RECT 16.695 112.005 16.865 112.195 ;
        RECT 20.375 112.005 20.545 112.195 ;
        RECT 21.295 112.025 21.465 112.215 ;
        RECT 21.755 112.025 21.925 112.215 ;
        RECT 24.510 112.055 24.630 112.165 ;
        RECT 25.435 112.025 25.605 112.215 ;
        RECT 27.740 112.005 27.910 112.195 ;
        RECT 29.125 112.050 29.285 112.160 ;
        RECT 30.035 112.005 30.205 112.195 ;
        RECT 30.955 112.025 31.125 112.215 ;
        RECT 32.790 112.055 32.910 112.165 ;
        RECT 33.255 112.025 33.425 112.215 ;
        RECT 37.390 112.055 37.510 112.165 ;
        RECT 11.955 111.195 13.325 112.005 ;
        RECT 13.335 111.195 14.705 112.005 ;
        RECT 14.715 111.095 16.545 112.005 ;
        RECT 16.665 111.325 20.130 112.005 ;
        RECT 20.235 111.325 27.545 112.005 ;
        RECT 19.210 111.095 20.130 111.325 ;
        RECT 23.750 111.105 24.660 111.325 ;
        RECT 26.195 111.095 27.545 111.325 ;
        RECT 27.595 111.095 28.945 112.005 ;
        RECT 29.895 111.325 37.205 112.005 ;
        RECT 38.310 111.975 38.480 112.195 ;
        RECT 40.615 112.165 40.785 112.215 ;
        RECT 43.375 112.195 43.545 112.215 ;
        RECT 40.610 112.055 40.785 112.165 ;
        RECT 40.615 112.025 40.785 112.055 ;
        RECT 41.075 112.025 41.245 112.195 ;
        RECT 43.375 112.025 43.550 112.195 ;
        RECT 41.080 112.005 41.245 112.025 ;
        RECT 43.380 112.005 43.550 112.025 ;
        RECT 45.215 112.005 45.385 112.195 ;
        RECT 46.595 112.005 46.765 112.195 ;
        RECT 51.195 112.025 51.365 112.215 ;
        RECT 52.115 112.005 52.285 112.195 ;
        RECT 53.960 112.165 54.130 112.245 ;
        RECT 56.090 112.215 57.025 112.245 ;
        RECT 57.035 112.215 64.345 112.895 ;
        RECT 64.395 112.215 65.745 113.125 ;
        RECT 65.775 112.215 67.145 113.025 ;
        RECT 67.165 112.215 68.515 113.125 ;
        RECT 68.575 112.895 69.925 113.125 ;
        RECT 71.460 112.895 72.370 113.115 ;
        RECT 68.575 112.215 75.885 112.895 ;
        RECT 76.365 112.300 76.795 113.085 ;
        RECT 76.815 112.215 82.325 113.025 ;
        RECT 82.335 112.215 86.005 113.025 ;
        RECT 86.015 112.215 87.385 112.995 ;
        RECT 87.880 112.895 89.225 113.125 ;
        RECT 87.395 112.215 89.225 112.895 ;
        RECT 89.235 112.215 90.605 113.025 ;
        RECT 53.950 112.055 54.130 112.165 ;
        RECT 53.960 112.025 54.130 112.055 ;
        RECT 54.420 112.005 54.590 112.195 ;
        RECT 57.175 112.025 57.345 112.215 ;
        RECT 58.555 112.005 58.725 112.195 ;
        RECT 60.390 112.055 60.510 112.165 ;
        RECT 63.155 112.005 63.325 112.195 ;
        RECT 64.075 112.005 64.245 112.195 ;
        RECT 64.540 112.025 64.710 112.215 ;
        RECT 65.915 112.025 66.085 112.215 ;
        RECT 67.765 112.050 67.925 112.160 ;
        RECT 68.215 112.025 68.385 112.215 ;
        RECT 71.895 112.005 72.065 112.195 ;
        RECT 72.355 112.005 72.525 112.195 ;
        RECT 74.655 112.005 74.825 112.195 ;
        RECT 75.575 112.025 75.745 112.215 ;
        RECT 76.030 112.055 76.150 112.165 ;
        RECT 76.955 112.025 77.125 112.215 ;
        RECT 78.335 112.005 78.505 112.195 ;
        RECT 82.475 112.025 82.645 112.215 ;
        RECT 86.155 112.025 86.325 112.215 ;
        RECT 87.535 112.025 87.705 112.215 ;
        RECT 88.915 112.005 89.085 112.195 ;
        RECT 90.295 112.005 90.465 112.215 ;
        RECT 39.510 111.975 40.465 112.005 ;
        RECT 33.410 111.105 34.320 111.325 ;
        RECT 35.855 111.095 37.205 111.325 ;
        RECT 37.725 111.135 38.155 111.920 ;
        RECT 38.185 111.295 40.465 111.975 ;
        RECT 41.080 111.325 42.915 112.005 ;
        RECT 39.510 111.095 40.465 111.295 ;
        RECT 41.985 111.095 42.915 111.325 ;
        RECT 43.235 111.095 45.065 112.005 ;
        RECT 45.085 111.095 46.435 112.005 ;
        RECT 46.455 111.195 51.965 112.005 ;
        RECT 51.975 111.195 53.805 112.005 ;
        RECT 54.275 111.325 58.370 112.005 ;
        RECT 54.760 111.095 58.370 111.325 ;
        RECT 58.415 111.195 60.245 112.005 ;
        RECT 60.715 111.095 63.465 112.005 ;
        RECT 63.485 111.135 63.915 111.920 ;
        RECT 63.935 111.325 67.605 112.005 ;
        RECT 66.675 111.095 67.605 111.325 ;
        RECT 68.630 111.325 72.095 112.005 ;
        RECT 68.630 111.095 69.550 111.325 ;
        RECT 72.215 111.095 74.505 112.005 ;
        RECT 74.515 111.195 78.185 112.005 ;
        RECT 78.195 111.325 85.505 112.005 ;
        RECT 81.710 111.105 82.620 111.325 ;
        RECT 84.155 111.095 85.505 111.325 ;
        RECT 85.650 111.325 89.115 112.005 ;
        RECT 85.650 111.095 86.570 111.325 ;
        RECT 89.235 111.195 90.605 112.005 ;
      LAYER nwell ;
        RECT 11.760 107.975 90.800 110.805 ;
      LAYER pwell ;
        RECT 11.955 106.775 13.325 107.585 ;
        RECT 16.850 107.455 17.760 107.675 ;
        RECT 19.295 107.455 20.645 107.685 ;
        RECT 13.335 106.775 20.645 107.455 ;
        RECT 20.695 106.775 22.525 107.685 ;
        RECT 22.845 107.455 23.775 107.685 ;
        RECT 22.845 106.775 24.680 107.455 ;
        RECT 24.845 106.860 25.275 107.645 ;
        RECT 27.585 107.485 28.940 107.685 ;
        RECT 26.260 107.455 28.940 107.485 ;
        RECT 29.435 107.485 30.390 107.685 ;
        RECT 26.260 106.805 29.425 107.455 ;
        RECT 27.585 106.775 29.425 106.805 ;
        RECT 29.435 106.805 31.715 107.485 ;
        RECT 29.435 106.775 30.390 106.805 ;
        RECT 12.095 106.565 12.265 106.775 ;
        RECT 13.475 106.725 13.645 106.775 ;
        RECT 13.470 106.615 13.645 106.725 ;
        RECT 13.475 106.585 13.645 106.615 ;
        RECT 13.940 106.565 14.110 106.755 ;
        RECT 18.995 106.565 19.165 106.755 ;
        RECT 19.465 106.610 19.625 106.720 ;
        RECT 20.370 106.565 20.540 106.755 ;
        RECT 20.840 106.585 21.010 106.775 ;
        RECT 24.515 106.755 24.680 106.775 ;
        RECT 21.765 106.565 21.935 106.755 ;
        RECT 23.130 106.615 23.250 106.725 ;
        RECT 24.515 106.585 24.685 106.755 ;
        RECT 24.970 106.565 25.140 106.755 ;
        RECT 25.435 106.565 25.605 106.755 ;
        RECT 29.115 106.585 29.285 106.775 ;
        RECT 30.035 106.565 30.205 106.755 ;
        RECT 30.495 106.565 30.665 106.755 ;
        RECT 31.420 106.585 31.590 106.805 ;
        RECT 31.735 106.775 33.565 107.585 ;
        RECT 34.055 106.775 35.405 107.685 ;
        RECT 35.415 107.485 36.360 107.685 ;
        RECT 37.695 107.485 38.625 107.685 ;
        RECT 35.415 107.005 38.625 107.485 ;
        RECT 38.730 107.455 39.650 107.685 ;
        RECT 43.455 107.595 44.405 107.685 ;
        RECT 35.415 106.805 38.485 107.005 ;
        RECT 35.415 106.775 36.360 106.805 ;
        RECT 31.875 106.585 32.045 106.775 ;
        RECT 33.710 106.615 33.830 106.725 ;
        RECT 34.170 106.585 34.340 106.775 ;
        RECT 38.315 106.585 38.485 106.805 ;
        RECT 38.730 106.775 42.195 107.455 ;
        RECT 42.475 106.775 44.405 107.595 ;
        RECT 44.615 106.775 48.285 107.585 ;
        RECT 49.665 107.455 50.585 107.685 ;
        RECT 48.295 106.775 50.585 107.455 ;
        RECT 50.605 106.860 51.035 107.645 ;
        RECT 51.055 106.775 60.160 107.455 ;
        RECT 60.255 106.775 63.925 107.585 ;
        RECT 64.865 106.775 66.215 107.685 ;
        RECT 66.235 106.775 67.605 107.585 ;
        RECT 67.615 107.485 68.565 107.685 ;
        RECT 69.895 107.485 70.825 107.685 ;
        RECT 72.170 107.485 73.125 107.685 ;
        RECT 67.615 107.005 70.825 107.485 ;
        RECT 67.615 106.805 70.680 107.005 ;
        RECT 70.845 106.805 73.125 107.485 ;
        RECT 67.615 106.775 68.550 106.805 ;
        RECT 41.995 106.755 42.165 106.775 ;
        RECT 42.475 106.755 42.625 106.775 ;
        RECT 40.615 106.565 40.785 106.755 ;
        RECT 41.990 106.585 42.165 106.755 ;
        RECT 41.990 106.565 42.160 106.585 ;
        RECT 42.455 106.565 42.625 106.755 ;
        RECT 44.755 106.585 44.925 106.775 ;
        RECT 48.435 106.585 48.605 106.775 ;
        RECT 49.825 106.610 49.985 106.720 ;
        RECT 51.195 106.585 51.365 106.775 ;
        RECT 53.955 106.565 54.125 106.755 ;
        RECT 54.410 106.615 54.530 106.725 ;
        RECT 54.875 106.565 55.045 106.755 ;
        RECT 57.175 106.565 57.345 106.755 ;
        RECT 60.395 106.585 60.565 106.775 ;
        RECT 60.855 106.565 61.025 106.755 ;
        RECT 64.080 106.565 64.250 106.755 ;
        RECT 64.995 106.585 65.165 106.775 ;
        RECT 65.915 106.565 66.085 106.755 ;
        RECT 66.375 106.585 66.545 106.775 ;
        RECT 70.510 106.585 70.680 106.805 ;
        RECT 70.970 106.585 71.140 106.805 ;
        RECT 72.170 106.775 73.125 106.805 ;
        RECT 73.135 106.775 75.325 107.685 ;
        RECT 76.365 106.860 76.795 107.645 ;
        RECT 76.815 107.005 78.650 107.685 ;
        RECT 76.960 106.775 78.650 107.005 ;
        RECT 79.115 106.775 80.485 107.585 ;
        RECT 80.495 107.455 81.425 107.685 ;
        RECT 80.495 106.775 84.395 107.455 ;
        RECT 84.635 106.775 86.005 107.585 ;
        RECT 86.015 106.775 87.385 107.555 ;
        RECT 87.395 106.775 89.225 107.585 ;
        RECT 89.235 106.775 90.605 107.585 ;
        RECT 100.400 107.200 106.500 116.990 ;
        RECT 100.400 107.170 106.510 107.200 ;
        RECT 71.430 106.615 71.550 106.725 ;
        RECT 71.900 106.565 72.070 106.755 ;
        RECT 73.280 106.585 73.450 106.775 ;
        RECT 75.585 106.620 75.745 106.730 ;
        RECT 76.960 106.585 77.130 106.775 ;
        RECT 77.410 106.565 77.580 106.755 ;
        RECT 79.255 106.565 79.425 106.775 ;
        RECT 79.715 106.565 79.885 106.755 ;
        RECT 80.910 106.585 81.080 106.775 ;
        RECT 83.395 106.565 83.565 106.755 ;
        RECT 84.775 106.585 84.945 106.775 ;
        RECT 86.155 106.585 86.325 106.775 ;
        RECT 87.535 106.585 87.705 106.775 ;
        RECT 87.995 106.565 88.165 106.755 ;
        RECT 88.465 106.610 88.625 106.720 ;
        RECT 90.295 106.565 90.465 106.775 ;
        RECT 100.600 106.770 101.760 107.170 ;
        RECT 11.955 105.755 13.325 106.565 ;
        RECT 13.795 105.655 17.465 106.565 ;
        RECT 17.475 105.885 19.305 106.565 ;
        RECT 17.475 105.655 18.820 105.885 ;
        RECT 20.255 105.655 21.605 106.565 ;
        RECT 21.615 105.785 22.985 106.565 ;
        RECT 23.455 105.655 25.285 106.565 ;
        RECT 25.295 105.755 26.665 106.565 ;
        RECT 26.770 105.885 30.235 106.565 ;
        RECT 30.355 105.885 37.665 106.565 ;
        RECT 26.770 105.655 27.690 105.885 ;
        RECT 33.870 105.665 34.780 105.885 ;
        RECT 36.315 105.655 37.665 105.885 ;
        RECT 37.725 105.695 38.155 106.480 ;
        RECT 38.185 105.655 40.915 106.565 ;
        RECT 40.955 105.655 42.305 106.565 ;
        RECT 42.315 105.885 49.625 106.565 ;
        RECT 45.830 105.665 46.740 105.885 ;
        RECT 48.275 105.655 49.625 105.885 ;
        RECT 50.690 105.885 54.155 106.565 ;
        RECT 54.735 105.885 57.025 106.565 ;
        RECT 57.145 105.885 60.610 106.565 ;
        RECT 50.690 105.655 51.610 105.885 ;
        RECT 56.105 105.655 57.025 105.885 ;
        RECT 59.690 105.655 60.610 105.885 ;
        RECT 60.715 105.755 63.465 106.565 ;
        RECT 63.485 105.695 63.915 106.480 ;
        RECT 63.935 105.655 65.765 106.565 ;
        RECT 65.775 105.755 71.285 106.565 ;
        RECT 71.755 105.885 74.030 106.565 ;
        RECT 72.660 105.655 74.030 105.885 ;
        RECT 74.250 105.655 77.725 106.565 ;
        RECT 77.735 105.885 79.565 106.565 ;
        RECT 77.735 105.655 79.080 105.885 ;
        RECT 79.575 105.755 83.245 106.565 ;
        RECT 83.255 105.755 84.625 106.565 ;
        RECT 84.730 105.885 88.195 106.565 ;
        RECT 84.730 105.655 85.650 105.885 ;
        RECT 89.235 105.755 90.605 106.565 ;
      LAYER nwell ;
        RECT 11.760 102.535 90.800 105.365 ;
      LAYER pwell ;
        RECT 103.720 105.090 106.510 107.170 ;
      LAYER nwell ;
        RECT 101.610 102.980 106.450 105.090 ;
        RECT 107.730 104.750 117.920 117.000 ;
      LAYER pwell ;
        RECT 120.330 107.200 126.430 116.990 ;
        RECT 120.330 107.170 126.440 107.200 ;
        RECT 120.530 106.770 121.690 107.170 ;
        RECT 123.650 105.090 126.440 107.170 ;
      LAYER nwell ;
        RECT 121.540 102.980 126.380 105.090 ;
        RECT 127.660 104.750 137.850 117.000 ;
      LAYER pwell ;
        RECT 140.360 107.200 146.460 116.990 ;
        RECT 140.360 107.170 146.470 107.200 ;
        RECT 140.560 106.770 141.720 107.170 ;
        RECT 143.680 105.090 146.470 107.170 ;
      LAYER nwell ;
        RECT 141.570 102.980 146.410 105.090 ;
        RECT 147.690 104.750 157.880 117.000 ;
      LAYER pwell ;
        RECT 11.955 101.335 13.325 102.145 ;
        RECT 13.335 101.335 15.165 102.015 ;
        RECT 16.115 101.335 17.465 102.245 ;
        RECT 20.130 102.015 21.050 102.245 ;
        RECT 17.585 101.335 21.050 102.015 ;
        RECT 21.715 101.335 24.825 102.245 ;
        RECT 24.845 101.420 25.275 102.205 ;
        RECT 28.810 102.015 29.720 102.235 ;
        RECT 31.255 102.015 32.605 102.245 ;
        RECT 25.295 101.335 32.605 102.015 ;
        RECT 32.655 101.335 36.325 102.145 ;
        RECT 36.795 101.335 38.145 102.245 ;
        RECT 38.635 101.335 41.845 102.245 ;
        RECT 41.855 101.335 45.355 102.245 ;
        RECT 45.535 101.335 49.205 102.145 ;
        RECT 49.225 101.335 50.575 102.245 ;
        RECT 50.605 101.420 51.035 102.205 ;
        RECT 52.015 102.015 53.365 102.245 ;
        RECT 54.900 102.015 55.810 102.235 ;
        RECT 59.335 102.015 60.265 102.245 ;
        RECT 63.960 102.015 65.305 102.245 ;
        RECT 52.015 101.335 59.325 102.015 ;
        RECT 59.335 101.335 63.235 102.015 ;
        RECT 63.475 101.335 65.305 102.015 ;
        RECT 65.315 101.335 66.665 102.245 ;
        RECT 66.695 101.335 70.365 102.145 ;
        RECT 71.295 101.335 72.645 102.245 ;
        RECT 72.675 101.335 75.885 102.245 ;
        RECT 76.365 101.420 76.795 102.205 ;
        RECT 76.815 101.335 78.645 102.145 ;
        RECT 82.630 102.015 83.540 102.235 ;
        RECT 85.075 102.015 86.425 102.245 ;
        RECT 79.115 101.335 86.425 102.015 ;
        RECT 86.475 101.335 89.225 102.145 ;
        RECT 89.235 101.335 90.605 102.145 ;
        RECT 12.095 101.125 12.265 101.335 ;
        RECT 13.475 101.125 13.645 101.335 ;
        RECT 15.325 101.180 15.485 101.290 ;
        RECT 16.230 101.145 16.400 101.335 ;
        RECT 17.615 101.145 17.785 101.335 ;
        RECT 21.290 101.175 21.410 101.285 ;
        RECT 21.755 101.145 21.925 101.335 ;
        RECT 24.055 101.125 24.225 101.315 ;
        RECT 24.510 101.125 24.680 101.315 ;
        RECT 25.435 101.145 25.605 101.335 ;
        RECT 25.895 101.125 26.065 101.315 ;
        RECT 31.415 101.125 31.585 101.315 ;
        RECT 32.795 101.145 32.965 101.335 ;
        RECT 36.470 101.175 36.590 101.285 ;
        RECT 36.945 101.170 37.105 101.280 ;
        RECT 37.860 101.145 38.030 101.335 ;
        RECT 38.315 101.285 38.485 101.315 ;
        RECT 38.310 101.175 38.485 101.285 ;
        RECT 38.315 101.125 38.485 101.175 ;
        RECT 38.765 101.145 38.935 101.335 ;
        RECT 45.220 101.315 45.355 101.335 ;
        RECT 41.070 101.175 41.190 101.285 ;
        RECT 41.810 101.125 41.980 101.315 ;
        RECT 45.220 101.145 45.390 101.315 ;
        RECT 45.675 101.125 45.845 101.335 ;
        RECT 50.275 101.145 50.445 101.335 ;
        RECT 51.205 101.180 51.365 101.290 ;
        RECT 55.790 101.125 55.960 101.315 ;
        RECT 56.255 101.125 56.425 101.315 ;
        RECT 59.015 101.145 59.185 101.335 ;
        RECT 59.750 101.145 59.920 101.335 ;
        RECT 63.615 101.145 63.785 101.335 ;
        RECT 64.350 101.125 64.520 101.315 ;
        RECT 65.460 101.145 65.630 101.335 ;
        RECT 66.835 101.145 67.005 101.335 ;
        RECT 68.215 101.125 68.385 101.315 ;
        RECT 70.050 101.175 70.170 101.285 ;
        RECT 70.525 101.180 70.685 101.290 ;
        RECT 72.360 101.145 72.530 101.335 ;
        RECT 75.575 101.315 75.745 101.335 ;
        RECT 73.275 101.125 73.445 101.315 ;
        RECT 75.570 101.145 75.745 101.315 ;
        RECT 76.030 101.175 76.150 101.285 ;
        RECT 76.955 101.145 77.125 101.335 ;
        RECT 75.570 101.125 75.740 101.145 ;
        RECT 11.955 100.315 13.325 101.125 ;
        RECT 13.335 100.445 20.645 101.125 ;
        RECT 16.850 100.225 17.760 100.445 ;
        RECT 19.295 100.215 20.645 100.445 ;
        RECT 20.695 100.445 24.365 101.125 ;
        RECT 20.695 100.215 21.625 100.445 ;
        RECT 24.395 100.215 25.745 101.125 ;
        RECT 25.755 100.315 31.265 101.125 ;
        RECT 31.275 100.315 36.785 101.125 ;
        RECT 37.725 100.255 38.155 101.040 ;
        RECT 38.175 100.315 40.925 101.125 ;
        RECT 41.395 100.445 45.295 101.125 ;
        RECT 45.535 100.445 52.845 101.125 ;
        RECT 41.395 100.215 42.325 100.445 ;
        RECT 49.050 100.225 49.960 100.445 ;
        RECT 51.495 100.215 52.845 100.445 ;
        RECT 52.990 100.215 56.105 101.125 ;
        RECT 56.115 100.445 63.425 101.125 ;
        RECT 59.630 100.225 60.540 100.445 ;
        RECT 62.075 100.215 63.425 100.445 ;
        RECT 63.485 100.255 63.915 101.040 ;
        RECT 63.935 100.445 67.835 101.125 ;
        RECT 63.935 100.215 64.865 100.445 ;
        RECT 68.075 100.315 69.905 101.125 ;
        RECT 70.505 100.215 73.505 101.125 ;
        RECT 73.675 100.215 75.885 101.125 ;
        RECT 75.895 101.095 76.850 101.125 ;
        RECT 77.880 101.095 78.050 101.315 ;
        RECT 78.340 101.125 78.510 101.315 ;
        RECT 78.790 101.175 78.910 101.285 ;
        RECT 79.255 101.145 79.425 101.335 ;
        RECT 80.630 101.175 80.750 101.285 ;
        RECT 81.370 101.125 81.540 101.315 ;
        RECT 85.235 101.125 85.405 101.315 ;
        RECT 86.615 101.145 86.785 101.335 ;
        RECT 88.910 101.175 89.030 101.285 ;
        RECT 90.295 101.125 90.465 101.335 ;
        RECT 75.895 100.415 78.175 101.095 ;
        RECT 78.195 100.445 80.470 101.125 ;
        RECT 75.895 100.215 76.850 100.415 ;
        RECT 79.100 100.215 80.470 100.445 ;
        RECT 80.955 100.445 84.855 101.125 ;
        RECT 80.955 100.215 81.885 100.445 ;
        RECT 85.095 100.315 88.765 101.125 ;
        RECT 89.235 100.315 90.605 101.125 ;
      LAYER nwell ;
        RECT 11.760 97.095 90.800 99.925 ;
      LAYER pwell ;
        RECT 11.955 95.895 13.325 96.705 ;
        RECT 13.335 95.895 17.005 96.705 ;
        RECT 17.015 95.895 18.845 96.805 ;
        RECT 18.950 96.575 19.870 96.805 ;
        RECT 18.950 95.895 22.415 96.575 ;
        RECT 22.535 95.895 24.365 96.705 ;
        RECT 24.845 95.980 25.275 96.765 ;
        RECT 25.295 95.895 30.805 96.705 ;
        RECT 30.815 95.895 32.645 96.705 ;
        RECT 36.170 96.575 37.080 96.795 ;
        RECT 38.615 96.575 39.965 96.805 ;
        RECT 32.655 95.895 39.965 96.575 ;
        RECT 40.110 96.575 41.030 96.805 ;
        RECT 40.110 95.895 43.575 96.575 ;
        RECT 43.695 95.895 46.445 96.705 ;
        RECT 46.455 96.575 47.385 96.805 ;
        RECT 46.455 95.895 50.355 96.575 ;
        RECT 50.605 95.980 51.035 96.765 ;
        RECT 51.055 96.575 51.985 96.805 ;
        RECT 51.055 95.895 54.955 96.575 ;
        RECT 55.195 95.895 58.865 96.705 ;
        RECT 58.875 95.895 60.245 96.705 ;
        RECT 62.910 96.575 63.830 96.805 ;
        RECT 60.365 95.895 63.830 96.575 ;
        RECT 63.935 95.895 65.765 96.705 ;
        RECT 65.775 96.575 66.695 96.805 ;
        RECT 65.775 95.895 68.065 96.575 ;
        RECT 68.075 95.895 69.425 96.805 ;
        RECT 69.455 95.895 72.205 96.705 ;
        RECT 74.010 96.605 74.965 96.805 ;
        RECT 72.685 95.925 74.965 96.605 ;
        RECT 12.095 95.685 12.265 95.895 ;
        RECT 13.475 95.685 13.645 95.895 ;
        RECT 15.130 95.685 15.300 95.875 ;
        RECT 17.160 95.705 17.330 95.895 ;
        RECT 18.990 95.735 19.110 95.845 ;
        RECT 11.955 94.875 13.325 95.685 ;
        RECT 13.335 94.875 14.705 95.685 ;
        RECT 14.715 95.005 18.615 95.685 ;
        RECT 19.455 95.655 19.625 95.875 ;
        RECT 22.215 95.685 22.385 95.895 ;
        RECT 22.675 95.705 22.845 95.895 ;
        RECT 24.510 95.735 24.630 95.845 ;
        RECT 24.975 95.685 25.145 95.875 ;
        RECT 25.435 95.705 25.605 95.895 ;
        RECT 30.955 95.705 31.125 95.895 ;
        RECT 32.795 95.705 32.965 95.895 ;
        RECT 33.990 95.685 34.160 95.875 ;
        RECT 38.310 95.735 38.430 95.845 ;
        RECT 39.050 95.685 39.220 95.875 ;
        RECT 42.915 95.685 43.085 95.875 ;
        RECT 43.375 95.705 43.545 95.895 ;
        RECT 43.835 95.705 44.005 95.895 ;
        RECT 45.215 95.685 45.385 95.875 ;
        RECT 46.870 95.705 47.040 95.895 ;
        RECT 50.735 95.685 50.905 95.875 ;
        RECT 51.470 95.705 51.640 95.895 ;
        RECT 53.490 95.735 53.610 95.845 ;
        RECT 55.335 95.705 55.505 95.895 ;
        RECT 59.015 95.705 59.185 95.895 ;
        RECT 60.395 95.705 60.565 95.895 ;
        RECT 60.855 95.685 61.025 95.875 ;
        RECT 61.315 95.685 61.485 95.875 ;
        RECT 63.150 95.735 63.270 95.845 ;
        RECT 64.075 95.705 64.245 95.895 ;
        RECT 67.755 95.875 67.925 95.895 ;
        RECT 66.835 95.685 67.005 95.875 ;
        RECT 67.290 95.735 67.410 95.845 ;
        RECT 67.745 95.705 67.925 95.875 ;
        RECT 68.220 95.705 68.390 95.895 ;
        RECT 69.595 95.705 69.765 95.895 ;
        RECT 67.745 95.685 67.915 95.705 ;
        RECT 70.975 95.685 71.145 95.875 ;
        RECT 72.350 95.735 72.470 95.845 ;
        RECT 20.655 95.655 22.035 95.685 ;
        RECT 14.715 94.775 15.645 95.005 ;
        RECT 19.330 94.975 22.035 95.655 ;
        RECT 20.655 94.775 22.035 94.975 ;
        RECT 22.075 94.875 24.825 95.685 ;
        RECT 24.835 95.005 32.565 95.685 ;
        RECT 28.350 94.785 29.260 95.005 ;
        RECT 30.795 94.775 32.565 95.005 ;
        RECT 33.575 95.005 37.475 95.685 ;
        RECT 33.575 94.775 34.505 95.005 ;
        RECT 37.725 94.815 38.155 95.600 ;
        RECT 38.635 95.005 42.535 95.685 ;
        RECT 42.775 95.005 45.065 95.685 ;
        RECT 38.635 94.775 39.565 95.005 ;
        RECT 44.145 94.775 45.065 95.005 ;
        RECT 45.075 94.875 50.585 95.685 ;
        RECT 50.595 94.875 53.345 95.685 ;
        RECT 53.855 95.005 61.165 95.685 ;
        RECT 53.855 94.775 55.205 95.005 ;
        RECT 56.740 94.785 57.650 95.005 ;
        RECT 61.175 94.875 63.005 95.685 ;
        RECT 63.485 94.815 63.915 95.600 ;
        RECT 63.935 94.775 67.145 95.685 ;
        RECT 67.615 94.775 70.825 95.685 ;
        RECT 70.835 94.875 72.665 95.685 ;
        RECT 72.810 95.655 72.980 95.925 ;
        RECT 74.010 95.895 74.965 95.925 ;
        RECT 74.975 95.895 76.345 96.705 ;
        RECT 76.365 95.980 76.795 96.765 ;
        RECT 80.935 96.575 81.865 96.805 ;
        RECT 77.965 95.895 81.865 96.575 ;
        RECT 81.875 95.895 87.385 96.705 ;
        RECT 87.395 95.895 89.225 96.705 ;
        RECT 89.235 95.895 90.605 96.705 ;
        RECT 75.115 95.705 75.285 95.895 ;
        RECT 76.965 95.740 77.125 95.850 ;
        RECT 77.425 95.730 77.585 95.840 ;
        RECT 75.120 95.685 75.285 95.705 ;
        RECT 78.335 95.685 78.505 95.875 ;
        RECT 81.280 95.705 81.450 95.895 ;
        RECT 81.555 95.685 81.725 95.875 ;
        RECT 82.015 95.705 82.185 95.895 ;
        RECT 87.075 95.685 87.245 95.875 ;
        RECT 87.535 95.705 87.705 95.895 ;
        RECT 88.910 95.735 89.030 95.845 ;
        RECT 90.295 95.685 90.465 95.895 ;
        RECT 74.010 95.655 74.965 95.685 ;
        RECT 72.685 94.975 74.965 95.655 ;
        RECT 75.120 95.005 76.955 95.685 ;
        RECT 74.010 94.775 74.965 94.975 ;
        RECT 76.025 94.775 76.955 95.005 ;
        RECT 78.195 94.775 81.405 95.685 ;
        RECT 81.415 94.875 86.925 95.685 ;
        RECT 86.935 94.875 88.765 95.685 ;
        RECT 89.235 94.875 90.605 95.685 ;
      LAYER nwell ;
        RECT 11.760 91.655 90.800 94.485 ;
        RECT 99.800 92.735 112.970 100.575 ;
      LAYER pwell ;
        RECT 134.270 96.400 158.480 102.920 ;
        RECT 11.955 90.455 13.325 91.265 ;
        RECT 16.850 91.135 17.760 91.355 ;
        RECT 19.295 91.135 21.065 91.365 ;
        RECT 23.445 91.135 24.365 91.365 ;
        RECT 13.335 90.455 21.065 91.135 ;
        RECT 22.075 90.455 24.365 91.135 ;
        RECT 24.845 90.540 25.275 91.325 ;
        RECT 25.755 91.135 26.685 91.365 ;
        RECT 25.755 90.455 29.655 91.135 ;
        RECT 29.895 90.455 35.405 91.265 ;
        RECT 35.415 90.455 39.085 91.265 ;
        RECT 41.750 91.135 42.670 91.365 ;
        RECT 39.205 90.455 42.670 91.135 ;
        RECT 42.775 90.455 44.605 91.265 ;
        RECT 47.795 91.165 48.745 91.365 ;
        RECT 45.075 90.485 48.745 91.165 ;
        RECT 12.095 90.245 12.265 90.455 ;
        RECT 13.475 90.245 13.645 90.455 ;
        RECT 15.310 90.295 15.430 90.405 ;
        RECT 11.955 89.435 13.325 90.245 ;
        RECT 13.335 89.435 15.165 90.245 ;
        RECT 15.635 90.215 16.590 90.245 ;
        RECT 17.620 90.215 17.790 90.435 ;
        RECT 18.075 90.245 18.245 90.435 ;
        RECT 21.305 90.300 21.465 90.410 ;
        RECT 22.215 90.265 22.385 90.455 ;
        RECT 25.435 90.405 25.605 90.435 ;
        RECT 24.510 90.295 24.630 90.405 ;
        RECT 25.430 90.295 25.605 90.405 ;
        RECT 25.435 90.245 25.605 90.295 ;
        RECT 26.170 90.265 26.340 90.455 ;
        RECT 27.735 90.245 27.905 90.435 ;
        RECT 30.035 90.265 30.205 90.455 ;
        RECT 30.495 90.245 30.665 90.435 ;
        RECT 35.555 90.265 35.725 90.455 ;
        RECT 38.590 90.245 38.760 90.435 ;
        RECT 39.235 90.265 39.405 90.455 ;
        RECT 42.455 90.245 42.625 90.435 ;
        RECT 42.915 90.265 43.085 90.455 ;
        RECT 44.300 90.245 44.470 90.435 ;
        RECT 44.750 90.295 44.870 90.405 ;
        RECT 45.220 90.265 45.390 90.485 ;
        RECT 47.795 90.455 48.745 90.485 ;
        RECT 48.755 90.455 50.585 91.265 ;
        RECT 50.605 90.540 51.035 91.325 ;
        RECT 51.055 90.455 56.565 91.265 ;
        RECT 56.575 90.455 62.085 91.265 ;
        RECT 62.095 90.455 65.765 91.265 ;
        RECT 65.875 90.455 68.065 91.365 ;
        RECT 68.075 90.455 69.905 91.265 ;
        RECT 71.285 91.135 72.205 91.365 ;
        RECT 69.915 90.455 72.205 91.135 ;
        RECT 72.215 90.455 75.885 91.265 ;
        RECT 76.365 90.540 76.795 91.325 ;
        RECT 76.815 90.455 79.025 91.365 ;
        RECT 79.125 90.455 80.475 91.365 ;
        RECT 80.495 90.455 84.165 91.265 ;
        RECT 84.175 90.455 85.545 91.265 ;
        RECT 85.650 91.135 86.570 91.365 ;
        RECT 85.650 90.455 89.115 91.135 ;
        RECT 89.235 90.455 90.605 91.265 ;
        RECT 48.895 90.265 49.065 90.455 ;
        RECT 15.635 89.535 17.915 90.215 ;
        RECT 17.935 89.565 25.245 90.245 ;
        RECT 25.295 89.565 27.585 90.245 ;
        RECT 15.635 89.335 16.590 89.535 ;
        RECT 21.450 89.345 22.360 89.565 ;
        RECT 23.895 89.335 25.245 89.565 ;
        RECT 26.665 89.335 27.585 89.565 ;
        RECT 27.595 89.435 30.345 90.245 ;
        RECT 30.355 89.565 37.665 90.245 ;
        RECT 33.870 89.345 34.780 89.565 ;
        RECT 36.315 89.335 37.665 89.565 ;
        RECT 37.725 89.375 38.155 90.160 ;
        RECT 38.175 89.565 42.075 90.245 ;
        RECT 38.175 89.335 39.105 89.565 ;
        RECT 42.315 89.435 44.145 90.245 ;
        RECT 44.155 89.335 47.630 90.245 ;
        RECT 47.835 90.215 48.770 90.245 ;
        RECT 50.730 90.215 50.900 90.435 ;
        RECT 51.195 90.265 51.365 90.455 ;
        RECT 53.495 90.245 53.665 90.435 ;
        RECT 53.955 90.245 54.125 90.435 ;
        RECT 55.795 90.245 55.965 90.435 ;
        RECT 56.715 90.265 56.885 90.455 ;
        RECT 62.235 90.265 62.405 90.455 ;
        RECT 63.150 90.295 63.270 90.405 ;
        RECT 64.080 90.245 64.250 90.435 ;
        RECT 67.750 90.400 67.920 90.455 ;
        RECT 67.750 90.290 67.925 90.400 ;
        RECT 67.750 90.265 67.920 90.290 ;
        RECT 68.215 90.265 68.385 90.455 ;
        RECT 68.675 90.245 68.845 90.435 ;
        RECT 70.055 90.265 70.225 90.455 ;
        RECT 71.440 90.245 71.610 90.435 ;
        RECT 72.355 90.265 72.525 90.455 ;
        RECT 73.275 90.245 73.445 90.435 ;
        RECT 76.030 90.295 76.150 90.405 ;
        RECT 76.495 90.245 76.665 90.435 ;
        RECT 76.960 90.265 77.130 90.455 ;
        RECT 79.710 90.295 79.830 90.405 ;
        RECT 80.175 90.245 80.345 90.455 ;
        RECT 80.635 90.265 80.805 90.455 ;
        RECT 84.315 90.265 84.485 90.455 ;
        RECT 87.535 90.245 87.705 90.435 ;
        RECT 88.915 90.265 89.085 90.455 ;
        RECT 90.295 90.245 90.465 90.455 ;
        RECT 47.835 90.015 50.900 90.215 ;
        RECT 47.835 89.535 51.045 90.015 ;
        RECT 47.835 89.335 48.785 89.535 ;
        RECT 50.115 89.335 51.045 89.535 ;
        RECT 51.055 89.565 53.805 90.245 ;
        RECT 51.055 89.335 51.985 89.565 ;
        RECT 53.815 89.435 55.645 90.245 ;
        RECT 55.655 89.565 62.965 90.245 ;
        RECT 59.170 89.345 60.080 89.565 ;
        RECT 61.615 89.335 62.965 89.565 ;
        RECT 63.485 89.375 63.915 90.160 ;
        RECT 63.935 89.335 67.605 90.245 ;
        RECT 68.535 89.565 71.285 90.245 ;
        RECT 70.355 89.335 71.285 89.565 ;
        RECT 71.295 89.335 73.125 90.245 ;
        RECT 73.135 89.435 75.885 90.245 ;
        RECT 76.355 89.335 79.565 90.245 ;
        RECT 80.035 89.565 87.345 90.245 ;
        RECT 87.395 89.565 89.225 90.245 ;
        RECT 83.550 89.345 84.460 89.565 ;
        RECT 85.995 89.335 87.345 89.565 ;
        RECT 87.880 89.335 89.225 89.565 ;
        RECT 89.235 89.435 90.605 90.245 ;
      LAYER nwell ;
        RECT 11.760 86.215 90.800 89.045 ;
      LAYER pwell ;
        RECT 99.810 88.235 112.980 92.025 ;
        RECT 11.955 85.015 13.325 85.825 ;
        RECT 13.335 85.015 17.005 85.825 ;
        RECT 17.015 85.015 18.385 85.825 ;
        RECT 19.445 85.695 20.375 85.925 ;
        RECT 18.540 85.015 20.375 85.695 ;
        RECT 20.895 85.835 21.845 85.925 ;
        RECT 20.895 85.015 22.825 85.835 ;
        RECT 23.465 85.015 24.815 85.925 ;
        RECT 24.845 85.100 25.275 85.885 ;
        RECT 29.730 85.695 30.640 85.915 ;
        RECT 32.175 85.695 33.945 85.925 ;
        RECT 26.215 85.015 33.945 85.695 ;
        RECT 34.035 85.015 37.705 85.825 ;
        RECT 38.730 85.695 39.650 85.925 ;
        RECT 42.315 85.725 43.245 85.925 ;
        RECT 44.575 85.725 45.525 85.925 ;
        RECT 38.730 85.015 42.195 85.695 ;
        RECT 42.315 85.245 45.525 85.725 ;
        RECT 42.460 85.045 45.525 85.245 ;
        RECT 12.095 84.805 12.265 85.015 ;
        RECT 13.475 84.805 13.645 85.015 ;
        RECT 17.155 84.825 17.325 85.015 ;
        RECT 18.540 84.995 18.705 85.015 ;
        RECT 22.675 84.995 22.825 85.015 ;
        RECT 18.535 84.825 18.705 84.995 ;
        RECT 18.995 84.805 19.165 84.995 ;
        RECT 22.675 84.825 22.845 84.995 ;
        RECT 23.130 84.855 23.250 84.965 ;
        RECT 23.595 84.825 23.765 85.015 ;
        RECT 24.515 84.805 24.685 84.995 ;
        RECT 25.445 84.860 25.605 84.970 ;
        RECT 26.355 84.965 26.525 85.015 ;
        RECT 26.350 84.855 26.525 84.965 ;
        RECT 26.355 84.825 26.525 84.855 ;
        RECT 27.090 84.805 27.260 84.995 ;
        RECT 30.955 84.805 31.125 84.995 ;
        RECT 34.175 84.825 34.345 85.015 ;
        RECT 36.475 84.805 36.645 84.995 ;
        RECT 37.865 84.860 38.025 84.970 ;
        RECT 38.315 84.805 38.485 84.995 ;
        RECT 41.995 84.825 42.165 85.015 ;
        RECT 42.460 84.825 42.630 85.045 ;
        RECT 44.590 85.015 45.525 85.045 ;
        RECT 46.455 85.695 47.385 85.925 ;
        RECT 46.455 85.015 49.205 85.695 ;
        RECT 49.215 85.015 50.585 85.825 ;
        RECT 50.605 85.100 51.035 85.885 ;
        RECT 51.055 85.695 51.985 85.925 ;
        RECT 59.170 85.695 60.080 85.915 ;
        RECT 61.615 85.695 62.965 85.925 ;
        RECT 51.055 85.015 54.955 85.695 ;
        RECT 55.655 85.015 62.965 85.695 ;
        RECT 63.015 85.015 66.225 85.925 ;
        RECT 66.545 85.695 67.475 85.925 ;
        RECT 66.545 85.015 68.380 85.695 ;
        RECT 68.535 85.015 69.885 85.925 ;
        RECT 69.915 85.015 71.285 85.825 ;
        RECT 71.295 85.015 73.125 85.925 ;
        RECT 75.105 85.695 76.035 85.925 ;
        RECT 74.200 85.015 76.035 85.695 ;
        RECT 76.365 85.100 76.795 85.885 ;
        RECT 76.965 85.015 80.620 85.925 ;
        RECT 81.875 85.695 82.805 85.925 ;
        RECT 81.875 85.015 85.775 85.695 ;
        RECT 86.015 85.015 87.385 85.795 ;
        RECT 87.395 85.015 89.225 85.825 ;
        RECT 89.235 85.015 90.605 85.825 ;
        RECT 45.685 84.860 45.845 84.970 ;
        RECT 11.955 83.995 13.325 84.805 ;
        RECT 13.335 83.995 18.845 84.805 ;
        RECT 18.855 83.995 24.365 84.805 ;
        RECT 24.375 83.995 26.205 84.805 ;
        RECT 26.675 84.125 30.575 84.805 ;
        RECT 26.675 83.895 27.605 84.125 ;
        RECT 30.815 83.995 36.325 84.805 ;
        RECT 36.335 83.995 37.705 84.805 ;
        RECT 37.725 83.935 38.155 84.720 ;
        RECT 38.175 84.125 45.485 84.805 ;
        RECT 41.690 83.905 42.600 84.125 ;
        RECT 44.135 83.895 45.485 84.125 ;
        RECT 45.535 84.775 46.480 84.805 ;
        RECT 47.970 84.775 48.140 84.995 ;
        RECT 48.430 84.855 48.550 84.965 ;
        RECT 48.895 84.805 49.065 85.015 ;
        RECT 49.355 84.825 49.525 85.015 ;
        RECT 51.470 84.825 51.640 85.015 ;
        RECT 55.330 84.855 55.450 84.965 ;
        RECT 55.795 84.825 55.965 85.015 ;
        RECT 59.475 84.805 59.645 84.995 ;
        RECT 59.935 84.805 60.105 84.995 ;
        RECT 63.145 84.825 63.315 85.015 ;
        RECT 68.215 84.995 68.380 85.015 ;
        RECT 64.085 84.850 64.245 84.960 ;
        RECT 45.535 84.095 48.285 84.775 ;
        RECT 48.755 84.125 56.065 84.805 ;
        RECT 45.535 83.895 46.480 84.095 ;
        RECT 52.270 83.905 53.180 84.125 ;
        RECT 54.715 83.895 56.065 84.125 ;
        RECT 56.210 84.125 59.675 84.805 ;
        RECT 56.210 83.895 57.130 84.125 ;
        RECT 59.795 83.995 63.465 84.805 ;
        RECT 65.000 84.775 65.170 84.995 ;
        RECT 68.215 84.825 68.385 84.995 ;
        RECT 69.600 84.825 69.770 85.015 ;
        RECT 70.055 84.825 70.225 85.015 ;
        RECT 70.515 84.805 70.685 84.995 ;
        RECT 70.975 84.805 71.145 84.995 ;
        RECT 71.440 84.825 71.610 85.015 ;
        RECT 74.200 84.995 74.365 85.015 ;
        RECT 76.965 84.995 77.125 85.015 ;
        RECT 73.285 84.860 73.445 84.970 ;
        RECT 74.195 84.825 74.365 84.995 ;
        RECT 75.575 84.805 75.745 84.995 ;
        RECT 76.035 84.805 76.205 84.995 ;
        RECT 76.955 84.825 77.125 84.995 ;
        RECT 81.105 84.860 81.265 84.970 ;
        RECT 81.555 84.805 81.725 84.995 ;
        RECT 82.290 84.825 82.460 85.015 ;
        RECT 84.315 84.805 84.485 84.995 ;
        RECT 86.155 84.825 86.325 85.015 ;
        RECT 87.535 84.825 87.705 85.015 ;
        RECT 88.915 84.805 89.085 84.995 ;
        RECT 90.295 84.805 90.465 85.015 ;
        RECT 67.130 84.775 68.065 84.805 ;
        RECT 63.485 83.935 63.915 84.720 ;
        RECT 65.000 84.575 68.065 84.775 ;
        RECT 64.855 84.095 68.065 84.575 ;
        RECT 64.855 83.895 65.785 84.095 ;
        RECT 67.115 83.895 68.065 84.095 ;
        RECT 68.075 84.125 70.825 84.805 ;
        RECT 68.075 83.895 69.005 84.125 ;
        RECT 70.835 83.995 73.585 84.805 ;
        RECT 73.595 84.125 75.885 84.805 ;
        RECT 73.595 83.895 74.515 84.125 ;
        RECT 75.895 83.995 81.405 84.805 ;
        RECT 81.415 83.995 84.165 84.805 ;
        RECT 84.175 84.025 85.545 84.805 ;
        RECT 85.650 84.125 89.115 84.805 ;
        RECT 85.650 83.895 86.570 84.125 ;
        RECT 89.235 83.995 90.605 84.805 ;
      LAYER nwell ;
        RECT 11.760 80.775 90.800 83.605 ;
      LAYER pwell ;
        RECT 99.810 80.745 113.660 87.965 ;
      LAYER nwell ;
        RECT 117.410 82.420 129.660 92.610 ;
      LAYER pwell ;
        RECT 127.210 81.190 129.320 81.200 ;
        RECT 15.835 80.395 16.785 80.485 ;
        RECT 11.955 79.575 13.325 80.385 ;
        RECT 13.335 79.575 15.165 80.385 ;
        RECT 15.835 79.575 17.765 80.395 ;
        RECT 17.935 79.575 19.285 80.485 ;
        RECT 19.315 79.575 20.665 80.485 ;
        RECT 21.615 80.285 22.545 80.485 ;
        RECT 23.880 80.285 24.825 80.485 ;
        RECT 21.615 79.805 24.825 80.285 ;
        RECT 21.755 79.605 24.825 79.805 ;
        RECT 24.845 79.660 25.275 80.445 ;
        RECT 12.095 79.365 12.265 79.575 ;
        RECT 13.475 79.385 13.645 79.575 ;
        RECT 17.615 79.555 17.765 79.575 ;
        RECT 14.395 79.365 14.565 79.555 ;
        RECT 15.310 79.415 15.430 79.525 ;
        RECT 17.615 79.385 17.785 79.555 ;
        RECT 19.000 79.385 19.170 79.575 ;
        RECT 19.460 79.385 19.630 79.575 ;
        RECT 20.845 79.420 21.005 79.530 ;
        RECT 21.755 79.365 21.925 79.605 ;
        RECT 23.880 79.575 24.825 79.605 ;
        RECT 25.295 79.575 26.665 80.385 ;
        RECT 26.675 80.255 27.605 80.485 ;
        RECT 26.675 79.575 30.575 80.255 ;
        RECT 30.815 79.575 36.325 80.385 ;
        RECT 40.455 80.255 41.385 80.485 ;
        RECT 37.485 79.575 41.385 80.255 ;
        RECT 41.395 79.575 43.225 80.385 ;
        RECT 43.330 80.255 44.250 80.485 ;
        RECT 49.570 80.255 50.490 80.485 ;
        RECT 43.330 79.575 46.795 80.255 ;
        RECT 47.025 79.575 50.490 80.255 ;
        RECT 50.605 79.660 51.035 80.445 ;
        RECT 51.055 80.255 51.975 80.485 ;
        RECT 53.355 80.255 54.285 80.485 ;
        RECT 51.055 79.575 53.345 80.255 ;
        RECT 53.355 79.575 57.255 80.255 ;
        RECT 57.495 79.575 63.005 80.385 ;
        RECT 65.670 80.255 66.590 80.485 ;
        RECT 68.065 80.255 68.985 80.485 ;
        RECT 63.125 79.575 66.590 80.255 ;
        RECT 66.695 79.575 68.985 80.255 ;
        RECT 68.995 79.575 71.745 80.385 ;
        RECT 72.365 79.575 76.020 80.485 ;
        RECT 76.365 79.660 76.795 80.445 ;
        RECT 76.815 79.575 80.025 80.485 ;
        RECT 83.550 80.255 84.460 80.475 ;
        RECT 85.995 80.255 87.345 80.485 ;
        RECT 87.880 80.255 89.225 80.485 ;
        RECT 80.035 79.575 87.345 80.255 ;
        RECT 87.395 79.575 89.225 80.255 ;
        RECT 89.235 79.575 90.605 80.385 ;
        RECT 11.955 78.555 13.325 79.365 ;
        RECT 14.255 78.685 21.565 79.365 ;
        RECT 17.770 78.465 18.680 78.685 ;
        RECT 20.215 78.455 21.565 78.685 ;
        RECT 21.615 78.555 23.445 79.365 ;
        RECT 23.595 79.335 23.765 79.555 ;
        RECT 25.435 79.385 25.605 79.575 ;
        RECT 26.810 79.415 26.930 79.525 ;
        RECT 27.090 79.385 27.260 79.575 ;
        RECT 27.275 79.365 27.445 79.555 ;
        RECT 30.955 79.385 31.125 79.575 ;
        RECT 35.095 79.365 35.265 79.555 ;
        RECT 36.485 79.420 36.645 79.530 ;
        RECT 38.315 79.365 38.485 79.555 ;
        RECT 40.800 79.385 40.970 79.575 ;
        RECT 41.535 79.385 41.705 79.575 ;
        RECT 45.670 79.415 45.790 79.525 ;
        RECT 46.595 79.385 46.765 79.575 ;
        RECT 47.055 79.385 47.225 79.575 ;
        RECT 53.035 79.365 53.205 79.575 ;
        RECT 53.495 79.365 53.665 79.555 ;
        RECT 53.770 79.385 53.940 79.575 ;
        RECT 57.635 79.385 57.805 79.575 ;
        RECT 63.155 79.365 63.325 79.575 ;
        RECT 64.075 79.365 64.245 79.555 ;
        RECT 66.835 79.385 67.005 79.575 ;
        RECT 67.300 79.365 67.470 79.555 ;
        RECT 69.135 79.385 69.305 79.575 ;
        RECT 72.365 79.555 72.525 79.575 ;
        RECT 70.525 79.410 70.685 79.520 ;
        RECT 71.890 79.415 72.010 79.525 ;
        RECT 72.355 79.385 72.525 79.555 ;
        RECT 73.735 79.365 73.905 79.555 ;
        RECT 76.495 79.365 76.665 79.555 ;
        RECT 76.955 79.365 77.125 79.575 ;
        RECT 80.175 79.385 80.345 79.575 ;
        RECT 80.635 79.365 80.805 79.555 ;
        RECT 82.290 79.365 82.460 79.555 ;
        RECT 86.155 79.365 86.325 79.555 ;
        RECT 87.535 79.365 87.705 79.575 ;
        RECT 90.295 79.365 90.465 79.575 ;
        RECT 25.720 79.335 26.665 79.365 ;
        RECT 23.595 79.135 26.665 79.335 ;
        RECT 23.455 78.655 26.665 79.135 ;
        RECT 27.135 78.685 34.865 79.365 ;
        RECT 23.455 78.455 24.385 78.655 ;
        RECT 25.720 78.455 26.665 78.655 ;
        RECT 30.650 78.465 31.560 78.685 ;
        RECT 33.095 78.455 34.865 78.685 ;
        RECT 34.955 78.555 37.705 79.365 ;
        RECT 37.725 78.495 38.155 79.280 ;
        RECT 38.175 78.685 45.485 79.365 ;
        RECT 41.690 78.465 42.600 78.685 ;
        RECT 44.135 78.455 45.485 78.685 ;
        RECT 46.035 78.685 53.345 79.365 ;
        RECT 46.035 78.455 47.385 78.685 ;
        RECT 48.920 78.465 49.830 78.685 ;
        RECT 53.355 78.555 56.105 79.365 ;
        RECT 56.155 78.685 63.465 79.365 ;
        RECT 56.155 78.455 57.505 78.685 ;
        RECT 59.040 78.465 59.950 78.685 ;
        RECT 63.485 78.495 63.915 79.280 ;
        RECT 64.015 78.455 67.015 79.365 ;
        RECT 67.155 78.455 70.075 79.365 ;
        RECT 71.305 78.455 74.035 79.365 ;
        RECT 74.065 78.455 76.795 79.365 ;
        RECT 76.815 78.555 80.485 79.365 ;
        RECT 80.495 78.555 81.865 79.365 ;
        RECT 81.875 78.685 85.775 79.365 ;
        RECT 81.875 78.455 82.805 78.685 ;
        RECT 86.015 78.585 87.385 79.365 ;
        RECT 87.395 78.555 89.225 79.365 ;
        RECT 89.235 78.555 90.605 79.365 ;
      LAYER nwell ;
        RECT 11.760 75.335 90.800 78.165 ;
      LAYER pwell ;
        RECT 11.955 74.135 13.325 74.945 ;
        RECT 13.335 74.135 15.165 74.945 ;
        RECT 15.485 74.815 16.415 75.045 ;
        RECT 17.935 74.845 18.865 75.045 ;
        RECT 20.195 74.845 21.145 75.045 ;
        RECT 15.485 74.135 17.320 74.815 ;
        RECT 17.935 74.365 21.145 74.845 ;
        RECT 21.615 74.845 22.545 75.045 ;
        RECT 23.880 74.845 24.825 75.045 ;
        RECT 21.615 74.365 24.825 74.845 ;
        RECT 12.095 73.925 12.265 74.135 ;
        RECT 13.475 74.085 13.645 74.135 ;
        RECT 17.155 74.115 17.320 74.135 ;
        RECT 18.080 74.165 21.145 74.365 ;
        RECT 13.470 73.975 13.645 74.085 ;
        RECT 13.475 73.945 13.645 73.975 ;
        RECT 14.210 73.925 14.380 74.115 ;
        RECT 17.155 73.945 17.325 74.115 ;
        RECT 17.610 73.975 17.730 74.085 ;
        RECT 18.080 73.945 18.250 74.165 ;
        RECT 20.210 74.135 21.145 74.165 ;
        RECT 21.755 74.165 24.825 74.365 ;
        RECT 24.845 74.220 25.275 75.005 ;
        RECT 18.350 73.925 18.520 74.115 ;
        RECT 21.290 73.975 21.410 74.085 ;
        RECT 21.755 73.945 21.925 74.165 ;
        RECT 23.880 74.135 24.825 74.165 ;
        RECT 25.295 74.135 27.125 74.945 ;
        RECT 31.110 74.815 32.020 75.035 ;
        RECT 33.555 74.815 35.325 75.045 ;
        RECT 27.595 74.135 35.325 74.815 ;
        RECT 35.415 74.135 39.085 74.945 ;
        RECT 40.935 74.815 41.865 75.045 ;
        RECT 45.075 74.815 46.005 75.045 ;
        RECT 39.560 74.135 40.925 74.815 ;
        RECT 40.935 74.135 44.835 74.815 ;
        RECT 45.075 74.135 48.975 74.815 ;
        RECT 49.215 74.135 50.585 74.945 ;
        RECT 50.605 74.220 51.035 75.005 ;
        RECT 51.055 74.815 51.985 75.045 ;
        RECT 55.695 74.815 57.045 75.045 ;
        RECT 58.580 74.815 59.490 75.035 ;
        RECT 65.670 74.815 66.590 75.045 ;
        RECT 51.055 74.135 54.955 74.815 ;
        RECT 55.695 74.135 63.005 74.815 ;
        RECT 63.125 74.135 66.590 74.815 ;
        RECT 66.695 74.135 69.905 75.045 ;
        RECT 71.055 74.955 72.005 75.045 ;
        RECT 70.075 74.135 72.005 74.955 ;
        RECT 72.215 74.135 73.565 75.045 ;
        RECT 74.540 74.815 75.885 75.045 ;
        RECT 74.055 74.135 75.885 74.815 ;
        RECT 76.365 74.220 76.795 75.005 ;
        RECT 76.815 74.135 79.565 74.945 ;
        RECT 83.550 74.815 84.460 75.035 ;
        RECT 85.995 74.815 87.345 75.045 ;
        RECT 87.880 74.815 89.225 75.045 ;
        RECT 80.035 74.135 87.345 74.815 ;
        RECT 87.395 74.135 89.225 74.815 ;
        RECT 89.235 74.135 90.605 74.945 ;
        RECT 99.810 74.755 110.700 80.745 ;
        RECT 117.420 78.410 129.320 81.190 ;
        RECT 117.420 76.450 127.240 78.410 ;
        RECT 117.420 75.290 127.640 76.450 ;
      LAYER nwell ;
        RECT 129.320 76.300 131.430 81.140 ;
        RECT 134.240 78.800 139.890 84.990 ;
      LAYER pwell ;
        RECT 134.230 75.340 139.880 78.440 ;
        RECT 117.420 75.090 127.240 75.290 ;
        RECT 22.225 73.970 22.385 74.080 ;
        RECT 25.435 73.945 25.605 74.135 ;
        RECT 26.540 73.925 26.710 74.115 ;
        RECT 27.275 74.085 27.445 74.115 ;
        RECT 27.270 73.975 27.445 74.085 ;
        RECT 27.275 73.925 27.445 73.975 ;
        RECT 27.735 73.945 27.905 74.135 ;
        RECT 32.335 73.925 32.505 74.115 ;
        RECT 35.555 73.945 35.725 74.135 ;
        RECT 38.325 73.970 38.485 74.080 ;
        RECT 39.235 73.925 39.405 74.115 ;
        RECT 41.350 73.945 41.520 74.135 ;
        RECT 44.295 73.925 44.465 74.115 ;
        RECT 45.490 73.945 45.660 74.135 ;
        RECT 47.055 73.925 47.225 74.115 ;
        RECT 49.355 73.945 49.525 74.135 ;
        RECT 51.470 73.945 51.640 74.135 ;
        RECT 54.690 73.925 54.860 74.115 ;
        RECT 55.330 73.975 55.450 74.085 ;
        RECT 61.775 73.925 61.945 74.115 ;
        RECT 62.235 73.925 62.405 74.115 ;
        RECT 62.695 73.945 62.865 74.135 ;
        RECT 63.155 73.945 63.325 74.135 ;
        RECT 64.075 73.945 64.245 74.115 ;
        RECT 66.835 73.945 67.005 74.135 ;
        RECT 70.075 74.115 70.225 74.135 ;
        RECT 68.220 73.925 68.390 74.115 ;
        RECT 69.600 73.925 69.770 74.115 ;
        RECT 70.055 73.945 70.225 74.115 ;
        RECT 70.970 73.925 71.140 74.115 ;
        RECT 71.445 73.970 71.605 74.080 ;
        RECT 72.355 73.925 72.525 74.115 ;
        RECT 73.280 73.945 73.450 74.135 ;
        RECT 73.730 73.975 73.850 74.085 ;
        RECT 74.195 73.945 74.365 74.135 ;
        RECT 76.030 73.975 76.150 74.085 ;
        RECT 76.955 73.945 77.125 74.135 ;
        RECT 78.790 73.925 78.960 74.115 ;
        RECT 79.255 73.925 79.425 74.115 ;
        RECT 79.710 73.975 79.830 74.085 ;
        RECT 80.175 73.945 80.345 74.135 ;
        RECT 81.090 73.975 81.210 74.085 ;
        RECT 81.830 73.925 82.000 74.115 ;
        RECT 87.535 73.945 87.705 74.135 ;
        RECT 88.915 73.925 89.085 74.115 ;
        RECT 90.295 73.925 90.465 74.135 ;
        RECT 11.955 73.115 13.325 73.925 ;
        RECT 13.795 73.245 17.695 73.925 ;
        RECT 17.935 73.245 21.835 73.925 ;
        RECT 23.225 73.245 27.125 73.925 ;
        RECT 27.135 73.245 31.950 73.925 ;
        RECT 13.795 73.015 14.725 73.245 ;
        RECT 17.935 73.015 18.865 73.245 ;
        RECT 26.195 73.015 27.125 73.245 ;
        RECT 32.195 73.115 37.705 73.925 ;
        RECT 37.725 73.055 38.155 73.840 ;
        RECT 39.095 73.245 43.910 73.925 ;
        RECT 44.155 73.115 46.905 73.925 ;
        RECT 46.915 73.245 54.225 73.925 ;
        RECT 50.430 73.025 51.340 73.245 ;
        RECT 52.875 73.015 54.225 73.245 ;
        RECT 54.275 73.245 58.175 73.925 ;
        RECT 58.510 73.245 61.975 73.925 ;
        RECT 54.275 73.015 55.205 73.245 ;
        RECT 58.510 73.015 59.430 73.245 ;
        RECT 62.095 73.115 63.465 73.925 ;
        RECT 63.485 73.055 63.915 73.840 ;
        RECT 64.340 73.245 66.765 73.925 ;
        RECT 67.155 73.015 68.505 73.925 ;
        RECT 68.535 73.015 69.885 73.925 ;
        RECT 69.935 73.015 71.285 73.925 ;
        RECT 72.215 73.015 75.425 73.925 ;
        RECT 75.630 73.015 79.105 73.925 ;
        RECT 79.115 73.115 80.945 73.925 ;
        RECT 81.415 73.245 85.315 73.925 ;
        RECT 85.650 73.245 89.115 73.925 ;
        RECT 81.415 73.015 82.345 73.245 ;
        RECT 85.650 73.015 86.570 73.245 ;
        RECT 89.235 73.115 90.605 73.925 ;
      LAYER nwell ;
        RECT 11.760 69.895 90.800 72.725 ;
      LAYER pwell ;
        RECT 11.955 68.695 13.325 69.505 ;
        RECT 16.850 69.375 17.760 69.595 ;
        RECT 19.295 69.375 21.065 69.605 ;
        RECT 13.335 68.695 21.065 69.375 ;
        RECT 21.155 68.695 24.825 69.505 ;
        RECT 24.845 68.780 25.275 69.565 ;
        RECT 28.810 69.375 29.720 69.595 ;
        RECT 31.255 69.375 33.025 69.605 ;
        RECT 25.295 68.695 33.025 69.375 ;
        RECT 33.115 68.695 34.945 69.505 ;
        RECT 34.955 69.375 35.885 69.605 ;
        RECT 42.610 69.375 43.520 69.595 ;
        RECT 45.055 69.375 46.405 69.605 ;
        RECT 34.955 68.695 38.855 69.375 ;
        RECT 39.095 68.695 46.405 69.375 ;
        RECT 46.455 69.375 47.385 69.605 ;
        RECT 46.455 68.695 50.355 69.375 ;
        RECT 50.605 68.780 51.035 69.565 ;
        RECT 51.150 69.375 52.070 69.605 ;
        RECT 51.150 68.695 54.615 69.375 ;
        RECT 54.735 68.695 58.405 69.505 ;
        RECT 67.050 69.375 67.970 69.605 ;
        RECT 59.335 68.695 64.150 69.375 ;
        RECT 64.505 68.695 67.970 69.375 ;
        RECT 68.275 69.515 69.225 69.605 ;
        RECT 68.275 68.695 70.205 69.515 ;
        RECT 70.385 68.695 71.735 69.605 ;
        RECT 71.775 68.695 73.125 69.605 ;
        RECT 74.470 69.405 75.425 69.605 ;
        RECT 73.145 68.725 75.425 69.405 ;
        RECT 76.365 68.780 76.795 69.565 ;
        RECT 12.095 68.485 12.265 68.695 ;
        RECT 13.475 68.505 13.645 68.695 ;
        RECT 14.855 68.485 15.025 68.675 ;
        RECT 15.325 68.530 15.485 68.640 ;
        RECT 16.235 68.485 16.405 68.675 ;
        RECT 21.295 68.505 21.465 68.695 ;
        RECT 25.435 68.505 25.605 68.695 ;
        RECT 27.460 68.485 27.630 68.675 ;
        RECT 28.195 68.485 28.365 68.675 ;
        RECT 33.255 68.505 33.425 68.695 ;
        RECT 33.715 68.485 33.885 68.675 ;
        RECT 35.370 68.505 35.540 68.695 ;
        RECT 37.390 68.535 37.510 68.645 ;
        RECT 38.310 68.535 38.430 68.645 ;
        RECT 39.235 68.505 39.405 68.695 ;
        RECT 41.995 68.485 42.165 68.675 ;
        RECT 45.225 68.485 45.395 68.675 ;
        RECT 45.675 68.485 45.845 68.675 ;
        RECT 46.870 68.505 47.040 68.695 ;
        RECT 50.275 68.485 50.445 68.675 ;
        RECT 50.745 68.530 50.905 68.640 ;
        RECT 51.930 68.485 52.100 68.675 ;
        RECT 54.415 68.505 54.585 68.695 ;
        RECT 54.875 68.505 55.045 68.695 ;
        RECT 58.565 68.540 58.725 68.650 ;
        RECT 59.475 68.505 59.645 68.695 ;
        RECT 62.695 68.485 62.865 68.675 ;
        RECT 63.150 68.535 63.270 68.645 ;
        RECT 64.350 68.485 64.520 68.675 ;
        RECT 64.535 68.505 64.705 68.695 ;
        RECT 70.055 68.675 70.205 68.695 ;
        RECT 71.435 68.675 71.605 68.695 ;
        RECT 68.215 68.485 68.385 68.675 ;
        RECT 70.055 68.505 70.225 68.675 ;
        RECT 70.970 68.535 71.090 68.645 ;
        RECT 71.430 68.505 71.605 68.675 ;
        RECT 71.890 68.505 72.060 68.695 ;
        RECT 73.270 68.505 73.440 68.725 ;
        RECT 74.470 68.695 75.425 68.725 ;
        RECT 77.735 68.695 80.945 69.605 ;
        RECT 80.955 68.695 83.705 69.505 ;
        RECT 83.715 69.375 85.060 69.605 ;
        RECT 85.650 69.375 86.570 69.605 ;
        RECT 83.715 68.695 85.545 69.375 ;
        RECT 85.650 68.695 89.115 69.375 ;
        RECT 89.235 68.695 90.605 69.505 ;
        RECT 76.950 68.650 77.120 68.675 ;
        RECT 75.585 68.540 75.745 68.650 ;
        RECT 76.950 68.540 77.125 68.650 ;
        RECT 11.955 67.675 13.325 68.485 ;
        RECT 13.335 67.805 15.165 68.485 ;
        RECT 16.095 67.805 23.825 68.485 ;
        RECT 24.145 67.805 28.045 68.485 ;
        RECT 13.335 67.575 14.680 67.805 ;
        RECT 19.610 67.585 20.520 67.805 ;
        RECT 22.055 67.575 23.825 67.805 ;
        RECT 27.115 67.575 28.045 67.805 ;
        RECT 28.055 67.675 33.565 68.485 ;
        RECT 33.575 67.675 37.245 68.485 ;
        RECT 37.725 67.615 38.155 68.400 ;
        RECT 38.730 67.805 42.195 68.485 ;
        RECT 38.730 67.575 39.650 67.805 ;
        RECT 42.315 67.575 45.525 68.485 ;
        RECT 45.535 67.675 46.905 68.485 ;
        RECT 47.010 67.805 50.475 68.485 ;
        RECT 51.515 67.805 55.415 68.485 ;
        RECT 55.695 67.805 63.005 68.485 ;
        RECT 47.010 67.575 47.930 67.805 ;
        RECT 51.515 67.575 52.445 67.805 ;
        RECT 55.695 67.575 57.045 67.805 ;
        RECT 58.580 67.585 59.490 67.805 ;
        RECT 63.485 67.615 63.915 68.400 ;
        RECT 63.935 67.805 67.835 68.485 ;
        RECT 63.935 67.575 64.865 67.805 ;
        RECT 68.075 67.675 70.825 68.485 ;
        RECT 71.430 68.455 71.600 68.505 ;
        RECT 76.950 68.485 77.120 68.540 ;
        RECT 77.415 68.485 77.585 68.675 ;
        RECT 77.875 68.505 78.045 68.695 ;
        RECT 80.635 68.485 80.805 68.675 ;
        RECT 81.095 68.505 81.265 68.695 ;
        RECT 85.235 68.505 85.405 68.695 ;
        RECT 88.915 68.485 89.085 68.695 ;
        RECT 90.295 68.485 90.465 68.695 ;
        RECT 72.630 68.455 73.585 68.485 ;
        RECT 71.305 67.775 73.585 68.455 ;
        RECT 72.630 67.575 73.585 67.775 ;
        RECT 73.790 67.575 77.265 68.485 ;
        RECT 77.275 67.575 80.485 68.485 ;
        RECT 80.495 67.805 87.805 68.485 ;
        RECT 84.010 67.585 84.920 67.805 ;
        RECT 86.455 67.575 87.805 67.805 ;
        RECT 87.855 67.705 89.225 68.485 ;
        RECT 89.235 67.675 90.605 68.485 ;
      LAYER nwell ;
        RECT 11.760 64.455 90.800 67.285 ;
      LAYER pwell ;
        RECT 11.955 63.255 13.325 64.065 ;
        RECT 13.335 63.935 14.680 64.165 ;
        RECT 15.175 63.935 16.520 64.165 ;
        RECT 13.335 63.255 15.165 63.935 ;
        RECT 15.175 63.255 17.005 63.935 ;
        RECT 17.015 63.255 18.385 64.065 ;
        RECT 18.395 63.935 19.740 64.165 ;
        RECT 18.395 63.255 20.225 63.935 ;
        RECT 20.235 63.255 23.905 64.065 ;
        RECT 24.845 63.340 25.275 64.125 ;
        RECT 25.295 63.255 28.770 64.165 ;
        RECT 30.025 63.935 30.955 64.165 ;
        RECT 29.120 63.255 30.955 63.935 ;
        RECT 31.275 63.255 33.105 64.065 ;
        RECT 36.630 63.935 37.540 64.155 ;
        RECT 39.075 63.935 40.425 64.165 ;
        RECT 33.115 63.255 40.425 63.935 ;
        RECT 40.475 63.255 43.225 64.065 ;
        RECT 43.235 63.935 44.165 64.165 ;
        RECT 43.235 63.255 47.135 63.935 ;
        RECT 47.845 63.255 50.585 63.935 ;
        RECT 50.605 63.340 51.035 64.125 ;
        RECT 54.570 63.935 55.480 64.155 ;
        RECT 57.015 63.935 58.365 64.165 ;
        RECT 51.055 63.255 58.365 63.935 ;
        RECT 58.510 63.935 59.430 64.165 ;
        RECT 64.750 63.935 65.670 64.165 ;
        RECT 58.510 63.255 61.975 63.935 ;
        RECT 62.205 63.255 65.670 63.935 ;
        RECT 65.775 63.255 67.605 64.165 ;
        RECT 75.105 63.935 76.035 64.165 ;
        RECT 68.535 63.255 73.350 63.935 ;
        RECT 74.200 63.255 76.035 63.935 ;
        RECT 76.365 63.340 76.795 64.125 ;
        RECT 76.815 63.255 78.645 64.065 ;
        RECT 81.310 63.935 82.230 64.165 ;
        RECT 78.765 63.255 82.230 63.935 ;
        RECT 82.335 63.935 83.265 64.165 ;
        RECT 87.880 63.935 89.225 64.165 ;
        RECT 82.335 63.255 86.235 63.935 ;
        RECT 87.395 63.255 89.225 63.935 ;
        RECT 89.235 63.255 90.605 64.065 ;
        RECT 12.095 63.045 12.265 63.255 ;
        RECT 13.475 63.045 13.645 63.235 ;
        RECT 14.855 63.065 15.025 63.255 ;
        RECT 16.695 63.065 16.865 63.255 ;
        RECT 14.860 63.045 15.025 63.065 ;
        RECT 17.155 63.045 17.325 63.255 ;
        RECT 19.915 63.065 20.085 63.255 ;
        RECT 20.375 63.065 20.545 63.255 ;
        RECT 22.700 63.065 22.870 63.235 ;
        RECT 22.700 63.045 22.810 63.065 ;
        RECT 23.135 63.045 23.305 63.235 ;
        RECT 24.065 63.100 24.225 63.210 ;
        RECT 25.440 63.065 25.610 63.255 ;
        RECT 29.120 63.235 29.285 63.255 ;
        RECT 29.115 63.065 29.285 63.235 ;
        RECT 30.495 63.045 30.665 63.235 ;
        RECT 31.415 63.065 31.585 63.255 ;
        RECT 33.255 63.065 33.425 63.255 ;
        RECT 38.315 63.045 38.485 63.235 ;
        RECT 40.615 63.065 40.785 63.255 ;
        RECT 41.075 63.045 41.245 63.235 ;
        RECT 43.650 63.065 43.820 63.255 ;
        RECT 47.510 63.095 47.630 63.205 ;
        RECT 48.435 63.045 48.605 63.235 ;
        RECT 50.275 63.065 50.445 63.255 ;
        RECT 51.195 63.065 51.365 63.255 ;
        RECT 53.680 63.045 53.850 63.235 ;
        RECT 54.415 63.045 54.585 63.235 ;
        RECT 61.775 63.065 61.945 63.255 ;
        RECT 62.235 63.065 62.405 63.255 ;
        RECT 63.155 63.045 63.325 63.235 ;
        RECT 66.835 63.045 67.005 63.235 ;
        RECT 67.290 63.065 67.460 63.255 ;
        RECT 68.675 63.235 68.845 63.255 ;
        RECT 74.200 63.235 74.365 63.255 ;
        RECT 67.765 63.100 67.925 63.210 ;
        RECT 68.220 63.045 68.390 63.235 ;
        RECT 68.675 63.065 68.850 63.235 ;
        RECT 73.730 63.095 73.850 63.205 ;
        RECT 74.195 63.065 74.365 63.235 ;
        RECT 76.955 63.065 77.125 63.255 ;
        RECT 78.795 63.065 78.965 63.255 ;
        RECT 68.680 63.045 68.850 63.065 ;
        RECT 79.710 63.045 79.880 63.235 ;
        RECT 81.105 63.090 81.265 63.200 ;
        RECT 82.290 63.045 82.460 63.235 ;
        RECT 82.750 63.065 82.920 63.255 ;
        RECT 86.625 63.100 86.785 63.210 ;
        RECT 87.075 63.045 87.245 63.235 ;
        RECT 87.535 63.045 87.705 63.255 ;
        RECT 90.295 63.045 90.465 63.255 ;
        RECT 11.955 62.235 13.325 63.045 ;
        RECT 13.335 62.235 14.705 63.045 ;
        RECT 14.860 62.365 16.695 63.045 ;
        RECT 15.765 62.135 16.695 62.365 ;
        RECT 17.015 62.235 18.385 63.045 ;
        RECT 18.395 62.365 22.810 63.045 ;
        RECT 22.995 62.365 30.305 63.045 ;
        RECT 30.355 62.365 37.665 63.045 ;
        RECT 18.395 62.135 22.325 62.365 ;
        RECT 26.510 62.145 27.420 62.365 ;
        RECT 28.955 62.135 30.305 62.365 ;
        RECT 33.870 62.145 34.780 62.365 ;
        RECT 36.315 62.135 37.665 62.365 ;
        RECT 37.725 62.175 38.155 62.960 ;
        RECT 38.175 62.235 40.925 63.045 ;
        RECT 40.935 62.365 48.245 63.045 ;
        RECT 44.450 62.145 45.360 62.365 ;
        RECT 46.895 62.135 48.245 62.365 ;
        RECT 48.295 62.235 50.125 63.045 ;
        RECT 50.365 62.365 54.265 63.045 ;
        RECT 53.335 62.135 54.265 62.365 ;
        RECT 54.275 62.235 56.105 63.045 ;
        RECT 56.155 62.365 63.465 63.045 ;
        RECT 56.155 62.135 57.505 62.365 ;
        RECT 59.040 62.145 59.950 62.365 ;
        RECT 63.485 62.175 63.915 62.960 ;
        RECT 63.935 62.135 67.145 63.045 ;
        RECT 67.155 62.135 68.505 63.045 ;
        RECT 68.535 62.135 79.545 63.045 ;
        RECT 79.595 62.135 80.945 63.045 ;
        RECT 81.875 62.365 85.775 63.045 ;
        RECT 81.875 62.135 82.805 62.365 ;
        RECT 86.015 62.265 87.385 63.045 ;
        RECT 87.395 62.365 89.225 63.045 ;
        RECT 87.880 62.135 89.225 62.365 ;
        RECT 89.235 62.235 90.605 63.045 ;
      LAYER nwell ;
        RECT 11.760 59.015 90.800 61.845 ;
      LAYER pwell ;
        RECT 11.955 57.815 13.325 58.625 ;
        RECT 13.335 58.495 14.680 58.725 ;
        RECT 18.690 58.495 19.600 58.715 ;
        RECT 21.135 58.495 22.485 58.725 ;
        RECT 13.335 57.815 15.165 58.495 ;
        RECT 15.175 57.815 22.485 58.495 ;
        RECT 22.535 57.815 24.365 58.625 ;
        RECT 24.845 57.900 25.275 58.685 ;
        RECT 26.345 58.495 27.275 58.725 ;
        RECT 25.440 57.815 27.275 58.495 ;
        RECT 28.250 57.815 31.725 58.725 ;
        RECT 31.735 57.815 33.565 58.625 ;
        RECT 37.090 58.495 38.000 58.715 ;
        RECT 39.535 58.495 40.885 58.725 ;
        RECT 33.575 57.815 40.885 58.495 ;
        RECT 40.935 58.495 41.865 58.725 ;
        RECT 48.735 58.495 49.665 58.725 ;
        RECT 40.935 57.815 44.835 58.495 ;
        RECT 45.765 57.815 49.665 58.495 ;
        RECT 50.605 57.900 51.035 58.685 ;
        RECT 51.055 57.815 54.725 58.625 ;
        RECT 54.735 58.495 55.665 58.725 ;
        RECT 54.735 57.815 58.635 58.495 ;
        RECT 58.875 57.815 64.385 58.625 ;
        RECT 64.395 57.815 67.605 58.725 ;
        RECT 67.635 57.815 68.985 58.725 ;
        RECT 68.995 57.815 71.915 58.725 ;
        RECT 72.365 57.815 76.020 58.725 ;
        RECT 76.365 57.900 76.795 58.685 ;
        RECT 76.815 57.815 80.025 58.725 ;
        RECT 84.010 58.495 84.920 58.715 ;
        RECT 86.455 58.495 87.805 58.725 ;
        RECT 80.495 57.815 87.805 58.495 ;
        RECT 87.855 57.815 89.225 58.595 ;
        RECT 89.235 57.815 90.605 58.625 ;
        RECT 12.095 57.605 12.265 57.815 ;
        RECT 14.855 57.795 15.025 57.815 ;
        RECT 13.475 57.605 13.645 57.795 ;
        RECT 14.855 57.625 15.030 57.795 ;
        RECT 15.315 57.625 15.485 57.815 ;
        RECT 14.860 57.605 15.030 57.625 ;
        RECT 18.540 57.605 18.710 57.795 ;
        RECT 22.675 57.625 22.845 57.815 ;
        RECT 25.440 57.795 25.605 57.815 ;
        RECT 24.510 57.655 24.630 57.765 ;
        RECT 24.985 57.605 25.155 57.795 ;
        RECT 25.435 57.625 25.605 57.795 ;
        RECT 27.730 57.655 27.850 57.765 ;
        RECT 28.650 57.605 28.820 57.795 ;
        RECT 29.115 57.605 29.285 57.795 ;
        RECT 31.410 57.625 31.580 57.815 ;
        RECT 31.875 57.625 32.045 57.815 ;
        RECT 33.715 57.625 33.885 57.815 ;
        RECT 36.475 57.605 36.645 57.795 ;
        RECT 38.590 57.605 38.760 57.795 ;
        RECT 41.350 57.625 41.520 57.815 ;
        RECT 45.210 57.655 45.330 57.765 ;
        RECT 45.675 57.605 45.845 57.795 ;
        RECT 46.125 57.605 46.295 57.795 ;
        RECT 49.080 57.625 49.250 57.815 ;
        RECT 49.355 57.605 49.525 57.795 ;
        RECT 49.825 57.660 49.985 57.770 ;
        RECT 51.195 57.625 51.365 57.815 ;
        RECT 51.470 57.605 51.640 57.795 ;
        RECT 55.150 57.625 55.320 57.815 ;
        RECT 58.555 57.605 58.725 57.795 ;
        RECT 59.015 57.765 59.185 57.815 ;
        RECT 59.010 57.655 59.185 57.765 ;
        RECT 59.015 57.625 59.185 57.655 ;
        RECT 62.695 57.605 62.865 57.795 ;
        RECT 63.150 57.655 63.270 57.765 ;
        RECT 64.075 57.605 64.245 57.795 ;
        RECT 67.295 57.625 67.465 57.815 ;
        RECT 67.750 57.625 67.920 57.815 ;
        RECT 69.140 57.795 69.310 57.815 ;
        RECT 72.365 57.795 72.525 57.815 ;
        RECT 69.130 57.625 69.310 57.795 ;
        RECT 69.130 57.605 69.300 57.625 ;
        RECT 70.970 57.605 71.140 57.795 ;
        RECT 71.445 57.650 71.605 57.760 ;
        RECT 72.355 57.625 72.525 57.795 ;
        RECT 75.570 57.605 75.740 57.795 ;
        RECT 76.955 57.625 77.125 57.815 ;
        RECT 78.335 57.625 78.505 57.795 ;
        RECT 78.790 57.655 78.910 57.765 ;
        RECT 78.335 57.605 78.355 57.625 ;
        RECT 79.255 57.605 79.425 57.795 ;
        RECT 80.170 57.655 80.290 57.765 ;
        RECT 80.635 57.625 80.805 57.815 ;
        RECT 86.625 57.650 86.785 57.760 ;
        RECT 87.535 57.605 87.705 57.795 ;
        RECT 88.915 57.625 89.085 57.815 ;
        RECT 90.295 57.605 90.465 57.815 ;
        RECT 11.955 56.795 13.325 57.605 ;
        RECT 13.335 56.795 14.705 57.605 ;
        RECT 14.715 56.695 18.190 57.605 ;
        RECT 18.395 56.695 21.870 57.605 ;
        RECT 22.075 56.695 25.285 57.605 ;
        RECT 25.490 56.695 28.965 57.605 ;
        RECT 28.975 56.925 36.285 57.605 ;
        RECT 32.490 56.705 33.400 56.925 ;
        RECT 34.935 56.695 36.285 56.925 ;
        RECT 36.335 56.795 37.705 57.605 ;
        RECT 37.725 56.735 38.155 57.520 ;
        RECT 38.175 56.925 42.075 57.605 ;
        RECT 42.410 56.925 45.875 57.605 ;
        RECT 38.175 56.695 39.105 56.925 ;
        RECT 42.410 56.695 43.330 56.925 ;
        RECT 45.995 56.695 49.205 57.605 ;
        RECT 49.215 56.795 51.045 57.605 ;
        RECT 51.055 56.925 54.955 57.605 ;
        RECT 55.290 56.925 58.755 57.605 ;
        RECT 59.430 56.925 62.895 57.605 ;
        RECT 51.055 56.695 51.985 56.925 ;
        RECT 55.290 56.695 56.210 56.925 ;
        RECT 59.430 56.695 60.350 56.925 ;
        RECT 63.485 56.735 63.915 57.520 ;
        RECT 64.045 56.925 67.510 57.605 ;
        RECT 66.590 56.695 67.510 56.925 ;
        RECT 67.615 56.695 69.445 57.605 ;
        RECT 69.455 56.695 71.285 57.605 ;
        RECT 72.300 56.925 75.885 57.605 ;
        RECT 74.965 56.695 75.885 56.925 ;
        RECT 75.905 56.925 78.355 57.605 ;
        RECT 79.115 56.925 86.425 57.605 ;
        RECT 87.395 56.925 89.225 57.605 ;
        RECT 75.905 56.695 77.865 56.925 ;
        RECT 82.630 56.705 83.540 56.925 ;
        RECT 85.075 56.695 86.425 56.925 ;
        RECT 87.880 56.695 89.225 56.925 ;
        RECT 89.235 56.795 90.605 57.605 ;
      LAYER nwell ;
        RECT 11.760 53.575 90.800 56.405 ;
      LAYER pwell ;
        RECT 11.955 52.375 13.325 53.185 ;
        RECT 14.385 53.055 15.315 53.285 ;
        RECT 19.150 53.055 20.060 53.275 ;
        RECT 21.595 53.055 22.945 53.285 ;
        RECT 13.480 52.375 15.315 53.055 ;
        RECT 15.635 52.375 22.945 53.055 ;
        RECT 22.995 52.375 24.825 53.185 ;
        RECT 24.845 52.460 25.275 53.245 ;
        RECT 25.295 52.375 30.110 53.055 ;
        RECT 30.355 52.375 33.565 53.285 ;
        RECT 33.575 52.375 39.085 53.185 ;
        RECT 39.095 52.375 44.605 53.185 ;
        RECT 44.615 52.375 47.365 53.185 ;
        RECT 47.375 52.375 50.585 53.285 ;
        RECT 50.605 52.460 51.035 53.245 ;
        RECT 55.490 53.055 56.400 53.275 ;
        RECT 57.935 53.055 59.285 53.285 ;
        RECT 51.975 52.375 59.285 53.055 ;
        RECT 59.375 53.055 60.725 53.285 ;
        RECT 62.260 53.055 63.170 53.275 ;
        RECT 66.735 53.055 68.085 53.285 ;
        RECT 69.620 53.055 70.530 53.275 ;
        RECT 59.375 52.375 66.685 53.055 ;
        RECT 66.735 52.375 74.045 53.055 ;
        RECT 74.075 52.375 75.425 53.285 ;
        RECT 76.365 52.460 76.795 53.245 ;
        RECT 76.910 53.055 77.830 53.285 ;
        RECT 80.955 53.055 81.885 53.285 ;
        RECT 85.190 53.055 86.110 53.285 ;
        RECT 76.910 52.375 80.375 53.055 ;
        RECT 80.955 52.375 84.855 53.055 ;
        RECT 85.190 52.375 88.655 53.055 ;
        RECT 89.235 52.375 90.605 53.185 ;
        RECT 12.095 52.165 12.265 52.375 ;
        RECT 13.480 52.355 13.645 52.375 ;
        RECT 13.475 52.185 13.645 52.355 ;
        RECT 14.855 52.165 15.025 52.355 ;
        RECT 15.775 52.185 15.945 52.375 ;
        RECT 16.695 52.165 16.865 52.355 ;
        RECT 17.155 52.165 17.325 52.355 ;
        RECT 22.670 52.215 22.790 52.325 ;
        RECT 23.135 52.185 23.305 52.375 ;
        RECT 25.435 52.185 25.605 52.375 ;
        RECT 23.140 52.165 23.305 52.185 ;
        RECT 30.035 52.165 30.205 52.355 ;
        RECT 30.495 52.185 30.665 52.355 ;
        RECT 30.500 52.165 30.665 52.185 ;
        RECT 32.795 52.165 32.965 52.355 ;
        RECT 33.265 52.185 33.435 52.375 ;
        RECT 33.715 52.185 33.885 52.375 ;
        RECT 37.395 52.185 37.565 52.355 ;
        RECT 38.310 52.215 38.430 52.325 ;
        RECT 38.765 52.165 38.935 52.355 ;
        RECT 39.235 52.185 39.405 52.375 ;
        RECT 41.990 52.215 42.110 52.325 ;
        RECT 42.455 52.165 42.625 52.355 ;
        RECT 44.755 52.185 44.925 52.375 ;
        RECT 47.505 52.185 47.675 52.375 ;
        RECT 49.815 52.165 49.985 52.355 ;
        RECT 51.205 52.220 51.365 52.330 ;
        RECT 52.115 52.185 52.285 52.375 ;
        RECT 57.450 52.165 57.620 52.355 ;
        RECT 61.315 52.165 61.485 52.355 ;
        RECT 63.150 52.215 63.270 52.325 ;
        RECT 64.075 52.165 64.245 52.355 ;
        RECT 66.375 52.185 66.545 52.375 ;
        RECT 69.595 52.165 69.765 52.355 ;
        RECT 73.735 52.185 73.905 52.375 ;
        RECT 74.190 52.185 74.360 52.375 ;
        RECT 75.115 52.165 75.285 52.355 ;
        RECT 75.585 52.220 75.745 52.330 ;
        RECT 76.955 52.165 77.125 52.355 ;
        RECT 78.335 52.165 78.505 52.355 ;
        RECT 80.175 52.185 80.345 52.375 ;
        RECT 80.630 52.215 80.750 52.325 ;
        RECT 81.370 52.185 81.540 52.375 ;
        RECT 83.855 52.165 84.025 52.355 ;
        RECT 87.530 52.215 87.650 52.325 ;
        RECT 88.455 52.185 88.625 52.375 ;
        RECT 88.915 52.325 89.085 52.355 ;
        RECT 88.910 52.215 89.085 52.325 ;
        RECT 88.915 52.165 89.085 52.215 ;
        RECT 90.295 52.165 90.465 52.375 ;
        RECT 11.955 51.355 13.325 52.165 ;
        RECT 13.335 51.485 15.165 52.165 ;
        RECT 15.175 51.485 17.005 52.165 ;
        RECT 13.335 51.255 14.680 51.485 ;
        RECT 15.175 51.255 16.520 51.485 ;
        RECT 17.015 51.355 22.525 52.165 ;
        RECT 23.140 51.485 24.975 52.165 ;
        RECT 25.530 51.485 30.345 52.165 ;
        RECT 30.500 51.485 32.335 52.165 ;
        RECT 24.045 51.255 24.975 51.485 ;
        RECT 31.405 51.255 32.335 51.485 ;
        RECT 32.655 51.355 34.485 52.165 ;
        RECT 34.875 51.485 37.300 52.165 ;
        RECT 37.725 51.295 38.155 52.080 ;
        RECT 38.635 51.255 41.845 52.165 ;
        RECT 42.315 51.485 49.625 52.165 ;
        RECT 49.675 51.485 56.985 52.165 ;
        RECT 45.830 51.265 46.740 51.485 ;
        RECT 48.275 51.255 49.625 51.485 ;
        RECT 53.190 51.265 54.100 51.485 ;
        RECT 55.635 51.255 56.985 51.485 ;
        RECT 57.035 51.485 60.935 52.165 ;
        RECT 57.035 51.255 57.965 51.485 ;
        RECT 61.175 51.355 63.005 52.165 ;
        RECT 63.485 51.295 63.915 52.080 ;
        RECT 63.935 51.355 69.445 52.165 ;
        RECT 69.455 51.355 74.965 52.165 ;
        RECT 74.975 51.355 76.805 52.165 ;
        RECT 76.825 51.255 78.175 52.165 ;
        RECT 78.195 51.355 83.705 52.165 ;
        RECT 83.715 51.355 87.385 52.165 ;
        RECT 87.855 51.385 89.225 52.165 ;
        RECT 89.235 51.355 90.605 52.165 ;
      LAYER nwell ;
        RECT 11.760 48.135 90.800 50.965 ;
      LAYER pwell ;
        RECT 11.955 46.935 13.325 47.745 ;
        RECT 13.335 47.615 14.680 47.845 ;
        RECT 13.335 46.935 15.165 47.615 ;
        RECT 16.290 46.935 19.765 47.845 ;
        RECT 19.775 47.615 21.120 47.845 ;
        RECT 19.775 46.935 21.605 47.615 ;
        RECT 21.615 46.935 24.365 47.745 ;
        RECT 24.845 47.020 25.275 47.805 ;
        RECT 25.950 46.935 29.425 47.845 ;
        RECT 32.950 47.615 33.860 47.835 ;
        RECT 35.395 47.615 36.745 47.845 ;
        RECT 40.310 47.615 41.220 47.835 ;
        RECT 42.755 47.615 44.105 47.845 ;
        RECT 29.435 46.935 36.745 47.615 ;
        RECT 36.795 46.935 44.105 47.615 ;
        RECT 44.155 47.615 45.085 47.845 ;
        RECT 44.155 46.935 48.055 47.615 ;
        RECT 48.295 46.935 50.125 47.745 ;
        RECT 50.605 47.020 51.035 47.805 ;
        RECT 51.150 47.615 52.070 47.845 ;
        RECT 56.075 47.645 57.485 47.845 ;
        RECT 51.150 46.935 54.615 47.615 ;
        RECT 54.750 46.965 57.485 47.645 ;
        RECT 12.095 46.725 12.265 46.935 ;
        RECT 13.475 46.725 13.645 46.915 ;
        RECT 14.855 46.745 15.025 46.935 ;
        RECT 15.325 46.780 15.485 46.890 ;
        RECT 14.860 46.725 15.025 46.745 ;
        RECT 17.155 46.725 17.325 46.915 ;
        RECT 19.450 46.745 19.620 46.935 ;
        RECT 21.295 46.745 21.465 46.935 ;
        RECT 21.755 46.745 21.925 46.935 ;
        RECT 24.515 46.885 24.685 46.915 ;
        RECT 24.510 46.775 24.685 46.885 ;
        RECT 25.430 46.775 25.550 46.885 ;
        RECT 24.515 46.745 24.685 46.775 ;
        RECT 29.110 46.745 29.280 46.935 ;
        RECT 29.575 46.745 29.745 46.935 ;
        RECT 24.520 46.725 24.685 46.745 ;
        RECT 30.030 46.725 30.200 46.915 ;
        RECT 30.495 46.725 30.665 46.915 ;
        RECT 36.935 46.745 37.105 46.935 ;
        RECT 38.315 46.725 38.485 46.915 ;
        RECT 44.570 46.745 44.740 46.935 ;
        RECT 46.595 46.725 46.765 46.915 ;
        RECT 47.055 46.725 47.225 46.915 ;
        RECT 48.435 46.745 48.605 46.935 ;
        RECT 49.820 46.725 49.990 46.915 ;
        RECT 50.270 46.775 50.390 46.885 ;
        RECT 53.495 46.725 53.665 46.915 ;
        RECT 54.415 46.745 54.585 46.935 ;
        RECT 54.875 46.745 55.045 46.965 ;
        RECT 56.090 46.935 57.485 46.965 ;
        RECT 57.495 46.935 59.325 47.615 ;
        RECT 59.335 46.935 60.705 47.745 ;
        RECT 60.715 46.935 63.925 47.845 ;
        RECT 64.595 47.615 68.525 47.845 ;
        RECT 64.110 46.935 68.525 47.615 ;
        RECT 68.535 46.935 71.745 47.845 ;
        RECT 72.065 47.615 72.995 47.845 ;
        RECT 72.065 46.935 73.900 47.615 ;
        RECT 74.055 46.935 75.885 47.745 ;
        RECT 76.365 47.020 76.795 47.805 ;
        RECT 77.010 46.935 80.485 47.845 ;
        RECT 80.495 46.935 86.005 47.745 ;
        RECT 86.015 46.935 88.765 47.745 ;
        RECT 89.235 46.935 90.605 47.745 ;
        RECT 55.335 46.725 55.505 46.915 ;
        RECT 57.635 46.745 57.805 46.935 ;
        RECT 58.105 46.770 58.265 46.880 ;
        RECT 59.475 46.745 59.645 46.935 ;
        RECT 60.850 46.725 61.020 46.915 ;
        RECT 61.315 46.725 61.485 46.915 ;
        RECT 63.150 46.775 63.270 46.885 ;
        RECT 63.615 46.745 63.785 46.935 ;
        RECT 64.110 46.915 64.220 46.935 ;
        RECT 64.050 46.745 64.245 46.915 ;
        RECT 67.295 46.745 67.465 46.915 ;
        RECT 64.075 46.725 64.245 46.745 ;
        RECT 67.755 46.725 67.925 46.915 ;
        RECT 68.675 46.745 68.845 46.935 ;
        RECT 73.735 46.915 73.900 46.935 ;
        RECT 72.815 46.725 72.985 46.915 ;
        RECT 73.735 46.745 73.905 46.915 ;
        RECT 74.195 46.745 74.365 46.935 ;
        RECT 80.170 46.915 80.340 46.935 ;
        RECT 76.030 46.775 76.150 46.885 ;
        RECT 80.170 46.745 80.345 46.915 ;
        RECT 80.635 46.745 80.805 46.935 ;
        RECT 80.175 46.725 80.345 46.745 ;
        RECT 85.695 46.725 85.865 46.915 ;
        RECT 86.155 46.745 86.325 46.935 ;
        RECT 87.535 46.725 87.705 46.915 ;
        RECT 88.910 46.775 89.030 46.885 ;
        RECT 90.295 46.725 90.465 46.935 ;
        RECT 11.955 45.915 13.325 46.725 ;
        RECT 13.335 45.915 14.705 46.725 ;
        RECT 14.860 46.045 16.695 46.725 ;
        RECT 17.015 46.045 24.325 46.725 ;
        RECT 24.520 46.045 26.355 46.725 ;
        RECT 15.765 45.815 16.695 46.045 ;
        RECT 20.530 45.825 21.440 46.045 ;
        RECT 22.975 45.815 24.325 46.045 ;
        RECT 25.425 45.815 26.355 46.045 ;
        RECT 26.870 45.815 30.345 46.725 ;
        RECT 30.355 46.045 37.665 46.725 ;
        RECT 33.870 45.825 34.780 46.045 ;
        RECT 36.315 45.815 37.665 46.045 ;
        RECT 37.725 45.855 38.155 46.640 ;
        RECT 38.175 46.045 42.990 46.725 ;
        RECT 43.330 46.045 46.795 46.725 ;
        RECT 46.915 46.045 49.655 46.725 ;
        RECT 43.330 45.815 44.250 46.045 ;
        RECT 49.680 45.815 53.265 46.725 ;
        RECT 53.355 45.915 55.185 46.725 ;
        RECT 55.195 45.915 57.285 46.725 ;
        RECT 58.975 45.815 61.165 46.725 ;
        RECT 61.175 45.915 63.005 46.725 ;
        RECT 63.485 45.855 63.915 46.640 ;
        RECT 63.935 45.915 65.765 46.725 ;
        RECT 65.775 46.045 67.140 46.725 ;
        RECT 67.615 46.045 72.430 46.725 ;
        RECT 72.675 46.045 79.985 46.725 ;
        RECT 76.190 45.825 77.100 46.045 ;
        RECT 78.635 45.815 79.985 46.045 ;
        RECT 80.035 45.915 85.545 46.725 ;
        RECT 85.555 45.915 87.385 46.725 ;
        RECT 87.395 46.045 89.225 46.725 ;
        RECT 87.880 45.815 89.225 46.045 ;
        RECT 89.235 45.915 90.605 46.725 ;
      LAYER nwell ;
        RECT 11.760 42.695 90.800 45.525 ;
      LAYER pwell ;
        RECT 11.955 41.495 13.325 42.305 ;
        RECT 16.850 42.175 17.760 42.395 ;
        RECT 19.295 42.175 20.645 42.405 ;
        RECT 13.335 41.495 20.645 42.175 ;
        RECT 20.695 42.175 22.040 42.405 ;
        RECT 20.695 41.495 22.525 42.175 ;
        RECT 22.535 41.495 24.365 42.305 ;
        RECT 24.845 41.580 25.275 42.365 ;
        RECT 25.295 41.495 28.505 42.405 ;
        RECT 28.530 42.175 29.900 42.405 ;
        RECT 28.530 41.495 30.805 42.175 ;
        RECT 30.825 41.495 32.175 42.405 ;
        RECT 32.195 41.495 37.705 42.305 ;
        RECT 38.175 42.175 39.105 42.405 ;
        RECT 46.750 42.175 47.660 42.395 ;
        RECT 49.195 42.175 50.545 42.405 ;
        RECT 38.175 41.495 42.075 42.175 ;
        RECT 43.235 41.495 50.545 42.175 ;
        RECT 50.605 41.580 51.035 42.365 ;
        RECT 51.065 41.495 52.415 42.405 ;
        RECT 55.950 42.175 56.860 42.395 ;
        RECT 58.395 42.175 59.745 42.405 ;
        RECT 64.230 42.175 65.140 42.395 ;
        RECT 66.675 42.175 68.025 42.405 ;
        RECT 52.435 41.495 59.745 42.175 ;
        RECT 60.715 41.495 68.025 42.175 ;
        RECT 69.190 41.495 72.665 42.405 ;
        RECT 73.725 42.175 74.655 42.405 ;
        RECT 72.820 41.495 74.655 42.175 ;
        RECT 74.975 41.495 76.345 42.305 ;
        RECT 76.365 41.580 76.795 42.365 ;
        RECT 80.330 42.175 81.240 42.395 ;
        RECT 82.775 42.175 84.125 42.405 ;
        RECT 76.815 41.495 84.125 42.175 ;
        RECT 84.175 41.495 87.845 42.305 ;
        RECT 87.855 41.495 89.225 42.305 ;
        RECT 89.235 41.495 90.605 42.305 ;
        RECT 12.095 41.285 12.265 41.495 ;
        RECT 13.475 41.305 13.645 41.495 ;
        RECT 14.400 41.285 14.570 41.475 ;
        RECT 19.915 41.305 20.085 41.475 ;
        RECT 19.915 41.285 20.080 41.305 ;
        RECT 20.375 41.285 20.545 41.475 ;
        RECT 22.215 41.305 22.385 41.495 ;
        RECT 22.675 41.305 22.845 41.495 ;
        RECT 23.595 41.285 23.765 41.475 ;
        RECT 24.510 41.335 24.630 41.445 ;
        RECT 27.270 41.335 27.390 41.445 ;
        RECT 27.740 41.285 27.910 41.475 ;
        RECT 28.205 41.305 28.375 41.495 ;
        RECT 29.115 41.285 29.285 41.475 ;
        RECT 30.490 41.305 30.660 41.495 ;
        RECT 30.955 41.305 31.125 41.495 ;
        RECT 32.335 41.305 32.505 41.495 ;
        RECT 32.335 41.285 32.485 41.305 ;
        RECT 32.795 41.285 32.965 41.475 ;
        RECT 36.475 41.285 36.645 41.475 ;
        RECT 37.850 41.335 37.970 41.445 ;
        RECT 38.315 41.285 38.485 41.475 ;
        RECT 38.590 41.305 38.760 41.495 ;
        RECT 40.145 41.285 40.315 41.475 ;
        RECT 42.465 41.340 42.625 41.450 ;
        RECT 43.375 41.285 43.545 41.495 ;
        RECT 46.130 41.335 46.250 41.445 ;
        RECT 46.870 41.285 47.040 41.475 ;
        RECT 51.195 41.305 51.365 41.495 ;
        RECT 52.575 41.305 52.745 41.495 ;
        RECT 11.955 40.475 13.325 41.285 ;
        RECT 14.255 40.375 17.730 41.285 ;
        RECT 18.245 40.605 20.080 41.285 ;
        RECT 18.245 40.375 19.175 40.605 ;
        RECT 20.235 40.375 23.445 41.285 ;
        RECT 23.455 40.475 27.125 41.285 ;
        RECT 27.595 40.375 28.945 41.285 ;
        RECT 28.975 40.475 30.345 41.285 ;
        RECT 30.555 40.465 32.485 41.285 ;
        RECT 32.655 40.475 36.325 41.285 ;
        RECT 36.335 40.475 37.705 41.285 ;
        RECT 30.555 40.375 31.505 40.465 ;
        RECT 37.725 40.415 38.155 41.200 ;
        RECT 38.175 40.475 40.005 41.285 ;
        RECT 40.015 40.375 43.225 41.285 ;
        RECT 43.235 40.475 45.985 41.285 ;
        RECT 46.455 40.605 50.355 41.285 ;
        RECT 50.595 41.255 51.990 41.285 ;
        RECT 53.035 41.255 53.205 41.475 ;
        RECT 53.490 41.335 53.610 41.445 ;
        RECT 54.875 41.285 55.045 41.475 ;
        RECT 59.935 41.285 60.105 41.475 ;
        RECT 60.395 41.305 60.565 41.475 ;
        RECT 60.855 41.305 61.025 41.495 ;
        RECT 63.150 41.335 63.270 41.445 ;
        RECT 60.425 41.285 60.565 41.305 ;
        RECT 64.080 41.285 64.250 41.475 ;
        RECT 67.750 41.335 67.870 41.445 ;
        RECT 68.215 41.305 68.385 41.475 ;
        RECT 68.220 41.285 68.385 41.305 ;
        RECT 70.520 41.285 70.690 41.475 ;
        RECT 72.350 41.305 72.520 41.495 ;
        RECT 72.820 41.475 72.985 41.495 ;
        RECT 72.815 41.305 72.985 41.475 ;
        RECT 72.835 41.285 72.985 41.305 ;
        RECT 75.115 41.285 75.285 41.495 ;
        RECT 76.955 41.305 77.125 41.495 ;
        RECT 82.010 41.285 82.180 41.475 ;
        RECT 83.385 41.285 83.555 41.475 ;
        RECT 83.855 41.285 84.025 41.475 ;
        RECT 84.315 41.305 84.485 41.495 ;
        RECT 87.995 41.305 88.165 41.495 ;
        RECT 90.295 41.285 90.465 41.495 ;
        RECT 46.455 40.375 47.385 40.605 ;
        RECT 50.595 40.575 53.330 41.255 ;
        RECT 50.595 40.375 52.005 40.575 ;
        RECT 53.825 40.375 55.175 41.285 ;
        RECT 55.430 40.605 60.245 41.285 ;
        RECT 60.425 40.465 62.995 41.285 ;
        RECT 61.405 40.375 62.995 40.465 ;
        RECT 63.485 40.415 63.915 41.200 ;
        RECT 63.935 40.375 67.410 41.285 ;
        RECT 68.220 40.605 70.055 41.285 ;
        RECT 69.125 40.375 70.055 40.605 ;
        RECT 70.375 40.375 72.565 41.285 ;
        RECT 72.835 40.465 74.765 41.285 ;
        RECT 74.975 40.475 78.645 41.285 ;
        RECT 73.815 40.375 74.765 40.465 ;
        RECT 78.850 40.375 82.325 41.285 ;
        RECT 82.335 40.505 83.705 41.285 ;
        RECT 83.715 40.475 89.225 41.285 ;
        RECT 89.235 40.475 90.605 41.285 ;
      LAYER nwell ;
        RECT 11.760 37.255 90.800 40.085 ;
      LAYER pwell ;
        RECT 11.955 36.055 13.325 36.865 ;
        RECT 13.335 36.055 16.085 36.865 ;
        RECT 20.070 36.735 20.980 36.955 ;
        RECT 22.515 36.735 23.865 36.965 ;
        RECT 16.555 36.055 23.865 36.735 ;
        RECT 24.845 36.140 25.275 36.925 ;
        RECT 25.605 36.735 26.535 36.965 ;
        RECT 25.605 36.055 27.440 36.735 ;
        RECT 28.710 36.055 32.185 36.965 ;
        RECT 32.295 36.055 34.485 36.965 ;
        RECT 34.495 36.055 36.325 36.865 ;
        RECT 36.375 36.735 37.725 36.965 ;
        RECT 39.260 36.735 40.170 36.955 ;
        RECT 36.375 36.055 43.685 36.735 ;
        RECT 43.695 36.055 47.170 36.965 ;
        RECT 47.375 36.055 50.125 36.865 ;
        RECT 50.605 36.140 51.035 36.925 ;
        RECT 51.055 36.055 53.805 36.865 ;
        RECT 53.815 36.735 54.745 36.965 ;
        RECT 58.050 36.735 58.970 36.965 ;
        RECT 53.815 36.055 57.715 36.735 ;
        RECT 58.050 36.055 61.515 36.735 ;
        RECT 61.635 36.055 63.465 36.735 ;
        RECT 63.475 36.055 68.985 36.865 ;
        RECT 68.995 36.055 72.665 36.865 ;
        RECT 72.675 36.055 74.045 36.865 ;
        RECT 75.105 36.735 76.035 36.965 ;
        RECT 74.200 36.055 76.035 36.735 ;
        RECT 76.365 36.140 76.795 36.925 ;
        RECT 77.930 36.055 81.405 36.965 ;
        RECT 84.930 36.735 85.840 36.955 ;
        RECT 87.375 36.735 88.725 36.965 ;
        RECT 81.415 36.055 88.725 36.735 ;
        RECT 89.235 36.055 90.605 36.865 ;
        RECT 12.095 35.845 12.265 36.055 ;
        RECT 13.475 35.845 13.645 36.055 ;
        RECT 16.230 35.895 16.350 36.005 ;
        RECT 16.695 35.865 16.865 36.055 ;
        RECT 27.275 36.035 27.440 36.055 ;
        RECT 19.005 35.890 19.165 36.000 ;
        RECT 19.920 35.845 20.090 36.035 ;
        RECT 23.595 35.845 23.765 36.035 ;
        RECT 24.065 35.900 24.225 36.010 ;
        RECT 25.435 35.845 25.605 36.035 ;
        RECT 27.275 35.865 27.445 36.035 ;
        RECT 27.745 35.900 27.905 36.010 ;
        RECT 27.280 35.845 27.445 35.865 ;
        RECT 29.575 35.845 29.745 36.035 ;
        RECT 31.870 35.865 32.040 36.055 ;
        RECT 34.170 35.865 34.340 36.055 ;
        RECT 34.635 35.865 34.805 36.055 ;
        RECT 36.945 35.890 37.105 36.000 ;
        RECT 38.315 35.845 38.485 36.035 ;
        RECT 41.535 35.865 41.705 36.035 ;
        RECT 43.375 35.865 43.545 36.055 ;
        RECT 43.840 36.035 44.010 36.055 ;
        RECT 43.835 35.865 44.010 36.035 ;
        RECT 47.515 35.865 47.685 36.055 ;
        RECT 51.195 36.035 51.365 36.055 ;
        RECT 41.540 35.845 41.705 35.865 ;
        RECT 43.835 35.845 44.005 35.865 ;
        RECT 49.355 35.845 49.525 36.035 ;
        RECT 50.270 35.895 50.390 36.005 ;
        RECT 51.195 35.865 51.370 36.035 ;
        RECT 54.230 35.865 54.400 36.055 ;
        RECT 51.200 35.845 51.370 35.865 ;
        RECT 54.875 35.845 55.045 36.035 ;
        RECT 56.255 35.845 56.425 36.035 ;
        RECT 61.315 35.865 61.485 36.055 ;
        RECT 61.775 35.865 61.945 36.055 ;
        RECT 63.615 35.865 63.785 36.055 ;
        RECT 64.075 35.845 64.245 36.035 ;
        RECT 67.750 35.895 67.870 36.005 ;
        RECT 69.135 35.865 69.305 36.055 ;
        RECT 70.515 35.865 70.685 36.035 ;
        RECT 70.515 35.845 70.655 35.865 ;
        RECT 70.980 35.845 71.150 36.035 ;
        RECT 72.815 35.865 72.985 36.055 ;
        RECT 74.200 36.035 74.365 36.055 ;
        RECT 73.275 35.845 73.445 36.035 ;
        RECT 74.195 35.865 74.365 36.035 ;
        RECT 75.110 35.895 75.230 36.005 ;
        RECT 75.575 35.865 75.745 36.035 ;
        RECT 76.965 35.900 77.125 36.010 ;
        RECT 75.580 35.845 75.745 35.865 ;
        RECT 80.635 35.845 80.805 36.035 ;
        RECT 81.090 36.000 81.260 36.055 ;
        RECT 81.090 35.890 81.265 36.000 ;
        RECT 81.090 35.865 81.260 35.890 ;
        RECT 81.555 35.865 81.725 36.055 ;
        RECT 82.015 35.845 82.185 36.035 ;
        RECT 88.910 35.895 89.030 36.005 ;
        RECT 90.295 35.845 90.465 36.055 ;
        RECT 11.955 35.035 13.325 35.845 ;
        RECT 13.335 35.035 18.845 35.845 ;
        RECT 19.775 34.935 23.250 35.845 ;
        RECT 23.455 35.165 25.285 35.845 ;
        RECT 23.940 34.935 25.285 35.165 ;
        RECT 25.295 35.035 27.125 35.845 ;
        RECT 27.280 35.165 29.115 35.845 ;
        RECT 29.435 35.165 36.745 35.845 ;
        RECT 28.185 34.935 29.115 35.165 ;
        RECT 32.950 34.945 33.860 35.165 ;
        RECT 35.395 34.935 36.745 35.165 ;
        RECT 37.725 34.975 38.155 35.760 ;
        RECT 38.175 34.935 41.385 35.845 ;
        RECT 41.540 35.165 43.375 35.845 ;
        RECT 42.445 34.935 43.375 35.165 ;
        RECT 43.695 35.035 49.205 35.845 ;
        RECT 49.215 35.035 51.045 35.845 ;
        RECT 51.060 34.935 54.645 35.845 ;
        RECT 54.735 35.035 56.105 35.845 ;
        RECT 56.115 35.165 63.425 35.845 ;
        RECT 59.630 34.945 60.540 35.165 ;
        RECT 62.075 34.935 63.425 35.165 ;
        RECT 63.485 34.975 63.915 35.760 ;
        RECT 63.935 35.035 67.605 35.845 ;
        RECT 68.085 35.025 70.655 35.845 ;
        RECT 68.085 34.935 69.675 35.025 ;
        RECT 70.835 34.935 73.025 35.845 ;
        RECT 73.135 35.035 74.965 35.845 ;
        RECT 75.580 35.165 77.415 35.845 ;
        RECT 76.485 34.935 77.415 35.165 ;
        RECT 77.735 34.935 80.945 35.845 ;
        RECT 81.875 35.165 89.185 35.845 ;
        RECT 85.390 34.945 86.300 35.165 ;
        RECT 87.835 34.935 89.185 35.165 ;
        RECT 89.235 35.035 90.605 35.845 ;
      LAYER nwell ;
        RECT 11.760 31.815 90.800 34.645 ;
      LAYER pwell ;
        RECT 11.955 30.615 13.325 31.425 ;
        RECT 13.335 31.295 14.680 31.525 ;
        RECT 15.945 31.295 16.875 31.525 ;
        RECT 13.335 30.615 15.165 31.295 ;
        RECT 15.945 30.615 17.780 31.295 ;
        RECT 17.935 30.615 19.765 31.425 ;
        RECT 20.235 30.615 23.710 31.525 ;
        RECT 24.845 30.700 25.275 31.485 ;
        RECT 25.295 30.615 30.805 31.425 ;
        RECT 30.815 30.615 36.325 31.425 ;
        RECT 36.335 30.615 41.845 31.425 ;
        RECT 43.825 31.295 44.755 31.525 ;
        RECT 42.920 30.615 44.755 31.295 ;
        RECT 45.075 30.615 46.905 31.425 ;
        RECT 47.375 30.615 50.585 31.525 ;
        RECT 50.605 30.700 51.035 31.485 ;
        RECT 51.055 30.615 52.425 31.425 ;
        RECT 52.630 30.615 56.105 31.525 ;
        RECT 56.425 31.295 57.355 31.525 ;
        RECT 61.930 31.295 62.840 31.515 ;
        RECT 64.375 31.295 65.725 31.525 ;
        RECT 56.425 30.615 58.260 31.295 ;
        RECT 58.415 30.615 65.725 31.295 ;
        RECT 66.085 31.295 67.015 31.525 ;
        RECT 71.590 31.295 72.500 31.515 ;
        RECT 74.035 31.295 75.385 31.525 ;
        RECT 66.085 30.615 67.920 31.295 ;
        RECT 68.075 30.615 75.385 31.295 ;
        RECT 76.365 30.700 76.795 31.485 ;
        RECT 78.325 31.295 79.255 31.525 ;
        RECT 77.420 30.615 79.255 31.295 ;
        RECT 79.575 30.615 85.085 31.425 ;
        RECT 85.095 30.615 86.925 31.425 ;
        RECT 87.880 31.295 89.225 31.525 ;
        RECT 87.395 30.615 89.225 31.295 ;
        RECT 89.235 30.615 90.605 31.425 ;
        RECT 12.095 30.405 12.265 30.615 ;
        RECT 13.470 30.455 13.590 30.565 ;
        RECT 13.940 30.405 14.110 30.595 ;
        RECT 14.855 30.425 15.025 30.615 ;
        RECT 17.615 30.595 17.780 30.615 ;
        RECT 15.310 30.455 15.430 30.565 ;
        RECT 17.615 30.405 17.785 30.595 ;
        RECT 18.075 30.425 18.245 30.615 ;
        RECT 19.910 30.455 20.030 30.565 ;
        RECT 20.380 30.425 20.550 30.615 ;
        RECT 24.065 30.460 24.225 30.570 ;
        RECT 25.435 30.425 25.605 30.615 ;
        RECT 26.815 30.425 26.985 30.595 ;
        RECT 27.270 30.455 27.390 30.565 ;
        RECT 26.815 30.405 26.980 30.425 ;
        RECT 27.740 30.405 27.910 30.595 ;
        RECT 30.955 30.425 31.125 30.615 ;
        RECT 31.410 30.455 31.530 30.565 ;
        RECT 35.090 30.405 35.260 30.595 ;
        RECT 35.555 30.425 35.725 30.595 ;
        RECT 36.475 30.425 36.645 30.615 ;
        RECT 42.920 30.595 43.085 30.615 ;
        RECT 35.560 30.405 35.725 30.425 ;
        RECT 38.315 30.405 38.485 30.595 ;
        RECT 41.075 30.405 41.245 30.595 ;
        RECT 42.005 30.460 42.165 30.570 ;
        RECT 42.915 30.425 43.085 30.595 ;
        RECT 45.215 30.425 45.385 30.615 ;
        RECT 47.050 30.455 47.170 30.565 ;
        RECT 47.515 30.425 47.685 30.615 ;
        RECT 48.435 30.405 48.605 30.595 ;
        RECT 49.815 30.405 49.985 30.595 ;
        RECT 51.195 30.425 51.365 30.615 ;
        RECT 55.790 30.425 55.960 30.615 ;
        RECT 58.095 30.595 58.260 30.615 ;
        RECT 57.170 30.455 57.290 30.565 ;
        RECT 57.640 30.405 57.810 30.595 ;
        RECT 58.095 30.425 58.265 30.595 ;
        RECT 58.555 30.425 58.725 30.615 ;
        RECT 67.755 30.595 67.920 30.615 ;
        RECT 63.155 30.425 63.325 30.595 ;
        RECT 64.085 30.450 64.245 30.560 ;
        RECT 63.155 30.405 63.320 30.425 ;
        RECT 67.755 30.405 67.925 30.595 ;
        RECT 68.215 30.425 68.385 30.615 ;
        RECT 77.420 30.595 77.585 30.615 ;
        RECT 71.430 30.405 71.600 30.595 ;
        RECT 71.895 30.405 72.065 30.595 ;
        RECT 73.730 30.455 73.850 30.565 ;
        RECT 74.195 30.405 74.365 30.595 ;
        RECT 75.585 30.460 75.745 30.570 ;
        RECT 76.950 30.455 77.070 30.565 ;
        RECT 77.415 30.425 77.585 30.595 ;
        RECT 79.715 30.425 79.885 30.615 ;
        RECT 84.315 30.405 84.485 30.595 ;
        RECT 84.775 30.405 84.945 30.595 ;
        RECT 85.235 30.425 85.405 30.615 ;
        RECT 87.070 30.455 87.190 30.565 ;
        RECT 87.535 30.425 87.705 30.615 ;
        RECT 88.465 30.450 88.625 30.560 ;
        RECT 90.295 30.405 90.465 30.615 ;
        RECT 11.955 29.595 13.325 30.405 ;
        RECT 13.795 29.495 17.270 30.405 ;
        RECT 17.475 29.725 24.785 30.405 ;
        RECT 20.990 29.505 21.900 29.725 ;
        RECT 23.435 29.495 24.785 29.725 ;
        RECT 25.145 29.725 26.980 30.405 ;
        RECT 25.145 29.495 26.075 29.725 ;
        RECT 27.595 29.495 31.070 30.405 ;
        RECT 31.930 29.495 35.405 30.405 ;
        RECT 35.560 29.725 37.395 30.405 ;
        RECT 36.465 29.495 37.395 29.725 ;
        RECT 37.725 29.535 38.155 30.320 ;
        RECT 38.175 29.595 40.925 30.405 ;
        RECT 40.935 29.725 48.245 30.405 ;
        RECT 44.450 29.505 45.360 29.725 ;
        RECT 46.895 29.495 48.245 29.725 ;
        RECT 48.295 29.595 49.665 30.405 ;
        RECT 49.675 29.725 56.985 30.405 ;
        RECT 53.190 29.505 54.100 29.725 ;
        RECT 55.635 29.495 56.985 29.725 ;
        RECT 57.495 29.495 60.970 30.405 ;
        RECT 61.485 29.725 63.320 30.405 ;
        RECT 61.485 29.495 62.415 29.725 ;
        RECT 63.485 29.535 63.915 30.320 ;
        RECT 64.855 29.495 68.065 30.405 ;
        RECT 68.270 29.495 71.745 30.405 ;
        RECT 71.755 29.595 73.585 30.405 ;
        RECT 74.055 29.725 81.365 30.405 ;
        RECT 77.570 29.505 78.480 29.725 ;
        RECT 80.015 29.495 81.365 29.725 ;
        RECT 81.415 29.495 84.625 30.405 ;
        RECT 84.635 29.595 88.305 30.405 ;
        RECT 89.235 29.595 90.605 30.405 ;
      LAYER nwell ;
        RECT 11.760 26.375 90.800 29.205 ;
      LAYER pwell ;
        RECT 11.955 25.175 13.325 25.985 ;
        RECT 16.850 25.855 17.760 26.075 ;
        RECT 19.295 25.855 20.645 26.085 ;
        RECT 13.335 25.175 20.645 25.855 ;
        RECT 20.695 25.175 23.905 26.085 ;
        RECT 24.845 25.260 25.275 26.045 ;
        RECT 25.295 25.175 26.665 25.985 ;
        RECT 30.190 25.855 31.100 26.075 ;
        RECT 32.635 25.855 33.985 26.085 ;
        RECT 37.550 25.855 38.460 26.075 ;
        RECT 39.995 25.855 41.345 26.085 ;
        RECT 26.675 25.175 33.985 25.855 ;
        RECT 34.035 25.175 41.345 25.855 ;
        RECT 42.315 25.175 45.790 26.085 ;
        RECT 45.995 25.175 47.825 25.985 ;
        RECT 49.345 25.855 50.275 26.085 ;
        RECT 48.440 25.175 50.275 25.855 ;
        RECT 50.605 25.260 51.035 26.045 ;
        RECT 51.055 25.175 54.530 26.085 ;
        RECT 54.735 25.175 56.565 25.985 ;
        RECT 56.575 25.855 57.920 26.085 ;
        RECT 56.575 25.175 58.405 25.855 ;
        RECT 58.415 25.175 63.925 25.985 ;
        RECT 63.935 25.175 69.445 25.985 ;
        RECT 69.455 25.175 73.125 25.985 ;
        RECT 75.105 25.855 76.035 26.085 ;
        RECT 74.200 25.175 76.035 25.855 ;
        RECT 76.365 25.260 76.795 26.045 ;
        RECT 76.815 25.175 80.290 26.085 ;
        RECT 80.495 25.175 81.865 25.985 ;
        RECT 85.390 25.855 86.300 26.075 ;
        RECT 87.835 25.855 89.185 26.085 ;
        RECT 81.875 25.175 89.185 25.855 ;
        RECT 89.235 25.175 90.605 25.985 ;
        RECT 12.095 24.965 12.265 25.175 ;
        RECT 13.475 24.985 13.645 25.175 ;
        RECT 14.855 24.965 15.025 25.155 ;
        RECT 15.315 24.965 15.485 25.155 ;
        RECT 18.075 24.965 18.245 25.155 ;
        RECT 19.915 24.965 20.085 25.155 ;
        RECT 20.385 25.010 20.545 25.120 ;
        RECT 20.835 24.985 21.005 25.175 ;
        RECT 21.295 24.965 21.465 25.155 ;
        RECT 24.065 25.020 24.225 25.130 ;
        RECT 24.515 24.965 24.685 25.155 ;
        RECT 25.435 24.985 25.605 25.175 ;
        RECT 26.365 25.010 26.525 25.120 ;
        RECT 26.815 24.985 26.985 25.175 ;
        RECT 27.275 24.985 27.445 25.155 ;
        RECT 27.280 24.965 27.445 24.985 ;
        RECT 29.575 24.965 29.745 25.155 ;
        RECT 34.175 24.985 34.345 25.175 ;
        RECT 35.095 24.965 35.265 25.155 ;
        RECT 38.315 24.965 38.485 25.155 ;
        RECT 40.155 24.965 40.325 25.155 ;
        RECT 41.545 25.020 41.705 25.130 ;
        RECT 42.460 24.985 42.630 25.175 ;
        RECT 43.375 24.965 43.545 25.155 ;
        RECT 44.755 24.965 44.925 25.155 ;
        RECT 46.135 24.985 46.305 25.175 ;
        RECT 48.440 25.155 48.605 25.175 ;
        RECT 47.975 25.125 48.145 25.155 ;
        RECT 47.970 25.015 48.145 25.125 ;
        RECT 47.975 24.965 48.145 25.015 ;
        RECT 48.435 24.985 48.605 25.155 ;
        RECT 51.200 24.985 51.370 25.175 ;
        RECT 53.495 24.965 53.665 25.155 ;
        RECT 54.875 24.985 55.045 25.175 ;
        RECT 57.170 25.015 57.290 25.125 ;
        RECT 57.640 24.965 57.810 25.155 ;
        RECT 58.095 24.985 58.265 25.175 ;
        RECT 58.555 24.985 58.725 25.175 ;
        RECT 63.155 24.985 63.325 25.155 ;
        RECT 64.075 24.985 64.245 25.175 ;
        RECT 63.155 24.965 63.320 24.985 ;
        RECT 66.835 24.965 67.005 25.155 ;
        RECT 67.300 24.965 67.470 25.155 ;
        RECT 69.595 24.985 69.765 25.175 ;
        RECT 74.200 25.155 74.365 25.175 ;
        RECT 72.815 24.985 72.985 25.155 ;
        RECT 72.815 24.965 72.980 24.985 ;
        RECT 73.275 24.965 73.445 25.155 ;
        RECT 74.195 24.985 74.365 25.155 ;
        RECT 75.110 25.015 75.230 25.125 ;
        RECT 76.960 24.985 77.130 25.175 ;
        RECT 78.335 24.965 78.505 25.155 ;
        RECT 80.635 24.985 80.805 25.175 ;
        RECT 82.015 25.155 82.185 25.175 ;
        RECT 82.010 24.985 82.185 25.155 ;
        RECT 82.010 24.965 82.180 24.985 ;
        RECT 82.475 24.965 82.645 25.155 ;
        RECT 83.855 24.965 84.025 25.155 ;
        RECT 85.695 24.965 85.865 25.155 ;
        RECT 88.915 24.965 89.085 25.155 ;
        RECT 90.295 24.965 90.465 25.175 ;
        RECT 11.955 24.155 13.325 24.965 ;
        RECT 13.335 24.285 15.165 24.965 ;
        RECT 13.335 24.055 14.680 24.285 ;
        RECT 15.175 24.155 16.545 24.965 ;
        RECT 16.555 24.285 18.385 24.965 ;
        RECT 18.395 24.285 20.225 24.965 ;
        RECT 16.555 24.055 17.900 24.285 ;
        RECT 18.395 24.055 19.740 24.285 ;
        RECT 21.155 24.055 24.365 24.965 ;
        RECT 24.375 24.285 26.205 24.965 ;
        RECT 27.280 24.285 29.115 24.965 ;
        RECT 24.860 24.055 26.205 24.285 ;
        RECT 28.185 24.055 29.115 24.285 ;
        RECT 29.435 24.155 34.945 24.965 ;
        RECT 34.955 24.155 37.705 24.965 ;
        RECT 37.725 24.095 38.155 24.880 ;
        RECT 38.175 24.155 40.005 24.965 ;
        RECT 40.015 24.055 43.225 24.965 ;
        RECT 43.235 24.155 44.605 24.965 ;
        RECT 44.615 24.055 47.825 24.965 ;
        RECT 47.835 24.155 53.345 24.965 ;
        RECT 53.355 24.155 57.025 24.965 ;
        RECT 57.495 24.055 60.970 24.965 ;
        RECT 61.485 24.285 63.320 24.965 ;
        RECT 61.485 24.055 62.415 24.285 ;
        RECT 63.485 24.095 63.915 24.880 ;
        RECT 63.935 24.055 67.145 24.965 ;
        RECT 67.155 24.055 70.630 24.965 ;
        RECT 71.145 24.285 72.980 24.965 ;
        RECT 71.145 24.055 72.075 24.285 ;
        RECT 73.135 24.155 74.965 24.965 ;
        RECT 75.435 24.055 78.645 24.965 ;
        RECT 78.850 24.055 82.325 24.965 ;
        RECT 82.335 24.155 83.705 24.965 ;
        RECT 83.715 24.285 85.545 24.965 ;
        RECT 85.555 24.285 87.385 24.965 ;
        RECT 84.200 24.055 85.545 24.285 ;
        RECT 86.040 24.055 87.385 24.285 ;
        RECT 87.395 24.285 89.225 24.965 ;
        RECT 87.395 24.055 88.740 24.285 ;
        RECT 89.235 24.155 90.605 24.965 ;
      LAYER nwell ;
        RECT 11.760 20.935 90.800 23.765 ;
      LAYER pwell ;
        RECT 11.955 19.735 13.325 20.545 ;
        RECT 13.795 19.735 17.270 20.645 ;
        RECT 18.395 20.415 19.740 20.645 ;
        RECT 18.395 19.735 20.225 20.415 ;
        RECT 20.235 19.735 23.710 20.645 ;
        RECT 24.845 19.820 25.275 20.605 ;
        RECT 25.950 19.735 29.425 20.645 ;
        RECT 29.630 19.735 33.105 20.645 ;
        RECT 36.630 20.415 37.540 20.635 ;
        RECT 39.075 20.415 40.425 20.645 ;
        RECT 33.115 19.735 40.425 20.415 ;
        RECT 41.395 19.735 44.870 20.645 ;
        RECT 45.075 19.735 46.905 20.545 ;
        RECT 46.915 19.735 50.390 20.645 ;
        RECT 50.605 19.820 51.035 20.605 ;
        RECT 51.055 19.735 52.885 20.545 ;
        RECT 53.355 19.735 56.830 20.645 ;
        RECT 60.550 20.415 61.460 20.635 ;
        RECT 62.995 20.415 64.345 20.645 ;
        RECT 67.910 20.415 68.820 20.635 ;
        RECT 70.355 20.415 71.705 20.645 ;
        RECT 57.035 19.735 64.345 20.415 ;
        RECT 64.395 19.735 71.705 20.415 ;
        RECT 71.755 19.735 75.230 20.645 ;
        RECT 76.365 19.820 76.795 20.605 ;
        RECT 77.470 19.735 80.945 20.645 ;
        RECT 81.150 19.735 84.625 20.645 ;
        RECT 85.120 20.415 86.465 20.645 ;
        RECT 86.960 20.415 88.305 20.645 ;
        RECT 84.635 19.735 86.465 20.415 ;
        RECT 86.475 19.735 88.305 20.415 ;
        RECT 89.235 19.735 90.605 20.545 ;
        RECT 12.095 19.525 12.265 19.735 ;
        RECT 13.470 19.680 13.590 19.685 ;
        RECT 13.470 19.575 13.645 19.680 ;
        RECT 13.485 19.570 13.645 19.575 ;
        RECT 13.940 19.545 14.110 19.735 ;
        RECT 14.395 19.545 14.565 19.715 ;
        RECT 14.400 19.525 14.565 19.545 ;
        RECT 16.695 19.525 16.865 19.715 ;
        RECT 17.625 19.580 17.785 19.690 ;
        RECT 18.075 19.525 18.245 19.715 ;
        RECT 19.915 19.545 20.085 19.735 ;
        RECT 20.380 19.545 20.550 19.735 ;
        RECT 24.065 19.580 24.225 19.690 ;
        RECT 25.435 19.685 25.605 19.715 ;
        RECT 25.430 19.575 25.605 19.685 ;
        RECT 25.435 19.545 25.605 19.575 ;
        RECT 25.440 19.525 25.605 19.545 ;
        RECT 27.735 19.525 27.905 19.715 ;
        RECT 29.110 19.545 29.280 19.735 ;
        RECT 32.790 19.545 32.960 19.735 ;
        RECT 33.255 19.545 33.425 19.735 ;
        RECT 36.935 19.545 37.105 19.715 ;
        RECT 37.390 19.575 37.510 19.685 ;
        RECT 38.310 19.575 38.430 19.685 ;
        RECT 40.625 19.580 40.785 19.690 ;
        RECT 41.540 19.545 41.710 19.735 ;
        RECT 45.215 19.545 45.385 19.735 ;
        RECT 36.935 19.525 37.100 19.545 ;
        RECT 45.675 19.525 45.845 19.715 ;
        RECT 46.130 19.575 46.250 19.685 ;
        RECT 46.595 19.525 46.765 19.715 ;
        RECT 47.060 19.545 47.230 19.735 ;
        RECT 51.195 19.545 51.365 19.735 ;
        RECT 53.030 19.575 53.150 19.685 ;
        RECT 53.500 19.545 53.670 19.735 ;
        RECT 53.955 19.525 54.125 19.715 ;
        RECT 57.175 19.545 57.345 19.735 ;
        RECT 63.155 19.545 63.325 19.715 ;
        RECT 64.535 19.545 64.705 19.735 ;
        RECT 63.155 19.525 63.320 19.545 ;
        RECT 66.835 19.525 67.005 19.715 ;
        RECT 67.295 19.525 67.465 19.715 ;
        RECT 68.675 19.525 68.845 19.715 ;
        RECT 71.900 19.545 72.070 19.735 ;
        RECT 75.585 19.580 75.745 19.690 ;
        RECT 76.035 19.545 76.205 19.715 ;
        RECT 76.950 19.575 77.070 19.685 ;
        RECT 76.040 19.525 76.205 19.545 ;
        RECT 78.335 19.525 78.505 19.715 ;
        RECT 79.715 19.525 79.885 19.715 ;
        RECT 80.630 19.545 80.800 19.735 ;
        RECT 84.310 19.545 84.480 19.735 ;
        RECT 84.775 19.545 84.945 19.735 ;
        RECT 86.615 19.545 86.785 19.735 ;
        RECT 87.075 19.525 87.245 19.715 ;
        RECT 88.465 19.580 88.625 19.690 ;
        RECT 88.910 19.575 89.030 19.685 ;
        RECT 90.295 19.525 90.465 19.735 ;
        RECT 11.955 18.715 13.325 19.525 ;
        RECT 14.400 18.845 16.235 19.525 ;
        RECT 15.305 18.615 16.235 18.845 ;
        RECT 16.555 18.715 17.925 19.525 ;
        RECT 17.935 18.845 25.245 19.525 ;
        RECT 25.440 18.845 27.275 19.525 ;
        RECT 27.595 18.845 34.905 19.525 ;
        RECT 21.450 18.625 22.360 18.845 ;
        RECT 23.895 18.615 25.245 18.845 ;
        RECT 26.345 18.615 27.275 18.845 ;
        RECT 31.110 18.625 32.020 18.845 ;
        RECT 33.555 18.615 34.905 18.845 ;
        RECT 35.265 18.845 37.100 19.525 ;
        RECT 35.265 18.615 36.195 18.845 ;
        RECT 37.725 18.655 38.155 19.440 ;
        RECT 38.675 18.845 45.985 19.525 ;
        RECT 46.455 18.845 53.765 19.525 ;
        RECT 53.815 18.845 61.125 19.525 ;
        RECT 38.675 18.615 40.025 18.845 ;
        RECT 41.560 18.625 42.470 18.845 ;
        RECT 49.970 18.625 50.880 18.845 ;
        RECT 52.415 18.615 53.765 18.845 ;
        RECT 57.330 18.625 58.240 18.845 ;
        RECT 59.775 18.615 61.125 18.845 ;
        RECT 61.485 18.845 63.320 19.525 ;
        RECT 61.485 18.615 62.415 18.845 ;
        RECT 63.485 18.655 63.915 19.440 ;
        RECT 63.935 18.615 67.145 19.525 ;
        RECT 67.155 18.715 68.525 19.525 ;
        RECT 68.535 18.845 75.845 19.525 ;
        RECT 76.040 18.845 77.875 19.525 ;
        RECT 72.050 18.625 72.960 18.845 ;
        RECT 74.495 18.615 75.845 18.845 ;
        RECT 76.945 18.615 77.875 18.845 ;
        RECT 78.195 18.715 79.565 19.525 ;
        RECT 79.575 18.845 86.885 19.525 ;
        RECT 86.935 18.845 88.765 19.525 ;
        RECT 83.090 18.625 84.000 18.845 ;
        RECT 85.535 18.615 86.885 18.845 ;
        RECT 87.420 18.615 88.765 18.845 ;
        RECT 89.235 18.715 90.605 19.525 ;
      LAYER nwell ;
        RECT 11.760 15.495 90.800 18.325 ;
      LAYER pwell ;
        RECT 11.955 14.295 13.325 15.105 ;
        RECT 16.850 14.975 17.760 15.195 ;
        RECT 19.295 14.975 20.645 15.205 ;
        RECT 13.335 14.295 20.645 14.975 ;
        RECT 21.925 14.975 22.855 15.205 ;
        RECT 21.925 14.295 23.760 14.975 ;
        RECT 24.845 14.380 25.275 15.165 ;
        RECT 26.215 14.975 27.560 15.205 ;
        RECT 28.515 14.975 29.860 15.205 ;
        RECT 30.355 14.975 31.700 15.205 ;
        RECT 32.195 14.975 33.540 15.205 ;
        RECT 34.035 14.975 35.380 15.205 ;
        RECT 35.875 14.975 37.220 15.205 ;
        RECT 26.215 14.295 28.045 14.975 ;
        RECT 28.515 14.295 30.345 14.975 ;
        RECT 30.355 14.295 32.185 14.975 ;
        RECT 32.195 14.295 34.025 14.975 ;
        RECT 34.035 14.295 35.865 14.975 ;
        RECT 35.875 14.295 37.705 14.975 ;
        RECT 37.725 14.380 38.155 15.165 ;
        RECT 39.095 14.295 42.305 15.205 ;
        RECT 43.365 14.975 44.295 15.205 ;
        RECT 42.460 14.295 44.295 14.975 ;
        RECT 44.615 14.975 45.960 15.205 ;
        RECT 46.940 14.975 48.285 15.205 ;
        RECT 49.345 14.975 50.275 15.205 ;
        RECT 44.615 14.295 46.445 14.975 ;
        RECT 46.455 14.295 48.285 14.975 ;
        RECT 48.440 14.295 50.275 14.975 ;
        RECT 50.605 14.380 51.035 15.165 ;
        RECT 51.975 14.975 53.320 15.205 ;
        RECT 51.975 14.295 53.805 14.975 ;
        RECT 53.815 14.295 55.185 15.105 ;
        RECT 55.195 14.975 56.540 15.205 ;
        RECT 55.195 14.295 57.025 14.975 ;
        RECT 57.035 14.295 58.405 15.105 ;
        RECT 58.900 14.975 60.245 15.205 ;
        RECT 58.415 14.295 60.245 14.975 ;
        RECT 60.255 14.295 61.625 15.105 ;
        RECT 61.635 14.975 62.980 15.205 ;
        RECT 61.635 14.295 63.465 14.975 ;
        RECT 63.485 14.380 63.915 15.165 ;
        RECT 64.855 14.975 66.200 15.205 ;
        RECT 64.855 14.295 66.685 14.975 ;
        RECT 66.695 14.295 68.065 15.105 ;
        RECT 68.075 14.975 69.420 15.205 ;
        RECT 68.075 14.295 69.905 14.975 ;
        RECT 69.915 14.295 71.285 15.105 ;
        RECT 71.780 14.975 73.125 15.205 ;
        RECT 71.295 14.295 73.125 14.975 ;
        RECT 73.135 14.295 74.505 15.105 ;
        RECT 74.515 14.975 75.860 15.205 ;
        RECT 74.515 14.295 76.345 14.975 ;
        RECT 76.365 14.380 76.795 15.165 ;
        RECT 77.865 14.975 78.795 15.205 ;
        RECT 80.165 14.975 81.095 15.205 ;
        RECT 85.390 14.975 86.300 15.195 ;
        RECT 87.835 14.975 89.185 15.205 ;
        RECT 76.960 14.295 78.795 14.975 ;
        RECT 79.260 14.295 81.095 14.975 ;
        RECT 81.875 14.295 89.185 14.975 ;
        RECT 89.235 14.295 90.605 15.105 ;
        RECT 12.095 14.105 12.265 14.295 ;
        RECT 13.475 14.105 13.645 14.295 ;
        RECT 23.595 14.275 23.760 14.295 ;
        RECT 20.845 14.140 21.005 14.250 ;
        RECT 23.595 14.105 23.765 14.275 ;
        RECT 24.065 14.140 24.225 14.250 ;
        RECT 25.445 14.140 25.605 14.250 ;
        RECT 27.735 14.105 27.905 14.295 ;
        RECT 28.190 14.135 28.310 14.245 ;
        RECT 30.035 14.105 30.205 14.295 ;
        RECT 31.875 14.105 32.045 14.295 ;
        RECT 33.715 14.105 33.885 14.295 ;
        RECT 35.555 14.105 35.725 14.295 ;
        RECT 37.395 14.105 37.565 14.295 ;
        RECT 38.325 14.140 38.485 14.250 ;
        RECT 39.235 14.105 39.405 14.295 ;
        RECT 42.460 14.275 42.625 14.295 ;
        RECT 42.455 14.105 42.625 14.275 ;
        RECT 46.135 14.105 46.305 14.295 ;
        RECT 46.595 14.105 46.765 14.295 ;
        RECT 48.440 14.275 48.605 14.295 ;
        RECT 48.435 14.105 48.605 14.275 ;
        RECT 51.205 14.140 51.365 14.250 ;
        RECT 53.495 14.105 53.665 14.295 ;
        RECT 53.955 14.105 54.125 14.295 ;
        RECT 56.715 14.105 56.885 14.295 ;
        RECT 57.175 14.105 57.345 14.295 ;
        RECT 58.555 14.105 58.725 14.295 ;
        RECT 60.395 14.105 60.565 14.295 ;
        RECT 63.155 14.105 63.325 14.295 ;
        RECT 64.085 14.140 64.245 14.250 ;
        RECT 66.375 14.105 66.545 14.295 ;
        RECT 66.835 14.105 67.005 14.295 ;
        RECT 69.595 14.105 69.765 14.295 ;
        RECT 70.055 14.105 70.225 14.295 ;
        RECT 71.435 14.105 71.605 14.295 ;
        RECT 73.275 14.105 73.445 14.295 ;
        RECT 76.035 14.105 76.205 14.295 ;
        RECT 76.960 14.275 77.125 14.295 ;
        RECT 79.260 14.275 79.425 14.295 ;
        RECT 76.955 14.105 77.125 14.275 ;
        RECT 79.255 14.105 79.425 14.275 ;
        RECT 81.550 14.135 81.670 14.245 ;
        RECT 82.015 14.105 82.185 14.295 ;
        RECT 90.295 14.105 90.465 14.295 ;
      LAYER li1 ;
        RECT 112.275 219.210 112.445 219.295 ;
        RECT 114.995 219.210 115.165 219.295 ;
        RECT 117.715 219.210 117.885 219.295 ;
        RECT 120.435 219.210 120.605 219.295 ;
        RECT 123.155 219.210 123.325 219.295 ;
        RECT 125.875 219.210 126.045 219.295 ;
        RECT 128.595 219.210 128.765 219.295 ;
        RECT 131.315 219.210 131.485 219.295 ;
        RECT 134.035 219.210 134.205 219.295 ;
        RECT 136.755 219.210 136.925 219.295 ;
        RECT 139.475 219.210 139.645 219.295 ;
        RECT 142.195 219.210 142.365 219.295 ;
        RECT 144.915 219.210 145.085 219.295 ;
        RECT 147.635 219.210 147.805 219.295 ;
        RECT 112.275 218.690 113.735 219.210 ;
        RECT 112.275 218.000 113.195 218.690 ;
        RECT 113.905 218.520 116.255 219.210 ;
        RECT 116.425 218.690 119.175 219.210 ;
        RECT 113.365 218.000 116.795 218.520 ;
        RECT 116.965 218.000 118.635 218.690 ;
        RECT 119.345 218.520 121.695 219.210 ;
        RECT 121.865 218.690 124.615 219.210 ;
        RECT 118.805 218.000 122.235 218.520 ;
        RECT 122.405 218.000 124.075 218.690 ;
        RECT 124.785 218.520 127.135 219.210 ;
        RECT 127.305 218.690 130.055 219.210 ;
        RECT 124.245 218.000 127.675 218.520 ;
        RECT 127.845 218.000 129.515 218.690 ;
        RECT 130.225 218.520 132.575 219.210 ;
        RECT 132.745 218.690 135.495 219.210 ;
        RECT 129.685 218.000 133.115 218.520 ;
        RECT 133.285 218.000 134.955 218.690 ;
        RECT 135.665 218.520 138.015 219.210 ;
        RECT 138.185 218.690 140.935 219.210 ;
        RECT 135.125 218.000 138.555 218.520 ;
        RECT 138.725 218.000 140.395 218.690 ;
        RECT 141.105 218.520 143.455 219.210 ;
        RECT 143.625 218.690 146.375 219.210 ;
        RECT 140.565 218.000 143.995 218.520 ;
        RECT 144.165 218.000 145.835 218.690 ;
        RECT 146.545 218.520 147.805 219.210 ;
        RECT 146.005 218.000 147.805 218.520 ;
        RECT 112.275 217.830 112.445 218.000 ;
        RECT 114.995 217.830 115.165 218.000 ;
        RECT 112.275 216.245 112.990 217.830 ;
        RECT 114.560 217.825 115.165 217.830 ;
        RECT 117.715 217.825 117.885 218.000 ;
        RECT 114.560 217.565 116.315 217.825 ;
        RECT 116.875 217.565 117.885 217.825 ;
        RECT 118.540 217.780 119.375 217.830 ;
        RECT 114.560 216.965 115.165 217.565 ;
        RECT 115.335 217.220 117.545 217.390 ;
        RECT 115.335 217.135 116.240 217.220 ;
        RECT 116.970 217.135 117.545 217.220 ;
        RECT 117.715 217.280 117.885 217.565 ;
        RECT 118.105 217.770 119.375 217.780 ;
        RECT 120.435 217.825 120.605 218.000 ;
        RECT 123.155 217.825 123.325 218.000 ;
        RECT 125.875 217.825 126.045 218.000 ;
        RECT 128.595 217.830 128.765 218.000 ;
        RECT 131.315 217.830 131.485 218.000 ;
        RECT 128.595 217.825 130.055 217.830 ;
        RECT 118.105 217.660 120.220 217.770 ;
        RECT 118.105 217.605 118.665 217.660 ;
        RECT 119.245 217.615 120.220 217.660 ;
        RECT 118.105 217.450 118.625 217.605 ;
        RECT 117.715 217.110 118.495 217.280 ;
        RECT 116.475 216.965 116.805 217.050 ;
        RECT 117.715 216.965 117.885 217.110 ;
        RECT 114.560 216.635 115.925 216.965 ;
        RECT 116.095 216.795 117.165 216.965 ;
        RECT 112.275 215.905 113.820 216.245 ;
        RECT 112.275 212.485 112.990 215.905 ;
        RECT 114.560 214.560 115.165 216.635 ;
        RECT 116.095 216.420 116.265 216.795 ;
        RECT 115.335 216.250 116.265 216.420 ;
        RECT 116.445 216.160 116.815 216.515 ;
        RECT 116.995 216.420 117.165 216.795 ;
        RECT 117.335 216.635 117.885 216.965 ;
        RECT 118.795 216.940 119.125 217.490 ;
        RECT 119.295 217.440 120.220 217.615 ;
        RECT 120.435 217.565 121.755 217.825 ;
        RECT 122.315 217.565 123.325 217.825 ;
        RECT 123.585 217.570 124.045 217.740 ;
        RECT 120.435 217.270 120.605 217.565 ;
        RECT 123.155 217.400 123.325 217.565 ;
        RECT 119.425 217.100 120.605 217.270 ;
        RECT 120.775 217.220 122.985 217.390 ;
        RECT 120.775 217.135 121.680 217.220 ;
        RECT 122.410 217.135 122.985 217.220 ;
        RECT 116.995 216.250 117.545 216.420 ;
        RECT 117.715 216.350 117.885 216.635 ;
        RECT 118.100 216.930 119.125 216.940 ;
        RECT 120.435 216.965 120.605 217.100 ;
        RECT 123.155 217.070 123.705 217.400 ;
        RECT 123.875 217.305 124.045 217.570 ;
        RECT 124.215 217.475 124.865 217.825 ;
        RECT 125.035 217.570 125.705 217.740 ;
        RECT 125.035 217.305 125.205 217.570 ;
        RECT 125.875 217.565 127.195 217.825 ;
        RECT 127.755 217.565 130.055 217.825 ;
        RECT 125.875 217.400 126.045 217.565 ;
        RECT 123.875 217.075 125.205 217.305 ;
        RECT 125.375 217.070 126.045 217.400 ;
        RECT 126.215 217.220 128.425 217.390 ;
        RECT 126.215 217.135 127.120 217.220 ;
        RECT 127.850 217.135 128.425 217.220 ;
        RECT 128.595 217.310 130.055 217.565 ;
        RECT 121.915 216.965 122.245 217.050 ;
        RECT 123.155 216.965 123.325 217.070 ;
        RECT 118.100 216.740 120.265 216.930 ;
        RECT 118.100 216.610 118.625 216.740 ;
        RECT 119.330 216.590 120.265 216.740 ;
        RECT 120.435 216.635 121.365 216.965 ;
        RECT 121.535 216.795 122.605 216.965 ;
        RECT 117.715 216.140 118.415 216.350 ;
        RECT 115.335 214.895 117.545 215.065 ;
        RECT 115.335 214.730 116.305 214.895 ;
        RECT 116.975 214.810 117.545 214.895 ;
        RECT 116.475 214.640 116.805 214.725 ;
        RECT 117.715 214.640 117.885 216.140 ;
        RECT 118.795 215.865 119.125 216.570 ;
        RECT 119.330 216.035 119.705 216.590 ;
        RECT 120.435 216.360 120.605 216.635 ;
        RECT 121.535 216.420 121.705 216.795 ;
        RECT 119.935 216.045 120.605 216.360 ;
        RECT 120.775 216.250 121.705 216.420 ;
        RECT 121.885 216.160 122.255 216.515 ;
        RECT 122.435 216.420 122.605 216.795 ;
        RECT 122.775 216.635 123.325 216.965 ;
        RECT 125.875 216.965 126.045 217.070 ;
        RECT 127.355 216.965 127.685 217.050 ;
        RECT 128.595 216.965 129.515 217.310 ;
        RECT 130.225 217.270 131.485 217.830 ;
        RECT 132.545 217.780 133.380 217.830 ;
        RECT 132.545 217.770 133.815 217.780 ;
        RECT 131.700 217.660 133.815 217.770 ;
        RECT 131.700 217.615 132.675 217.660 ;
        RECT 131.700 217.440 132.625 217.615 ;
        RECT 133.255 217.605 133.815 217.660 ;
        RECT 130.225 217.140 132.495 217.270 ;
        RECT 123.585 216.715 125.705 216.900 ;
        RECT 123.155 216.460 123.325 216.635 ;
        RECT 125.875 216.635 126.805 216.965 ;
        RECT 126.975 216.795 128.045 216.965 ;
        RECT 122.435 216.250 122.985 216.420 ;
        RECT 123.155 216.210 123.785 216.460 ;
        RECT 123.955 216.265 124.905 216.545 ;
        RECT 125.875 216.475 126.045 216.635 ;
        RECT 125.415 216.210 126.045 216.475 ;
        RECT 126.975 216.420 127.145 216.795 ;
        RECT 126.215 216.250 127.145 216.420 ;
        RECT 118.165 215.695 120.135 215.865 ;
        RECT 118.165 215.080 118.335 215.695 ;
        RECT 118.505 215.205 119.795 215.525 ;
        RECT 118.505 215.060 118.835 215.205 ;
        RECT 114.560 214.425 116.305 214.560 ;
        RECT 116.475 214.470 117.145 214.640 ;
        RECT 113.310 214.390 116.305 214.425 ;
        RECT 113.310 214.075 115.165 214.390 ;
        RECT 116.475 214.220 116.805 214.245 ;
        RECT 114.560 212.485 115.165 214.075 ;
        RECT 112.275 212.310 112.445 212.485 ;
        RECT 114.995 212.310 115.165 212.485 ;
        RECT 112.275 210.660 113.735 212.310 ;
        RECT 113.905 212.020 115.165 212.310 ;
        RECT 115.335 214.050 116.805 214.220 ;
        RECT 115.335 212.360 115.505 214.050 ;
        RECT 116.975 213.885 117.145 214.470 ;
        RECT 117.315 214.325 117.885 214.640 ;
        RECT 118.165 214.675 118.335 214.910 ;
        RECT 119.045 214.845 119.765 215.035 ;
        RECT 119.965 214.980 120.135 215.695 ;
        RECT 119.935 214.675 120.265 214.755 ;
        RECT 118.165 214.505 120.265 214.675 ;
        RECT 117.315 214.310 118.385 214.325 ;
        RECT 117.715 213.955 118.385 214.310 ;
        RECT 118.565 214.045 118.865 214.505 ;
        RECT 120.435 214.500 120.605 216.045 ;
        RECT 120.775 214.670 121.455 214.955 ;
        RECT 120.435 214.335 121.065 214.500 ;
        RECT 119.045 214.165 119.375 214.335 ;
        RECT 119.635 214.230 121.065 214.335 ;
        RECT 119.635 214.165 120.605 214.230 ;
        RECT 116.975 213.880 117.545 213.885 ;
        RECT 115.675 213.710 117.545 213.880 ;
        RECT 115.675 212.755 115.845 213.710 ;
        RECT 116.015 213.370 116.985 213.540 ;
        RECT 116.015 212.720 116.185 213.370 ;
        RECT 117.180 213.355 117.545 213.710 ;
        RECT 117.205 213.165 117.375 213.170 ;
        RECT 116.385 212.890 117.545 213.165 ;
        RECT 116.015 212.530 117.545 212.720 ;
        RECT 115.335 212.190 116.360 212.360 ;
        RECT 117.715 212.350 117.885 213.955 ;
        RECT 118.565 213.845 118.895 214.045 ;
        RECT 119.115 213.995 119.375 214.165 ;
        RECT 119.115 213.825 120.160 213.995 ;
        RECT 119.115 213.635 119.285 213.825 ;
        RECT 118.165 213.465 119.285 213.635 ;
        RECT 118.165 212.960 118.335 213.465 ;
        RECT 119.455 213.295 119.820 213.655 ;
        RECT 118.535 213.125 119.820 213.295 ;
        RECT 118.535 212.770 118.755 213.125 ;
        RECT 118.165 212.600 118.335 212.765 ;
        RECT 118.925 212.715 119.520 212.955 ;
        RECT 119.990 212.890 120.160 213.825 ;
        RECT 118.165 212.545 118.605 212.600 ;
        RECT 119.710 212.545 120.265 212.680 ;
        RECT 118.165 212.430 120.265 212.545 ;
        RECT 120.435 212.440 120.605 214.165 ;
        RECT 121.235 214.210 121.455 214.670 ;
        RECT 121.625 214.380 122.185 215.070 ;
        RECT 122.355 214.670 122.985 214.955 ;
        RECT 122.355 214.210 122.525 214.670 ;
        RECT 123.155 214.515 123.325 216.210 ;
        RECT 123.915 216.040 125.280 216.095 ;
        RECT 123.605 215.925 125.705 216.040 ;
        RECT 123.605 215.870 124.045 215.925 ;
        RECT 123.605 215.705 123.775 215.870 ;
        RECT 125.150 215.790 125.705 215.925 ;
        RECT 123.605 215.005 123.775 215.510 ;
        RECT 123.975 215.345 124.195 215.700 ;
        RECT 124.365 215.515 124.960 215.755 ;
        RECT 123.975 215.175 125.260 215.345 ;
        RECT 123.605 214.835 124.725 215.005 ;
        RECT 124.555 214.645 124.725 214.835 ;
        RECT 124.895 214.815 125.260 215.175 ;
        RECT 125.430 214.645 125.600 215.580 ;
        RECT 123.155 214.500 123.825 214.515 ;
        RECT 122.695 214.230 123.825 214.500 ;
        RECT 121.235 214.000 122.525 214.210 ;
        RECT 123.155 214.145 123.825 214.230 ;
        RECT 124.005 214.425 124.335 214.625 ;
        RECT 124.555 214.475 125.600 214.645 ;
        RECT 125.875 215.020 126.045 216.210 ;
        RECT 127.325 216.160 127.695 216.515 ;
        RECT 127.875 216.420 128.045 216.795 ;
        RECT 128.215 216.635 129.515 216.965 ;
        RECT 128.595 216.620 129.515 216.635 ;
        RECT 129.685 217.100 132.495 217.140 ;
        RECT 129.685 216.620 131.485 217.100 ;
        RECT 132.795 216.940 133.125 217.490 ;
        RECT 133.295 217.450 133.815 217.605 ;
        RECT 134.035 217.400 134.205 218.000 ;
        RECT 136.755 217.825 136.925 218.000 ;
        RECT 139.475 217.825 139.645 218.000 ;
        RECT 142.195 217.830 142.365 218.000 ;
        RECT 144.915 217.830 145.085 218.000 ;
        RECT 147.635 217.830 147.805 218.000 ;
        RECT 134.375 217.655 136.585 217.825 ;
        RECT 134.375 217.570 134.945 217.655 ;
        RECT 135.615 217.490 136.585 217.655 ;
        RECT 136.755 217.565 138.075 217.825 ;
        RECT 138.635 217.565 139.645 217.825 ;
        RECT 139.905 217.570 140.365 217.740 ;
        RECT 135.115 217.400 135.445 217.485 ;
        RECT 134.035 217.280 134.605 217.400 ;
        RECT 133.425 217.110 134.605 217.280 ;
        RECT 134.035 217.070 134.605 217.110 ;
        RECT 134.775 217.230 135.445 217.400 ;
        RECT 136.755 217.320 136.925 217.565 ;
        RECT 139.475 217.400 139.645 217.565 ;
        RECT 132.795 216.930 133.820 216.940 ;
        RECT 127.875 216.250 128.425 216.420 ;
        RECT 128.595 215.880 128.765 216.620 ;
        RECT 128.935 216.050 129.565 216.335 ;
        RECT 128.595 215.610 129.225 215.880 ;
        RECT 126.215 215.355 128.425 215.525 ;
        RECT 126.215 215.190 127.185 215.355 ;
        RECT 127.855 215.270 128.425 215.355 ;
        RECT 127.355 215.100 127.685 215.185 ;
        RECT 128.595 215.100 128.765 215.610 ;
        RECT 129.395 215.590 129.565 216.050 ;
        RECT 129.735 215.760 130.295 216.450 ;
        RECT 131.315 216.360 131.485 216.620 ;
        RECT 131.655 216.740 133.820 216.930 ;
        RECT 131.655 216.590 132.590 216.740 ;
        RECT 133.295 216.610 133.820 216.740 ;
        RECT 130.465 216.050 131.145 216.335 ;
        RECT 130.465 215.590 130.685 216.050 ;
        RECT 131.315 216.045 131.985 216.360 ;
        RECT 131.315 215.880 131.485 216.045 ;
        RECT 132.215 216.035 132.590 216.590 ;
        RECT 130.855 215.610 131.485 215.880 ;
        RECT 132.795 215.865 133.125 216.570 ;
        RECT 134.035 216.350 134.205 217.070 ;
        RECT 134.775 216.645 134.945 217.230 ;
        RECT 135.615 217.150 136.925 217.320 ;
        RECT 135.115 216.980 135.445 217.005 ;
        RECT 135.115 216.810 136.585 216.980 ;
        RECT 133.505 216.140 134.205 216.350 ;
        RECT 129.395 215.380 130.685 215.590 ;
        RECT 125.875 214.850 127.185 215.020 ;
        RECT 127.355 214.930 128.025 215.100 ;
        RECT 120.775 213.430 122.985 213.830 ;
        RECT 120.775 212.960 121.455 213.240 ;
        RECT 121.235 212.565 121.455 212.960 ;
        RECT 121.625 212.735 122.185 213.430 ;
        RECT 122.355 212.960 122.985 213.240 ;
        RECT 122.355 212.565 122.525 212.960 ;
        RECT 118.475 212.375 119.840 212.430 ;
        RECT 113.905 211.850 115.925 212.020 ;
        RECT 113.905 210.930 115.165 211.850 ;
        RECT 115.515 211.440 115.925 211.615 ;
        RECT 116.170 211.610 116.360 212.190 ;
        RECT 116.735 211.620 116.905 212.330 ;
        RECT 117.180 212.260 117.885 212.350 ;
        RECT 120.435 212.260 121.065 212.440 ;
        RECT 117.180 212.010 118.345 212.260 ;
        RECT 117.180 211.840 117.885 212.010 ;
        RECT 118.515 211.925 119.465 212.205 ;
        RECT 119.975 212.115 121.065 212.260 ;
        RECT 121.235 212.115 122.525 212.565 ;
        RECT 123.155 212.440 123.325 214.145 ;
        RECT 124.005 213.965 124.305 214.425 ;
        RECT 124.555 214.305 124.815 214.475 ;
        RECT 125.875 214.305 126.045 214.850 ;
        RECT 127.355 214.680 127.685 214.705 ;
        RECT 124.485 214.135 124.815 214.305 ;
        RECT 125.075 214.135 126.045 214.305 ;
        RECT 123.605 213.795 125.705 213.965 ;
        RECT 123.605 213.560 123.775 213.795 ;
        RECT 125.375 213.715 125.705 213.795 ;
        RECT 124.485 213.435 125.205 213.625 ;
        RECT 123.605 212.775 123.775 213.390 ;
        RECT 123.945 213.265 124.275 213.410 ;
        RECT 123.945 212.945 125.235 213.265 ;
        RECT 125.405 212.775 125.575 213.490 ;
        RECT 123.605 212.605 125.575 212.775 ;
        RECT 122.695 212.330 123.325 212.440 ;
        RECT 122.695 212.120 123.855 212.330 ;
        RECT 122.695 212.115 123.325 212.120 ;
        RECT 119.975 211.995 120.605 212.115 ;
        RECT 121.915 212.010 122.245 212.115 ;
        RECT 116.735 211.440 117.510 211.620 ;
        RECT 115.515 211.375 117.510 211.440 ;
        RECT 117.715 211.400 117.885 211.840 ;
        RECT 118.145 211.570 120.265 211.755 ;
        RECT 120.435 211.400 120.605 211.995 ;
        RECT 120.775 211.840 121.745 211.945 ;
        RECT 122.415 211.840 122.985 211.945 ;
        RECT 120.775 211.560 122.985 211.840 ;
        RECT 115.515 211.100 116.905 211.375 ;
        RECT 117.715 211.070 118.265 211.400 ;
        RECT 118.435 211.165 119.765 211.395 ;
        RECT 117.715 210.930 117.885 211.070 ;
        RECT 112.275 208.800 113.215 210.660 ;
        RECT 113.905 210.490 116.255 210.930 ;
        RECT 113.385 209.110 116.255 210.490 ;
        RECT 116.425 210.470 117.885 210.930 ;
        RECT 118.435 210.900 118.605 211.165 ;
        RECT 118.145 210.730 118.605 210.900 ;
        RECT 118.775 210.645 119.425 210.995 ;
        RECT 119.595 210.900 119.765 211.165 ;
        RECT 119.935 211.070 120.605 211.400 ;
        RECT 119.595 210.730 120.265 210.900 ;
        RECT 120.435 210.470 120.605 211.070 ;
        RECT 123.155 211.360 123.325 212.115 ;
        RECT 124.235 211.900 124.565 212.605 ;
        RECT 125.875 212.480 126.045 214.135 ;
        RECT 126.215 214.510 127.685 214.680 ;
        RECT 126.215 212.820 126.385 214.510 ;
        RECT 127.855 214.345 128.025 214.930 ;
        RECT 128.195 214.770 128.765 215.100 ;
        RECT 128.935 214.810 131.145 215.210 ;
        RECT 127.855 214.340 128.425 214.345 ;
        RECT 126.555 214.170 128.425 214.340 ;
        RECT 126.555 213.215 126.725 214.170 ;
        RECT 126.895 213.830 127.865 214.000 ;
        RECT 126.895 213.180 127.065 213.830 ;
        RECT 128.060 213.815 128.425 214.170 ;
        RECT 128.595 213.820 128.765 214.770 ;
        RECT 128.935 214.340 129.565 214.620 ;
        RECT 129.395 213.945 129.565 214.340 ;
        RECT 129.735 214.115 130.295 214.810 ;
        RECT 130.465 214.340 131.145 214.620 ;
        RECT 130.465 213.945 130.685 214.340 ;
        RECT 128.085 213.625 128.255 213.630 ;
        RECT 127.265 213.350 128.425 213.625 ;
        RECT 128.595 213.495 129.225 213.820 ;
        RECT 129.395 213.495 130.685 213.945 ;
        RECT 131.315 214.335 131.485 215.610 ;
        RECT 131.785 215.695 133.755 215.865 ;
        RECT 131.785 214.980 131.955 215.695 ;
        RECT 132.125 215.205 133.415 215.525 ;
        RECT 133.085 215.060 133.415 215.205 ;
        RECT 133.585 215.080 133.755 215.695 ;
        RECT 134.035 215.110 134.205 216.140 ;
        RECT 134.375 216.640 134.945 216.645 ;
        RECT 134.375 216.470 136.245 216.640 ;
        RECT 134.375 216.115 134.740 216.470 ;
        RECT 134.935 216.130 135.905 216.300 ;
        RECT 134.545 215.925 134.715 215.930 ;
        RECT 134.375 215.650 135.535 215.925 ;
        RECT 135.735 215.480 135.905 216.130 ;
        RECT 136.075 215.515 136.245 216.470 ;
        RECT 134.375 215.290 135.905 215.480 ;
        RECT 136.415 215.120 136.585 216.810 ;
        RECT 132.155 214.845 132.875 215.035 ;
        RECT 131.655 214.675 131.985 214.755 ;
        RECT 133.585 214.675 133.755 214.910 ;
        RECT 131.655 214.505 133.755 214.675 ;
        RECT 134.035 214.600 134.740 215.110 ;
        RECT 131.315 214.165 132.285 214.335 ;
        RECT 132.545 214.165 132.875 214.335 ;
        RECT 131.315 213.820 131.485 214.165 ;
        RECT 132.545 213.995 132.805 214.165 ;
        RECT 133.055 214.045 133.355 214.505 ;
        RECT 134.035 214.325 134.205 214.600 ;
        RECT 135.015 214.380 135.185 215.090 ;
        RECT 130.855 213.495 131.485 213.820 ;
        RECT 126.895 212.990 128.425 213.180 ;
        RECT 126.215 212.650 127.240 212.820 ;
        RECT 128.595 212.810 128.765 213.495 ;
        RECT 129.675 213.390 130.005 213.495 ;
        RECT 128.935 213.220 129.505 213.325 ;
        RECT 130.175 213.220 131.145 213.325 ;
        RECT 128.935 212.940 131.145 213.220 ;
        RECT 124.770 211.880 125.145 212.435 ;
        RECT 125.875 212.425 126.805 212.480 ;
        RECT 125.375 212.310 126.805 212.425 ;
        RECT 125.375 212.110 126.045 212.310 ;
        RECT 123.540 211.730 124.065 211.860 ;
        RECT 124.770 211.730 125.705 211.880 ;
        RECT 123.540 211.540 125.705 211.730 ;
        RECT 123.540 211.530 124.565 211.540 ;
        RECT 123.155 211.190 123.935 211.360 ;
        RECT 123.155 210.470 123.325 211.190 ;
        RECT 123.545 210.865 124.065 211.020 ;
        RECT 124.235 210.980 124.565 211.530 ;
        RECT 125.875 211.370 126.045 212.110 ;
        RECT 126.395 211.900 126.805 212.075 ;
        RECT 127.050 212.070 127.240 212.650 ;
        RECT 127.615 212.080 127.785 212.790 ;
        RECT 128.060 212.300 128.765 212.810 ;
        RECT 128.935 212.490 131.145 212.770 ;
        RECT 128.935 212.385 129.505 212.490 ;
        RECT 130.175 212.385 131.145 212.490 ;
        RECT 128.595 212.215 128.765 212.300 ;
        RECT 129.675 212.215 130.005 212.320 ;
        RECT 131.315 212.260 131.485 213.495 ;
        RECT 131.760 213.825 132.805 213.995 ;
        RECT 133.025 213.845 133.355 214.045 ;
        RECT 133.535 213.955 134.205 214.325 ;
        RECT 134.410 214.200 135.185 214.380 ;
        RECT 135.560 214.950 136.585 215.120 ;
        RECT 136.755 216.965 136.925 217.150 ;
        RECT 137.095 217.220 139.305 217.390 ;
        RECT 137.095 217.135 138.000 217.220 ;
        RECT 138.730 217.135 139.305 217.220 ;
        RECT 139.475 217.070 140.025 217.400 ;
        RECT 140.195 217.305 140.365 217.570 ;
        RECT 140.535 217.475 141.185 217.825 ;
        RECT 141.355 217.570 142.025 217.740 ;
        RECT 141.355 217.305 141.525 217.570 ;
        RECT 142.195 217.400 143.455 217.830 ;
        RECT 140.195 217.075 141.525 217.305 ;
        RECT 141.695 217.070 143.455 217.400 ;
        RECT 138.235 216.965 138.565 217.050 ;
        RECT 139.475 216.965 139.645 217.070 ;
        RECT 136.755 216.635 137.685 216.965 ;
        RECT 137.855 216.795 138.925 216.965 ;
        RECT 136.755 215.480 136.925 216.635 ;
        RECT 137.855 216.420 138.025 216.795 ;
        RECT 137.095 216.250 138.025 216.420 ;
        RECT 138.205 216.160 138.575 216.515 ;
        RECT 138.755 216.420 138.925 216.795 ;
        RECT 139.095 216.635 139.645 216.965 ;
        RECT 139.905 216.715 142.025 216.900 ;
        RECT 139.475 216.460 139.645 216.635 ;
        RECT 138.755 216.250 139.305 216.420 ;
        RECT 139.475 216.210 140.105 216.460 ;
        RECT 140.275 216.265 141.225 216.545 ;
        RECT 142.195 216.475 143.455 217.070 ;
        RECT 141.735 216.210 143.455 216.475 ;
        RECT 137.095 215.815 139.305 215.985 ;
        RECT 137.095 215.650 138.065 215.815 ;
        RECT 138.735 215.730 139.305 215.815 ;
        RECT 138.235 215.560 138.565 215.645 ;
        RECT 139.475 215.560 139.645 216.210 ;
        RECT 140.235 216.040 141.600 216.095 ;
        RECT 139.925 215.925 142.025 216.040 ;
        RECT 139.925 215.870 140.365 215.925 ;
        RECT 139.925 215.705 140.095 215.870 ;
        RECT 141.470 215.790 142.025 215.925 ;
        RECT 142.195 216.010 143.455 216.210 ;
        RECT 143.625 216.245 145.630 217.830 ;
        RECT 143.625 216.180 146.460 216.245 ;
        RECT 136.755 215.310 138.065 215.480 ;
        RECT 138.235 215.390 138.905 215.560 ;
        RECT 135.560 214.370 135.750 214.950 ;
        RECT 136.755 214.780 136.925 215.310 ;
        RECT 138.235 215.140 138.565 215.165 ;
        RECT 135.995 214.610 136.925 214.780 ;
        RECT 135.995 214.200 136.405 214.375 ;
        RECT 134.410 214.135 136.405 214.200 ;
        RECT 131.760 212.890 131.930 213.825 ;
        RECT 132.100 213.295 132.465 213.655 ;
        RECT 132.635 213.635 132.805 213.825 ;
        RECT 132.635 213.465 133.755 213.635 ;
        RECT 132.100 213.125 133.385 213.295 ;
        RECT 132.400 212.715 132.995 212.955 ;
        RECT 133.165 212.770 133.385 213.125 ;
        RECT 133.585 212.960 133.755 213.465 ;
        RECT 134.035 213.260 134.205 213.955 ;
        RECT 135.015 213.860 136.405 214.135 ;
        RECT 134.465 213.430 134.925 213.600 ;
        RECT 134.035 212.930 134.585 213.260 ;
        RECT 134.755 213.165 134.925 213.430 ;
        RECT 135.095 213.335 135.745 213.685 ;
        RECT 135.915 213.430 136.585 213.600 ;
        RECT 135.915 213.165 136.085 213.430 ;
        RECT 136.755 213.260 136.925 214.610 ;
        RECT 134.755 212.935 136.085 213.165 ;
        RECT 136.255 212.940 136.925 213.260 ;
        RECT 137.095 214.970 138.565 215.140 ;
        RECT 137.095 213.280 137.265 214.970 ;
        RECT 138.735 214.805 138.905 215.390 ;
        RECT 139.075 215.230 139.645 215.560 ;
        RECT 138.735 214.800 139.305 214.805 ;
        RECT 137.435 214.630 139.305 214.800 ;
        RECT 137.435 213.675 137.605 214.630 ;
        RECT 137.775 214.290 138.745 214.460 ;
        RECT 137.775 213.640 137.945 214.290 ;
        RECT 138.940 214.275 139.305 214.630 ;
        RECT 139.475 214.515 139.645 215.230 ;
        RECT 139.925 215.005 140.095 215.510 ;
        RECT 140.295 215.345 140.515 215.700 ;
        RECT 140.685 215.515 141.280 215.755 ;
        RECT 140.295 215.175 141.580 215.345 ;
        RECT 139.925 214.835 141.045 215.005 ;
        RECT 140.875 214.645 141.045 214.835 ;
        RECT 141.215 214.815 141.580 215.175 ;
        RECT 141.750 214.645 141.920 215.580 ;
        RECT 139.475 214.145 140.145 214.515 ;
        RECT 140.325 214.425 140.655 214.625 ;
        RECT 140.875 214.475 141.920 214.645 ;
        RECT 138.965 214.085 139.135 214.090 ;
        RECT 138.145 213.810 139.305 214.085 ;
        RECT 137.775 213.450 139.305 213.640 ;
        RECT 137.095 213.110 138.120 213.280 ;
        RECT 139.475 213.270 139.645 214.145 ;
        RECT 140.325 213.965 140.625 214.425 ;
        RECT 140.875 214.305 141.135 214.475 ;
        RECT 142.195 214.320 143.975 216.010 ;
        RECT 144.145 215.905 146.460 216.180 ;
        RECT 144.145 214.320 145.630 215.905 ;
        RECT 147.200 214.425 147.805 217.830 ;
        RECT 142.195 214.305 142.365 214.320 ;
        RECT 140.805 214.135 141.135 214.305 ;
        RECT 141.395 214.135 142.365 214.305 ;
        RECT 139.925 213.795 142.025 213.965 ;
        RECT 139.925 213.560 140.095 213.795 ;
        RECT 141.695 213.715 142.025 213.795 ;
        RECT 140.805 213.435 141.525 213.625 ;
        RECT 136.255 212.930 137.685 212.940 ;
        RECT 131.655 212.545 132.210 212.680 ;
        RECT 133.585 212.600 133.755 212.765 ;
        RECT 133.315 212.545 133.755 212.600 ;
        RECT 131.655 212.430 133.755 212.545 ;
        RECT 132.080 212.375 133.445 212.430 ;
        RECT 134.035 212.320 134.205 212.930 ;
        RECT 136.755 212.770 137.685 212.930 ;
        RECT 134.465 212.575 136.585 212.760 ;
        RECT 134.035 212.260 134.665 212.320 ;
        RECT 131.315 212.215 131.945 212.260 ;
        RECT 127.615 211.900 128.390 212.080 ;
        RECT 126.395 211.835 128.390 211.900 ;
        RECT 128.595 211.890 129.225 212.215 ;
        RECT 126.395 211.560 127.785 211.835 ;
        RECT 124.865 211.200 126.045 211.370 ;
        RECT 123.545 210.810 124.105 210.865 ;
        RECT 124.735 210.855 125.660 211.030 ;
        RECT 124.685 210.810 125.660 210.855 ;
        RECT 123.545 210.700 125.660 210.810 ;
        RECT 125.875 210.960 126.045 211.200 ;
        RECT 126.215 211.130 126.885 211.300 ;
        RECT 123.545 210.690 124.815 210.700 ;
        RECT 123.980 210.640 124.815 210.690 ;
        RECT 125.875 210.630 126.545 210.960 ;
        RECT 126.715 210.865 126.885 211.130 ;
        RECT 127.055 211.035 127.705 211.385 ;
        RECT 127.875 211.130 128.335 211.300 ;
        RECT 127.875 210.865 128.045 211.130 ;
        RECT 128.595 210.960 128.765 211.890 ;
        RECT 129.395 211.765 130.685 212.215 ;
        RECT 130.855 211.995 131.945 212.215 ;
        RECT 130.855 211.890 131.485 211.995 ;
        RECT 132.455 211.925 133.405 212.205 ;
        RECT 133.575 212.070 134.665 212.260 ;
        RECT 134.835 212.125 135.785 212.405 ;
        RECT 136.755 212.335 136.925 212.770 ;
        RECT 136.295 212.070 136.925 212.335 ;
        RECT 133.575 212.010 134.205 212.070 ;
        RECT 129.395 211.370 129.565 211.765 ;
        RECT 128.935 211.090 129.565 211.370 ;
        RECT 126.715 210.635 128.045 210.865 ;
        RECT 128.215 210.630 128.765 210.960 ;
        RECT 129.735 210.900 130.295 211.595 ;
        RECT 130.465 211.370 130.685 211.765 ;
        RECT 131.315 211.400 131.485 211.890 ;
        RECT 131.655 211.570 133.775 211.755 ;
        RECT 134.035 211.400 134.205 212.010 ;
        RECT 134.795 211.900 136.160 211.955 ;
        RECT 134.485 211.785 136.585 211.900 ;
        RECT 134.485 211.730 134.925 211.785 ;
        RECT 134.485 211.565 134.655 211.730 ;
        RECT 136.030 211.650 136.585 211.785 ;
        RECT 136.755 211.850 136.925 212.070 ;
        RECT 137.275 212.360 137.685 212.535 ;
        RECT 137.930 212.530 138.120 213.110 ;
        RECT 138.495 212.540 138.665 213.250 ;
        RECT 138.940 212.760 139.645 213.270 ;
        RECT 138.495 212.360 139.270 212.540 ;
        RECT 137.275 212.295 139.270 212.360 ;
        RECT 139.475 212.330 139.645 212.760 ;
        RECT 139.925 212.775 140.095 213.390 ;
        RECT 140.265 213.265 140.595 213.410 ;
        RECT 140.265 212.945 141.555 213.265 ;
        RECT 141.725 212.775 141.895 213.490 ;
        RECT 139.925 212.605 141.895 212.775 ;
        RECT 142.195 213.130 142.365 214.135 ;
        RECT 143.425 213.640 144.260 213.690 ;
        RECT 143.425 213.630 144.695 213.640 ;
        RECT 142.580 213.520 144.695 213.630 ;
        RECT 142.580 213.475 143.555 213.520 ;
        RECT 142.580 213.300 143.505 213.475 ;
        RECT 144.135 213.465 144.695 213.520 ;
        RECT 142.195 212.960 143.375 213.130 ;
        RECT 137.275 212.020 138.665 212.295 ;
        RECT 139.475 212.120 140.175 212.330 ;
        RECT 139.475 211.850 139.645 212.120 ;
        RECT 140.555 211.900 140.885 212.605 ;
        RECT 141.090 211.880 141.465 212.435 ;
        RECT 142.195 212.425 142.365 212.960 ;
        RECT 143.675 212.800 144.005 213.350 ;
        RECT 144.175 213.310 144.695 213.465 ;
        RECT 144.915 213.140 145.630 214.320 ;
        RECT 145.950 214.075 147.805 214.425 ;
        RECT 144.305 212.970 145.630 213.140 ;
        RECT 143.675 212.790 144.700 212.800 ;
        RECT 142.535 212.600 144.700 212.790 ;
        RECT 142.535 212.450 143.470 212.600 ;
        RECT 144.175 212.470 144.700 212.600 ;
        RECT 144.915 212.485 145.630 212.970 ;
        RECT 147.200 212.485 147.805 214.075 ;
        RECT 141.695 212.220 142.365 212.425 ;
        RECT 141.695 212.110 142.865 212.220 ;
        RECT 142.195 211.905 142.865 212.110 ;
        RECT 130.465 211.090 131.145 211.370 ;
        RECT 131.315 211.070 131.985 211.400 ;
        RECT 132.155 211.165 133.485 211.395 ;
        RECT 125.875 210.470 126.045 210.630 ;
        RECT 116.425 209.280 119.175 210.470 ;
        RECT 113.385 208.800 116.775 209.110 ;
        RECT 112.275 207.695 112.445 208.800 ;
        RECT 112.615 207.910 113.165 208.080 ;
        RECT 112.275 207.365 112.825 207.695 ;
        RECT 112.995 207.535 113.165 207.910 ;
        RECT 113.345 207.815 113.715 208.170 ;
        RECT 113.895 207.910 114.825 208.080 ;
        RECT 113.895 207.535 114.065 207.910 ;
        RECT 114.995 207.695 116.775 208.800 ;
        RECT 112.995 207.365 114.065 207.535 ;
        RECT 114.235 207.420 116.775 207.695 ;
        RECT 116.945 208.820 119.175 209.280 ;
        RECT 119.345 209.900 120.605 210.470 ;
        RECT 120.775 210.070 121.455 210.355 ;
        RECT 119.345 209.630 121.065 209.900 ;
        RECT 116.945 207.420 118.655 208.820 ;
        RECT 119.345 208.650 120.605 209.630 ;
        RECT 121.235 209.610 121.455 210.070 ;
        RECT 121.625 209.780 122.185 210.470 ;
        RECT 122.355 210.070 122.985 210.355 ;
        RECT 122.355 209.610 122.525 210.070 ;
        RECT 123.155 209.900 124.615 210.470 ;
        RECT 122.695 209.630 124.615 209.900 ;
        RECT 121.235 209.400 122.525 209.610 ;
        RECT 120.775 208.830 122.985 209.230 ;
        RECT 114.235 207.365 115.165 207.420 ;
        RECT 112.275 206.765 112.445 207.365 ;
        RECT 113.355 207.280 113.685 207.365 ;
        RECT 114.995 207.250 115.165 207.365 ;
        RECT 117.715 207.250 118.655 207.420 ;
        RECT 112.615 207.110 113.190 207.195 ;
        RECT 113.920 207.110 114.825 207.195 ;
        RECT 112.615 206.940 114.825 207.110 ;
        RECT 114.995 206.765 116.255 207.250 ;
        RECT 112.275 206.505 113.285 206.765 ;
        RECT 113.845 206.560 116.255 206.765 ;
        RECT 116.425 206.960 118.655 207.250 ;
        RECT 118.825 207.840 120.605 208.650 ;
        RECT 120.775 208.360 121.455 208.640 ;
        RECT 121.235 207.965 121.455 208.360 ;
        RECT 121.625 208.135 122.185 208.830 ;
        RECT 123.155 208.820 124.615 209.630 ;
        RECT 124.785 210.035 126.045 210.470 ;
        RECT 126.215 210.275 128.335 210.460 ;
        RECT 124.785 209.770 126.505 210.035 ;
        RECT 127.015 209.825 127.965 210.105 ;
        RECT 128.595 210.100 128.765 210.630 ;
        RECT 128.935 210.500 131.145 210.900 ;
        RECT 131.315 210.470 131.485 211.070 ;
        RECT 132.155 210.900 132.325 211.165 ;
        RECT 131.655 210.730 132.325 210.900 ;
        RECT 132.495 210.645 133.145 210.995 ;
        RECT 133.315 210.900 133.485 211.165 ;
        RECT 133.655 211.070 134.205 211.400 ;
        RECT 133.315 210.730 133.775 210.900 ;
        RECT 134.035 210.470 134.205 211.070 ;
        RECT 134.485 210.865 134.655 211.370 ;
        RECT 134.855 211.205 135.075 211.560 ;
        RECT 135.245 211.375 135.840 211.615 ;
        RECT 134.855 211.035 136.140 211.205 ;
        RECT 134.485 210.695 135.605 210.865 ;
        RECT 135.435 210.505 135.605 210.695 ;
        RECT 135.775 210.675 136.140 211.035 ;
        RECT 136.310 210.505 136.480 211.440 ;
        RECT 129.395 210.120 130.685 210.330 ;
        RECT 128.595 210.020 129.225 210.100 ;
        RECT 128.135 209.830 129.225 210.020 ;
        RECT 128.135 209.770 128.765 209.830 ;
        RECT 122.355 208.360 122.985 208.640 ;
        RECT 122.355 207.965 122.525 208.360 ;
        RECT 118.825 207.515 121.065 207.840 ;
        RECT 121.235 207.515 122.525 207.965 ;
        RECT 123.155 207.840 124.095 208.820 ;
        RECT 124.785 208.650 126.045 209.770 ;
        RECT 126.640 209.600 128.005 209.655 ;
        RECT 126.215 209.485 128.315 209.600 ;
        RECT 126.215 209.350 126.770 209.485 ;
        RECT 127.875 209.430 128.315 209.485 ;
        RECT 122.695 207.515 124.095 207.840 ;
        RECT 118.825 206.960 120.605 207.515 ;
        RECT 121.915 207.410 122.245 207.515 ;
        RECT 120.775 207.240 121.745 207.345 ;
        RECT 122.415 207.240 122.985 207.345 ;
        RECT 120.775 206.960 122.985 207.240 ;
        RECT 123.155 206.960 124.095 207.515 ;
        RECT 124.265 207.865 126.045 208.650 ;
        RECT 126.320 208.205 126.490 209.140 ;
        RECT 126.960 209.075 127.555 209.315 ;
        RECT 128.145 209.265 128.315 209.430 ;
        RECT 127.725 208.905 127.945 209.260 ;
        RECT 128.595 209.090 128.765 209.770 ;
        RECT 129.395 209.660 129.565 210.120 ;
        RECT 128.935 209.375 129.565 209.660 ;
        RECT 129.735 209.260 130.295 209.950 ;
        RECT 130.465 209.660 130.685 210.120 ;
        RECT 131.315 210.100 132.575 210.470 ;
        RECT 130.855 209.830 132.575 210.100 ;
        RECT 130.465 209.375 131.145 209.660 ;
        RECT 131.315 209.090 132.575 209.830 ;
        RECT 132.745 210.375 134.205 210.470 ;
        RECT 132.745 210.005 134.705 210.375 ;
        RECT 134.885 210.285 135.215 210.485 ;
        RECT 135.435 210.335 136.480 210.505 ;
        RECT 136.755 211.160 138.015 211.850 ;
        RECT 138.185 211.360 139.645 211.850 ;
        RECT 139.860 211.730 140.385 211.860 ;
        RECT 141.090 211.730 142.025 211.880 ;
        RECT 139.860 211.540 142.025 211.730 ;
        RECT 139.860 211.530 140.885 211.540 ;
        RECT 138.185 211.330 140.255 211.360 ;
        RECT 138.725 211.190 140.255 211.330 ;
        RECT 136.755 210.640 138.555 211.160 ;
        RECT 138.725 210.640 139.645 211.190 ;
        RECT 139.865 210.865 140.385 211.020 ;
        RECT 140.555 210.980 140.885 211.530 ;
        RECT 142.195 211.370 142.365 211.905 ;
        RECT 143.095 211.895 143.470 212.450 ;
        RECT 143.675 211.725 144.005 212.430 ;
        RECT 144.915 212.210 145.085 212.485 ;
        RECT 144.385 212.000 145.085 212.210 ;
        RECT 141.185 211.200 142.365 211.370 ;
        RECT 139.865 210.810 140.425 210.865 ;
        RECT 141.055 210.855 141.980 211.030 ;
        RECT 141.005 210.810 141.980 210.855 ;
        RECT 139.865 210.700 141.980 210.810 ;
        RECT 139.865 210.690 141.135 210.700 ;
        RECT 140.300 210.640 141.135 210.690 ;
        RECT 136.755 210.380 136.925 210.640 ;
        RECT 139.475 210.380 139.645 210.640 ;
        RECT 132.745 209.260 134.205 210.005 ;
        RECT 134.885 209.825 135.185 210.285 ;
        RECT 135.435 210.165 135.695 210.335 ;
        RECT 136.755 210.165 137.670 210.380 ;
        RECT 135.365 209.995 135.695 210.165 ;
        RECT 135.955 210.110 137.670 210.165 ;
        RECT 135.955 209.995 136.925 210.110 ;
        RECT 134.485 209.655 136.585 209.825 ;
        RECT 134.485 209.420 134.655 209.655 ;
        RECT 136.255 209.575 136.585 209.655 ;
        RECT 135.365 209.295 136.085 209.485 ;
        RECT 136.755 209.480 136.925 209.995 ;
        RECT 137.840 209.940 138.825 210.380 ;
        RECT 138.995 210.080 139.645 210.380 ;
        RECT 139.815 210.190 142.025 210.470 ;
        RECT 139.815 210.085 140.385 210.190 ;
        RECT 141.055 210.085 142.025 210.190 ;
        RECT 142.195 210.195 142.365 211.200 ;
        RECT 142.665 211.555 144.635 211.725 ;
        RECT 142.665 210.840 142.835 211.555 ;
        RECT 143.005 211.065 144.295 211.385 ;
        RECT 143.965 210.920 144.295 211.065 ;
        RECT 144.465 210.940 144.635 211.555 ;
        RECT 144.915 210.915 145.085 212.000 ;
        RECT 145.255 211.130 145.805 211.300 ;
        RECT 143.035 210.705 143.755 210.895 ;
        RECT 142.535 210.535 142.865 210.615 ;
        RECT 144.465 210.535 144.635 210.770 ;
        RECT 142.535 210.365 144.635 210.535 ;
        RECT 144.915 210.585 145.465 210.915 ;
        RECT 145.635 210.755 145.805 211.130 ;
        RECT 145.985 211.035 146.355 211.390 ;
        RECT 146.535 211.130 147.465 211.300 ;
        RECT 146.535 210.755 146.705 211.130 ;
        RECT 147.635 210.915 147.805 212.485 ;
        RECT 145.635 210.585 146.705 210.755 ;
        RECT 146.875 210.585 147.805 210.915 ;
        RECT 137.100 209.910 138.825 209.940 ;
        RECT 139.475 209.915 139.645 210.080 ;
        RECT 142.195 210.025 143.165 210.195 ;
        RECT 143.425 210.025 143.755 210.195 ;
        RECT 140.555 209.915 140.885 210.020 ;
        RECT 142.195 209.915 142.365 210.025 ;
        RECT 137.100 209.650 139.280 209.910 ;
        RECT 126.660 208.735 127.945 208.905 ;
        RECT 126.660 208.375 127.025 208.735 ;
        RECT 128.145 208.565 128.315 209.070 ;
        RECT 127.195 208.395 128.315 208.565 ;
        RECT 127.195 208.205 127.365 208.395 ;
        RECT 126.320 208.035 127.365 208.205 ;
        RECT 127.105 207.865 127.365 208.035 ;
        RECT 127.585 207.985 127.915 208.185 ;
        RECT 128.595 208.075 130.055 209.090 ;
        RECT 124.265 207.695 126.845 207.865 ;
        RECT 127.105 207.695 127.435 207.865 ;
        RECT 124.265 206.960 126.045 207.695 ;
        RECT 127.615 207.525 127.915 207.985 ;
        RECT 128.095 207.880 130.055 208.075 ;
        RECT 130.225 207.880 133.095 209.090 ;
        RECT 133.265 208.190 134.205 209.260 ;
        RECT 134.485 208.635 134.655 209.250 ;
        RECT 134.825 209.125 135.155 209.270 ;
        RECT 134.825 208.805 136.115 209.125 ;
        RECT 136.285 208.635 136.455 209.350 ;
        RECT 134.485 208.465 136.455 208.635 ;
        RECT 136.755 209.225 137.655 209.480 ;
        RECT 136.755 208.610 136.930 209.225 ;
        RECT 137.840 209.215 138.825 209.650 ;
        RECT 139.475 209.590 140.105 209.915 ;
        RECT 139.475 209.480 139.645 209.590 ;
        RECT 138.995 209.220 139.645 209.480 ;
        RECT 137.840 209.040 138.065 209.215 ;
        RECT 137.100 208.780 138.065 209.040 ;
        RECT 133.265 207.980 134.735 208.190 ;
        RECT 133.265 207.880 134.205 207.980 ;
        RECT 128.095 207.705 129.535 207.880 ;
        RECT 130.225 207.710 131.485 207.880 ;
        RECT 126.215 207.355 128.315 207.525 ;
        RECT 126.215 207.275 126.545 207.355 ;
        RECT 116.425 206.730 117.885 206.960 ;
        RECT 113.845 206.505 116.795 206.560 ;
        RECT 112.275 206.330 112.445 206.505 ;
        RECT 114.995 206.330 116.795 206.505 ;
        RECT 112.275 206.040 113.170 206.330 ;
        RECT 113.830 206.040 116.795 206.330 ;
        RECT 116.965 206.330 117.885 206.730 ;
        RECT 120.435 206.330 120.605 206.960 ;
        RECT 116.965 206.040 118.610 206.330 ;
        RECT 119.270 206.040 120.605 206.330 ;
        RECT 120.955 206.515 122.345 206.790 ;
        RECT 120.955 206.450 122.950 206.515 ;
        RECT 120.955 206.275 121.365 206.450 ;
        RECT 112.275 205.405 112.445 206.040 ;
        RECT 114.995 205.405 115.165 206.040 ;
        RECT 117.715 205.870 117.885 206.040 ;
        RECT 120.435 205.870 121.365 206.040 ;
        RECT 116.225 205.820 117.060 205.870 ;
        RECT 116.225 205.810 117.495 205.820 ;
        RECT 115.380 205.700 117.495 205.810 ;
        RECT 115.380 205.655 116.355 205.700 ;
        RECT 115.380 205.480 116.305 205.655 ;
        RECT 116.935 205.645 117.495 205.700 ;
        RECT 112.275 205.145 113.285 205.405 ;
        RECT 113.845 205.310 115.165 205.405 ;
        RECT 113.845 205.145 116.175 205.310 ;
        RECT 112.275 204.545 112.445 205.145 ;
        RECT 114.995 205.140 116.175 205.145 ;
        RECT 112.615 204.800 114.825 204.970 ;
        RECT 112.615 204.715 113.190 204.800 ;
        RECT 113.920 204.715 114.825 204.800 ;
        RECT 113.355 204.545 113.685 204.630 ;
        RECT 114.995 204.545 115.165 205.140 ;
        RECT 116.475 204.980 116.805 205.530 ;
        RECT 116.975 205.490 117.495 205.645 ;
        RECT 117.715 205.565 118.395 205.870 ;
        RECT 117.715 205.320 117.885 205.565 ;
        RECT 118.565 205.555 119.125 205.870 ;
        RECT 120.435 205.860 120.605 205.870 ;
        RECT 119.625 205.565 120.605 205.860 ;
        RECT 121.610 205.700 121.800 206.280 ;
        RECT 117.105 205.150 117.885 205.320 ;
        RECT 116.475 204.970 117.500 204.980 ;
        RECT 115.335 204.780 117.500 204.970 ;
        RECT 115.335 204.630 116.270 204.780 ;
        RECT 116.975 204.650 117.500 204.780 ;
        RECT 117.715 204.965 117.885 205.150 ;
        RECT 118.065 205.140 120.265 205.385 ;
        RECT 118.065 205.135 119.125 205.140 ;
        RECT 117.715 204.705 118.410 204.965 ;
        RECT 112.275 204.215 112.825 204.545 ;
        RECT 112.995 204.375 114.065 204.545 ;
        RECT 112.275 203.140 112.445 204.215 ;
        RECT 112.995 204.000 113.165 204.375 ;
        RECT 112.615 203.830 113.165 204.000 ;
        RECT 113.345 203.740 113.715 204.095 ;
        RECT 113.895 204.000 114.065 204.375 ;
        RECT 114.235 204.400 115.165 204.545 ;
        RECT 114.235 204.215 115.665 204.400 ;
        RECT 114.995 204.085 115.665 204.215 ;
        RECT 113.895 203.830 114.825 204.000 ;
        RECT 112.705 203.310 113.165 203.480 ;
        RECT 112.275 202.810 112.825 203.140 ;
        RECT 112.995 203.045 113.165 203.310 ;
        RECT 113.335 203.215 113.985 203.565 ;
        RECT 114.155 203.310 114.825 203.480 ;
        RECT 114.155 203.045 114.325 203.310 ;
        RECT 114.995 203.140 115.165 204.085 ;
        RECT 115.895 204.075 116.270 204.630 ;
        RECT 116.475 203.905 116.805 204.610 ;
        RECT 117.715 204.390 117.885 204.705 ;
        RECT 118.875 204.525 119.125 205.135 ;
        RECT 120.435 204.965 120.605 205.565 ;
        RECT 119.625 204.705 120.605 204.965 ;
        RECT 117.185 204.180 117.885 204.390 ;
        RECT 118.065 204.275 120.260 204.525 ;
        RECT 117.715 204.105 117.885 204.180 ;
        RECT 112.995 202.815 114.325 203.045 ;
        RECT 114.495 202.810 115.165 203.140 ;
        RECT 115.465 203.735 117.435 203.905 ;
        RECT 115.465 203.020 115.635 203.735 ;
        RECT 115.805 203.245 117.095 203.565 ;
        RECT 116.765 203.100 117.095 203.245 ;
        RECT 117.265 203.120 117.435 203.735 ;
        RECT 117.715 203.845 118.445 204.105 ;
        RECT 117.715 203.245 117.885 203.845 ;
        RECT 118.080 203.415 118.705 203.675 ;
        RECT 115.835 202.885 116.555 203.075 ;
        RECT 117.715 202.985 118.365 203.245 ;
        RECT 112.275 202.200 112.445 202.810 ;
        RECT 112.705 202.455 114.825 202.640 ;
        RECT 114.995 202.375 115.165 202.810 ;
        RECT 115.335 202.715 115.665 202.795 ;
        RECT 117.265 202.715 117.435 202.950 ;
        RECT 115.335 202.545 117.435 202.715 ;
        RECT 11.950 201.785 90.610 201.955 ;
        RECT 112.275 201.950 112.905 202.200 ;
        RECT 113.075 202.005 114.025 202.285 ;
        RECT 114.995 202.215 115.965 202.375 ;
        RECT 114.535 202.205 115.965 202.215 ;
        RECT 116.225 202.205 116.555 202.375 ;
        RECT 114.535 201.950 115.165 202.205 ;
        RECT 116.225 202.035 116.485 202.205 ;
        RECT 116.735 202.085 117.035 202.545 ;
        RECT 117.715 202.385 117.885 202.985 ;
        RECT 118.535 202.815 118.705 203.415 ;
        RECT 118.080 202.555 118.705 202.815 ;
        RECT 117.715 202.365 118.365 202.385 ;
        RECT 12.035 200.695 13.245 201.785 ;
        RECT 13.415 201.350 18.760 201.785 ;
        RECT 18.935 201.350 24.280 201.785 ;
        RECT 12.035 199.985 12.555 200.525 ;
        RECT 12.725 200.155 13.245 200.695 ;
        RECT 12.035 199.235 13.245 199.985 ;
        RECT 15.000 199.780 15.340 200.610 ;
        RECT 16.820 200.100 17.170 201.350 ;
        RECT 20.520 199.780 20.860 200.610 ;
        RECT 22.340 200.100 22.690 201.350 ;
        RECT 24.915 200.620 25.205 201.785 ;
        RECT 25.375 201.350 30.720 201.785 ;
        RECT 30.895 201.350 36.240 201.785 ;
        RECT 13.415 199.235 18.760 199.780 ;
        RECT 18.935 199.235 24.280 199.780 ;
        RECT 24.915 199.235 25.205 199.960 ;
        RECT 26.960 199.780 27.300 200.610 ;
        RECT 28.780 200.100 29.130 201.350 ;
        RECT 32.480 199.780 32.820 200.610 ;
        RECT 34.300 200.100 34.650 201.350 ;
        RECT 36.415 200.695 37.625 201.785 ;
        RECT 36.415 199.985 36.935 200.525 ;
        RECT 37.105 200.155 37.625 200.695 ;
        RECT 37.795 200.620 38.085 201.785 ;
        RECT 38.255 201.350 43.600 201.785 ;
        RECT 43.775 201.350 49.120 201.785 ;
        RECT 25.375 199.235 30.720 199.780 ;
        RECT 30.895 199.235 36.240 199.780 ;
        RECT 36.415 199.235 37.625 199.985 ;
        RECT 37.795 199.235 38.085 199.960 ;
        RECT 39.840 199.780 40.180 200.610 ;
        RECT 41.660 200.100 42.010 201.350 ;
        RECT 45.360 199.780 45.700 200.610 ;
        RECT 47.180 200.100 47.530 201.350 ;
        RECT 49.295 200.695 50.505 201.785 ;
        RECT 49.295 199.985 49.815 200.525 ;
        RECT 49.985 200.155 50.505 200.695 ;
        RECT 50.675 200.620 50.965 201.785 ;
        RECT 51.135 201.350 56.480 201.785 ;
        RECT 38.255 199.235 43.600 199.780 ;
        RECT 43.775 199.235 49.120 199.780 ;
        RECT 49.295 199.235 50.505 199.985 ;
        RECT 50.675 199.235 50.965 199.960 ;
        RECT 52.720 199.780 53.060 200.610 ;
        RECT 54.540 200.100 54.890 201.350 ;
        RECT 56.655 200.915 56.930 201.615 ;
        RECT 57.100 201.240 57.355 201.785 ;
        RECT 57.525 201.275 58.005 201.615 ;
        RECT 58.180 201.230 58.785 201.785 ;
        RECT 58.170 201.130 58.785 201.230 ;
        RECT 58.170 201.105 58.355 201.130 ;
        RECT 56.655 199.885 56.825 200.915 ;
        RECT 57.100 200.785 57.855 201.035 ;
        RECT 58.025 200.860 58.355 201.105 ;
        RECT 57.100 200.750 57.870 200.785 ;
        RECT 57.100 200.740 57.885 200.750 ;
        RECT 56.995 200.725 57.890 200.740 ;
        RECT 56.995 200.710 57.910 200.725 ;
        RECT 56.995 200.700 57.930 200.710 ;
        RECT 56.995 200.690 57.955 200.700 ;
        RECT 56.995 200.660 58.025 200.690 ;
        RECT 56.995 200.630 58.045 200.660 ;
        RECT 56.995 200.600 58.065 200.630 ;
        RECT 56.995 200.575 58.095 200.600 ;
        RECT 56.995 200.540 58.130 200.575 ;
        RECT 56.995 200.535 58.160 200.540 ;
        RECT 56.995 200.140 57.225 200.535 ;
        RECT 57.770 200.530 58.160 200.535 ;
        RECT 57.795 200.520 58.160 200.530 ;
        RECT 57.810 200.515 58.160 200.520 ;
        RECT 57.825 200.510 58.160 200.515 ;
        RECT 58.525 200.510 58.785 200.960 ;
        RECT 58.955 200.695 61.545 201.785 ;
        RECT 57.825 200.505 58.785 200.510 ;
        RECT 57.835 200.495 58.785 200.505 ;
        RECT 57.845 200.490 58.785 200.495 ;
        RECT 57.855 200.480 58.785 200.490 ;
        RECT 57.860 200.470 58.785 200.480 ;
        RECT 57.865 200.465 58.785 200.470 ;
        RECT 57.875 200.450 58.785 200.465 ;
        RECT 57.880 200.435 58.785 200.450 ;
        RECT 57.890 200.410 58.785 200.435 ;
        RECT 57.395 199.940 57.725 200.365 ;
        RECT 51.135 199.235 56.480 199.780 ;
        RECT 56.655 199.405 56.915 199.885 ;
        RECT 57.085 199.235 57.335 199.775 ;
        RECT 57.505 199.455 57.725 199.940 ;
        RECT 57.895 200.340 58.785 200.410 ;
        RECT 57.895 199.615 58.065 200.340 ;
        RECT 58.235 199.785 58.785 200.170 ;
        RECT 58.955 200.005 60.165 200.525 ;
        RECT 60.335 200.175 61.545 200.695 ;
        RECT 61.805 200.855 61.975 201.615 ;
        RECT 62.155 201.025 62.485 201.785 ;
        RECT 61.805 200.685 62.470 200.855 ;
        RECT 62.655 200.710 62.925 201.615 ;
        RECT 62.300 200.540 62.470 200.685 ;
        RECT 61.735 200.135 62.065 200.505 ;
        RECT 62.300 200.210 62.585 200.540 ;
        RECT 57.895 199.445 58.785 199.615 ;
        RECT 58.955 199.235 61.545 200.005 ;
        RECT 62.300 199.955 62.470 200.210 ;
        RECT 61.805 199.785 62.470 199.955 ;
        RECT 62.755 199.910 62.925 200.710 ;
        RECT 63.555 200.620 63.845 201.785 ;
        RECT 64.015 201.350 69.360 201.785 ;
        RECT 61.805 199.405 61.975 199.785 ;
        RECT 62.155 199.235 62.485 199.615 ;
        RECT 62.665 199.405 62.925 199.910 ;
        RECT 63.555 199.235 63.845 199.960 ;
        RECT 65.600 199.780 65.940 200.610 ;
        RECT 67.420 200.100 67.770 201.350 ;
        RECT 69.535 200.695 71.205 201.785 ;
        RECT 69.535 200.005 70.285 200.525 ;
        RECT 70.455 200.175 71.205 200.695 ;
        RECT 71.375 200.710 71.645 201.615 ;
        RECT 71.815 201.025 72.145 201.785 ;
        RECT 72.325 200.855 72.495 201.615 ;
        RECT 64.015 199.235 69.360 199.780 ;
        RECT 69.535 199.235 71.205 200.005 ;
        RECT 71.375 199.910 71.545 200.710 ;
        RECT 71.830 200.685 72.495 200.855 ;
        RECT 72.755 200.695 76.265 201.785 ;
        RECT 71.830 200.540 72.000 200.685 ;
        RECT 71.715 200.210 72.000 200.540 ;
        RECT 71.830 199.955 72.000 200.210 ;
        RECT 72.235 200.135 72.565 200.505 ;
        RECT 72.755 200.005 74.405 200.525 ;
        RECT 74.575 200.175 76.265 200.695 ;
        RECT 76.435 200.620 76.725 201.785 ;
        RECT 76.895 201.350 82.240 201.785 ;
        RECT 82.415 201.350 87.760 201.785 ;
        RECT 71.375 199.405 71.635 199.910 ;
        RECT 71.830 199.785 72.495 199.955 ;
        RECT 71.815 199.235 72.145 199.615 ;
        RECT 72.325 199.405 72.495 199.785 ;
        RECT 72.755 199.235 76.265 200.005 ;
        RECT 76.435 199.235 76.725 199.960 ;
        RECT 78.480 199.780 78.820 200.610 ;
        RECT 80.300 200.100 80.650 201.350 ;
        RECT 84.000 199.780 84.340 200.610 ;
        RECT 85.820 200.100 86.170 201.350 ;
        RECT 87.935 200.695 89.145 201.785 ;
        RECT 87.935 199.985 88.455 200.525 ;
        RECT 88.625 200.155 89.145 200.695 ;
        RECT 89.315 200.695 90.525 201.785 ;
        RECT 89.315 200.155 89.835 200.695 ;
        RECT 90.005 199.985 90.525 200.525 ;
        RECT 76.895 199.235 82.240 199.780 ;
        RECT 82.415 199.235 87.760 199.780 ;
        RECT 87.935 199.235 89.145 199.985 ;
        RECT 89.315 199.235 90.525 199.985 ;
        RECT 112.275 200.255 112.445 201.950 ;
        RECT 113.035 201.780 114.400 201.835 ;
        RECT 112.725 201.665 114.825 201.780 ;
        RECT 112.725 201.610 113.165 201.665 ;
        RECT 112.725 201.445 112.895 201.610 ;
        RECT 114.270 201.530 114.825 201.665 ;
        RECT 112.725 200.745 112.895 201.250 ;
        RECT 113.095 201.085 113.315 201.440 ;
        RECT 113.485 201.255 114.080 201.495 ;
        RECT 113.095 200.915 114.380 201.085 ;
        RECT 112.725 200.575 113.845 200.745 ;
        RECT 113.675 200.385 113.845 200.575 ;
        RECT 114.015 200.555 114.380 200.915 ;
        RECT 114.550 200.385 114.720 201.320 ;
        RECT 112.275 199.885 112.945 200.255 ;
        RECT 113.125 200.165 113.455 200.365 ;
        RECT 113.675 200.215 114.720 200.385 ;
        RECT 114.995 200.300 115.165 201.950 ;
        RECT 115.440 201.865 116.485 202.035 ;
        RECT 116.705 201.885 117.035 202.085 ;
        RECT 117.215 202.125 118.365 202.365 ;
        RECT 117.215 201.995 117.885 202.125 ;
        RECT 115.440 200.930 115.610 201.865 ;
        RECT 115.780 201.335 116.145 201.695 ;
        RECT 116.315 201.675 116.485 201.865 ;
        RECT 116.315 201.505 117.435 201.675 ;
        RECT 115.780 201.165 117.065 201.335 ;
        RECT 116.080 200.755 116.675 200.995 ;
        RECT 116.845 200.810 117.065 201.165 ;
        RECT 117.265 201.000 117.435 201.505 ;
        RECT 117.715 201.525 117.885 201.995 ;
        RECT 118.535 201.955 118.705 202.555 ;
        RECT 118.080 201.695 118.705 201.955 ;
        RECT 117.715 201.280 118.365 201.525 ;
        RECT 115.335 200.585 115.890 200.720 ;
        RECT 117.265 200.640 117.435 200.805 ;
        RECT 116.995 200.585 117.435 200.640 ;
        RECT 115.335 200.470 117.435 200.585 ;
        RECT 117.715 200.665 117.885 201.280 ;
        RECT 118.535 201.110 118.705 201.695 ;
        RECT 118.080 200.835 118.705 201.110 ;
        RECT 115.760 200.415 117.125 200.470 ;
        RECT 117.715 200.420 118.365 200.665 ;
        RECT 117.715 200.300 117.885 200.420 ;
        RECT 11.950 199.065 90.610 199.235 ;
        RECT 12.035 198.315 13.245 199.065 ;
        RECT 13.415 198.520 18.760 199.065 ;
        RECT 18.935 198.520 24.280 199.065 ;
        RECT 24.455 198.520 29.800 199.065 ;
        RECT 29.975 198.520 35.320 199.065 ;
        RECT 12.035 197.775 12.555 198.315 ;
        RECT 12.725 197.605 13.245 198.145 ;
        RECT 15.000 197.690 15.340 198.520 ;
        RECT 12.035 196.515 13.245 197.605 ;
        RECT 16.820 196.950 17.170 198.200 ;
        RECT 20.520 197.690 20.860 198.520 ;
        RECT 22.340 196.950 22.690 198.200 ;
        RECT 26.040 197.690 26.380 198.520 ;
        RECT 27.860 196.950 28.210 198.200 ;
        RECT 31.560 197.690 31.900 198.520 ;
        RECT 35.495 198.295 37.165 199.065 ;
        RECT 37.795 198.340 38.085 199.065 ;
        RECT 38.255 198.295 40.845 199.065 ;
        RECT 33.380 196.950 33.730 198.200 ;
        RECT 35.495 197.775 36.245 198.295 ;
        RECT 36.415 197.605 37.165 198.125 ;
        RECT 38.255 197.775 39.465 198.295 ;
        RECT 41.025 198.255 41.295 199.065 ;
        RECT 41.465 198.255 41.795 198.895 ;
        RECT 41.965 198.255 42.205 199.065 ;
        RECT 42.395 198.685 43.285 198.855 ;
        RECT 13.415 196.515 18.760 196.950 ;
        RECT 18.935 196.515 24.280 196.950 ;
        RECT 24.455 196.515 29.800 196.950 ;
        RECT 29.975 196.515 35.320 196.950 ;
        RECT 35.495 196.515 37.165 197.605 ;
        RECT 37.795 196.515 38.085 197.680 ;
        RECT 39.635 197.605 40.845 198.125 ;
        RECT 41.015 197.825 41.365 198.075 ;
        RECT 41.535 197.655 41.705 198.255 ;
        RECT 42.395 198.130 42.945 198.515 ;
        RECT 41.875 197.825 42.225 198.075 ;
        RECT 43.115 197.960 43.285 198.685 ;
        RECT 42.395 197.890 43.285 197.960 ;
        RECT 43.455 198.360 43.675 198.845 ;
        RECT 43.845 198.525 44.095 199.065 ;
        RECT 44.265 198.415 44.525 198.895 ;
        RECT 43.455 197.935 43.785 198.360 ;
        RECT 42.395 197.865 43.290 197.890 ;
        RECT 42.395 197.850 43.300 197.865 ;
        RECT 42.395 197.835 43.305 197.850 ;
        RECT 42.395 197.830 43.315 197.835 ;
        RECT 42.395 197.820 43.320 197.830 ;
        RECT 42.395 197.810 43.325 197.820 ;
        RECT 42.395 197.805 43.335 197.810 ;
        RECT 42.395 197.795 43.345 197.805 ;
        RECT 42.395 197.790 43.355 197.795 ;
        RECT 38.255 196.515 40.845 197.605 ;
        RECT 41.025 196.515 41.355 197.655 ;
        RECT 41.535 197.485 42.215 197.655 ;
        RECT 41.885 196.700 42.215 197.485 ;
        RECT 42.395 197.340 42.655 197.790 ;
        RECT 43.020 197.785 43.355 197.790 ;
        RECT 43.020 197.780 43.370 197.785 ;
        RECT 43.020 197.770 43.385 197.780 ;
        RECT 43.020 197.765 43.410 197.770 ;
        RECT 43.955 197.765 44.185 198.160 ;
        RECT 43.020 197.760 44.185 197.765 ;
        RECT 43.050 197.725 44.185 197.760 ;
        RECT 43.085 197.700 44.185 197.725 ;
        RECT 43.115 197.670 44.185 197.700 ;
        RECT 43.135 197.640 44.185 197.670 ;
        RECT 43.155 197.610 44.185 197.640 ;
        RECT 43.225 197.600 44.185 197.610 ;
        RECT 43.250 197.590 44.185 197.600 ;
        RECT 43.270 197.575 44.185 197.590 ;
        RECT 43.290 197.560 44.185 197.575 ;
        RECT 43.295 197.550 44.080 197.560 ;
        RECT 43.310 197.515 44.080 197.550 ;
        RECT 42.825 197.195 43.155 197.440 ;
        RECT 43.325 197.265 44.080 197.515 ;
        RECT 44.355 197.385 44.525 198.415 ;
        RECT 44.785 198.515 44.955 198.805 ;
        RECT 45.125 198.685 45.455 199.065 ;
        RECT 44.785 198.345 45.450 198.515 ;
        RECT 44.700 197.525 45.050 198.175 ;
        RECT 42.825 197.170 43.010 197.195 ;
        RECT 42.395 197.070 43.010 197.170 ;
        RECT 42.395 196.515 43.000 197.070 ;
        RECT 43.175 196.685 43.655 197.025 ;
        RECT 43.825 196.515 44.080 197.060 ;
        RECT 44.250 196.685 44.525 197.385 ;
        RECT 45.220 197.355 45.450 198.345 ;
        RECT 44.785 197.185 45.450 197.355 ;
        RECT 44.785 196.685 44.955 197.185 ;
        RECT 45.125 196.515 45.455 197.015 ;
        RECT 45.625 196.685 45.810 198.805 ;
        RECT 46.065 198.605 46.315 199.065 ;
        RECT 46.485 198.615 46.820 198.785 ;
        RECT 47.015 198.615 47.690 198.785 ;
        RECT 46.485 198.475 46.655 198.615 ;
        RECT 45.980 197.485 46.260 198.435 ;
        RECT 46.430 198.345 46.655 198.475 ;
        RECT 46.430 197.240 46.600 198.345 ;
        RECT 46.825 198.195 47.350 198.415 ;
        RECT 46.770 197.430 47.010 198.025 ;
        RECT 47.180 197.495 47.350 198.195 ;
        RECT 47.520 197.835 47.690 198.615 ;
        RECT 48.010 198.565 48.380 199.065 ;
        RECT 48.560 198.615 48.965 198.785 ;
        RECT 49.135 198.615 49.920 198.785 ;
        RECT 48.560 198.385 48.730 198.615 ;
        RECT 47.900 198.085 48.730 198.385 ;
        RECT 49.115 198.115 49.580 198.445 ;
        RECT 47.900 198.055 48.100 198.085 ;
        RECT 48.220 197.835 48.390 197.905 ;
        RECT 47.520 197.665 48.390 197.835 ;
        RECT 47.880 197.575 48.390 197.665 ;
        RECT 46.430 197.110 46.735 197.240 ;
        RECT 47.180 197.130 47.710 197.495 ;
        RECT 46.050 196.515 46.315 196.975 ;
        RECT 46.485 196.685 46.735 197.110 ;
        RECT 47.880 196.960 48.050 197.575 ;
        RECT 46.945 196.790 48.050 196.960 ;
        RECT 48.220 196.515 48.390 197.315 ;
        RECT 48.560 197.015 48.730 198.085 ;
        RECT 48.900 197.185 49.090 197.905 ;
        RECT 49.260 197.155 49.580 198.115 ;
        RECT 49.750 198.155 49.920 198.615 ;
        RECT 50.195 198.535 50.405 199.065 ;
        RECT 50.665 198.325 50.995 198.850 ;
        RECT 51.165 198.455 51.335 199.065 ;
        RECT 51.505 198.410 51.835 198.845 ;
        RECT 51.505 198.325 51.885 198.410 ;
        RECT 50.795 198.155 50.995 198.325 ;
        RECT 51.660 198.285 51.885 198.325 ;
        RECT 49.750 197.825 50.625 198.155 ;
        RECT 50.795 197.825 51.545 198.155 ;
        RECT 48.560 196.685 48.810 197.015 ;
        RECT 49.750 196.985 49.920 197.825 ;
        RECT 50.795 197.620 50.985 197.825 ;
        RECT 51.715 197.705 51.885 198.285 ;
        RECT 52.055 198.295 55.565 199.065 ;
        RECT 55.825 198.515 55.995 198.805 ;
        RECT 56.165 198.685 56.495 199.065 ;
        RECT 55.825 198.345 56.490 198.515 ;
        RECT 52.055 197.775 53.705 198.295 ;
        RECT 51.670 197.655 51.885 197.705 ;
        RECT 50.090 197.245 50.985 197.620 ;
        RECT 51.495 197.575 51.885 197.655 ;
        RECT 53.875 197.605 55.565 198.125 ;
        RECT 49.035 196.815 49.920 196.985 ;
        RECT 50.100 196.515 50.415 197.015 ;
        RECT 50.645 196.685 50.985 197.245 ;
        RECT 51.155 196.515 51.325 197.525 ;
        RECT 51.495 196.730 51.825 197.575 ;
        RECT 52.055 196.515 55.565 197.605 ;
        RECT 55.740 197.525 56.090 198.175 ;
        RECT 56.260 197.355 56.490 198.345 ;
        RECT 55.825 197.185 56.490 197.355 ;
        RECT 55.825 196.685 55.995 197.185 ;
        RECT 56.165 196.515 56.495 197.015 ;
        RECT 56.665 196.685 56.850 198.805 ;
        RECT 57.105 198.605 57.355 199.065 ;
        RECT 57.525 198.615 57.860 198.785 ;
        RECT 58.055 198.615 58.730 198.785 ;
        RECT 57.525 198.475 57.695 198.615 ;
        RECT 57.020 197.485 57.300 198.435 ;
        RECT 57.470 198.345 57.695 198.475 ;
        RECT 57.470 197.240 57.640 198.345 ;
        RECT 57.865 198.195 58.390 198.415 ;
        RECT 57.810 197.430 58.050 198.025 ;
        RECT 58.220 197.495 58.390 198.195 ;
        RECT 58.560 197.835 58.730 198.615 ;
        RECT 59.050 198.565 59.420 199.065 ;
        RECT 59.600 198.615 60.005 198.785 ;
        RECT 60.175 198.615 60.960 198.785 ;
        RECT 59.600 198.385 59.770 198.615 ;
        RECT 58.940 198.085 59.770 198.385 ;
        RECT 60.155 198.115 60.620 198.445 ;
        RECT 58.940 198.055 59.140 198.085 ;
        RECT 59.260 197.835 59.430 197.905 ;
        RECT 58.560 197.665 59.430 197.835 ;
        RECT 58.920 197.575 59.430 197.665 ;
        RECT 57.470 197.110 57.775 197.240 ;
        RECT 58.220 197.130 58.750 197.495 ;
        RECT 57.090 196.515 57.355 196.975 ;
        RECT 57.525 196.685 57.775 197.110 ;
        RECT 58.920 196.960 59.090 197.575 ;
        RECT 57.985 196.790 59.090 196.960 ;
        RECT 59.260 196.515 59.430 197.315 ;
        RECT 59.600 197.015 59.770 198.085 ;
        RECT 59.940 197.185 60.130 197.905 ;
        RECT 60.300 197.155 60.620 198.115 ;
        RECT 60.790 198.155 60.960 198.615 ;
        RECT 61.235 198.535 61.445 199.065 ;
        RECT 61.705 198.325 62.035 198.850 ;
        RECT 62.205 198.455 62.375 199.065 ;
        RECT 62.545 198.410 62.875 198.845 ;
        RECT 62.545 198.325 62.925 198.410 ;
        RECT 63.555 198.340 63.845 199.065 ;
        RECT 61.835 198.155 62.035 198.325 ;
        RECT 62.700 198.285 62.925 198.325 ;
        RECT 60.790 197.825 61.665 198.155 ;
        RECT 61.835 197.825 62.585 198.155 ;
        RECT 59.600 196.685 59.850 197.015 ;
        RECT 60.790 196.985 60.960 197.825 ;
        RECT 61.835 197.620 62.025 197.825 ;
        RECT 62.755 197.705 62.925 198.285 ;
        RECT 64.015 198.295 65.685 199.065 ;
        RECT 66.365 198.410 66.695 198.845 ;
        RECT 66.865 198.455 67.035 199.065 ;
        RECT 66.315 198.325 66.695 198.410 ;
        RECT 67.205 198.325 67.535 198.850 ;
        RECT 67.795 198.535 68.005 199.065 ;
        RECT 68.280 198.615 69.065 198.785 ;
        RECT 69.235 198.615 69.640 198.785 ;
        RECT 64.015 197.775 64.765 198.295 ;
        RECT 66.315 198.285 66.540 198.325 ;
        RECT 62.710 197.655 62.925 197.705 ;
        RECT 61.130 197.245 62.025 197.620 ;
        RECT 62.535 197.575 62.925 197.655 ;
        RECT 60.075 196.815 60.960 196.985 ;
        RECT 61.140 196.515 61.455 197.015 ;
        RECT 61.685 196.685 62.025 197.245 ;
        RECT 62.195 196.515 62.365 197.525 ;
        RECT 62.535 196.730 62.865 197.575 ;
        RECT 63.555 196.515 63.845 197.680 ;
        RECT 64.935 197.605 65.685 198.125 ;
        RECT 64.015 196.515 65.685 197.605 ;
        RECT 66.315 197.705 66.485 198.285 ;
        RECT 67.205 198.155 67.405 198.325 ;
        RECT 68.280 198.155 68.450 198.615 ;
        RECT 66.655 197.825 67.405 198.155 ;
        RECT 67.575 197.825 68.450 198.155 ;
        RECT 66.315 197.655 66.530 197.705 ;
        RECT 66.315 197.575 66.705 197.655 ;
        RECT 66.375 196.730 66.705 197.575 ;
        RECT 67.215 197.620 67.405 197.825 ;
        RECT 66.875 196.515 67.045 197.525 ;
        RECT 67.215 197.245 68.110 197.620 ;
        RECT 67.215 196.685 67.555 197.245 ;
        RECT 67.785 196.515 68.100 197.015 ;
        RECT 68.280 196.985 68.450 197.825 ;
        RECT 68.620 198.115 69.085 198.445 ;
        RECT 69.470 198.385 69.640 198.615 ;
        RECT 69.820 198.565 70.190 199.065 ;
        RECT 70.510 198.615 71.185 198.785 ;
        RECT 71.380 198.615 71.715 198.785 ;
        RECT 68.620 197.155 68.940 198.115 ;
        RECT 69.470 198.085 70.300 198.385 ;
        RECT 69.110 197.185 69.300 197.905 ;
        RECT 69.470 197.015 69.640 198.085 ;
        RECT 70.100 198.055 70.300 198.085 ;
        RECT 69.810 197.835 69.980 197.905 ;
        RECT 70.510 197.835 70.680 198.615 ;
        RECT 71.545 198.475 71.715 198.615 ;
        RECT 71.885 198.605 72.135 199.065 ;
        RECT 69.810 197.665 70.680 197.835 ;
        RECT 70.850 198.195 71.375 198.415 ;
        RECT 71.545 198.345 71.770 198.475 ;
        RECT 69.810 197.575 70.320 197.665 ;
        RECT 68.280 196.815 69.165 196.985 ;
        RECT 69.390 196.685 69.640 197.015 ;
        RECT 69.810 196.515 69.980 197.315 ;
        RECT 70.150 196.960 70.320 197.575 ;
        RECT 70.850 197.495 71.020 198.195 ;
        RECT 70.490 197.130 71.020 197.495 ;
        RECT 71.190 197.430 71.430 198.025 ;
        RECT 71.600 197.240 71.770 198.345 ;
        RECT 71.940 197.485 72.220 198.435 ;
        RECT 71.465 197.110 71.770 197.240 ;
        RECT 70.150 196.790 71.255 196.960 ;
        RECT 71.465 196.685 71.715 197.110 ;
        RECT 71.885 196.515 72.150 196.975 ;
        RECT 72.390 196.685 72.575 198.805 ;
        RECT 72.745 198.685 73.075 199.065 ;
        RECT 73.245 198.515 73.415 198.805 ;
        RECT 73.675 198.520 79.020 199.065 ;
        RECT 79.195 198.520 84.540 199.065 ;
        RECT 72.750 198.345 73.415 198.515 ;
        RECT 72.750 197.355 72.980 198.345 ;
        RECT 73.150 197.525 73.500 198.175 ;
        RECT 75.260 197.690 75.600 198.520 ;
        RECT 72.750 197.185 73.415 197.355 ;
        RECT 72.745 196.515 73.075 197.015 ;
        RECT 73.245 196.685 73.415 197.185 ;
        RECT 77.080 196.950 77.430 198.200 ;
        RECT 80.780 197.690 81.120 198.520 ;
        RECT 84.715 198.295 88.225 199.065 ;
        RECT 89.315 198.315 90.525 199.065 ;
        RECT 82.600 196.950 82.950 198.200 ;
        RECT 84.715 197.775 86.365 198.295 ;
        RECT 86.535 197.605 88.225 198.125 ;
        RECT 73.675 196.515 79.020 196.950 ;
        RECT 79.195 196.515 84.540 196.950 ;
        RECT 84.715 196.515 88.225 197.605 ;
        RECT 89.315 197.605 89.835 198.145 ;
        RECT 90.005 197.775 90.525 198.315 ;
        RECT 112.275 198.070 112.445 199.885 ;
        RECT 113.125 199.705 113.425 200.165 ;
        RECT 113.675 200.045 113.935 200.215 ;
        RECT 114.995 200.045 115.625 200.300 ;
        RECT 113.605 199.875 113.935 200.045 ;
        RECT 114.195 200.035 115.625 200.045 ;
        RECT 114.195 199.875 115.165 200.035 ;
        RECT 116.135 199.965 117.085 200.245 ;
        RECT 117.255 200.050 117.885 200.300 ;
        RECT 118.535 200.250 118.705 200.835 ;
        RECT 112.725 199.535 114.825 199.705 ;
        RECT 112.725 199.300 112.895 199.535 ;
        RECT 114.495 199.455 114.825 199.535 ;
        RECT 114.995 199.440 115.165 199.875 ;
        RECT 117.715 199.810 117.885 200.050 ;
        RECT 118.080 199.990 118.705 200.250 ;
        RECT 115.335 199.610 117.455 199.795 ;
        RECT 117.715 199.560 118.365 199.810 ;
        RECT 117.715 199.440 117.885 199.560 ;
        RECT 113.605 199.175 114.325 199.365 ;
        RECT 112.725 198.515 112.895 199.130 ;
        RECT 113.065 199.005 113.395 199.150 ;
        RECT 113.065 198.685 114.355 199.005 ;
        RECT 114.525 198.515 114.695 199.230 ;
        RECT 112.725 198.345 114.695 198.515 ;
        RECT 114.995 199.110 115.665 199.440 ;
        RECT 115.835 199.205 117.165 199.435 ;
        RECT 112.275 197.860 112.975 198.070 ;
        RECT 89.315 196.515 90.525 197.605 ;
        RECT 112.275 197.100 112.445 197.860 ;
        RECT 113.355 197.640 113.685 198.345 ;
        RECT 113.890 197.620 114.265 198.175 ;
        RECT 114.995 198.165 115.165 199.110 ;
        RECT 115.835 198.940 116.005 199.205 ;
        RECT 115.335 198.770 116.005 198.940 ;
        RECT 116.175 198.685 116.825 199.035 ;
        RECT 116.995 198.940 117.165 199.205 ;
        RECT 117.335 199.110 117.885 199.440 ;
        RECT 118.535 199.390 118.705 199.990 ;
        RECT 118.080 199.130 118.705 199.390 ;
        RECT 117.715 198.950 117.885 199.110 ;
        RECT 116.995 198.770 117.455 198.940 ;
        RECT 117.715 198.700 118.365 198.950 ;
        RECT 115.335 198.335 117.545 198.505 ;
        RECT 115.335 198.170 116.305 198.335 ;
        RECT 116.975 198.250 117.545 198.335 ;
        RECT 114.495 198.000 115.165 198.165 ;
        RECT 116.475 198.080 116.805 198.165 ;
        RECT 117.715 198.090 117.885 198.700 ;
        RECT 118.535 198.530 118.705 199.130 ;
        RECT 118.080 198.270 118.705 198.530 ;
        RECT 118.535 198.095 118.705 198.270 ;
        RECT 118.875 198.265 119.125 204.275 ;
        RECT 120.435 204.105 120.605 204.705 ;
        RECT 119.635 203.845 120.605 204.105 ;
        RECT 119.295 203.415 120.260 203.675 ;
        RECT 120.430 203.500 120.605 203.845 ;
        RECT 120.775 205.530 121.800 205.700 ;
        RECT 122.175 206.270 122.950 206.450 ;
        RECT 123.155 206.330 123.325 206.960 ;
        RECT 125.875 206.330 126.045 206.960 ;
        RECT 122.175 205.560 122.345 206.270 ;
        RECT 123.155 206.050 124.050 206.330 ;
        RECT 122.620 206.040 124.050 206.050 ;
        RECT 124.710 206.040 126.045 206.330 ;
        RECT 126.345 206.335 126.515 207.050 ;
        RECT 126.715 206.995 127.435 207.185 ;
        RECT 128.145 207.120 128.315 207.355 ;
        RECT 127.645 206.825 127.975 206.970 ;
        RECT 126.685 206.505 127.975 206.825 ;
        RECT 128.145 206.335 128.315 206.950 ;
        RECT 126.345 206.165 128.315 206.335 ;
        RECT 128.595 206.500 129.535 207.705 ;
        RECT 129.705 207.240 131.485 207.710 ;
        RECT 134.035 207.250 134.205 207.880 ;
        RECT 135.115 207.760 135.445 208.465 ;
        RECT 136.755 208.365 137.655 208.610 ;
        RECT 135.650 207.740 136.025 208.295 ;
        RECT 136.755 208.285 136.930 208.365 ;
        RECT 136.255 207.970 136.930 208.285 ;
        RECT 137.825 208.180 138.065 208.780 ;
        RECT 136.755 207.750 136.930 207.970 ;
        RECT 137.100 207.920 138.065 208.180 ;
        RECT 134.420 207.590 134.945 207.720 ;
        RECT 135.650 207.590 136.585 207.740 ;
        RECT 134.420 207.400 136.585 207.590 ;
        RECT 136.755 207.505 137.655 207.750 ;
        RECT 134.420 207.390 135.445 207.400 ;
        RECT 129.705 206.945 132.295 207.240 ;
        RECT 129.705 206.500 131.485 206.945 ;
        RECT 132.795 206.935 133.355 207.250 ;
        RECT 133.525 207.220 134.205 207.250 ;
        RECT 133.525 207.050 134.815 207.220 ;
        RECT 133.525 206.945 134.205 207.050 ;
        RECT 131.655 206.520 133.855 206.765 ;
        RECT 128.595 206.330 128.765 206.500 ;
        RECT 131.315 206.345 131.485 206.500 ;
        RECT 132.795 206.515 133.855 206.520 ;
        RECT 131.315 206.330 132.295 206.345 ;
        RECT 122.620 205.540 123.325 206.040 ;
        RECT 125.875 205.985 126.045 206.040 ;
        RECT 123.585 205.610 124.045 205.780 ;
        RECT 120.775 203.840 120.945 205.530 ;
        RECT 123.155 205.440 123.325 205.540 ;
        RECT 121.455 205.170 122.985 205.360 ;
        RECT 121.115 204.180 121.285 205.135 ;
        RECT 121.455 204.520 121.625 205.170 ;
        RECT 123.155 205.110 123.705 205.440 ;
        RECT 123.875 205.345 124.045 205.610 ;
        RECT 124.215 205.515 124.865 205.865 ;
        RECT 125.035 205.610 125.705 205.780 ;
        RECT 125.875 205.670 126.545 205.985 ;
        RECT 125.035 205.345 125.205 205.610 ;
        RECT 125.875 205.440 126.045 205.670 ;
        RECT 126.775 205.440 127.150 205.995 ;
        RECT 127.355 205.460 127.685 206.165 ;
        RECT 128.595 206.040 129.490 206.330 ;
        RECT 130.150 206.085 132.295 206.330 ;
        RECT 130.150 206.040 131.485 206.085 ;
        RECT 128.595 205.890 128.765 206.040 ;
        RECT 128.065 205.860 128.765 205.890 ;
        RECT 128.065 205.680 129.575 205.860 ;
        RECT 128.595 205.590 129.575 205.680 ;
        RECT 123.875 205.115 125.205 205.345 ;
        RECT 125.375 205.110 126.045 205.440 ;
        RECT 121.825 204.725 122.985 205.000 ;
        RECT 121.965 204.720 122.135 204.725 ;
        RECT 121.455 204.350 122.425 204.520 ;
        RECT 122.620 204.180 122.985 204.535 ;
        RECT 121.115 204.010 122.985 204.180 ;
        RECT 122.415 204.005 122.985 204.010 ;
        RECT 123.155 204.500 123.325 205.110 ;
        RECT 123.585 204.755 125.705 204.940 ;
        RECT 125.875 204.930 126.045 205.110 ;
        RECT 126.215 205.290 127.150 205.440 ;
        RECT 127.855 205.290 128.380 205.420 ;
        RECT 126.215 205.100 128.380 205.290 ;
        RECT 127.355 205.090 128.380 205.100 ;
        RECT 125.875 204.760 127.055 204.930 ;
        RECT 123.155 204.250 123.785 204.500 ;
        RECT 123.955 204.305 124.905 204.585 ;
        RECT 125.875 204.515 126.045 204.760 ;
        RECT 125.415 204.250 126.045 204.515 ;
        RECT 126.260 204.415 127.185 204.590 ;
        RECT 127.355 204.540 127.685 205.090 ;
        RECT 128.595 204.920 128.765 205.590 ;
        RECT 129.755 205.520 130.005 205.870 ;
        RECT 131.315 205.860 131.485 206.040 ;
        RECT 132.795 205.905 133.045 206.515 ;
        RECT 134.035 206.345 134.205 206.945 ;
        RECT 134.425 206.725 134.945 206.880 ;
        RECT 135.115 206.840 135.445 207.390 ;
        RECT 136.755 207.230 136.930 207.505 ;
        RECT 137.825 207.320 138.065 207.920 ;
        RECT 135.745 207.060 136.930 207.230 ;
        RECT 137.100 207.060 138.065 207.320 ;
        RECT 136.755 206.890 136.930 207.060 ;
        RECT 134.425 206.670 134.985 206.725 ;
        RECT 135.615 206.715 136.540 206.890 ;
        RECT 135.565 206.670 136.540 206.715 ;
        RECT 134.425 206.560 136.540 206.670 ;
        RECT 136.755 206.645 137.655 206.890 ;
        RECT 134.425 206.550 135.695 206.560 ;
        RECT 134.860 206.500 135.695 206.550 ;
        RECT 133.510 206.330 134.205 206.345 ;
        RECT 136.755 206.330 136.930 206.645 ;
        RECT 137.825 206.475 138.065 207.060 ;
        RECT 133.510 206.085 134.930 206.330 ;
        RECT 134.035 206.040 134.930 206.085 ;
        RECT 135.590 206.045 136.930 206.330 ;
        RECT 137.100 206.215 138.065 206.475 ;
        RECT 135.590 206.040 137.655 206.045 ;
        RECT 130.175 205.530 131.485 205.860 ;
        RECT 131.660 205.655 133.855 205.905 ;
        RECT 131.315 205.485 131.485 205.530 ;
        RECT 128.935 205.350 129.575 205.420 ;
        RECT 128.935 205.180 130.345 205.350 ;
        RECT 128.935 205.090 129.575 205.180 ;
        RECT 127.985 204.750 129.575 204.920 ;
        RECT 128.595 204.680 129.575 204.750 ;
        RECT 127.855 204.425 128.375 204.580 ;
        RECT 126.260 204.370 127.235 204.415 ;
        RECT 127.815 204.370 128.375 204.425 ;
        RECT 126.260 204.260 128.375 204.370 ;
        RECT 120.775 203.670 122.245 203.840 ;
        RECT 121.915 203.645 122.245 203.670 ;
        RECT 119.295 202.815 119.535 203.415 ;
        RECT 120.430 203.330 121.745 203.500 ;
        RECT 122.415 203.420 122.585 204.005 ;
        RECT 123.155 203.580 123.325 204.250 ;
        RECT 123.915 204.080 125.280 204.135 ;
        RECT 123.605 203.965 125.705 204.080 ;
        RECT 123.605 203.910 124.045 203.965 ;
        RECT 123.605 203.745 123.775 203.910 ;
        RECT 125.150 203.830 125.705 203.965 ;
        RECT 120.430 203.245 120.605 203.330 ;
        RECT 119.705 202.985 120.605 203.245 ;
        RECT 121.915 203.250 122.585 203.420 ;
        RECT 122.755 203.250 123.325 203.580 ;
        RECT 121.915 203.165 122.245 203.250 ;
        RECT 119.295 202.555 120.260 202.815 ;
        RECT 120.430 202.650 120.605 202.985 ;
        RECT 120.775 202.995 121.745 203.160 ;
        RECT 122.415 202.995 122.985 203.080 ;
        RECT 120.775 202.825 122.985 202.995 ;
        RECT 123.155 202.650 123.325 203.250 ;
        RECT 123.605 203.045 123.775 203.550 ;
        RECT 123.975 203.385 124.195 203.740 ;
        RECT 124.365 203.555 124.960 203.795 ;
        RECT 123.975 203.215 125.260 203.385 ;
        RECT 123.605 202.875 124.725 203.045 ;
        RECT 124.555 202.685 124.725 202.875 ;
        RECT 124.895 202.855 125.260 203.215 ;
        RECT 125.430 202.685 125.600 203.620 ;
        RECT 119.295 201.955 119.535 202.555 ;
        RECT 120.430 202.385 121.695 202.650 ;
        RECT 119.705 202.125 121.695 202.385 ;
        RECT 119.295 201.695 120.260 201.955 ;
        RECT 120.430 201.730 121.695 202.125 ;
        RECT 121.865 202.555 123.325 202.650 ;
        RECT 121.865 202.185 123.825 202.555 ;
        RECT 124.005 202.465 124.335 202.665 ;
        RECT 124.555 202.515 125.600 202.685 ;
        RECT 125.875 203.520 126.045 204.250 ;
        RECT 127.105 204.250 128.375 204.260 ;
        RECT 127.105 204.200 127.940 204.250 ;
        RECT 126.215 203.855 128.425 204.025 ;
        RECT 126.215 203.690 127.185 203.855 ;
        RECT 127.855 203.770 128.425 203.855 ;
        RECT 128.595 203.890 128.765 204.680 ;
        RECT 129.755 204.660 130.005 205.010 ;
        RECT 130.175 205.000 130.345 205.180 ;
        RECT 131.315 205.225 132.285 205.485 ;
        RECT 130.175 204.670 131.130 205.000 ;
        RECT 131.315 204.625 131.490 205.225 ;
        RECT 131.660 204.795 132.625 205.055 ;
        RECT 128.935 204.060 129.585 204.390 ;
        RECT 127.355 203.600 127.685 203.685 ;
        RECT 128.595 203.600 129.225 203.890 ;
        RECT 125.875 203.350 127.185 203.520 ;
        RECT 127.355 203.430 128.025 203.600 ;
        RECT 121.865 201.900 123.325 202.185 ;
        RECT 124.005 202.005 124.305 202.465 ;
        RECT 124.555 202.345 124.815 202.515 ;
        RECT 125.875 202.345 126.045 203.350 ;
        RECT 127.355 203.180 127.685 203.205 ;
        RECT 124.485 202.175 124.815 202.345 ;
        RECT 125.075 202.175 126.045 202.345 ;
        RECT 119.295 201.095 119.535 201.695 ;
        RECT 120.430 201.525 122.215 201.730 ;
        RECT 119.705 201.265 122.215 201.525 ;
        RECT 119.295 200.835 120.260 201.095 ;
        RECT 120.430 200.980 122.215 201.265 ;
        RECT 122.385 200.980 123.325 201.900 ;
        RECT 123.605 201.835 125.705 202.005 ;
        RECT 123.605 201.600 123.775 201.835 ;
        RECT 125.375 201.755 125.705 201.835 ;
        RECT 124.485 201.475 125.205 201.665 ;
        RECT 119.295 200.250 119.535 200.835 ;
        RECT 120.430 200.665 120.605 200.980 ;
        RECT 119.705 200.420 120.605 200.665 ;
        RECT 120.775 200.550 121.445 200.720 ;
        RECT 120.430 200.380 120.605 200.420 ;
        RECT 119.295 199.990 120.260 200.250 ;
        RECT 120.430 200.050 121.105 200.380 ;
        RECT 121.275 200.285 121.445 200.550 ;
        RECT 121.615 200.455 122.265 200.805 ;
        RECT 122.435 200.550 122.895 200.720 ;
        RECT 122.435 200.285 122.605 200.550 ;
        RECT 123.155 200.380 123.325 200.980 ;
        RECT 123.605 200.815 123.775 201.430 ;
        RECT 123.945 201.305 124.275 201.450 ;
        RECT 123.945 200.985 125.235 201.305 ;
        RECT 125.405 200.815 125.575 201.530 ;
        RECT 123.605 200.645 125.575 200.815 ;
        RECT 125.875 200.980 126.045 202.175 ;
        RECT 126.215 203.010 127.685 203.180 ;
        RECT 126.215 201.320 126.385 203.010 ;
        RECT 127.855 202.845 128.025 203.430 ;
        RECT 128.195 203.560 129.225 203.600 ;
        RECT 128.195 203.270 128.765 203.560 ;
        RECT 129.415 203.345 129.585 204.060 ;
        RECT 129.755 203.920 130.005 204.430 ;
        RECT 131.315 204.370 132.215 204.625 ;
        RECT 130.195 204.365 132.215 204.370 ;
        RECT 130.195 204.040 131.490 204.365 ;
        RECT 132.385 204.195 132.625 204.795 ;
        RECT 131.315 203.765 131.490 204.040 ;
        RECT 131.660 203.935 132.625 204.195 ;
        RECT 127.855 202.840 128.425 202.845 ;
        RECT 126.555 202.670 128.425 202.840 ;
        RECT 126.555 201.715 126.725 202.670 ;
        RECT 126.895 202.330 127.865 202.500 ;
        RECT 126.895 201.680 127.065 202.330 ;
        RECT 128.060 202.315 128.425 202.670 ;
        RECT 128.595 202.815 128.765 203.270 ;
        RECT 128.935 203.015 129.585 203.345 ;
        RECT 129.755 203.340 131.070 203.710 ;
        RECT 131.315 203.505 132.215 203.765 ;
        RECT 128.595 202.485 129.225 202.815 ;
        RECT 127.405 202.125 127.575 202.130 ;
        RECT 127.265 201.850 128.425 202.125 ;
        RECT 126.895 201.490 128.425 201.680 ;
        RECT 128.595 201.320 128.765 202.485 ;
        RECT 129.415 202.260 129.585 203.015 ;
        RECT 129.755 202.840 131.070 203.170 ;
        RECT 131.315 202.905 131.490 203.505 ;
        RECT 132.385 203.335 132.625 203.935 ;
        RECT 131.660 203.075 132.625 203.335 ;
        RECT 131.315 202.645 132.215 202.905 ;
        RECT 129.755 202.300 131.070 202.630 ;
        RECT 129.095 202.090 129.585 202.260 ;
        RECT 128.950 201.590 129.585 201.920 ;
        RECT 129.755 201.710 129.965 202.130 ;
        RECT 131.315 202.045 131.490 202.645 ;
        RECT 132.385 202.475 132.625 203.075 ;
        RECT 131.660 202.215 132.625 202.475 ;
        RECT 130.135 201.780 131.145 202.030 ;
        RECT 131.315 201.800 132.215 202.045 ;
        RECT 129.395 201.540 129.585 201.590 ;
        RECT 130.135 201.540 130.425 201.780 ;
        RECT 131.315 201.610 131.490 201.800 ;
        RECT 132.385 201.630 132.625 202.215 ;
        RECT 126.215 201.150 127.240 201.320 ;
        RECT 128.595 201.310 129.225 201.320 ;
        RECT 125.875 200.810 126.805 200.980 ;
        RECT 121.275 200.055 122.605 200.285 ;
        RECT 122.775 200.370 123.325 200.380 ;
        RECT 122.775 200.160 123.855 200.370 ;
        RECT 122.775 200.050 123.325 200.160 ;
        RECT 119.295 199.390 119.535 199.990 ;
        RECT 120.430 199.805 120.605 200.050 ;
        RECT 119.705 199.560 120.605 199.805 ;
        RECT 120.775 199.695 122.895 199.880 ;
        RECT 120.430 199.455 120.605 199.560 ;
        RECT 119.295 199.130 120.260 199.390 ;
        RECT 120.430 199.190 121.065 199.455 ;
        RECT 121.575 199.245 122.525 199.525 ;
        RECT 123.155 199.440 123.325 200.050 ;
        RECT 124.235 199.940 124.565 200.645 ;
        RECT 124.770 199.920 125.145 200.475 ;
        RECT 125.875 200.465 126.045 200.810 ;
        RECT 125.375 200.150 126.045 200.465 ;
        RECT 123.540 199.770 124.065 199.900 ;
        RECT 124.770 199.770 125.705 199.920 ;
        RECT 123.540 199.580 125.705 199.770 ;
        RECT 123.540 199.570 124.565 199.580 ;
        RECT 122.695 199.400 123.325 199.440 ;
        RECT 122.695 199.230 123.935 199.400 ;
        RECT 122.695 199.190 123.325 199.230 ;
        RECT 119.295 198.530 119.535 199.130 ;
        RECT 120.430 198.945 120.605 199.190 ;
        RECT 121.200 199.020 122.565 199.075 ;
        RECT 119.705 198.700 120.605 198.945 ;
        RECT 120.775 198.905 122.875 199.020 ;
        RECT 120.775 198.770 121.330 198.905 ;
        RECT 122.435 198.850 122.875 198.905 ;
        RECT 119.295 198.270 120.260 198.530 ;
        RECT 119.295 198.095 119.520 198.270 ;
        RECT 117.715 198.080 118.365 198.090 ;
        RECT 114.495 197.850 116.305 198.000 ;
        RECT 116.475 197.910 117.145 198.080 ;
        RECT 114.995 197.830 116.305 197.850 ;
        RECT 112.660 197.470 113.185 197.600 ;
        RECT 113.890 197.470 114.825 197.620 ;
        RECT 112.660 197.280 114.825 197.470 ;
        RECT 112.660 197.270 113.685 197.280 ;
        RECT 112.275 196.930 113.055 197.100 ;
        RECT 11.950 196.345 90.610 196.515 ;
        RECT 12.035 195.255 13.245 196.345 ;
        RECT 13.415 195.910 18.760 196.345 ;
        RECT 18.935 195.910 24.280 196.345 ;
        RECT 12.035 194.545 12.555 195.085 ;
        RECT 12.725 194.715 13.245 195.255 ;
        RECT 12.035 193.795 13.245 194.545 ;
        RECT 15.000 194.340 15.340 195.170 ;
        RECT 16.820 194.660 17.170 195.910 ;
        RECT 20.520 194.340 20.860 195.170 ;
        RECT 22.340 194.660 22.690 195.910 ;
        RECT 24.915 195.180 25.205 196.345 ;
        RECT 25.375 195.910 30.720 196.345 ;
        RECT 30.895 195.910 36.240 196.345 ;
        RECT 13.415 193.795 18.760 194.340 ;
        RECT 18.935 193.795 24.280 194.340 ;
        RECT 24.915 193.795 25.205 194.520 ;
        RECT 26.960 194.340 27.300 195.170 ;
        RECT 28.780 194.660 29.130 195.910 ;
        RECT 32.480 194.340 32.820 195.170 ;
        RECT 34.300 194.660 34.650 195.910 ;
        RECT 36.965 195.675 37.135 196.175 ;
        RECT 37.305 195.845 37.635 196.345 ;
        RECT 36.965 195.505 37.630 195.675 ;
        RECT 36.880 194.685 37.230 195.335 ;
        RECT 37.400 194.515 37.630 195.505 ;
        RECT 36.965 194.345 37.630 194.515 ;
        RECT 25.375 193.795 30.720 194.340 ;
        RECT 30.895 193.795 36.240 194.340 ;
        RECT 36.965 194.055 37.135 194.345 ;
        RECT 37.305 193.795 37.635 194.175 ;
        RECT 37.805 194.055 37.990 196.175 ;
        RECT 38.230 195.885 38.495 196.345 ;
        RECT 38.665 195.750 38.915 196.175 ;
        RECT 39.125 195.900 40.230 196.070 ;
        RECT 38.610 195.620 38.915 195.750 ;
        RECT 38.160 194.425 38.440 195.375 ;
        RECT 38.610 194.515 38.780 195.620 ;
        RECT 38.950 194.835 39.190 195.430 ;
        RECT 39.360 195.365 39.890 195.730 ;
        RECT 39.360 194.665 39.530 195.365 ;
        RECT 40.060 195.285 40.230 195.900 ;
        RECT 40.400 195.545 40.570 196.345 ;
        RECT 40.740 195.845 40.990 196.175 ;
        RECT 41.215 195.875 42.100 196.045 ;
        RECT 40.060 195.195 40.570 195.285 ;
        RECT 38.610 194.385 38.835 194.515 ;
        RECT 39.005 194.445 39.530 194.665 ;
        RECT 39.700 195.025 40.570 195.195 ;
        RECT 38.245 193.795 38.495 194.255 ;
        RECT 38.665 194.245 38.835 194.385 ;
        RECT 39.700 194.245 39.870 195.025 ;
        RECT 40.400 194.955 40.570 195.025 ;
        RECT 40.080 194.775 40.280 194.805 ;
        RECT 40.740 194.775 40.910 195.845 ;
        RECT 41.080 194.955 41.270 195.675 ;
        RECT 40.080 194.475 40.910 194.775 ;
        RECT 41.440 194.745 41.760 195.705 ;
        RECT 38.665 194.075 39.000 194.245 ;
        RECT 39.195 194.075 39.870 194.245 ;
        RECT 40.190 193.795 40.560 194.295 ;
        RECT 40.740 194.245 40.910 194.475 ;
        RECT 41.295 194.415 41.760 194.745 ;
        RECT 41.930 195.035 42.100 195.875 ;
        RECT 42.280 195.845 42.595 196.345 ;
        RECT 42.825 195.615 43.165 196.175 ;
        RECT 42.270 195.240 43.165 195.615 ;
        RECT 43.335 195.335 43.505 196.345 ;
        RECT 42.975 195.035 43.165 195.240 ;
        RECT 43.675 195.285 44.005 196.130 ;
        RECT 44.695 195.475 44.970 196.175 ;
        RECT 45.140 195.800 45.395 196.345 ;
        RECT 45.565 195.835 46.045 196.175 ;
        RECT 46.220 195.790 46.825 196.345 ;
        RECT 46.210 195.690 46.825 195.790 ;
        RECT 46.210 195.665 46.395 195.690 ;
        RECT 43.675 195.205 44.065 195.285 ;
        RECT 43.850 195.155 44.065 195.205 ;
        RECT 41.930 194.705 42.805 195.035 ;
        RECT 42.975 194.705 43.725 195.035 ;
        RECT 41.930 194.245 42.100 194.705 ;
        RECT 42.975 194.535 43.175 194.705 ;
        RECT 43.895 194.575 44.065 195.155 ;
        RECT 43.840 194.535 44.065 194.575 ;
        RECT 40.740 194.075 41.145 194.245 ;
        RECT 41.315 194.075 42.100 194.245 ;
        RECT 42.375 193.795 42.585 194.325 ;
        RECT 42.845 194.010 43.175 194.535 ;
        RECT 43.685 194.450 44.065 194.535 ;
        RECT 43.345 193.795 43.515 194.405 ;
        RECT 43.685 194.015 44.015 194.450 ;
        RECT 44.695 194.445 44.865 195.475 ;
        RECT 45.140 195.345 45.895 195.595 ;
        RECT 46.065 195.420 46.395 195.665 ;
        RECT 45.140 195.310 45.910 195.345 ;
        RECT 45.140 195.300 45.925 195.310 ;
        RECT 45.035 195.285 45.930 195.300 ;
        RECT 45.035 195.270 45.950 195.285 ;
        RECT 45.035 195.260 45.970 195.270 ;
        RECT 45.035 195.250 45.995 195.260 ;
        RECT 45.035 195.220 46.065 195.250 ;
        RECT 45.035 195.190 46.085 195.220 ;
        RECT 45.035 195.160 46.105 195.190 ;
        RECT 45.035 195.135 46.135 195.160 ;
        RECT 45.035 195.100 46.170 195.135 ;
        RECT 45.035 195.095 46.200 195.100 ;
        RECT 45.035 194.700 45.265 195.095 ;
        RECT 45.810 195.090 46.200 195.095 ;
        RECT 45.835 195.080 46.200 195.090 ;
        RECT 45.850 195.075 46.200 195.080 ;
        RECT 45.865 195.070 46.200 195.075 ;
        RECT 46.565 195.070 46.825 195.520 ;
        RECT 47.005 195.375 47.335 196.160 ;
        RECT 47.005 195.205 47.685 195.375 ;
        RECT 47.865 195.205 48.195 196.345 ;
        RECT 48.375 195.790 48.980 196.345 ;
        RECT 49.155 195.835 49.635 196.175 ;
        RECT 49.805 195.800 50.060 196.345 ;
        RECT 48.375 195.690 48.990 195.790 ;
        RECT 48.805 195.665 48.990 195.690 ;
        RECT 45.865 195.065 46.825 195.070 ;
        RECT 45.875 195.055 46.825 195.065 ;
        RECT 45.885 195.050 46.825 195.055 ;
        RECT 45.895 195.040 46.825 195.050 ;
        RECT 45.900 195.030 46.825 195.040 ;
        RECT 45.905 195.025 46.825 195.030 ;
        RECT 45.915 195.010 46.825 195.025 ;
        RECT 45.920 194.995 46.825 195.010 ;
        RECT 45.930 194.970 46.825 194.995 ;
        RECT 45.435 194.500 45.765 194.925 ;
        RECT 44.695 193.965 44.955 194.445 ;
        RECT 45.125 193.795 45.375 194.335 ;
        RECT 45.545 194.015 45.765 194.500 ;
        RECT 45.935 194.900 46.825 194.970 ;
        RECT 45.935 194.175 46.105 194.900 ;
        RECT 46.995 194.785 47.345 195.035 ;
        RECT 46.275 194.345 46.825 194.730 ;
        RECT 47.515 194.605 47.685 195.205 ;
        RECT 48.375 195.070 48.635 195.520 ;
        RECT 48.805 195.420 49.135 195.665 ;
        RECT 49.305 195.345 50.060 195.595 ;
        RECT 50.230 195.475 50.505 196.175 ;
        RECT 49.290 195.310 50.060 195.345 ;
        RECT 49.275 195.300 50.060 195.310 ;
        RECT 49.270 195.285 50.165 195.300 ;
        RECT 49.250 195.270 50.165 195.285 ;
        RECT 49.230 195.260 50.165 195.270 ;
        RECT 49.205 195.250 50.165 195.260 ;
        RECT 49.135 195.220 50.165 195.250 ;
        RECT 49.115 195.190 50.165 195.220 ;
        RECT 49.095 195.160 50.165 195.190 ;
        RECT 49.065 195.135 50.165 195.160 ;
        RECT 49.030 195.100 50.165 195.135 ;
        RECT 49.000 195.095 50.165 195.100 ;
        RECT 49.000 195.090 49.390 195.095 ;
        RECT 49.000 195.080 49.365 195.090 ;
        RECT 49.000 195.075 49.350 195.080 ;
        RECT 49.000 195.070 49.335 195.075 ;
        RECT 48.375 195.065 49.335 195.070 ;
        RECT 48.375 195.055 49.325 195.065 ;
        RECT 48.375 195.050 49.315 195.055 ;
        RECT 48.375 195.040 49.305 195.050 ;
        RECT 47.855 194.785 48.205 195.035 ;
        RECT 48.375 195.030 49.300 195.040 ;
        RECT 48.375 195.025 49.295 195.030 ;
        RECT 48.375 195.010 49.285 195.025 ;
        RECT 48.375 194.995 49.280 195.010 ;
        RECT 48.375 194.970 49.270 194.995 ;
        RECT 48.375 194.900 49.265 194.970 ;
        RECT 45.935 194.005 46.825 194.175 ;
        RECT 47.015 193.795 47.255 194.605 ;
        RECT 47.425 193.965 47.755 194.605 ;
        RECT 47.925 193.795 48.195 194.605 ;
        RECT 48.375 194.345 48.925 194.730 ;
        RECT 49.095 194.175 49.265 194.900 ;
        RECT 48.375 194.005 49.265 194.175 ;
        RECT 49.435 194.500 49.765 194.925 ;
        RECT 49.935 194.700 50.165 195.095 ;
        RECT 49.435 194.015 49.655 194.500 ;
        RECT 50.335 194.445 50.505 195.475 ;
        RECT 50.675 195.180 50.965 196.345 ;
        RECT 51.225 195.675 51.395 196.175 ;
        RECT 51.565 195.845 51.895 196.345 ;
        RECT 51.225 195.505 51.890 195.675 ;
        RECT 51.140 194.685 51.490 195.335 ;
        RECT 49.825 193.795 50.075 194.335 ;
        RECT 50.245 193.965 50.505 194.445 ;
        RECT 50.675 193.795 50.965 194.520 ;
        RECT 51.660 194.515 51.890 195.505 ;
        RECT 51.225 194.345 51.890 194.515 ;
        RECT 51.225 194.055 51.395 194.345 ;
        RECT 51.565 193.795 51.895 194.175 ;
        RECT 52.065 194.055 52.250 196.175 ;
        RECT 52.490 195.885 52.755 196.345 ;
        RECT 52.925 195.750 53.175 196.175 ;
        RECT 53.385 195.900 54.490 196.070 ;
        RECT 52.870 195.620 53.175 195.750 ;
        RECT 52.420 194.425 52.700 195.375 ;
        RECT 52.870 194.515 53.040 195.620 ;
        RECT 53.210 194.835 53.450 195.430 ;
        RECT 53.620 195.365 54.150 195.730 ;
        RECT 53.620 194.665 53.790 195.365 ;
        RECT 54.320 195.285 54.490 195.900 ;
        RECT 54.660 195.545 54.830 196.345 ;
        RECT 55.000 195.845 55.250 196.175 ;
        RECT 55.475 195.875 56.360 196.045 ;
        RECT 54.320 195.195 54.830 195.285 ;
        RECT 52.870 194.385 53.095 194.515 ;
        RECT 53.265 194.445 53.790 194.665 ;
        RECT 53.960 195.025 54.830 195.195 ;
        RECT 52.505 193.795 52.755 194.255 ;
        RECT 52.925 194.245 53.095 194.385 ;
        RECT 53.960 194.245 54.130 195.025 ;
        RECT 54.660 194.955 54.830 195.025 ;
        RECT 54.340 194.775 54.540 194.805 ;
        RECT 55.000 194.775 55.170 195.845 ;
        RECT 55.340 194.955 55.530 195.675 ;
        RECT 54.340 194.475 55.170 194.775 ;
        RECT 55.700 194.745 56.020 195.705 ;
        RECT 52.925 194.075 53.260 194.245 ;
        RECT 53.455 194.075 54.130 194.245 ;
        RECT 54.450 193.795 54.820 194.295 ;
        RECT 55.000 194.245 55.170 194.475 ;
        RECT 55.555 194.415 56.020 194.745 ;
        RECT 56.190 195.035 56.360 195.875 ;
        RECT 56.540 195.845 56.855 196.345 ;
        RECT 57.085 195.615 57.425 196.175 ;
        RECT 56.530 195.240 57.425 195.615 ;
        RECT 57.595 195.335 57.765 196.345 ;
        RECT 57.235 195.035 57.425 195.240 ;
        RECT 57.935 195.285 58.265 196.130 ;
        RECT 57.935 195.205 58.325 195.285 ;
        RECT 59.425 195.205 59.755 196.345 ;
        RECT 60.285 195.375 60.615 196.160 ;
        RECT 59.935 195.205 60.615 195.375 ;
        RECT 61.725 195.205 62.055 196.345 ;
        RECT 62.585 195.375 62.915 196.160 ;
        RECT 62.235 195.205 62.915 195.375 ;
        RECT 63.095 195.255 64.305 196.345 ;
        RECT 58.110 195.155 58.325 195.205 ;
        RECT 56.190 194.705 57.065 195.035 ;
        RECT 57.235 194.705 57.985 195.035 ;
        RECT 56.190 194.245 56.360 194.705 ;
        RECT 57.235 194.535 57.435 194.705 ;
        RECT 58.155 194.575 58.325 195.155 ;
        RECT 59.415 194.785 59.765 195.035 ;
        RECT 59.935 194.605 60.105 195.205 ;
        RECT 60.275 194.785 60.625 195.035 ;
        RECT 61.715 194.785 62.065 195.035 ;
        RECT 62.235 194.605 62.405 195.205 ;
        RECT 62.575 194.785 62.925 195.035 ;
        RECT 58.100 194.535 58.325 194.575 ;
        RECT 55.000 194.075 55.405 194.245 ;
        RECT 55.575 194.075 56.360 194.245 ;
        RECT 56.635 193.795 56.845 194.325 ;
        RECT 57.105 194.010 57.435 194.535 ;
        RECT 57.945 194.450 58.325 194.535 ;
        RECT 57.605 193.795 57.775 194.405 ;
        RECT 57.945 194.015 58.275 194.450 ;
        RECT 59.425 193.795 59.695 194.605 ;
        RECT 59.865 193.965 60.195 194.605 ;
        RECT 60.365 193.795 60.605 194.605 ;
        RECT 61.725 193.795 61.995 194.605 ;
        RECT 62.165 193.965 62.495 194.605 ;
        RECT 62.665 193.795 62.905 194.605 ;
        RECT 63.095 194.545 63.615 195.085 ;
        RECT 63.785 194.715 64.305 195.255 ;
        RECT 64.485 195.205 64.815 196.345 ;
        RECT 65.345 195.375 65.675 196.160 ;
        RECT 65.855 195.790 66.460 196.345 ;
        RECT 66.635 195.835 67.115 196.175 ;
        RECT 67.285 195.800 67.540 196.345 ;
        RECT 65.855 195.690 66.470 195.790 ;
        RECT 66.285 195.665 66.470 195.690 ;
        RECT 64.995 195.205 65.675 195.375 ;
        RECT 64.475 194.785 64.825 195.035 ;
        RECT 64.995 194.605 65.165 195.205 ;
        RECT 65.855 195.070 66.115 195.520 ;
        RECT 66.285 195.420 66.615 195.665 ;
        RECT 66.785 195.345 67.540 195.595 ;
        RECT 67.710 195.475 67.985 196.175 ;
        RECT 66.770 195.310 67.540 195.345 ;
        RECT 66.755 195.300 67.540 195.310 ;
        RECT 66.750 195.285 67.645 195.300 ;
        RECT 66.730 195.270 67.645 195.285 ;
        RECT 66.710 195.260 67.645 195.270 ;
        RECT 66.685 195.250 67.645 195.260 ;
        RECT 66.615 195.220 67.645 195.250 ;
        RECT 66.595 195.190 67.645 195.220 ;
        RECT 66.575 195.160 67.645 195.190 ;
        RECT 66.545 195.135 67.645 195.160 ;
        RECT 66.510 195.100 67.645 195.135 ;
        RECT 66.480 195.095 67.645 195.100 ;
        RECT 66.480 195.090 66.870 195.095 ;
        RECT 66.480 195.080 66.845 195.090 ;
        RECT 66.480 195.075 66.830 195.080 ;
        RECT 66.480 195.070 66.815 195.075 ;
        RECT 65.855 195.065 66.815 195.070 ;
        RECT 65.855 195.055 66.805 195.065 ;
        RECT 65.855 195.050 66.795 195.055 ;
        RECT 65.855 195.040 66.785 195.050 ;
        RECT 65.335 194.785 65.685 195.035 ;
        RECT 65.855 195.030 66.780 195.040 ;
        RECT 65.855 195.025 66.775 195.030 ;
        RECT 65.855 195.010 66.765 195.025 ;
        RECT 65.855 194.995 66.760 195.010 ;
        RECT 65.855 194.970 66.750 194.995 ;
        RECT 65.855 194.900 66.745 194.970 ;
        RECT 63.095 193.795 64.305 194.545 ;
        RECT 64.485 193.795 64.755 194.605 ;
        RECT 64.925 193.965 65.255 194.605 ;
        RECT 65.425 193.795 65.665 194.605 ;
        RECT 65.855 194.345 66.405 194.730 ;
        RECT 66.575 194.175 66.745 194.900 ;
        RECT 65.855 194.005 66.745 194.175 ;
        RECT 66.915 194.500 67.245 194.925 ;
        RECT 67.415 194.700 67.645 195.095 ;
        RECT 66.915 194.015 67.135 194.500 ;
        RECT 67.815 194.445 67.985 195.475 ;
        RECT 69.135 195.285 69.465 196.130 ;
        RECT 69.635 195.335 69.805 196.345 ;
        RECT 69.975 195.615 70.315 196.175 ;
        RECT 70.545 195.845 70.860 196.345 ;
        RECT 71.040 195.875 71.925 196.045 ;
        RECT 69.075 195.205 69.465 195.285 ;
        RECT 69.975 195.240 70.870 195.615 ;
        RECT 69.075 195.155 69.290 195.205 ;
        RECT 69.075 194.575 69.245 195.155 ;
        RECT 69.975 195.035 70.165 195.240 ;
        RECT 71.040 195.035 71.210 195.875 ;
        RECT 72.150 195.845 72.400 196.175 ;
        RECT 69.415 194.705 70.165 195.035 ;
        RECT 70.335 194.705 71.210 195.035 ;
        RECT 69.075 194.535 69.300 194.575 ;
        RECT 69.965 194.535 70.165 194.705 ;
        RECT 69.075 194.450 69.455 194.535 ;
        RECT 67.305 193.795 67.555 194.335 ;
        RECT 67.725 193.965 67.985 194.445 ;
        RECT 69.125 194.015 69.455 194.450 ;
        RECT 69.625 193.795 69.795 194.405 ;
        RECT 69.965 194.010 70.295 194.535 ;
        RECT 70.555 193.795 70.765 194.325 ;
        RECT 71.040 194.245 71.210 194.705 ;
        RECT 71.380 194.745 71.700 195.705 ;
        RECT 71.870 194.955 72.060 195.675 ;
        RECT 72.230 194.775 72.400 195.845 ;
        RECT 72.570 195.545 72.740 196.345 ;
        RECT 72.910 195.900 74.015 196.070 ;
        RECT 72.910 195.285 73.080 195.900 ;
        RECT 74.225 195.750 74.475 196.175 ;
        RECT 74.645 195.885 74.910 196.345 ;
        RECT 73.250 195.365 73.780 195.730 ;
        RECT 74.225 195.620 74.530 195.750 ;
        RECT 72.570 195.195 73.080 195.285 ;
        RECT 72.570 195.025 73.440 195.195 ;
        RECT 72.570 194.955 72.740 195.025 ;
        RECT 72.860 194.775 73.060 194.805 ;
        RECT 71.380 194.415 71.845 194.745 ;
        RECT 72.230 194.475 73.060 194.775 ;
        RECT 72.230 194.245 72.400 194.475 ;
        RECT 71.040 194.075 71.825 194.245 ;
        RECT 71.995 194.075 72.400 194.245 ;
        RECT 72.580 193.795 72.950 194.295 ;
        RECT 73.270 194.245 73.440 195.025 ;
        RECT 73.610 194.665 73.780 195.365 ;
        RECT 73.950 194.835 74.190 195.430 ;
        RECT 73.610 194.445 74.135 194.665 ;
        RECT 74.360 194.515 74.530 195.620 ;
        RECT 74.305 194.385 74.530 194.515 ;
        RECT 74.700 194.425 74.980 195.375 ;
        RECT 74.305 194.245 74.475 194.385 ;
        RECT 73.270 194.075 73.945 194.245 ;
        RECT 74.140 194.075 74.475 194.245 ;
        RECT 74.645 193.795 74.895 194.255 ;
        RECT 75.150 194.055 75.335 196.175 ;
        RECT 75.505 195.845 75.835 196.345 ;
        RECT 76.005 195.675 76.175 196.175 ;
        RECT 75.510 195.505 76.175 195.675 ;
        RECT 75.510 194.515 75.740 195.505 ;
        RECT 75.910 194.685 76.260 195.335 ;
        RECT 76.435 195.180 76.725 196.345 ;
        RECT 76.895 195.910 82.240 196.345 ;
        RECT 82.415 195.910 87.760 196.345 ;
        RECT 75.510 194.345 76.175 194.515 ;
        RECT 75.505 193.795 75.835 194.175 ;
        RECT 76.005 194.055 76.175 194.345 ;
        RECT 76.435 193.795 76.725 194.520 ;
        RECT 78.480 194.340 78.820 195.170 ;
        RECT 80.300 194.660 80.650 195.910 ;
        RECT 84.000 194.340 84.340 195.170 ;
        RECT 85.820 194.660 86.170 195.910 ;
        RECT 87.935 195.255 89.145 196.345 ;
        RECT 87.935 194.545 88.455 195.085 ;
        RECT 88.625 194.715 89.145 195.255 ;
        RECT 89.315 195.255 90.525 196.345 ;
        RECT 112.275 196.205 112.445 196.930 ;
        RECT 112.665 196.605 113.185 196.760 ;
        RECT 113.355 196.720 113.685 197.270 ;
        RECT 114.995 197.110 115.165 197.830 ;
        RECT 116.475 197.660 116.805 197.685 ;
        RECT 113.985 196.940 115.165 197.110 ;
        RECT 112.665 196.550 113.225 196.605 ;
        RECT 113.855 196.595 114.780 196.770 ;
        RECT 113.805 196.550 114.780 196.595 ;
        RECT 112.665 196.440 114.780 196.550 ;
        RECT 112.665 196.430 113.935 196.440 ;
        RECT 113.100 196.380 113.935 196.430 ;
        RECT 114.995 196.205 115.165 196.940 ;
        RECT 112.275 195.945 113.285 196.205 ;
        RECT 113.845 195.945 115.165 196.205 ;
        RECT 112.275 195.345 112.445 195.945 ;
        RECT 112.615 195.600 114.825 195.770 ;
        RECT 112.615 195.515 113.190 195.600 ;
        RECT 113.920 195.515 114.825 195.600 ;
        RECT 114.995 195.460 115.165 195.945 ;
        RECT 115.335 197.490 116.805 197.660 ;
        RECT 115.335 195.800 115.505 197.490 ;
        RECT 116.975 197.325 117.145 197.910 ;
        RECT 117.315 197.830 118.365 198.080 ;
        RECT 117.315 197.750 117.885 197.830 ;
        RECT 116.975 197.320 117.545 197.325 ;
        RECT 115.675 197.150 117.545 197.320 ;
        RECT 115.675 196.195 115.845 197.150 ;
        RECT 116.015 196.810 116.985 196.980 ;
        RECT 116.015 196.160 116.185 196.810 ;
        RECT 117.180 196.795 117.545 197.150 ;
        RECT 117.715 197.230 117.885 197.750 ;
        RECT 118.535 197.660 119.520 198.095 ;
        RECT 120.430 198.085 120.605 198.700 ;
        RECT 119.705 197.830 120.605 198.085 ;
        RECT 118.080 197.400 120.260 197.660 ;
        RECT 118.535 197.370 120.260 197.400 ;
        RECT 117.715 196.930 118.365 197.230 ;
        RECT 118.535 196.930 119.520 197.370 ;
        RECT 120.435 197.285 120.605 197.830 ;
        RECT 120.880 197.625 121.050 198.560 ;
        RECT 121.520 198.495 122.115 198.735 ;
        RECT 122.705 198.685 122.875 198.850 ;
        RECT 122.285 198.325 122.505 198.680 ;
        RECT 123.155 198.500 123.325 199.190 ;
        RECT 123.545 198.905 124.065 199.060 ;
        RECT 124.235 199.020 124.565 199.570 ;
        RECT 125.875 199.410 126.045 200.150 ;
        RECT 126.395 200.400 126.805 200.575 ;
        RECT 127.050 200.570 127.240 201.150 ;
        RECT 127.615 200.580 127.785 201.290 ;
        RECT 128.060 201.150 129.225 201.310 ;
        RECT 129.395 201.280 130.425 201.540 ;
        RECT 130.595 201.280 131.490 201.610 ;
        RECT 131.660 201.370 132.625 201.630 ;
        RECT 129.395 201.170 129.965 201.280 ;
        RECT 128.060 200.800 128.765 201.150 ;
        RECT 129.755 200.960 129.965 201.170 ;
        RECT 131.315 201.185 131.490 201.280 ;
        RECT 127.615 200.400 128.390 200.580 ;
        RECT 126.395 200.335 128.390 200.400 ;
        RECT 126.395 200.060 127.785 200.335 ;
        RECT 126.215 199.610 128.425 199.890 ;
        RECT 126.215 199.505 127.185 199.610 ;
        RECT 127.855 199.505 128.425 199.610 ;
        RECT 128.595 199.795 128.765 200.800 ;
        RECT 128.935 200.790 129.565 200.860 ;
        RECT 130.135 200.790 131.145 201.045 ;
        RECT 128.935 200.520 131.145 200.790 ;
        RECT 131.315 200.940 132.215 201.185 ;
        RECT 128.935 200.070 131.145 200.350 ;
        RECT 128.935 199.965 129.505 200.070 ;
        RECT 130.175 199.965 131.145 200.070 ;
        RECT 131.315 200.325 131.490 200.940 ;
        RECT 132.385 200.770 132.625 201.370 ;
        RECT 131.660 200.510 132.625 200.770 ;
        RECT 131.315 200.080 132.215 200.325 ;
        RECT 129.675 199.795 130.005 199.900 ;
        RECT 131.315 199.795 131.490 200.080 ;
        RECT 132.385 199.910 132.625 200.510 ;
        RECT 128.595 199.470 129.225 199.795 ;
        RECT 124.865 199.335 126.045 199.410 ;
        RECT 127.355 199.335 127.685 199.440 ;
        RECT 128.595 199.335 128.765 199.470 ;
        RECT 124.865 199.240 126.505 199.335 ;
        RECT 123.545 198.850 124.105 198.905 ;
        RECT 124.735 198.895 125.660 199.070 ;
        RECT 124.685 198.850 125.660 198.895 ;
        RECT 123.545 198.740 125.660 198.850 ;
        RECT 125.875 199.010 126.505 199.240 ;
        RECT 123.545 198.730 124.815 198.740 ;
        RECT 123.980 198.680 124.815 198.730 ;
        RECT 121.220 198.155 122.505 198.325 ;
        RECT 121.220 197.795 121.585 198.155 ;
        RECT 122.705 197.985 122.875 198.490 ;
        RECT 121.755 197.815 122.875 197.985 ;
        RECT 123.155 198.170 123.830 198.500 ;
        RECT 124.685 198.445 124.855 198.450 ;
        RECT 121.755 197.625 121.925 197.815 ;
        RECT 120.880 197.455 121.925 197.625 ;
        RECT 121.665 197.285 121.925 197.455 ;
        RECT 122.145 197.405 122.475 197.605 ;
        RECT 123.155 197.495 123.325 198.170 ;
        RECT 124.005 198.145 124.855 198.445 ;
        RECT 125.025 198.250 125.685 198.420 ;
        RECT 123.520 197.975 123.895 198.000 ;
        RECT 125.025 197.975 125.255 198.250 ;
        RECT 125.875 198.080 126.045 199.010 ;
        RECT 126.675 198.885 127.965 199.335 ;
        RECT 128.135 199.010 128.765 199.335 ;
        RECT 126.675 198.490 126.895 198.885 ;
        RECT 126.215 198.210 126.895 198.490 ;
        RECT 123.520 197.760 125.255 197.975 ;
        RECT 120.435 197.200 121.405 197.285 ;
        RECT 119.690 197.115 121.405 197.200 ;
        RECT 121.665 197.115 121.995 197.285 ;
        RECT 119.690 196.930 120.605 197.115 ;
        RECT 122.175 196.945 122.475 197.405 ;
        RECT 122.655 197.125 123.325 197.495 ;
        RECT 124.045 197.740 125.255 197.760 ;
        RECT 125.425 197.750 126.045 198.080 ;
        RECT 127.065 198.020 127.625 198.715 ;
        RECT 127.795 198.490 127.965 198.885 ;
        RECT 127.795 198.210 128.425 198.490 ;
        RECT 123.510 197.310 123.850 197.480 ;
        RECT 124.045 197.420 124.375 197.740 ;
        RECT 117.715 196.670 117.885 196.930 ;
        RECT 120.435 196.670 120.605 196.930 ;
        RECT 120.775 196.775 122.875 196.945 ;
        RECT 120.775 196.695 121.105 196.775 ;
        RECT 116.525 196.605 116.695 196.610 ;
        RECT 116.385 196.330 117.545 196.605 ;
        RECT 116.015 195.970 117.545 196.160 ;
        RECT 117.715 196.150 119.175 196.670 ;
        RECT 115.335 195.630 116.360 195.800 ;
        RECT 117.715 195.790 118.635 196.150 ;
        RECT 119.345 195.980 120.605 196.670 ;
        RECT 113.355 195.345 113.685 195.430 ;
        RECT 114.995 195.345 115.925 195.460 ;
        RECT 89.315 194.715 89.835 195.255 ;
        RECT 90.005 194.545 90.525 195.085 ;
        RECT 76.895 193.795 82.240 194.340 ;
        RECT 82.415 193.795 87.760 194.340 ;
        RECT 87.935 193.795 89.145 194.545 ;
        RECT 89.315 193.795 90.525 194.545 ;
        RECT 112.275 195.015 112.825 195.345 ;
        RECT 112.995 195.175 114.065 195.345 ;
        RECT 11.950 193.625 90.610 193.795 ;
        RECT 12.035 192.875 13.245 193.625 ;
        RECT 13.415 193.080 18.760 193.625 ;
        RECT 18.935 193.080 24.280 193.625 ;
        RECT 24.455 193.080 29.800 193.625 ;
        RECT 29.975 193.080 35.320 193.625 ;
        RECT 12.035 192.335 12.555 192.875 ;
        RECT 12.725 192.165 13.245 192.705 ;
        RECT 15.000 192.250 15.340 193.080 ;
        RECT 12.035 191.075 13.245 192.165 ;
        RECT 16.820 191.510 17.170 192.760 ;
        RECT 20.520 192.250 20.860 193.080 ;
        RECT 22.340 191.510 22.690 192.760 ;
        RECT 26.040 192.250 26.380 193.080 ;
        RECT 27.860 191.510 28.210 192.760 ;
        RECT 31.560 192.250 31.900 193.080 ;
        RECT 35.495 192.855 37.165 193.625 ;
        RECT 37.795 192.900 38.085 193.625 ;
        RECT 38.255 192.875 39.465 193.625 ;
        RECT 39.635 192.975 39.895 193.455 ;
        RECT 40.065 193.085 40.315 193.625 ;
        RECT 33.380 191.510 33.730 192.760 ;
        RECT 35.495 192.335 36.245 192.855 ;
        RECT 36.415 192.165 37.165 192.685 ;
        RECT 38.255 192.335 38.775 192.875 ;
        RECT 13.415 191.075 18.760 191.510 ;
        RECT 18.935 191.075 24.280 191.510 ;
        RECT 24.455 191.075 29.800 191.510 ;
        RECT 29.975 191.075 35.320 191.510 ;
        RECT 35.495 191.075 37.165 192.165 ;
        RECT 37.795 191.075 38.085 192.240 ;
        RECT 38.945 192.165 39.465 192.705 ;
        RECT 38.255 191.075 39.465 192.165 ;
        RECT 39.635 191.945 39.805 192.975 ;
        RECT 40.485 192.920 40.705 193.405 ;
        RECT 39.975 192.325 40.205 192.720 ;
        RECT 40.375 192.495 40.705 192.920 ;
        RECT 40.875 193.245 41.765 193.415 ;
        RECT 40.875 192.520 41.045 193.245 ;
        RECT 41.215 192.690 41.765 193.075 ;
        RECT 41.955 192.815 42.195 193.625 ;
        RECT 42.365 192.815 42.695 193.455 ;
        RECT 42.865 192.815 43.135 193.625 ;
        RECT 43.400 193.125 43.895 193.455 ;
        RECT 40.875 192.450 41.765 192.520 ;
        RECT 40.870 192.425 41.765 192.450 ;
        RECT 40.860 192.410 41.765 192.425 ;
        RECT 40.855 192.395 41.765 192.410 ;
        RECT 40.845 192.390 41.765 192.395 ;
        RECT 40.840 192.380 41.765 192.390 ;
        RECT 41.935 192.385 42.285 192.635 ;
        RECT 40.835 192.370 41.765 192.380 ;
        RECT 40.825 192.365 41.765 192.370 ;
        RECT 40.815 192.355 41.765 192.365 ;
        RECT 40.805 192.350 41.765 192.355 ;
        RECT 40.805 192.345 41.140 192.350 ;
        RECT 40.790 192.340 41.140 192.345 ;
        RECT 40.775 192.330 41.140 192.340 ;
        RECT 40.750 192.325 41.140 192.330 ;
        RECT 39.975 192.320 41.140 192.325 ;
        RECT 39.975 192.285 41.110 192.320 ;
        RECT 39.975 192.260 41.075 192.285 ;
        RECT 39.975 192.230 41.045 192.260 ;
        RECT 39.975 192.200 41.025 192.230 ;
        RECT 39.975 192.170 41.005 192.200 ;
        RECT 39.975 192.160 40.935 192.170 ;
        RECT 39.975 192.150 40.910 192.160 ;
        RECT 39.975 192.135 40.890 192.150 ;
        RECT 39.975 192.120 40.870 192.135 ;
        RECT 40.080 192.110 40.865 192.120 ;
        RECT 40.080 192.075 40.850 192.110 ;
        RECT 39.635 191.245 39.910 191.945 ;
        RECT 40.080 191.825 40.835 192.075 ;
        RECT 41.005 191.755 41.335 192.000 ;
        RECT 41.505 191.900 41.765 192.350 ;
        RECT 42.455 192.215 42.625 192.815 ;
        RECT 42.795 192.385 43.145 192.635 ;
        RECT 41.945 192.045 42.625 192.215 ;
        RECT 41.150 191.730 41.335 191.755 ;
        RECT 41.150 191.630 41.765 191.730 ;
        RECT 40.080 191.075 40.335 191.620 ;
        RECT 40.505 191.245 40.985 191.585 ;
        RECT 41.160 191.075 41.765 191.630 ;
        RECT 41.945 191.260 42.275 192.045 ;
        RECT 42.805 191.075 43.135 192.215 ;
        RECT 43.315 191.635 43.555 192.945 ;
        RECT 43.725 192.215 43.895 193.125 ;
        RECT 44.115 192.385 44.465 193.350 ;
        RECT 44.645 192.385 44.945 193.355 ;
        RECT 45.125 192.385 45.405 193.355 ;
        RECT 45.585 192.825 45.855 193.625 ;
        RECT 46.025 192.905 46.365 193.415 ;
        RECT 46.560 193.235 46.890 193.625 ;
        RECT 47.060 193.065 47.285 193.445 ;
        RECT 45.600 192.385 45.930 192.635 ;
        RECT 45.600 192.215 45.915 192.385 ;
        RECT 43.725 192.045 45.915 192.215 ;
        RECT 43.320 191.075 43.655 191.455 ;
        RECT 43.825 191.245 44.075 192.045 ;
        RECT 44.295 191.075 44.625 191.795 ;
        RECT 44.810 191.245 45.060 192.045 ;
        RECT 45.525 191.075 45.855 191.875 ;
        RECT 46.105 191.505 46.365 192.905 ;
        RECT 46.545 192.385 46.785 193.035 ;
        RECT 46.955 192.885 47.285 193.065 ;
        RECT 46.955 192.215 47.130 192.885 ;
        RECT 47.485 192.715 47.715 193.335 ;
        RECT 47.895 192.895 48.195 193.625 ;
        RECT 48.375 192.790 48.665 193.625 ;
        RECT 48.835 193.225 49.790 193.395 ;
        RECT 50.205 193.235 50.535 193.625 ;
        RECT 47.300 192.385 47.715 192.715 ;
        RECT 47.895 192.385 48.190 192.715 ;
        RECT 48.835 192.345 49.005 193.225 ;
        RECT 50.705 193.055 50.875 193.375 ;
        RECT 51.045 193.235 51.375 193.625 ;
        RECT 51.595 193.080 56.940 193.625 ;
        RECT 49.175 192.885 51.425 193.055 ;
        RECT 49.175 192.385 49.405 192.885 ;
        RECT 49.575 192.465 49.950 192.635 ;
        RECT 46.025 191.245 46.365 191.505 ;
        RECT 46.545 192.025 47.130 192.215 ;
        RECT 46.545 191.255 46.820 192.025 ;
        RECT 47.300 191.855 48.195 192.185 ;
        RECT 46.990 191.685 48.195 191.855 ;
        RECT 46.990 191.255 47.320 191.685 ;
        RECT 47.490 191.075 47.685 191.515 ;
        RECT 47.865 191.255 48.195 191.685 ;
        RECT 48.375 192.175 49.005 192.345 ;
        RECT 49.780 192.265 49.950 192.465 ;
        RECT 50.120 192.435 50.670 192.635 ;
        RECT 50.840 192.265 51.085 192.715 ;
        RECT 48.375 191.245 48.695 192.175 ;
        RECT 49.780 192.095 51.085 192.265 ;
        RECT 51.255 191.925 51.425 192.885 ;
        RECT 53.180 192.250 53.520 193.080 ;
        RECT 57.115 192.855 60.625 193.625 ;
        RECT 60.855 193.145 61.135 193.625 ;
        RECT 61.305 192.975 61.565 193.365 ;
        RECT 61.740 193.145 61.995 193.625 ;
        RECT 62.165 192.975 62.460 193.365 ;
        RECT 62.640 193.145 62.915 193.625 ;
        RECT 63.085 193.125 63.385 193.455 ;
        RECT 48.875 191.755 50.115 191.925 ;
        RECT 48.875 191.245 49.275 191.755 ;
        RECT 49.445 191.075 49.615 191.585 ;
        RECT 49.785 191.245 50.115 191.755 ;
        RECT 50.285 191.075 50.455 191.925 ;
        RECT 51.045 191.245 51.425 191.925 ;
        RECT 55.000 191.510 55.350 192.760 ;
        RECT 57.115 192.335 58.765 192.855 ;
        RECT 60.810 192.805 62.460 192.975 ;
        RECT 58.935 192.165 60.625 192.685 ;
        RECT 51.595 191.075 56.940 191.510 ;
        RECT 57.115 191.075 60.625 192.165 ;
        RECT 60.810 192.295 61.215 192.805 ;
        RECT 61.385 192.465 62.525 192.635 ;
        RECT 60.810 192.125 61.565 192.295 ;
        RECT 60.850 191.075 61.135 191.945 ;
        RECT 61.305 191.875 61.565 192.125 ;
        RECT 62.355 192.215 62.525 192.465 ;
        RECT 62.695 192.385 63.045 192.955 ;
        RECT 63.215 192.215 63.385 193.125 ;
        RECT 63.555 192.900 63.845 193.625 ;
        RECT 64.100 193.125 64.595 193.455 ;
        RECT 62.355 192.045 63.385 192.215 ;
        RECT 61.305 191.705 62.425 191.875 ;
        RECT 61.305 191.245 61.565 191.705 ;
        RECT 61.740 191.075 61.995 191.535 ;
        RECT 62.165 191.245 62.425 191.705 ;
        RECT 62.595 191.075 62.905 191.875 ;
        RECT 63.075 191.245 63.385 192.045 ;
        RECT 63.555 191.075 63.845 192.240 ;
        RECT 64.015 191.635 64.255 192.945 ;
        RECT 64.425 192.215 64.595 193.125 ;
        RECT 64.815 192.385 65.165 193.350 ;
        RECT 65.345 192.385 65.645 193.355 ;
        RECT 65.825 192.385 66.105 193.355 ;
        RECT 66.285 192.825 66.555 193.625 ;
        RECT 66.725 192.905 67.065 193.415 ;
        RECT 67.260 193.235 67.590 193.625 ;
        RECT 67.760 193.065 67.985 193.445 ;
        RECT 66.300 192.385 66.630 192.635 ;
        RECT 66.300 192.215 66.615 192.385 ;
        RECT 64.425 192.045 66.615 192.215 ;
        RECT 64.020 191.075 64.355 191.455 ;
        RECT 64.525 191.245 64.775 192.045 ;
        RECT 64.995 191.075 65.325 191.795 ;
        RECT 65.510 191.245 65.760 192.045 ;
        RECT 66.225 191.075 66.555 191.875 ;
        RECT 66.805 191.505 67.065 192.905 ;
        RECT 67.245 192.385 67.485 193.035 ;
        RECT 67.655 192.885 67.985 193.065 ;
        RECT 67.655 192.215 67.830 192.885 ;
        RECT 68.185 192.715 68.415 193.335 ;
        RECT 68.595 192.895 68.895 193.625 ;
        RECT 69.160 193.125 69.655 193.455 ;
        RECT 68.000 192.385 68.415 192.715 ;
        RECT 68.595 192.385 68.890 192.715 ;
        RECT 66.725 191.245 67.065 191.505 ;
        RECT 67.245 192.025 67.830 192.215 ;
        RECT 67.245 191.255 67.520 192.025 ;
        RECT 68.000 191.855 68.895 192.185 ;
        RECT 67.690 191.685 68.895 191.855 ;
        RECT 67.690 191.255 68.020 191.685 ;
        RECT 68.190 191.075 68.385 191.515 ;
        RECT 68.565 191.255 68.895 191.685 ;
        RECT 69.075 191.635 69.315 192.945 ;
        RECT 69.485 192.215 69.655 193.125 ;
        RECT 69.875 192.385 70.225 193.350 ;
        RECT 70.405 192.385 70.705 193.355 ;
        RECT 70.885 192.385 71.165 193.355 ;
        RECT 71.345 192.825 71.615 193.625 ;
        RECT 71.785 192.905 72.125 193.415 ;
        RECT 72.460 193.115 72.700 193.625 ;
        RECT 72.880 193.115 73.160 193.445 ;
        RECT 73.390 193.115 73.605 193.625 ;
        RECT 71.360 192.385 71.690 192.635 ;
        RECT 71.360 192.215 71.675 192.385 ;
        RECT 69.485 192.045 71.675 192.215 ;
        RECT 69.080 191.075 69.415 191.455 ;
        RECT 69.585 191.245 69.835 192.045 ;
        RECT 70.055 191.075 70.385 191.795 ;
        RECT 70.570 191.245 70.820 192.045 ;
        RECT 71.285 191.075 71.615 191.875 ;
        RECT 71.865 191.505 72.125 192.905 ;
        RECT 72.355 192.385 72.710 192.945 ;
        RECT 72.880 192.215 73.050 193.115 ;
        RECT 73.220 192.385 73.485 192.945 ;
        RECT 73.775 192.885 74.390 193.455 ;
        RECT 74.595 193.080 79.940 193.625 ;
        RECT 80.115 193.080 85.460 193.625 ;
        RECT 73.735 192.215 73.905 192.715 ;
        RECT 72.480 192.045 73.905 192.215 ;
        RECT 72.480 191.870 72.870 192.045 ;
        RECT 71.785 191.245 72.125 191.505 ;
        RECT 73.355 191.075 73.685 191.875 ;
        RECT 74.075 191.865 74.390 192.885 ;
        RECT 76.180 192.250 76.520 193.080 ;
        RECT 73.855 191.245 74.390 191.865 ;
        RECT 78.000 191.510 78.350 192.760 ;
        RECT 81.700 192.250 82.040 193.080 ;
        RECT 85.635 192.855 89.145 193.625 ;
        RECT 89.315 192.875 90.525 193.625 ;
        RECT 83.520 191.510 83.870 192.760 ;
        RECT 85.635 192.335 87.285 192.855 ;
        RECT 87.455 192.165 89.145 192.685 ;
        RECT 74.595 191.075 79.940 191.510 ;
        RECT 80.115 191.075 85.460 191.510 ;
        RECT 85.635 191.075 89.145 192.165 ;
        RECT 89.315 192.165 89.835 192.705 ;
        RECT 90.005 192.335 90.525 192.875 ;
        RECT 112.275 193.450 112.445 195.015 ;
        RECT 112.995 194.800 113.165 195.175 ;
        RECT 112.615 194.630 113.165 194.800 ;
        RECT 113.345 194.540 113.715 194.895 ;
        RECT 113.895 194.800 114.065 195.175 ;
        RECT 114.235 195.290 115.925 195.345 ;
        RECT 114.235 195.015 115.165 195.290 ;
        RECT 113.895 194.630 114.825 194.800 ;
        RECT 114.995 193.450 115.165 195.015 ;
        RECT 115.515 194.880 115.925 195.055 ;
        RECT 116.170 195.050 116.360 195.630 ;
        RECT 116.735 195.060 116.905 195.770 ;
        RECT 117.180 195.460 118.635 195.790 ;
        RECT 118.805 195.460 120.605 195.980 ;
        RECT 120.905 195.755 121.075 196.470 ;
        RECT 121.275 196.415 121.995 196.605 ;
        RECT 122.705 196.540 122.875 196.775 ;
        RECT 123.155 196.720 123.325 197.125 ;
        RECT 123.655 197.250 123.850 197.310 ;
        RECT 124.545 197.265 125.660 197.550 ;
        RECT 124.545 197.250 124.715 197.265 ;
        RECT 123.655 197.080 124.715 197.250 ;
        RECT 125.875 197.220 126.045 197.750 ;
        RECT 126.215 197.620 128.425 198.020 ;
        RECT 128.595 197.680 128.765 199.010 ;
        RECT 129.395 199.345 130.685 199.795 ;
        RECT 130.855 199.470 131.490 199.795 ;
        RECT 131.660 199.650 132.625 199.910 ;
        RECT 129.395 198.950 129.565 199.345 ;
        RECT 128.935 198.670 129.565 198.950 ;
        RECT 129.735 198.480 130.295 199.175 ;
        RECT 130.465 198.950 130.685 199.345 ;
        RECT 131.315 199.465 131.490 199.470 ;
        RECT 132.400 199.475 132.625 199.650 ;
        RECT 132.795 199.645 133.045 205.655 ;
        RECT 134.035 205.485 134.205 206.040 ;
        RECT 134.465 205.610 134.925 205.780 ;
        RECT 133.475 205.440 134.205 205.485 ;
        RECT 133.475 205.225 134.585 205.440 ;
        RECT 134.035 205.110 134.585 205.225 ;
        RECT 134.755 205.345 134.925 205.610 ;
        RECT 135.095 205.515 135.745 205.865 ;
        RECT 136.755 205.785 137.655 206.040 ;
        RECT 135.915 205.610 136.585 205.780 ;
        RECT 135.915 205.345 136.085 205.610 ;
        RECT 136.755 205.440 136.930 205.785 ;
        RECT 137.825 205.615 138.065 206.215 ;
        RECT 134.755 205.115 136.085 205.345 ;
        RECT 136.255 205.185 136.930 205.440 ;
        RECT 137.100 205.355 138.065 205.615 ;
        RECT 136.255 205.110 137.655 205.185 ;
        RECT 133.215 204.795 133.840 205.055 ;
        RECT 133.215 204.195 133.385 204.795 ;
        RECT 134.035 204.625 134.205 205.110 ;
        RECT 134.465 204.755 136.585 204.940 ;
        RECT 136.755 204.925 137.655 205.110 ;
        RECT 133.555 204.500 134.205 204.625 ;
        RECT 133.555 204.365 134.665 204.500 ;
        RECT 134.035 204.250 134.665 204.365 ;
        RECT 134.835 204.305 135.785 204.585 ;
        RECT 136.755 204.515 136.930 204.925 ;
        RECT 137.825 204.755 138.065 205.355 ;
        RECT 136.295 204.325 136.930 204.515 ;
        RECT 137.100 204.495 138.065 204.755 ;
        RECT 136.295 204.250 137.655 204.325 ;
        RECT 133.215 203.935 133.840 204.195 ;
        RECT 133.215 203.335 133.385 203.935 ;
        RECT 134.035 203.765 134.205 204.250 ;
        RECT 134.795 204.080 136.160 204.135 ;
        RECT 133.555 203.505 134.205 203.765 ;
        RECT 134.485 203.965 136.585 204.080 ;
        RECT 134.485 203.910 134.925 203.965 ;
        RECT 134.485 203.745 134.655 203.910 ;
        RECT 136.030 203.830 136.585 203.965 ;
        RECT 136.755 204.065 137.655 204.250 ;
        RECT 133.215 203.075 133.840 203.335 ;
        RECT 133.215 202.490 133.385 203.075 ;
        RECT 134.035 202.905 134.205 203.505 ;
        RECT 133.555 202.660 134.205 202.905 ;
        RECT 134.485 203.045 134.655 203.550 ;
        RECT 134.855 203.385 135.075 203.740 ;
        RECT 135.245 203.555 135.840 203.795 ;
        RECT 134.855 203.215 136.140 203.385 ;
        RECT 134.485 202.875 135.605 203.045 ;
        RECT 135.435 202.685 135.605 202.875 ;
        RECT 135.775 202.855 136.140 203.215 ;
        RECT 136.310 202.685 136.480 203.620 ;
        RECT 134.035 202.555 134.205 202.660 ;
        RECT 133.215 202.215 133.840 202.490 ;
        RECT 133.215 201.630 133.385 202.215 ;
        RECT 134.035 202.185 134.705 202.555 ;
        RECT 134.885 202.465 135.215 202.665 ;
        RECT 135.435 202.515 136.480 202.685 ;
        RECT 136.755 203.465 136.930 204.065 ;
        RECT 137.825 203.895 138.065 204.495 ;
        RECT 137.100 203.635 138.065 203.895 ;
        RECT 136.755 203.205 137.725 203.465 ;
        RECT 136.755 202.605 136.925 203.205 ;
        RECT 138.235 203.035 138.485 209.045 ;
        RECT 138.655 209.040 138.825 209.215 ;
        RECT 138.655 208.780 139.280 209.040 ;
        RECT 138.655 208.180 138.825 208.780 ;
        RECT 139.475 208.610 139.645 209.220 ;
        RECT 140.275 209.465 141.565 209.915 ;
        RECT 141.735 209.590 142.365 209.915 ;
        RECT 143.425 209.855 143.685 210.025 ;
        RECT 143.935 209.905 144.235 210.365 ;
        RECT 144.915 210.185 145.085 210.585 ;
        RECT 145.995 210.500 146.325 210.585 ;
        RECT 140.275 209.070 140.445 209.465 ;
        RECT 139.815 208.790 140.445 209.070 ;
        RECT 138.995 208.360 139.645 208.610 ;
        RECT 140.615 208.600 141.175 209.295 ;
        RECT 141.345 209.070 141.565 209.465 ;
        RECT 141.345 208.790 142.025 209.070 ;
        RECT 138.655 207.920 139.280 208.180 ;
        RECT 138.655 207.320 138.825 207.920 ;
        RECT 139.475 207.800 139.645 208.360 ;
        RECT 139.815 208.200 142.025 208.600 ;
        RECT 142.195 208.120 142.365 209.590 ;
        RECT 142.640 209.685 143.685 209.855 ;
        RECT 143.905 209.705 144.235 209.905 ;
        RECT 144.415 209.985 145.085 210.185 ;
        RECT 145.255 210.330 145.830 210.415 ;
        RECT 146.560 210.330 147.465 210.415 ;
        RECT 145.255 210.160 147.465 210.330 ;
        RECT 147.635 209.985 147.805 210.585 ;
        RECT 144.415 209.815 145.925 209.985 ;
        RECT 144.915 209.725 145.925 209.815 ;
        RECT 146.485 209.725 147.805 209.985 ;
        RECT 142.640 208.750 142.810 209.685 ;
        RECT 142.980 209.155 143.345 209.515 ;
        RECT 143.515 209.495 143.685 209.685 ;
        RECT 143.515 209.325 144.635 209.495 ;
        RECT 142.980 208.985 144.265 209.155 ;
        RECT 143.280 208.575 143.875 208.815 ;
        RECT 144.045 208.630 144.265 208.985 ;
        RECT 144.465 208.820 144.635 209.325 ;
        RECT 142.535 208.405 143.090 208.540 ;
        RECT 144.465 208.460 144.635 208.625 ;
        RECT 144.195 208.405 144.635 208.460 ;
        RECT 142.535 208.290 144.635 208.405 ;
        RECT 144.915 208.490 145.085 209.725 ;
        RECT 145.255 209.380 146.665 209.550 ;
        RECT 147.635 209.540 147.805 209.725 ;
        RECT 145.255 209.060 145.825 209.380 ;
        RECT 145.255 208.660 145.825 208.890 ;
        RECT 145.995 208.805 146.325 209.210 ;
        RECT 146.495 209.030 146.665 209.380 ;
        RECT 146.835 209.210 147.805 209.540 ;
        RECT 146.495 208.780 147.465 209.030 ;
        RECT 142.960 208.235 144.325 208.290 ;
        RECT 144.915 208.120 145.485 208.490 ;
        RECT 140.275 207.820 141.565 208.030 ;
        RECT 139.475 207.750 140.105 207.800 ;
        RECT 138.995 207.530 140.105 207.750 ;
        RECT 138.995 207.500 139.645 207.530 ;
        RECT 138.655 207.060 139.280 207.320 ;
        RECT 138.655 206.475 138.825 207.060 ;
        RECT 139.475 206.890 139.645 207.500 ;
        RECT 140.275 207.360 140.445 207.820 ;
        RECT 139.815 207.075 140.445 207.360 ;
        RECT 140.615 206.960 141.175 207.650 ;
        RECT 141.345 207.360 141.565 207.820 ;
        RECT 142.195 207.855 142.825 208.120 ;
        RECT 144.455 208.070 145.485 208.120 ;
        RECT 142.195 207.800 142.365 207.855 ;
        RECT 141.735 207.530 142.365 207.800 ;
        RECT 143.335 207.785 144.285 208.065 ;
        RECT 144.455 207.870 145.085 208.070 ;
        RECT 145.655 207.900 145.825 208.660 ;
        RECT 145.995 208.340 147.125 208.590 ;
        RECT 141.345 207.075 142.025 207.360 ;
        RECT 142.195 207.260 142.365 207.530 ;
        RECT 142.535 207.430 144.655 207.615 ;
        RECT 144.915 207.560 145.085 207.870 ;
        RECT 145.255 207.730 145.825 207.900 ;
        RECT 145.995 207.940 147.125 208.140 ;
        RECT 145.995 207.895 146.325 207.940 ;
        RECT 147.295 207.770 147.465 208.780 ;
        RECT 144.915 207.260 145.825 207.560 ;
        RECT 145.995 207.320 146.275 207.710 ;
        RECT 146.445 207.600 147.465 207.770 ;
        RECT 138.995 206.645 139.645 206.890 ;
        RECT 138.655 206.200 139.280 206.475 ;
        RECT 139.475 206.330 139.645 206.645 ;
        RECT 142.195 206.930 142.865 207.260 ;
        RECT 143.035 207.025 144.365 207.255 ;
        RECT 142.195 206.330 142.365 206.930 ;
        RECT 143.035 206.760 143.205 207.025 ;
        RECT 142.535 206.590 143.205 206.760 ;
        RECT 143.375 206.505 144.025 206.855 ;
        RECT 144.195 206.760 144.365 207.025 ;
        RECT 144.535 207.110 145.825 207.260 ;
        RECT 146.445 207.150 146.615 207.600 ;
        RECT 147.635 207.430 147.805 209.210 ;
        RECT 144.535 206.930 145.085 207.110 ;
        RECT 145.995 206.980 146.615 207.150 ;
        RECT 146.785 207.115 147.805 207.430 ;
        RECT 144.195 206.590 144.655 206.760 ;
        RECT 138.655 205.615 138.825 206.200 ;
        RECT 139.475 206.040 140.370 206.330 ;
        RECT 141.030 206.040 142.365 206.330 ;
        RECT 144.915 206.330 145.085 206.930 ;
        RECT 145.265 206.810 145.825 206.940 ;
        RECT 146.835 206.810 147.465 206.940 ;
        RECT 145.265 206.500 147.465 206.810 ;
        RECT 147.635 206.330 147.805 207.115 ;
        RECT 142.535 206.070 143.205 206.240 ;
        RECT 139.475 206.030 139.645 206.040 ;
        RECT 138.995 205.785 139.645 206.030 ;
        RECT 142.195 205.900 142.365 206.040 ;
        RECT 138.655 205.355 139.280 205.615 ;
        RECT 139.475 205.440 139.645 205.785 ;
        RECT 139.815 205.695 142.025 205.865 ;
        RECT 139.815 205.610 140.385 205.695 ;
        RECT 141.055 205.530 142.025 205.695 ;
        RECT 142.195 205.570 142.865 205.900 ;
        RECT 143.035 205.805 143.205 206.070 ;
        RECT 143.375 205.975 144.025 206.325 ;
        RECT 144.195 206.070 144.655 206.240 ;
        RECT 144.195 205.805 144.365 206.070 ;
        RECT 144.915 206.040 145.810 206.330 ;
        RECT 146.470 206.040 147.805 206.330 ;
        RECT 144.915 205.900 145.085 206.040 ;
        RECT 143.035 205.575 144.365 205.805 ;
        RECT 144.535 205.570 145.085 205.900 ;
        RECT 140.555 205.440 140.885 205.525 ;
        RECT 138.655 204.755 138.825 205.355 ;
        RECT 139.475 205.185 140.045 205.440 ;
        RECT 138.995 205.110 140.045 205.185 ;
        RECT 140.215 205.270 140.885 205.440 ;
        RECT 142.195 205.360 142.365 205.570 ;
        RECT 138.995 204.925 139.645 205.110 ;
        RECT 138.655 204.495 139.280 204.755 ;
        RECT 138.655 203.895 138.825 204.495 ;
        RECT 139.475 204.325 139.645 204.925 ;
        RECT 140.215 204.685 140.385 205.270 ;
        RECT 141.055 205.190 142.365 205.360 ;
        RECT 142.535 205.215 144.655 205.400 ;
        RECT 140.555 205.020 140.885 205.045 ;
        RECT 140.555 204.850 142.025 205.020 ;
        RECT 138.995 204.065 139.645 204.325 ;
        RECT 139.815 204.680 140.385 204.685 ;
        RECT 139.815 204.510 141.685 204.680 ;
        RECT 139.815 204.155 140.180 204.510 ;
        RECT 140.375 204.170 141.345 204.340 ;
        RECT 138.655 203.635 139.280 203.895 ;
        RECT 139.475 203.465 139.645 204.065 ;
        RECT 140.665 203.965 140.835 203.970 ;
        RECT 139.815 203.690 140.975 203.965 ;
        RECT 141.175 203.520 141.345 204.170 ;
        RECT 141.515 203.555 141.685 204.510 ;
        RECT 138.915 203.205 139.645 203.465 ;
        RECT 139.815 203.330 141.345 203.520 ;
        RECT 139.475 203.150 139.645 203.205 ;
        RECT 141.855 203.160 142.025 204.850 ;
        RECT 137.100 202.785 139.295 203.035 ;
        RECT 134.035 202.045 134.205 202.185 ;
        RECT 133.555 201.800 134.205 202.045 ;
        RECT 134.885 202.005 135.185 202.465 ;
        RECT 135.435 202.345 135.695 202.515 ;
        RECT 136.755 202.345 137.735 202.605 ;
        RECT 135.365 202.175 135.695 202.345 ;
        RECT 135.955 202.175 136.925 202.345 ;
        RECT 133.215 201.370 133.840 201.630 ;
        RECT 133.215 200.770 133.385 201.370 ;
        RECT 134.035 201.190 134.205 201.800 ;
        RECT 134.485 201.835 136.585 202.005 ;
        RECT 134.485 201.600 134.655 201.835 ;
        RECT 136.255 201.755 136.585 201.835 ;
        RECT 136.755 201.745 136.925 202.175 ;
        RECT 138.235 202.175 138.485 202.785 ;
        RECT 139.475 202.640 140.180 203.150 ;
        RECT 139.475 202.605 139.645 202.640 ;
        RECT 138.950 202.345 139.645 202.605 ;
        RECT 140.455 202.420 140.625 203.130 ;
        RECT 138.235 202.170 139.295 202.175 ;
        RECT 137.095 201.925 139.295 202.170 ;
        RECT 135.365 201.475 136.085 201.665 ;
        RECT 133.555 200.940 134.205 201.190 ;
        RECT 133.215 200.510 133.840 200.770 ;
        RECT 133.215 199.910 133.385 200.510 ;
        RECT 134.035 200.370 134.205 200.940 ;
        RECT 134.485 200.815 134.655 201.430 ;
        RECT 134.825 201.305 135.155 201.450 ;
        RECT 134.825 200.985 136.115 201.305 ;
        RECT 136.285 200.815 136.455 201.530 ;
        RECT 134.485 200.645 136.455 200.815 ;
        RECT 136.755 201.450 137.735 201.745 ;
        RECT 136.755 200.715 136.925 201.450 ;
        RECT 138.235 201.440 138.795 201.755 ;
        RECT 139.475 201.745 139.645 202.345 ;
        RECT 139.850 202.240 140.625 202.420 ;
        RECT 141.000 202.990 142.025 203.160 ;
        RECT 142.195 204.975 142.365 205.190 ;
        RECT 142.195 204.710 142.825 204.975 ;
        RECT 143.335 204.765 144.285 205.045 ;
        RECT 144.915 204.960 145.085 205.570 ;
        RECT 144.455 204.710 145.085 204.960 ;
        RECT 141.000 202.410 141.190 202.990 ;
        RECT 142.195 202.820 142.365 204.710 ;
        RECT 142.960 204.540 144.325 204.595 ;
        RECT 142.535 204.425 144.635 204.540 ;
        RECT 142.535 204.290 143.090 204.425 ;
        RECT 144.195 204.370 144.635 204.425 ;
        RECT 142.640 203.145 142.810 204.080 ;
        RECT 143.280 204.015 143.875 204.255 ;
        RECT 144.465 204.205 144.635 204.370 ;
        RECT 144.915 204.380 145.085 204.710 ;
        RECT 145.255 204.550 145.885 204.835 ;
        RECT 144.045 203.845 144.265 204.200 ;
        RECT 144.915 204.110 145.545 204.380 ;
        RECT 142.980 203.675 144.265 203.845 ;
        RECT 142.980 203.315 143.345 203.675 ;
        RECT 144.465 203.505 144.635 204.010 ;
        RECT 143.515 203.335 144.635 203.505 ;
        RECT 143.515 203.145 143.685 203.335 ;
        RECT 142.640 202.975 143.685 203.145 ;
        RECT 141.435 202.805 142.365 202.820 ;
        RECT 143.425 202.805 143.685 202.975 ;
        RECT 143.905 202.925 144.235 203.125 ;
        RECT 144.915 203.015 145.085 204.110 ;
        RECT 145.715 204.090 145.885 204.550 ;
        RECT 146.055 204.260 146.615 204.950 ;
        RECT 146.785 204.550 147.465 204.835 ;
        RECT 146.785 204.090 147.005 204.550 ;
        RECT 147.635 204.380 147.805 206.040 ;
        RECT 147.175 204.110 147.805 204.380 ;
        RECT 145.715 203.880 147.005 204.090 ;
        RECT 145.255 203.310 147.465 203.710 ;
        RECT 141.435 202.650 143.165 202.805 ;
        RECT 142.195 202.635 143.165 202.650 ;
        RECT 143.425 202.635 143.755 202.805 ;
        RECT 141.435 202.240 141.845 202.415 ;
        RECT 139.850 202.175 141.845 202.240 ;
        RECT 140.455 201.900 141.845 202.175 ;
        RECT 138.965 201.440 139.645 201.745 ;
        RECT 137.095 200.990 139.305 201.270 ;
        RECT 137.095 200.885 138.065 200.990 ;
        RECT 138.735 200.885 139.305 200.990 ;
        RECT 139.475 201.105 139.645 201.440 ;
        RECT 139.475 200.865 140.155 201.105 ;
        RECT 138.235 200.715 138.565 200.820 ;
        RECT 139.475 200.715 139.645 200.865 ;
        RECT 140.325 200.855 140.885 201.210 ;
        RECT 134.035 200.330 134.735 200.370 ;
        RECT 133.555 200.160 134.735 200.330 ;
        RECT 133.555 200.080 134.205 200.160 ;
        RECT 133.215 199.650 133.840 199.910 ;
        RECT 133.215 199.475 133.385 199.650 ;
        RECT 131.315 199.210 132.215 199.465 ;
        RECT 130.465 198.670 131.145 198.950 ;
        RECT 131.315 198.580 131.485 199.210 ;
        RECT 132.400 199.040 133.385 199.475 ;
        RECT 134.035 199.470 134.205 200.080 ;
        RECT 135.115 199.940 135.445 200.645 ;
        RECT 135.650 199.920 136.025 200.475 ;
        RECT 136.755 200.465 137.385 200.715 ;
        RECT 136.255 200.390 137.385 200.465 ;
        RECT 136.255 200.150 136.925 200.390 ;
        RECT 134.420 199.770 134.945 199.900 ;
        RECT 135.650 199.770 136.585 199.920 ;
        RECT 134.420 199.580 136.585 199.770 ;
        RECT 134.420 199.570 135.445 199.580 ;
        RECT 133.555 199.400 134.205 199.470 ;
        RECT 133.555 199.230 134.815 199.400 ;
        RECT 133.555 199.210 134.205 199.230 ;
        RECT 131.660 198.780 133.840 199.040 ;
        RECT 131.660 198.750 133.385 198.780 ;
        RECT 128.935 198.080 131.145 198.480 ;
        RECT 131.315 198.310 132.230 198.580 ;
        RECT 132.400 198.310 133.385 198.750 ;
        RECT 134.035 198.610 134.205 199.210 ;
        RECT 134.425 198.905 134.945 199.060 ;
        RECT 135.115 199.020 135.445 199.570 ;
        RECT 136.755 199.410 136.925 200.150 ;
        RECT 137.555 200.265 138.845 200.715 ;
        RECT 139.015 200.390 139.645 200.715 ;
        RECT 141.055 200.695 141.400 201.085 ;
        RECT 142.195 200.925 142.365 202.635 ;
        RECT 143.935 202.465 144.235 202.925 ;
        RECT 144.415 202.645 145.085 203.015 ;
        RECT 145.255 202.840 145.885 203.120 ;
        RECT 142.535 202.295 144.635 202.465 ;
        RECT 142.535 202.215 142.865 202.295 ;
        RECT 142.665 201.275 142.835 201.990 ;
        RECT 143.035 201.935 143.755 202.125 ;
        RECT 144.465 202.060 144.635 202.295 ;
        RECT 144.915 202.320 145.085 202.645 ;
        RECT 145.715 202.445 145.885 202.840 ;
        RECT 146.055 202.615 146.615 203.310 ;
        RECT 146.785 202.840 147.465 203.120 ;
        RECT 146.785 202.445 147.005 202.840 ;
        RECT 144.915 201.995 145.545 202.320 ;
        RECT 145.715 201.995 147.005 202.445 ;
        RECT 147.635 202.320 147.805 204.110 ;
        RECT 147.175 201.995 147.805 202.320 ;
        RECT 143.965 201.765 144.295 201.910 ;
        RECT 143.005 201.445 144.295 201.765 ;
        RECT 144.465 201.275 144.635 201.890 ;
        RECT 142.665 201.105 144.635 201.275 ;
        RECT 141.055 200.685 141.225 200.695 ;
        RECT 139.825 200.515 141.225 200.685 ;
        RECT 139.825 200.405 140.155 200.515 ;
        RECT 137.555 199.870 137.775 200.265 ;
        RECT 137.095 199.590 137.775 199.870 ;
        RECT 135.745 199.240 136.925 199.410 ;
        RECT 137.945 199.400 138.505 200.095 ;
        RECT 138.675 199.870 138.845 200.265 ;
        RECT 139.475 200.175 139.645 200.390 ;
        RECT 139.475 199.960 140.155 200.175 ;
        RECT 140.325 200.080 140.885 200.345 ;
        RECT 138.675 199.590 139.305 199.870 ;
        RECT 134.425 198.850 134.985 198.905 ;
        RECT 135.615 198.895 136.540 199.070 ;
        RECT 135.565 198.850 136.540 198.895 ;
        RECT 134.425 198.740 136.540 198.850 ;
        RECT 134.425 198.730 135.695 198.740 ;
        RECT 134.860 198.680 135.695 198.730 ;
        RECT 133.555 198.310 134.205 198.610 ;
        RECT 129.395 197.700 130.685 197.910 ;
        RECT 126.675 197.240 127.965 197.450 ;
        RECT 122.205 196.245 122.535 196.390 ;
        RECT 121.245 195.925 122.535 196.245 ;
        RECT 122.705 195.755 122.875 196.370 ;
        RECT 120.905 195.585 122.875 195.755 ;
        RECT 123.155 196.320 123.820 196.720 ;
        RECT 124.185 196.690 124.715 197.080 ;
        RECT 123.155 195.730 123.325 196.320 ;
        RECT 124.185 196.260 124.565 196.690 ;
        RECT 124.885 196.395 125.195 197.090 ;
        RECT 125.875 197.085 126.505 197.220 ;
        RECT 125.405 196.950 126.505 197.085 ;
        RECT 125.405 196.400 126.045 196.950 ;
        RECT 126.675 196.780 126.895 197.240 ;
        RECT 126.215 196.495 126.895 196.780 ;
        RECT 123.495 196.090 124.015 196.150 ;
        RECT 124.820 196.090 125.605 196.220 ;
        RECT 123.495 195.915 125.605 196.090 ;
        RECT 125.875 196.210 126.045 196.400 ;
        RECT 127.065 196.380 127.625 197.070 ;
        RECT 127.795 196.780 127.965 197.240 ;
        RECT 128.595 197.410 129.225 197.680 ;
        RECT 128.595 197.220 128.765 197.410 ;
        RECT 129.395 197.240 129.565 197.700 ;
        RECT 128.135 196.950 128.765 197.220 ;
        RECT 128.935 196.955 129.565 197.240 ;
        RECT 127.795 196.495 128.425 196.780 ;
        RECT 128.595 196.670 128.765 196.950 ;
        RECT 129.735 196.840 130.295 197.530 ;
        RECT 130.465 197.240 130.685 197.700 ;
        RECT 131.315 197.680 131.485 198.310 ;
        RECT 134.035 198.050 134.205 198.310 ;
        RECT 136.755 198.600 136.925 199.240 ;
        RECT 137.095 199.000 139.305 199.400 ;
        RECT 139.475 198.910 139.645 199.960 ;
        RECT 141.055 199.830 141.225 200.515 ;
        RECT 142.195 200.610 142.865 200.925 ;
        RECT 142.195 200.210 142.365 200.610 ;
        RECT 143.095 200.380 143.470 200.935 ;
        RECT 143.675 200.400 144.005 201.105 ;
        RECT 144.915 200.830 145.085 201.995 ;
        RECT 145.995 201.890 146.325 201.995 ;
        RECT 145.255 201.720 145.825 201.825 ;
        RECT 146.495 201.720 147.465 201.825 ;
        RECT 145.255 201.440 147.465 201.720 ;
        RECT 144.385 200.620 145.085 200.830 ;
        RECT 141.395 199.880 142.365 200.210 ;
        RECT 142.535 200.230 143.470 200.380 ;
        RECT 144.175 200.230 144.700 200.360 ;
        RECT 142.535 200.040 144.700 200.230 ;
        RECT 139.815 199.490 140.385 199.790 ;
        RECT 140.555 199.660 141.225 199.830 ;
        RECT 142.195 199.870 142.365 199.880 ;
        RECT 143.675 200.030 144.700 200.040 ;
        RECT 144.915 200.345 145.085 200.620 ;
        RECT 147.635 200.345 147.805 201.995 ;
        RECT 144.915 200.085 145.925 200.345 ;
        RECT 146.485 200.085 147.805 200.345 ;
        RECT 141.405 199.490 142.025 199.710 ;
        RECT 139.815 199.175 142.025 199.490 ;
        RECT 142.195 199.700 143.375 199.870 ;
        RECT 142.195 198.910 142.365 199.700 ;
        RECT 142.580 199.355 143.505 199.530 ;
        RECT 143.675 199.480 144.005 200.030 ;
        RECT 144.915 199.860 145.085 200.085 ;
        RECT 144.305 199.690 145.085 199.860 ;
        RECT 144.175 199.365 144.695 199.520 ;
        RECT 142.580 199.310 143.555 199.355 ;
        RECT 144.135 199.310 144.695 199.365 ;
        RECT 142.580 199.200 144.695 199.310 ;
        RECT 143.425 199.190 144.695 199.200 ;
        RECT 144.915 199.485 145.085 199.690 ;
        RECT 145.255 199.740 147.465 199.910 ;
        RECT 145.255 199.655 145.830 199.740 ;
        RECT 146.560 199.655 147.465 199.740 ;
        RECT 145.995 199.485 146.325 199.570 ;
        RECT 147.635 199.485 147.805 200.085 ;
        RECT 143.425 199.140 144.260 199.190 ;
        RECT 144.915 199.155 145.465 199.485 ;
        RECT 145.635 199.315 146.705 199.485 ;
        RECT 137.555 198.620 138.845 198.830 ;
        RECT 136.755 198.330 137.385 198.600 ;
        RECT 136.755 198.050 136.925 198.330 ;
        RECT 137.555 198.160 137.775 198.620 ;
        RECT 130.855 197.495 131.485 197.680 ;
        RECT 131.655 197.770 133.865 198.050 ;
        RECT 131.655 197.665 132.625 197.770 ;
        RECT 133.295 197.665 133.865 197.770 ;
        RECT 134.035 197.780 134.840 198.050 ;
        RECT 135.800 197.780 136.925 198.050 ;
        RECT 137.095 197.875 137.775 198.160 ;
        RECT 132.795 197.495 133.125 197.600 ;
        RECT 134.035 197.495 134.205 197.780 ;
        RECT 130.855 197.410 131.945 197.495 ;
        RECT 130.465 196.955 131.145 197.240 ;
        RECT 131.315 197.170 131.945 197.410 ;
        RECT 131.315 196.670 131.485 197.170 ;
        RECT 128.595 196.210 130.055 196.670 ;
        RECT 125.875 195.730 127.135 196.210 ;
        RECT 117.180 195.280 117.885 195.460 ;
        RECT 116.735 194.880 117.510 195.060 ;
        RECT 115.515 194.815 117.510 194.880 ;
        RECT 117.715 194.850 117.885 195.280 ;
        RECT 120.435 195.405 120.605 195.460 ;
        RECT 118.055 195.030 118.605 195.200 ;
        RECT 115.515 194.540 116.905 194.815 ;
        RECT 117.715 194.520 118.265 194.850 ;
        RECT 118.435 194.705 118.605 195.030 ;
        RECT 118.785 194.940 119.155 195.270 ;
        RECT 119.335 195.030 120.265 195.200 ;
        RECT 120.435 195.090 121.105 195.405 ;
        RECT 119.335 194.705 119.505 195.030 ;
        RECT 120.435 194.850 120.605 195.090 ;
        RECT 121.335 194.860 121.710 195.415 ;
        RECT 121.915 194.880 122.245 195.585 ;
        RECT 123.155 195.460 123.960 195.730 ;
        RECT 124.920 195.460 127.135 195.730 ;
        RECT 123.155 195.310 123.325 195.460 ;
        RECT 122.625 195.290 123.325 195.310 ;
        RECT 125.875 195.290 127.135 195.460 ;
        RECT 122.625 195.100 124.615 195.290 ;
        RECT 118.435 194.535 119.505 194.705 ;
        RECT 117.715 193.470 117.885 194.520 ;
        RECT 118.860 194.420 119.190 194.535 ;
        RECT 119.675 194.520 120.605 194.850 ;
        RECT 120.775 194.710 121.710 194.860 ;
        RECT 122.415 194.710 122.940 194.840 ;
        RECT 120.775 194.520 122.940 194.710 ;
        RECT 120.435 194.350 120.605 194.520 ;
        RECT 121.915 194.510 122.940 194.520 ;
        RECT 118.055 194.250 118.560 194.340 ;
        RECT 119.360 194.250 120.265 194.350 ;
        RECT 118.055 194.080 120.265 194.250 ;
        RECT 120.435 194.180 121.615 194.350 ;
        RECT 118.055 193.650 118.605 193.820 ;
        RECT 117.715 193.450 118.265 193.470 ;
        RECT 112.275 193.160 113.170 193.450 ;
        RECT 113.830 193.160 116.330 193.450 ;
        RECT 116.990 193.160 118.265 193.450 ;
        RECT 89.315 191.075 90.525 192.165 ;
        RECT 112.275 191.595 112.445 193.160 ;
        RECT 114.995 192.435 115.165 193.160 ;
        RECT 117.715 193.140 118.265 193.160 ;
        RECT 118.435 193.325 118.605 193.650 ;
        RECT 118.785 193.560 119.155 193.890 ;
        RECT 119.335 193.650 120.265 193.820 ;
        RECT 119.335 193.325 119.505 193.650 ;
        RECT 120.435 193.470 120.605 194.180 ;
        RECT 120.820 193.835 121.745 194.010 ;
        RECT 121.915 193.960 122.245 194.510 ;
        RECT 123.155 194.340 124.615 195.100 ;
        RECT 122.545 194.170 124.615 194.340 ;
        RECT 123.155 194.080 124.615 194.170 ;
        RECT 124.785 194.830 127.135 195.290 ;
        RECT 127.305 196.150 130.055 196.210 ;
        RECT 127.305 195.460 129.515 196.150 ;
        RECT 130.225 195.980 131.485 196.670 ;
        RECT 132.115 197.045 133.405 197.495 ;
        RECT 133.575 197.190 134.205 197.495 ;
        RECT 134.375 197.420 136.485 197.595 ;
        RECT 134.375 197.360 134.895 197.420 ;
        RECT 135.700 197.290 136.485 197.420 ;
        RECT 136.755 197.590 136.925 197.780 ;
        RECT 137.945 197.760 138.505 198.450 ;
        RECT 138.675 198.160 138.845 198.620 ;
        RECT 139.475 198.700 140.465 198.910 ;
        RECT 141.055 198.700 142.365 198.910 ;
        RECT 139.475 198.600 139.645 198.700 ;
        RECT 139.015 198.330 139.645 198.600 ;
        RECT 138.675 197.875 139.305 198.160 ;
        RECT 139.475 198.030 139.645 198.330 ;
        RECT 139.815 198.280 142.025 198.530 ;
        RECT 139.815 198.200 140.445 198.280 ;
        RECT 141.045 198.200 142.025 198.280 ;
        RECT 142.195 198.230 142.365 198.700 ;
        RECT 142.535 198.620 144.745 198.935 ;
        RECT 142.535 198.400 143.155 198.620 ;
        RECT 143.335 198.280 144.005 198.450 ;
        RECT 144.175 198.320 144.745 198.620 ;
        RECT 139.475 197.800 140.465 198.030 ;
        RECT 139.475 197.590 139.645 197.800 ;
        RECT 140.635 197.780 140.885 198.110 ;
        RECT 142.195 198.030 143.165 198.230 ;
        RECT 141.055 197.900 143.165 198.030 ;
        RECT 141.055 197.800 142.365 197.900 ;
        RECT 133.575 197.170 134.700 197.190 ;
        RECT 132.115 196.650 132.335 197.045 ;
        RECT 131.655 196.370 132.335 196.650 ;
        RECT 132.505 196.180 133.065 196.875 ;
        RECT 133.235 196.650 133.405 197.045 ;
        RECT 134.035 196.790 134.700 197.170 ;
        RECT 135.065 196.820 135.445 197.250 ;
        RECT 133.235 196.370 133.865 196.650 ;
        RECT 129.685 195.460 131.485 195.980 ;
        RECT 131.655 195.780 133.865 196.180 ;
        RECT 127.305 195.000 128.765 195.460 ;
        RECT 131.315 195.380 131.485 195.460 ;
        RECT 132.115 195.400 133.405 195.610 ;
        RECT 129.095 195.120 131.145 195.290 ;
        RECT 129.095 195.015 129.440 195.120 ;
        RECT 130.175 195.015 131.145 195.120 ;
        RECT 131.315 195.110 131.945 195.380 ;
        RECT 122.415 193.845 122.935 194.000 ;
        RECT 120.820 193.790 121.795 193.835 ;
        RECT 122.375 193.790 122.935 193.845 ;
        RECT 120.820 193.680 122.935 193.790 ;
        RECT 121.665 193.670 122.935 193.680 ;
        RECT 121.665 193.620 122.500 193.670 ;
        RECT 118.435 193.155 119.505 193.325 ;
        RECT 119.675 193.450 120.605 193.470 ;
        RECT 123.155 193.450 124.095 194.080 ;
        RECT 124.785 193.910 127.655 194.830 ;
        RECT 119.675 193.160 121.770 193.450 ;
        RECT 122.430 193.160 124.095 193.450 ;
        RECT 115.335 192.710 117.545 192.990 ;
        RECT 115.335 192.605 116.305 192.710 ;
        RECT 116.975 192.605 117.545 192.710 ;
        RECT 116.475 192.435 116.805 192.540 ;
        RECT 117.715 192.435 117.885 193.140 ;
        RECT 118.860 193.040 119.190 193.155 ;
        RECT 119.675 193.140 120.605 193.160 ;
        RECT 118.055 192.870 118.560 192.960 ;
        RECT 119.360 192.870 120.265 192.970 ;
        RECT 118.055 192.700 120.265 192.870 ;
        RECT 114.995 192.110 115.625 192.435 ;
        RECT 112.615 191.810 113.165 191.980 ;
        RECT 112.275 191.265 112.825 191.595 ;
        RECT 112.995 191.435 113.165 191.810 ;
        RECT 113.345 191.715 113.715 192.070 ;
        RECT 113.895 191.810 114.825 191.980 ;
        RECT 113.895 191.435 114.065 191.810 ;
        RECT 114.995 191.595 115.165 192.110 ;
        RECT 112.995 191.265 114.065 191.435 ;
        RECT 114.235 191.265 115.165 191.595 ;
        RECT 115.795 191.985 117.085 192.435 ;
        RECT 117.255 192.110 117.885 192.435 ;
        RECT 118.055 192.270 118.605 192.440 ;
        RECT 115.795 191.590 116.015 191.985 ;
        RECT 115.335 191.310 116.015 191.590 ;
        RECT 11.950 190.905 90.610 191.075 ;
        RECT 12.035 189.815 13.245 190.905 ;
        RECT 13.415 190.470 18.760 190.905 ;
        RECT 18.935 190.470 24.280 190.905 ;
        RECT 12.035 189.105 12.555 189.645 ;
        RECT 12.725 189.275 13.245 189.815 ;
        RECT 12.035 188.355 13.245 189.105 ;
        RECT 15.000 188.900 15.340 189.730 ;
        RECT 16.820 189.220 17.170 190.470 ;
        RECT 20.520 188.900 20.860 189.730 ;
        RECT 22.340 189.220 22.690 190.470 ;
        RECT 24.915 189.740 25.205 190.905 ;
        RECT 25.375 190.470 30.720 190.905 ;
        RECT 30.895 190.470 36.240 190.905 ;
        RECT 13.415 188.355 18.760 188.900 ;
        RECT 18.935 188.355 24.280 188.900 ;
        RECT 24.915 188.355 25.205 189.080 ;
        RECT 26.960 188.900 27.300 189.730 ;
        RECT 28.780 189.220 29.130 190.470 ;
        RECT 32.480 188.900 32.820 189.730 ;
        RECT 34.300 189.220 34.650 190.470 ;
        RECT 36.415 189.815 39.925 190.905 ;
        RECT 36.415 189.125 38.065 189.645 ;
        RECT 38.235 189.295 39.925 189.815 ;
        RECT 40.095 190.035 40.370 190.735 ;
        RECT 40.540 190.360 40.795 190.905 ;
        RECT 40.965 190.395 41.445 190.735 ;
        RECT 41.620 190.350 42.225 190.905 ;
        RECT 42.395 190.470 47.740 190.905 ;
        RECT 41.610 190.250 42.225 190.350 ;
        RECT 41.610 190.225 41.795 190.250 ;
        RECT 25.375 188.355 30.720 188.900 ;
        RECT 30.895 188.355 36.240 188.900 ;
        RECT 36.415 188.355 39.925 189.125 ;
        RECT 40.095 189.005 40.265 190.035 ;
        RECT 40.540 189.905 41.295 190.155 ;
        RECT 41.465 189.980 41.795 190.225 ;
        RECT 40.540 189.870 41.310 189.905 ;
        RECT 40.540 189.860 41.325 189.870 ;
        RECT 40.435 189.845 41.330 189.860 ;
        RECT 40.435 189.830 41.350 189.845 ;
        RECT 40.435 189.820 41.370 189.830 ;
        RECT 40.435 189.810 41.395 189.820 ;
        RECT 40.435 189.780 41.465 189.810 ;
        RECT 40.435 189.750 41.485 189.780 ;
        RECT 40.435 189.720 41.505 189.750 ;
        RECT 40.435 189.695 41.535 189.720 ;
        RECT 40.435 189.660 41.570 189.695 ;
        RECT 40.435 189.655 41.600 189.660 ;
        RECT 40.435 189.260 40.665 189.655 ;
        RECT 41.210 189.650 41.600 189.655 ;
        RECT 41.235 189.640 41.600 189.650 ;
        RECT 41.250 189.635 41.600 189.640 ;
        RECT 41.265 189.630 41.600 189.635 ;
        RECT 41.965 189.630 42.225 190.080 ;
        RECT 41.265 189.625 42.225 189.630 ;
        RECT 41.275 189.615 42.225 189.625 ;
        RECT 41.285 189.610 42.225 189.615 ;
        RECT 41.295 189.600 42.225 189.610 ;
        RECT 41.300 189.590 42.225 189.600 ;
        RECT 41.305 189.585 42.225 189.590 ;
        RECT 41.315 189.570 42.225 189.585 ;
        RECT 41.320 189.555 42.225 189.570 ;
        RECT 41.330 189.530 42.225 189.555 ;
        RECT 40.835 189.060 41.165 189.485 ;
        RECT 40.095 188.525 40.355 189.005 ;
        RECT 40.525 188.355 40.775 188.895 ;
        RECT 40.945 188.575 41.165 189.060 ;
        RECT 41.335 189.460 42.225 189.530 ;
        RECT 41.335 188.735 41.505 189.460 ;
        RECT 41.675 188.905 42.225 189.290 ;
        RECT 43.980 188.900 44.320 189.730 ;
        RECT 45.800 189.220 46.150 190.470 ;
        RECT 47.915 189.815 50.505 190.905 ;
        RECT 47.915 189.125 49.125 189.645 ;
        RECT 49.295 189.295 50.505 189.815 ;
        RECT 50.675 189.740 50.965 190.905 ;
        RECT 51.135 189.815 54.645 190.905 ;
        RECT 51.135 189.125 52.785 189.645 ;
        RECT 52.955 189.295 54.645 189.815 ;
        RECT 55.745 190.295 56.075 190.725 ;
        RECT 56.255 190.465 56.450 190.905 ;
        RECT 56.620 190.295 56.950 190.725 ;
        RECT 55.745 190.125 56.950 190.295 ;
        RECT 55.745 189.795 56.640 190.125 ;
        RECT 57.120 189.955 57.395 190.725 ;
        RECT 56.810 189.765 57.395 189.955 ;
        RECT 55.750 189.265 56.045 189.595 ;
        RECT 56.225 189.265 56.640 189.595 ;
        RECT 41.335 188.565 42.225 188.735 ;
        RECT 42.395 188.355 47.740 188.900 ;
        RECT 47.915 188.355 50.505 189.125 ;
        RECT 50.675 188.355 50.965 189.080 ;
        RECT 51.135 188.355 54.645 189.125 ;
        RECT 55.745 188.355 56.045 189.085 ;
        RECT 56.225 188.645 56.455 189.265 ;
        RECT 56.810 189.095 56.985 189.765 ;
        RECT 56.655 188.915 56.985 189.095 ;
        RECT 57.155 188.945 57.395 189.595 ;
        RECT 56.655 188.535 56.880 188.915 ;
        RECT 57.050 188.355 57.380 188.745 ;
        RECT 57.575 188.635 57.855 190.735 ;
        RECT 58.045 190.145 58.830 190.905 ;
        RECT 59.225 190.075 59.610 190.735 ;
        RECT 59.225 189.975 59.635 190.075 ;
        RECT 58.025 189.765 59.635 189.975 ;
        RECT 59.935 189.885 60.135 190.675 ;
        RECT 58.025 189.165 58.300 189.765 ;
        RECT 59.805 189.715 60.135 189.885 ;
        RECT 60.305 189.725 60.625 190.905 ;
        RECT 59.805 189.595 59.985 189.715 ;
        RECT 58.470 189.345 58.825 189.595 ;
        RECT 59.020 189.545 59.485 189.595 ;
        RECT 59.015 189.375 59.485 189.545 ;
        RECT 59.020 189.345 59.485 189.375 ;
        RECT 59.655 189.345 59.985 189.595 ;
        RECT 60.160 189.345 60.625 189.545 ;
        RECT 60.795 189.300 61.075 190.735 ;
        RECT 61.245 190.130 61.955 190.905 ;
        RECT 62.125 189.960 62.455 190.735 ;
        RECT 61.305 189.745 62.455 189.960 ;
        RECT 58.025 188.985 59.275 189.165 ;
        RECT 58.910 188.915 59.275 188.985 ;
        RECT 59.445 188.965 60.625 189.135 ;
        RECT 58.085 188.355 58.255 188.815 ;
        RECT 59.445 188.745 59.775 188.965 ;
        RECT 58.525 188.565 59.775 188.745 ;
        RECT 59.945 188.355 60.115 188.795 ;
        RECT 60.285 188.550 60.625 188.965 ;
        RECT 60.795 188.525 61.135 189.300 ;
        RECT 61.305 189.175 61.590 189.745 ;
        RECT 61.775 189.345 62.245 189.575 ;
        RECT 62.650 189.545 62.865 190.660 ;
        RECT 63.045 190.185 63.375 190.905 ;
        RECT 64.015 190.035 64.290 190.735 ;
        RECT 64.460 190.360 64.715 190.905 ;
        RECT 64.885 190.395 65.365 190.735 ;
        RECT 65.540 190.350 66.145 190.905 ;
        RECT 65.530 190.250 66.145 190.350 ;
        RECT 65.530 190.225 65.715 190.250 ;
        RECT 63.155 189.545 63.385 189.885 ;
        RECT 62.415 189.365 62.865 189.545 ;
        RECT 62.415 189.345 62.745 189.365 ;
        RECT 63.055 189.345 63.385 189.545 ;
        RECT 61.305 188.985 62.015 189.175 ;
        RECT 61.715 188.845 62.015 188.985 ;
        RECT 62.205 188.985 63.385 189.175 ;
        RECT 62.205 188.905 62.535 188.985 ;
        RECT 61.715 188.835 62.030 188.845 ;
        RECT 61.715 188.825 62.040 188.835 ;
        RECT 61.715 188.820 62.050 188.825 ;
        RECT 61.305 188.355 61.475 188.815 ;
        RECT 61.715 188.810 62.055 188.820 ;
        RECT 61.715 188.805 62.060 188.810 ;
        RECT 61.715 188.795 62.065 188.805 ;
        RECT 61.715 188.790 62.070 188.795 ;
        RECT 61.715 188.525 62.075 188.790 ;
        RECT 62.705 188.355 62.875 188.815 ;
        RECT 63.045 188.525 63.385 188.985 ;
        RECT 64.015 189.005 64.185 190.035 ;
        RECT 64.460 189.905 65.215 190.155 ;
        RECT 65.385 189.980 65.715 190.225 ;
        RECT 64.460 189.870 65.230 189.905 ;
        RECT 64.460 189.860 65.245 189.870 ;
        RECT 64.355 189.845 65.250 189.860 ;
        RECT 64.355 189.830 65.270 189.845 ;
        RECT 64.355 189.820 65.290 189.830 ;
        RECT 64.355 189.810 65.315 189.820 ;
        RECT 64.355 189.780 65.385 189.810 ;
        RECT 64.355 189.750 65.405 189.780 ;
        RECT 64.355 189.720 65.425 189.750 ;
        RECT 64.355 189.695 65.455 189.720 ;
        RECT 64.355 189.660 65.490 189.695 ;
        RECT 64.355 189.655 65.520 189.660 ;
        RECT 64.355 189.260 64.585 189.655 ;
        RECT 65.130 189.650 65.520 189.655 ;
        RECT 65.155 189.640 65.520 189.650 ;
        RECT 65.170 189.635 65.520 189.640 ;
        RECT 65.185 189.630 65.520 189.635 ;
        RECT 65.885 189.630 66.145 190.080 ;
        RECT 66.315 189.815 68.905 190.905 ;
        RECT 65.185 189.625 66.145 189.630 ;
        RECT 65.195 189.615 66.145 189.625 ;
        RECT 65.205 189.610 66.145 189.615 ;
        RECT 65.215 189.600 66.145 189.610 ;
        RECT 65.220 189.590 66.145 189.600 ;
        RECT 65.225 189.585 66.145 189.590 ;
        RECT 65.235 189.570 66.145 189.585 ;
        RECT 65.240 189.555 66.145 189.570 ;
        RECT 65.250 189.530 66.145 189.555 ;
        RECT 64.755 189.060 65.085 189.485 ;
        RECT 64.015 188.525 64.275 189.005 ;
        RECT 64.445 188.355 64.695 188.895 ;
        RECT 64.865 188.575 65.085 189.060 ;
        RECT 65.255 189.460 66.145 189.530 ;
        RECT 65.255 188.735 65.425 189.460 ;
        RECT 65.595 188.905 66.145 189.290 ;
        RECT 66.315 189.125 67.525 189.645 ;
        RECT 67.695 189.295 68.905 189.815 ;
        RECT 69.535 189.765 69.815 190.905 ;
        RECT 69.985 189.755 70.315 190.735 ;
        RECT 70.485 189.765 70.745 190.905 ;
        RECT 70.915 190.470 76.260 190.905 ;
        RECT 69.545 189.325 69.880 189.595 ;
        RECT 70.050 189.155 70.220 189.755 ;
        RECT 70.390 189.345 70.725 189.595 ;
        RECT 65.255 188.565 66.145 188.735 ;
        RECT 66.315 188.355 68.905 189.125 ;
        RECT 69.535 188.355 69.845 189.155 ;
        RECT 70.050 188.525 70.745 189.155 ;
        RECT 72.500 188.900 72.840 189.730 ;
        RECT 74.320 189.220 74.670 190.470 ;
        RECT 76.435 189.740 76.725 190.905 ;
        RECT 76.895 190.470 82.240 190.905 ;
        RECT 82.415 190.470 87.760 190.905 ;
        RECT 70.915 188.355 76.260 188.900 ;
        RECT 76.435 188.355 76.725 189.080 ;
        RECT 78.480 188.900 78.820 189.730 ;
        RECT 80.300 189.220 80.650 190.470 ;
        RECT 84.000 188.900 84.340 189.730 ;
        RECT 85.820 189.220 86.170 190.470 ;
        RECT 87.935 189.815 89.145 190.905 ;
        RECT 87.935 189.105 88.455 189.645 ;
        RECT 88.625 189.275 89.145 189.815 ;
        RECT 89.315 189.815 90.525 190.905 ;
        RECT 112.275 190.665 112.445 191.265 ;
        RECT 113.355 191.180 113.685 191.265 ;
        RECT 112.615 191.010 113.190 191.095 ;
        RECT 113.920 191.010 114.825 191.095 ;
        RECT 112.615 190.840 114.825 191.010 ;
        RECT 114.995 190.665 115.165 191.265 ;
        RECT 116.185 191.120 116.745 191.815 ;
        RECT 116.915 191.590 117.085 191.985 ;
        RECT 117.715 192.090 117.885 192.110 ;
        RECT 117.715 191.760 118.265 192.090 ;
        RECT 118.435 191.945 118.605 192.270 ;
        RECT 118.785 192.180 119.155 192.510 ;
        RECT 120.435 192.480 120.605 193.140 ;
        RECT 120.775 192.815 122.985 192.985 ;
        RECT 120.775 192.650 121.745 192.815 ;
        RECT 122.415 192.730 122.985 192.815 ;
        RECT 123.155 192.700 124.095 193.160 ;
        RECT 124.265 193.620 127.655 193.910 ;
        RECT 127.825 194.825 128.765 195.000 ;
        RECT 129.675 194.845 130.005 194.950 ;
        RECT 127.825 194.445 129.165 194.825 ;
        RECT 129.335 194.675 130.345 194.845 ;
        RECT 131.315 194.805 131.485 195.110 ;
        RECT 132.115 194.940 132.335 195.400 ;
        RECT 127.825 193.935 128.765 194.445 ;
        RECT 129.335 194.275 129.505 194.675 ;
        RECT 128.985 194.105 129.505 194.275 ;
        RECT 129.675 194.125 130.005 194.505 ;
        RECT 130.175 194.355 130.345 194.675 ;
        RECT 130.515 194.525 131.485 194.805 ;
        RECT 131.655 194.655 132.335 194.940 ;
        RECT 132.505 194.540 133.065 195.230 ;
        RECT 133.235 194.940 133.405 195.400 ;
        RECT 134.035 195.380 134.205 196.790 ;
        RECT 135.065 196.430 135.595 196.820 ;
        RECT 134.535 196.260 135.595 196.430 ;
        RECT 135.765 196.420 136.075 197.115 ;
        RECT 136.755 197.110 138.015 197.590 ;
        RECT 136.285 196.900 138.015 197.110 ;
        RECT 138.185 197.160 139.645 197.590 ;
        RECT 139.905 197.330 140.365 197.500 ;
        RECT 138.185 197.070 140.025 197.160 ;
        RECT 136.285 196.425 138.555 196.900 ;
        RECT 134.535 196.200 134.730 196.260 ;
        RECT 134.390 196.030 134.730 196.200 ;
        RECT 135.425 196.245 135.595 196.260 ;
        RECT 136.755 196.380 138.555 196.425 ;
        RECT 138.725 196.830 140.025 197.070 ;
        RECT 140.195 197.065 140.365 197.330 ;
        RECT 140.535 197.235 141.185 197.585 ;
        RECT 141.355 197.330 142.025 197.500 ;
        RECT 141.355 197.065 141.525 197.330 ;
        RECT 142.195 197.160 142.365 197.800 ;
        RECT 143.335 197.595 143.505 198.280 ;
        RECT 144.915 198.150 145.085 199.155 ;
        RECT 145.635 198.940 145.805 199.315 ;
        RECT 145.255 198.770 145.805 198.940 ;
        RECT 145.985 198.680 146.355 199.035 ;
        RECT 146.535 198.940 146.705 199.315 ;
        RECT 146.875 199.155 147.805 199.485 ;
        RECT 146.535 198.770 147.465 198.940 ;
        RECT 143.675 197.765 144.235 198.030 ;
        RECT 144.405 197.940 145.085 198.150 ;
        RECT 145.255 198.110 145.885 198.395 ;
        RECT 144.405 197.935 145.545 197.940 ;
        RECT 144.405 197.595 144.735 197.705 ;
        RECT 143.335 197.425 144.735 197.595 ;
        RECT 144.915 197.670 145.545 197.935 ;
        RECT 143.335 197.415 143.505 197.425 ;
        RECT 140.195 196.835 141.525 197.065 ;
        RECT 141.695 196.830 142.365 197.160 ;
        RECT 143.160 197.025 143.505 197.415 ;
        RECT 143.675 196.900 144.235 197.255 ;
        RECT 144.915 197.245 145.085 197.670 ;
        RECT 145.715 197.650 145.885 198.110 ;
        RECT 146.055 197.820 146.615 198.510 ;
        RECT 146.785 198.110 147.465 198.395 ;
        RECT 146.785 197.650 147.005 198.110 ;
        RECT 147.635 197.940 147.805 199.155 ;
        RECT 147.175 197.670 147.805 197.940 ;
        RECT 145.715 197.440 147.005 197.650 ;
        RECT 144.405 197.005 145.085 197.245 ;
        RECT 138.725 196.380 139.645 196.830 ;
        RECT 139.905 196.475 142.025 196.660 ;
        RECT 134.925 195.770 135.255 196.090 ;
        RECT 135.425 195.960 136.540 196.245 ;
        RECT 134.925 195.750 136.135 195.770 ;
        RECT 136.755 195.760 136.925 196.380 ;
        RECT 139.475 196.220 139.645 196.380 ;
        RECT 134.400 195.535 136.135 195.750 ;
        RECT 134.400 195.510 134.775 195.535 ;
        RECT 133.575 195.340 134.205 195.380 ;
        RECT 133.575 195.110 134.710 195.340 ;
        RECT 134.035 195.010 134.710 195.110 ;
        RECT 134.885 195.065 135.735 195.365 ;
        RECT 135.905 195.260 136.135 195.535 ;
        RECT 136.305 195.430 136.925 195.760 ;
        RECT 135.905 195.090 136.565 195.260 ;
        RECT 134.885 195.060 135.055 195.065 ;
        RECT 133.235 194.655 133.865 194.940 ;
        RECT 130.175 194.185 130.635 194.355 ;
        RECT 127.825 193.620 129.165 193.935 ;
        RECT 124.265 193.450 126.045 193.620 ;
        RECT 128.595 193.605 129.165 193.620 ;
        RECT 128.595 193.450 128.765 193.605 ;
        RECT 124.265 193.160 127.210 193.450 ;
        RECT 127.870 193.160 128.765 193.450 ;
        RECT 129.335 193.430 129.505 194.105 ;
        RECT 128.985 193.260 129.505 193.430 ;
        RECT 129.675 193.215 130.295 193.955 ;
        RECT 124.265 192.700 126.045 193.160 ;
        RECT 128.595 193.060 128.765 193.160 ;
        RECT 121.915 192.560 122.245 192.645 ;
        RECT 123.155 192.560 123.325 192.700 ;
        RECT 119.335 192.270 120.265 192.440 ;
        RECT 120.435 192.310 121.745 192.480 ;
        RECT 121.915 192.390 122.585 192.560 ;
        RECT 119.335 191.945 119.505 192.270 ;
        RECT 120.435 192.090 120.605 192.310 ;
        RECT 121.915 192.140 122.245 192.165 ;
        RECT 118.435 191.775 119.505 191.945 ;
        RECT 116.915 191.310 117.545 191.590 ;
        RECT 115.335 190.720 117.545 191.120 ;
        RECT 112.275 190.405 113.285 190.665 ;
        RECT 113.845 190.405 115.165 190.665 ;
        RECT 117.715 190.710 117.885 191.760 ;
        RECT 118.860 191.660 119.190 191.775 ;
        RECT 119.675 191.760 120.605 192.090 ;
        RECT 118.055 191.490 118.560 191.580 ;
        RECT 119.360 191.490 120.265 191.590 ;
        RECT 118.055 191.320 120.265 191.490 ;
        RECT 118.055 190.890 118.605 191.060 ;
        RECT 89.315 189.275 89.835 189.815 ;
        RECT 112.275 189.790 112.445 190.405 ;
        RECT 114.995 190.320 115.165 190.405 ;
        RECT 115.795 190.340 117.085 190.550 ;
        RECT 112.615 190.050 114.825 190.230 ;
        RECT 112.615 189.970 113.120 190.050 ;
        RECT 113.920 189.960 114.825 190.050 ;
        RECT 114.995 190.050 115.625 190.320 ;
        RECT 90.005 189.105 90.525 189.645 ;
        RECT 76.895 188.355 82.240 188.900 ;
        RECT 82.415 188.355 87.760 188.900 ;
        RECT 87.935 188.355 89.145 189.105 ;
        RECT 89.315 188.355 90.525 189.105 ;
        RECT 112.275 189.460 112.825 189.790 ;
        RECT 113.420 189.775 113.750 189.880 ;
        RECT 114.995 189.790 115.165 190.050 ;
        RECT 115.795 189.880 116.015 190.340 ;
        RECT 112.995 189.605 114.065 189.775 ;
        RECT 11.950 188.185 90.610 188.355 ;
        RECT 12.035 187.435 13.245 188.185 ;
        RECT 13.415 187.640 18.760 188.185 ;
        RECT 12.035 186.895 12.555 187.435 ;
        RECT 12.725 186.725 13.245 187.265 ;
        RECT 15.000 186.810 15.340 187.640 ;
        RECT 18.935 187.435 20.145 188.185 ;
        RECT 20.315 187.535 20.575 188.015 ;
        RECT 20.745 187.645 20.995 188.185 ;
        RECT 12.035 185.635 13.245 186.725 ;
        RECT 16.820 186.070 17.170 187.320 ;
        RECT 18.935 186.895 19.455 187.435 ;
        RECT 19.625 186.725 20.145 187.265 ;
        RECT 13.415 185.635 18.760 186.070 ;
        RECT 18.935 185.635 20.145 186.725 ;
        RECT 20.315 186.505 20.485 187.535 ;
        RECT 21.165 187.480 21.385 187.965 ;
        RECT 20.655 186.885 20.885 187.280 ;
        RECT 21.055 187.055 21.385 187.480 ;
        RECT 21.555 187.805 22.445 187.975 ;
        RECT 21.555 187.080 21.725 187.805 ;
        RECT 21.895 187.250 22.445 187.635 ;
        RECT 22.615 187.415 26.125 188.185 ;
        RECT 26.385 187.635 26.555 187.925 ;
        RECT 26.725 187.805 27.055 188.185 ;
        RECT 26.385 187.465 27.050 187.635 ;
        RECT 21.555 187.010 22.445 187.080 ;
        RECT 21.550 186.985 22.445 187.010 ;
        RECT 21.540 186.970 22.445 186.985 ;
        RECT 21.535 186.955 22.445 186.970 ;
        RECT 21.525 186.950 22.445 186.955 ;
        RECT 21.520 186.940 22.445 186.950 ;
        RECT 21.515 186.930 22.445 186.940 ;
        RECT 21.505 186.925 22.445 186.930 ;
        RECT 21.495 186.915 22.445 186.925 ;
        RECT 21.485 186.910 22.445 186.915 ;
        RECT 21.485 186.905 21.820 186.910 ;
        RECT 21.470 186.900 21.820 186.905 ;
        RECT 21.455 186.890 21.820 186.900 ;
        RECT 21.430 186.885 21.820 186.890 ;
        RECT 20.655 186.880 21.820 186.885 ;
        RECT 20.655 186.845 21.790 186.880 ;
        RECT 20.655 186.820 21.755 186.845 ;
        RECT 20.655 186.790 21.725 186.820 ;
        RECT 20.655 186.760 21.705 186.790 ;
        RECT 20.655 186.730 21.685 186.760 ;
        RECT 20.655 186.720 21.615 186.730 ;
        RECT 20.655 186.710 21.590 186.720 ;
        RECT 20.655 186.695 21.570 186.710 ;
        RECT 20.655 186.680 21.550 186.695 ;
        RECT 20.760 186.670 21.545 186.680 ;
        RECT 20.760 186.635 21.530 186.670 ;
        RECT 20.315 185.805 20.590 186.505 ;
        RECT 20.760 186.385 21.515 186.635 ;
        RECT 21.685 186.315 22.015 186.560 ;
        RECT 22.185 186.460 22.445 186.910 ;
        RECT 22.615 186.895 24.265 187.415 ;
        RECT 24.435 186.725 26.125 187.245 ;
        RECT 21.830 186.290 22.015 186.315 ;
        RECT 21.830 186.190 22.445 186.290 ;
        RECT 20.760 185.635 21.015 186.180 ;
        RECT 21.185 185.805 21.665 186.145 ;
        RECT 21.840 185.635 22.445 186.190 ;
        RECT 22.615 185.635 26.125 186.725 ;
        RECT 26.300 186.645 26.650 187.295 ;
        RECT 26.820 186.475 27.050 187.465 ;
        RECT 26.385 186.305 27.050 186.475 ;
        RECT 26.385 185.805 26.555 186.305 ;
        RECT 26.725 185.635 27.055 186.135 ;
        RECT 27.225 185.805 27.410 187.925 ;
        RECT 27.665 187.725 27.915 188.185 ;
        RECT 28.085 187.735 28.420 187.905 ;
        RECT 28.615 187.735 29.290 187.905 ;
        RECT 28.085 187.595 28.255 187.735 ;
        RECT 27.580 186.605 27.860 187.555 ;
        RECT 28.030 187.465 28.255 187.595 ;
        RECT 28.030 186.360 28.200 187.465 ;
        RECT 28.425 187.315 28.950 187.535 ;
        RECT 28.370 186.550 28.610 187.145 ;
        RECT 28.780 186.615 28.950 187.315 ;
        RECT 29.120 186.955 29.290 187.735 ;
        RECT 29.610 187.685 29.980 188.185 ;
        RECT 30.160 187.735 30.565 187.905 ;
        RECT 30.735 187.735 31.520 187.905 ;
        RECT 30.160 187.505 30.330 187.735 ;
        RECT 29.500 187.205 30.330 187.505 ;
        RECT 30.715 187.235 31.180 187.565 ;
        RECT 29.500 187.175 29.700 187.205 ;
        RECT 29.820 186.955 29.990 187.025 ;
        RECT 29.120 186.785 29.990 186.955 ;
        RECT 29.480 186.695 29.990 186.785 ;
        RECT 28.030 186.230 28.335 186.360 ;
        RECT 28.780 186.250 29.310 186.615 ;
        RECT 27.650 185.635 27.915 186.095 ;
        RECT 28.085 185.805 28.335 186.230 ;
        RECT 29.480 186.080 29.650 186.695 ;
        RECT 28.545 185.910 29.650 186.080 ;
        RECT 29.820 185.635 29.990 186.435 ;
        RECT 30.160 186.135 30.330 187.205 ;
        RECT 30.500 186.305 30.690 187.025 ;
        RECT 30.860 186.275 31.180 187.235 ;
        RECT 31.350 187.275 31.520 187.735 ;
        RECT 31.795 187.655 32.005 188.185 ;
        RECT 32.265 187.445 32.595 187.970 ;
        RECT 32.765 187.575 32.935 188.185 ;
        RECT 33.105 187.530 33.435 187.965 ;
        RECT 33.105 187.445 33.485 187.530 ;
        RECT 32.395 187.275 32.595 187.445 ;
        RECT 33.260 187.405 33.485 187.445 ;
        RECT 31.350 186.945 32.225 187.275 ;
        RECT 32.395 186.945 33.145 187.275 ;
        RECT 30.160 185.805 30.410 186.135 ;
        RECT 31.350 186.105 31.520 186.945 ;
        RECT 32.395 186.740 32.585 186.945 ;
        RECT 33.315 186.825 33.485 187.405 ;
        RECT 33.655 187.415 37.165 188.185 ;
        RECT 37.795 187.460 38.085 188.185 ;
        RECT 38.345 187.635 38.515 187.925 ;
        RECT 38.685 187.805 39.015 188.185 ;
        RECT 38.345 187.465 39.010 187.635 ;
        RECT 33.655 186.895 35.305 187.415 ;
        RECT 33.270 186.775 33.485 186.825 ;
        RECT 31.690 186.365 32.585 186.740 ;
        RECT 33.095 186.695 33.485 186.775 ;
        RECT 35.475 186.725 37.165 187.245 ;
        RECT 30.635 185.935 31.520 186.105 ;
        RECT 31.700 185.635 32.015 186.135 ;
        RECT 32.245 185.805 32.585 186.365 ;
        RECT 32.755 185.635 32.925 186.645 ;
        RECT 33.095 185.850 33.425 186.695 ;
        RECT 33.655 185.635 37.165 186.725 ;
        RECT 37.795 185.635 38.085 186.800 ;
        RECT 38.260 186.645 38.610 187.295 ;
        RECT 38.780 186.475 39.010 187.465 ;
        RECT 38.345 186.305 39.010 186.475 ;
        RECT 38.345 185.805 38.515 186.305 ;
        RECT 38.685 185.635 39.015 186.135 ;
        RECT 39.185 185.805 39.370 187.925 ;
        RECT 39.625 187.725 39.875 188.185 ;
        RECT 40.045 187.735 40.380 187.905 ;
        RECT 40.575 187.735 41.250 187.905 ;
        RECT 40.045 187.595 40.215 187.735 ;
        RECT 39.540 186.605 39.820 187.555 ;
        RECT 39.990 187.465 40.215 187.595 ;
        RECT 39.990 186.360 40.160 187.465 ;
        RECT 40.385 187.315 40.910 187.535 ;
        RECT 40.330 186.550 40.570 187.145 ;
        RECT 40.740 186.615 40.910 187.315 ;
        RECT 41.080 186.955 41.250 187.735 ;
        RECT 41.570 187.685 41.940 188.185 ;
        RECT 42.120 187.735 42.525 187.905 ;
        RECT 42.695 187.735 43.480 187.905 ;
        RECT 42.120 187.505 42.290 187.735 ;
        RECT 41.460 187.205 42.290 187.505 ;
        RECT 42.675 187.235 43.140 187.565 ;
        RECT 41.460 187.175 41.660 187.205 ;
        RECT 41.780 186.955 41.950 187.025 ;
        RECT 41.080 186.785 41.950 186.955 ;
        RECT 41.440 186.695 41.950 186.785 ;
        RECT 39.990 186.230 40.295 186.360 ;
        RECT 40.740 186.250 41.270 186.615 ;
        RECT 39.610 185.635 39.875 186.095 ;
        RECT 40.045 185.805 40.295 186.230 ;
        RECT 41.440 186.080 41.610 186.695 ;
        RECT 40.505 185.910 41.610 186.080 ;
        RECT 41.780 185.635 41.950 186.435 ;
        RECT 42.120 186.135 42.290 187.205 ;
        RECT 42.460 186.305 42.650 187.025 ;
        RECT 42.820 186.275 43.140 187.235 ;
        RECT 43.310 187.275 43.480 187.735 ;
        RECT 43.755 187.655 43.965 188.185 ;
        RECT 44.225 187.445 44.555 187.970 ;
        RECT 44.725 187.575 44.895 188.185 ;
        RECT 45.065 187.530 45.395 187.965 ;
        RECT 45.615 187.640 50.960 188.185 ;
        RECT 45.065 187.445 45.445 187.530 ;
        RECT 44.355 187.275 44.555 187.445 ;
        RECT 45.220 187.405 45.445 187.445 ;
        RECT 43.310 186.945 44.185 187.275 ;
        RECT 44.355 186.945 45.105 187.275 ;
        RECT 42.120 185.805 42.370 186.135 ;
        RECT 43.310 186.105 43.480 186.945 ;
        RECT 44.355 186.740 44.545 186.945 ;
        RECT 45.275 186.825 45.445 187.405 ;
        RECT 45.230 186.775 45.445 186.825 ;
        RECT 47.200 186.810 47.540 187.640 ;
        RECT 51.135 187.415 54.645 188.185 ;
        RECT 55.285 187.455 55.585 188.185 ;
        RECT 43.650 186.365 44.545 186.740 ;
        RECT 45.055 186.695 45.445 186.775 ;
        RECT 42.595 185.935 43.480 186.105 ;
        RECT 43.660 185.635 43.975 186.135 ;
        RECT 44.205 185.805 44.545 186.365 ;
        RECT 44.715 185.635 44.885 186.645 ;
        RECT 45.055 185.850 45.385 186.695 ;
        RECT 49.020 186.070 49.370 187.320 ;
        RECT 51.135 186.895 52.785 187.415 ;
        RECT 55.765 187.275 55.995 187.895 ;
        RECT 56.195 187.625 56.420 188.005 ;
        RECT 56.590 187.795 56.920 188.185 ;
        RECT 56.195 187.445 56.525 187.625 ;
        RECT 52.955 186.725 54.645 187.245 ;
        RECT 55.290 186.945 55.585 187.275 ;
        RECT 55.765 186.945 56.180 187.275 ;
        RECT 56.350 186.775 56.525 187.445 ;
        RECT 56.695 186.945 56.935 187.595 ;
        RECT 57.115 187.415 58.785 188.185 ;
        RECT 59.420 187.655 59.710 188.005 ;
        RECT 59.905 187.825 60.235 188.185 ;
        RECT 60.405 187.655 60.635 187.960 ;
        RECT 59.420 187.485 60.635 187.655 ;
        RECT 57.115 186.895 57.865 187.415 ;
        RECT 60.825 187.315 60.995 187.880 ;
        RECT 45.615 185.635 50.960 186.070 ;
        RECT 51.135 185.635 54.645 186.725 ;
        RECT 55.285 186.415 56.180 186.745 ;
        RECT 56.350 186.585 56.935 186.775 ;
        RECT 58.035 186.725 58.785 187.245 ;
        RECT 59.480 187.165 59.740 187.275 ;
        RECT 59.475 186.995 59.740 187.165 ;
        RECT 59.480 186.945 59.740 186.995 ;
        RECT 59.920 186.945 60.305 187.275 ;
        RECT 60.475 187.145 60.995 187.315 ;
        RECT 61.255 187.415 62.925 188.185 ;
        RECT 63.555 187.460 63.845 188.185 ;
        RECT 64.015 187.640 69.360 188.185 ;
        RECT 69.535 187.640 74.880 188.185 ;
        RECT 75.055 187.640 80.400 188.185 ;
        RECT 80.575 187.640 85.920 188.185 ;
        RECT 55.285 186.245 56.490 186.415 ;
        RECT 55.285 185.815 55.615 186.245 ;
        RECT 55.795 185.635 55.990 186.075 ;
        RECT 56.160 185.815 56.490 186.245 ;
        RECT 56.660 185.815 56.935 186.585 ;
        RECT 57.115 185.635 58.785 186.725 ;
        RECT 59.420 185.635 59.740 186.775 ;
        RECT 59.920 185.895 60.115 186.945 ;
        RECT 60.475 186.765 60.645 187.145 ;
        RECT 60.295 186.485 60.645 186.765 ;
        RECT 60.835 186.615 61.080 186.975 ;
        RECT 61.255 186.895 62.005 187.415 ;
        RECT 62.175 186.725 62.925 187.245 ;
        RECT 65.600 186.810 65.940 187.640 ;
        RECT 60.295 185.805 60.625 186.485 ;
        RECT 60.825 185.635 61.080 186.435 ;
        RECT 61.255 185.635 62.925 186.725 ;
        RECT 63.555 185.635 63.845 186.800 ;
        RECT 67.420 186.070 67.770 187.320 ;
        RECT 71.120 186.810 71.460 187.640 ;
        RECT 72.940 186.070 73.290 187.320 ;
        RECT 76.640 186.810 76.980 187.640 ;
        RECT 78.460 186.070 78.810 187.320 ;
        RECT 82.160 186.810 82.500 187.640 ;
        RECT 86.095 187.415 88.685 188.185 ;
        RECT 89.315 187.435 90.525 188.185 ;
        RECT 83.980 186.070 84.330 187.320 ;
        RECT 86.095 186.895 87.305 187.415 ;
        RECT 87.475 186.725 88.685 187.245 ;
        RECT 64.015 185.635 69.360 186.070 ;
        RECT 69.535 185.635 74.880 186.070 ;
        RECT 75.055 185.635 80.400 186.070 ;
        RECT 80.575 185.635 85.920 186.070 ;
        RECT 86.095 185.635 88.685 186.725 ;
        RECT 89.315 186.725 89.835 187.265 ;
        RECT 90.005 186.895 90.525 187.435 ;
        RECT 112.275 187.925 112.445 189.460 ;
        RECT 112.995 189.280 113.165 189.605 ;
        RECT 112.615 189.110 113.165 189.280 ;
        RECT 113.345 189.040 113.715 189.380 ;
        RECT 113.895 189.280 114.065 189.605 ;
        RECT 114.235 189.460 115.165 189.790 ;
        RECT 115.335 189.595 116.015 189.880 ;
        RECT 116.185 189.480 116.745 190.170 ;
        RECT 116.915 189.880 117.085 190.340 ;
        RECT 117.715 190.380 118.265 190.710 ;
        RECT 118.435 190.565 118.605 190.890 ;
        RECT 118.785 190.800 119.155 191.130 ;
        RECT 119.335 190.890 120.265 191.060 ;
        RECT 119.335 190.565 119.505 190.890 ;
        RECT 120.435 190.710 120.605 191.760 ;
        RECT 118.435 190.395 119.505 190.565 ;
        RECT 117.715 190.320 117.885 190.380 ;
        RECT 117.255 190.050 117.885 190.320 ;
        RECT 118.860 190.280 119.190 190.395 ;
        RECT 119.675 190.380 120.605 190.710 ;
        RECT 116.915 189.595 117.545 189.880 ;
        RECT 117.715 189.760 117.885 190.050 ;
        RECT 118.055 190.110 118.560 190.200 ;
        RECT 119.360 190.110 120.265 190.210 ;
        RECT 118.055 189.940 120.265 190.110 ;
        RECT 120.435 189.940 120.605 190.380 ;
        RECT 120.775 191.970 122.245 192.140 ;
        RECT 120.775 190.280 120.945 191.970 ;
        RECT 122.415 191.805 122.585 192.390 ;
        RECT 122.755 192.230 123.325 192.560 ;
        RECT 122.415 191.800 122.985 191.805 ;
        RECT 121.115 191.630 122.985 191.800 ;
        RECT 121.115 190.675 121.285 191.630 ;
        RECT 121.455 191.290 122.425 191.460 ;
        RECT 121.455 190.640 121.625 191.290 ;
        RECT 122.620 191.275 122.985 191.630 ;
        RECT 123.155 191.500 123.325 192.230 ;
        RECT 123.495 191.670 124.125 191.955 ;
        RECT 123.155 191.230 123.785 191.500 ;
        RECT 122.645 191.085 122.815 191.090 ;
        RECT 121.825 190.810 122.985 191.085 ;
        RECT 121.455 190.450 122.985 190.640 ;
        RECT 120.775 190.110 121.800 190.280 ;
        RECT 123.155 190.270 123.325 191.230 ;
        RECT 123.955 191.210 124.125 191.670 ;
        RECT 124.295 191.380 124.855 192.070 ;
        RECT 125.025 191.670 125.705 191.955 ;
        RECT 125.875 191.700 126.045 192.700 ;
        RECT 126.685 192.690 128.025 192.815 ;
        RECT 126.255 192.645 128.025 192.690 ;
        RECT 128.595 192.730 129.265 193.060 ;
        RECT 130.465 193.045 130.635 194.185 ;
        RECT 128.595 192.660 128.765 192.730 ;
        RECT 126.255 192.360 126.855 192.645 ;
        RECT 127.025 192.230 127.685 192.475 ;
        RECT 126.265 191.930 126.855 192.180 ;
        RECT 127.855 192.160 128.025 192.645 ;
        RECT 128.195 192.330 128.765 192.660 ;
        RECT 129.675 192.535 130.005 192.945 ;
        RECT 130.175 192.725 130.635 193.045 ;
        RECT 125.025 191.210 125.245 191.670 ;
        RECT 125.875 191.500 126.515 191.700 ;
        RECT 125.415 191.370 126.515 191.500 ;
        RECT 125.415 191.230 126.045 191.370 ;
        RECT 123.955 191.000 125.245 191.210 ;
        RECT 123.495 190.430 125.705 190.830 ;
        RECT 125.875 190.700 126.045 191.230 ;
        RECT 126.685 191.140 126.855 191.930 ;
        RECT 127.025 191.750 127.685 192.015 ;
        RECT 127.855 191.830 128.365 192.160 ;
        RECT 128.595 192.120 128.765 192.330 ;
        RECT 128.985 192.530 130.005 192.535 ;
        RECT 128.985 192.290 130.600 192.530 ;
        RECT 130.805 192.305 131.095 194.355 ;
        RECT 131.315 193.450 131.485 194.525 ;
        RECT 134.035 193.450 134.205 195.010 ;
        RECT 136.755 194.380 136.925 195.430 ;
        RECT 137.145 194.550 137.435 196.205 ;
        RECT 137.605 195.885 138.065 196.205 ;
        RECT 137.605 194.785 137.775 195.885 ;
        RECT 138.235 195.855 138.805 196.205 ;
        RECT 139.475 196.200 140.105 196.220 ;
        RECT 138.975 195.970 140.105 196.200 ;
        RECT 140.275 196.025 141.225 196.305 ;
        RECT 142.195 196.235 142.365 196.830 ;
        RECT 142.535 196.410 143.465 196.580 ;
        RECT 141.735 196.195 142.365 196.235 ;
        RECT 141.735 195.970 143.125 196.195 ;
        RECT 138.975 195.870 139.645 195.970 ;
        RECT 137.945 194.975 138.565 195.685 ;
        RECT 138.735 195.500 139.255 195.670 ;
        RECT 137.605 194.615 138.065 194.785 ;
        RECT 136.755 194.100 137.725 194.380 ;
        RECT 137.895 194.230 138.065 194.615 ;
        RECT 138.235 194.400 138.565 194.805 ;
        RECT 138.735 194.800 138.905 195.500 ;
        RECT 139.475 195.300 139.645 195.870 ;
        RECT 142.195 195.865 143.125 195.970 ;
        RECT 143.295 196.035 143.465 196.410 ;
        RECT 143.645 196.315 144.015 196.670 ;
        RECT 144.195 196.410 144.745 196.580 ;
        RECT 144.195 196.035 144.365 196.410 ;
        RECT 144.915 196.195 145.085 197.005 ;
        RECT 145.255 196.870 147.465 197.270 ;
        RECT 145.255 196.400 145.885 196.680 ;
        RECT 143.295 195.865 144.365 196.035 ;
        RECT 144.535 195.880 145.085 196.195 ;
        RECT 145.715 196.005 145.885 196.400 ;
        RECT 146.055 196.175 146.615 196.870 ;
        RECT 146.785 196.400 147.465 196.680 ;
        RECT 146.785 196.005 147.005 196.400 ;
        RECT 144.535 195.865 145.545 195.880 ;
        RECT 140.235 195.800 141.600 195.855 ;
        RECT 139.925 195.685 142.025 195.800 ;
        RECT 139.925 195.630 140.365 195.685 ;
        RECT 139.925 195.465 140.095 195.630 ;
        RECT 141.470 195.550 142.025 195.685 ;
        RECT 139.075 194.970 139.645 195.300 ;
        RECT 138.735 194.630 139.255 194.800 ;
        RECT 138.735 194.230 138.905 194.630 ;
        RECT 139.475 194.460 139.645 194.970 ;
        RECT 139.925 194.765 140.095 195.270 ;
        RECT 140.295 195.105 140.515 195.460 ;
        RECT 140.685 195.275 141.280 195.515 ;
        RECT 140.295 194.935 141.580 195.105 ;
        RECT 139.925 194.595 141.045 194.765 ;
        RECT 134.385 193.600 136.585 193.910 ;
        RECT 134.385 193.470 134.945 193.600 ;
        RECT 135.955 193.470 136.585 193.600 ;
        RECT 131.315 193.160 132.650 193.450 ;
        RECT 133.310 193.300 134.205 193.450 ;
        RECT 136.755 193.450 136.925 194.100 ;
        RECT 137.895 194.060 138.905 194.230 ;
        RECT 139.075 194.275 139.645 194.460 ;
        RECT 140.875 194.405 141.045 194.595 ;
        RECT 141.215 194.575 141.580 194.935 ;
        RECT 141.750 194.405 141.920 195.340 ;
        RECT 139.075 194.080 140.145 194.275 ;
        RECT 138.235 193.960 138.565 194.060 ;
        RECT 139.475 193.905 140.145 194.080 ;
        RECT 140.325 194.185 140.655 194.385 ;
        RECT 140.875 194.235 141.920 194.405 ;
        RECT 142.195 195.265 142.365 195.865 ;
        RECT 143.675 195.780 144.005 195.865 ;
        RECT 142.535 195.610 143.440 195.695 ;
        RECT 144.170 195.610 144.745 195.695 ;
        RECT 142.535 195.440 144.745 195.610 ;
        RECT 144.915 195.555 145.545 195.865 ;
        RECT 145.715 195.555 147.005 196.005 ;
        RECT 147.635 195.880 147.805 197.670 ;
        RECT 147.175 195.555 147.805 195.880 ;
        RECT 144.915 195.265 145.085 195.555 ;
        RECT 145.995 195.450 146.325 195.555 ;
        RECT 142.195 195.005 143.515 195.265 ;
        RECT 144.075 195.005 145.085 195.265 ;
        RECT 142.195 194.790 142.365 195.005 ;
        RECT 142.195 194.560 143.505 194.790 ;
        RECT 137.095 193.790 138.065 193.890 ;
        RECT 138.800 193.790 139.145 193.890 ;
        RECT 137.095 193.620 139.145 193.790 ;
        RECT 139.475 193.450 139.645 193.905 ;
        RECT 140.325 193.725 140.625 194.185 ;
        RECT 140.875 194.065 141.135 194.235 ;
        RECT 142.195 194.065 142.365 194.560 ;
        RECT 143.675 194.480 143.925 194.810 ;
        RECT 144.915 194.790 145.085 195.005 ;
        RECT 145.255 195.280 145.825 195.385 ;
        RECT 146.495 195.280 147.465 195.385 ;
        RECT 145.255 195.000 147.465 195.280 ;
        RECT 144.095 194.560 145.085 194.790 ;
        RECT 145.255 194.570 145.805 194.740 ;
        RECT 144.915 194.390 145.085 194.560 ;
        RECT 140.805 193.895 141.135 194.065 ;
        RECT 141.395 193.895 142.365 194.065 ;
        RECT 142.535 194.310 143.515 194.390 ;
        RECT 144.115 194.310 144.745 194.390 ;
        RECT 142.535 194.060 144.745 194.310 ;
        RECT 144.915 194.060 145.465 194.390 ;
        RECT 145.635 194.245 145.805 194.570 ;
        RECT 145.985 194.470 146.355 194.810 ;
        RECT 146.535 194.570 147.465 194.750 ;
        RECT 146.535 194.245 146.705 194.570 ;
        RECT 147.635 194.390 147.805 195.555 ;
        RECT 145.635 194.075 146.705 194.245 ;
        RECT 142.195 193.890 142.365 193.895 ;
        RECT 144.915 193.890 145.085 194.060 ;
        RECT 146.060 193.970 146.390 194.075 ;
        RECT 146.875 194.060 147.805 194.390 ;
        RECT 133.310 193.160 134.945 193.300 ;
        RECT 135.115 193.260 135.735 193.430 ;
        RECT 136.755 193.295 138.090 193.450 ;
        RECT 131.315 192.120 131.485 193.160 ;
        RECT 127.025 191.270 127.685 191.555 ;
        RECT 126.265 190.890 126.855 191.140 ;
        RECT 127.025 190.880 127.685 191.095 ;
        RECT 127.355 190.790 127.685 190.880 ;
        RECT 125.875 190.450 127.185 190.700 ;
        RECT 127.855 190.620 128.025 191.830 ;
        RECT 128.595 191.780 129.265 192.120 ;
        RECT 129.435 191.780 130.005 192.120 ;
        RECT 130.240 191.780 131.485 192.120 ;
        RECT 131.705 191.800 131.995 192.990 ;
        RECT 132.165 192.645 132.625 192.970 ;
        RECT 132.795 192.645 133.125 192.990 ;
        RECT 133.295 192.720 133.815 192.975 ;
        RECT 134.035 192.850 134.945 193.160 ;
        RECT 132.165 191.970 132.335 192.645 ;
        RECT 132.505 192.280 133.125 192.475 ;
        RECT 132.165 191.800 132.625 191.970 ;
        RECT 128.595 191.590 128.765 191.780 ;
        RECT 131.315 191.630 131.485 191.780 ;
        RECT 128.595 191.350 129.575 191.590 ;
        RECT 128.595 190.780 128.765 191.350 ;
        RECT 129.755 191.260 130.005 191.610 ;
        RECT 130.175 191.270 131.130 191.600 ;
        RECT 131.315 191.350 132.285 191.630 ;
        RECT 132.455 191.480 132.625 191.800 ;
        RECT 132.795 191.650 133.125 192.280 ;
        RECT 133.295 192.050 133.465 192.720 ;
        RECT 134.035 192.550 134.205 192.850 ;
        RECT 135.115 192.700 135.395 193.090 ;
        RECT 135.565 192.810 135.735 193.260 ;
        RECT 135.905 193.160 138.090 193.295 ;
        RECT 138.750 193.160 139.645 193.450 ;
        RECT 139.925 193.555 142.025 193.725 ;
        RECT 139.925 193.320 140.095 193.555 ;
        RECT 141.695 193.475 142.025 193.555 ;
        RECT 142.195 193.680 143.505 193.890 ;
        RECT 144.095 193.680 145.085 193.890 ;
        RECT 142.195 193.450 142.365 193.680 ;
        RECT 144.915 193.450 145.085 193.680 ;
        RECT 145.255 193.800 145.760 193.880 ;
        RECT 146.560 193.800 147.465 193.890 ;
        RECT 145.255 193.620 147.465 193.800 ;
        RECT 147.635 193.450 147.805 194.060 ;
        RECT 140.805 193.195 141.525 193.385 ;
        RECT 135.905 192.980 136.925 193.160 ;
        RECT 133.635 192.340 134.205 192.550 ;
        RECT 134.375 192.510 134.945 192.680 ;
        RECT 135.565 192.640 136.585 192.810 ;
        RECT 133.635 192.220 134.605 192.340 ;
        RECT 133.295 191.880 133.815 192.050 ;
        RECT 134.035 191.920 134.605 192.220 ;
        RECT 133.295 191.480 133.465 191.880 ;
        RECT 134.035 191.710 134.205 191.920 ;
        RECT 134.775 191.750 134.945 192.510 ;
        RECT 135.115 192.470 135.445 192.515 ;
        RECT 135.115 192.270 136.245 192.470 ;
        RECT 135.115 191.820 136.245 192.070 ;
        RECT 128.935 191.090 129.575 191.180 ;
        RECT 130.175 191.090 130.345 191.270 ;
        RECT 128.935 190.920 130.345 191.090 ;
        RECT 128.935 190.850 129.575 190.920 ;
        RECT 127.355 190.450 128.025 190.620 ;
        RECT 128.195 190.680 128.765 190.780 ;
        RECT 128.195 190.450 129.575 190.680 ;
        RECT 120.435 189.770 121.365 189.940 ;
        RECT 117.715 189.490 118.695 189.760 ;
        RECT 113.895 189.100 114.825 189.280 ;
        RECT 114.995 188.380 115.165 189.460 ;
        RECT 117.715 188.820 117.885 189.490 ;
        RECT 118.875 189.420 119.125 189.770 ;
        RECT 120.435 189.760 120.605 189.770 ;
        RECT 119.295 189.430 120.605 189.760 ;
        RECT 118.055 189.250 118.695 189.320 ;
        RECT 118.055 189.080 119.465 189.250 ;
        RECT 118.055 188.990 118.695 189.080 ;
        RECT 117.715 188.580 118.695 188.820 ;
        RECT 114.995 188.050 115.885 188.380 ;
        RECT 116.185 188.160 116.725 188.390 ;
        RECT 116.525 188.060 116.725 188.160 ;
        RECT 116.895 188.050 117.545 188.390 ;
        RECT 112.275 187.590 112.950 187.925 ;
        RECT 89.315 185.635 90.525 186.725 ;
        RECT 112.275 186.165 112.445 187.590 ;
        RECT 113.125 187.570 113.975 187.870 ;
        RECT 114.145 187.670 114.805 187.840 ;
        RECT 112.640 187.400 113.015 187.420 ;
        RECT 114.145 187.400 114.375 187.670 ;
        RECT 114.995 187.500 115.165 188.050 ;
        RECT 115.410 187.750 116.705 187.870 ;
        RECT 115.410 187.655 116.725 187.750 ;
        RECT 112.640 187.180 114.375 187.400 ;
        RECT 113.165 187.165 114.375 187.180 ;
        RECT 114.545 187.170 115.165 187.500 ;
        RECT 112.630 186.730 112.970 186.900 ;
        RECT 113.165 186.865 113.495 187.165 ;
        RECT 112.775 186.695 112.970 186.730 ;
        RECT 113.665 186.710 114.780 186.995 ;
        RECT 114.995 186.960 115.165 187.170 ;
        RECT 115.335 187.130 116.325 187.460 ;
        RECT 116.525 187.420 116.725 187.655 ;
        RECT 116.895 187.540 117.085 188.050 ;
        RECT 117.715 187.880 117.885 188.580 ;
        RECT 118.875 188.560 119.125 188.910 ;
        RECT 119.295 188.900 119.465 189.080 ;
        RECT 119.295 188.570 120.250 188.900 ;
        RECT 120.435 188.410 120.605 189.430 ;
        RECT 120.955 189.360 121.365 189.535 ;
        RECT 121.610 189.530 121.800 190.110 ;
        RECT 122.175 189.540 122.345 190.250 ;
        RECT 122.620 189.760 123.325 190.270 ;
        RECT 123.495 189.960 124.125 190.240 ;
        RECT 122.175 189.360 122.950 189.540 ;
        RECT 120.955 189.295 122.950 189.360 ;
        RECT 123.155 189.440 123.325 189.760 ;
        RECT 123.955 189.565 124.125 189.960 ;
        RECT 124.295 189.735 124.855 190.430 ;
        RECT 125.025 189.960 125.705 190.240 ;
        RECT 125.025 189.565 125.245 189.960 ;
        RECT 120.955 189.020 122.345 189.295 ;
        RECT 123.155 189.115 123.785 189.440 ;
        RECT 123.955 189.115 125.245 189.565 ;
        RECT 125.875 189.440 126.045 190.450 ;
        RECT 127.355 190.310 127.685 190.450 ;
        RECT 128.595 190.410 129.575 190.450 ;
        RECT 126.255 190.140 127.105 190.280 ;
        RECT 127.870 190.140 128.380 190.280 ;
        RECT 126.255 189.950 128.380 190.140 ;
        RECT 125.415 189.115 126.045 189.440 ;
        RECT 120.775 188.590 121.705 188.760 ;
        RECT 118.250 188.135 120.265 188.390 ;
        RECT 118.250 188.030 118.625 188.135 ;
        RECT 119.280 188.050 120.265 188.135 ;
        RECT 120.435 188.080 121.365 188.410 ;
        RECT 121.535 188.265 121.705 188.590 ;
        RECT 121.885 188.500 122.255 188.830 ;
        RECT 122.435 188.590 122.985 188.760 ;
        RECT 122.435 188.265 122.605 188.590 ;
        RECT 123.155 188.410 123.325 189.115 ;
        RECT 124.235 189.010 124.565 189.115 ;
        RECT 123.495 188.840 124.065 188.945 ;
        RECT 124.735 188.840 125.705 188.945 ;
        RECT 123.495 188.560 125.705 188.840 ;
        RECT 125.875 188.635 126.045 189.115 ;
        RECT 128.595 189.790 128.765 190.410 ;
        RECT 129.755 190.400 130.005 190.750 ;
        RECT 131.315 190.740 131.485 191.350 ;
        RECT 132.455 191.310 133.465 191.480 ;
        RECT 133.635 191.330 134.205 191.710 ;
        RECT 134.375 191.520 134.945 191.750 ;
        RECT 136.415 191.630 136.585 192.640 ;
        RECT 132.795 191.205 133.125 191.310 ;
        RECT 131.655 191.035 132.625 191.140 ;
        RECT 133.360 191.035 133.705 191.140 ;
        RECT 131.655 190.865 133.705 191.035 ;
        RECT 130.175 190.690 131.485 190.740 ;
        RECT 134.035 190.690 134.205 191.330 ;
        RECT 134.375 191.030 134.945 191.350 ;
        RECT 135.115 191.200 135.445 191.605 ;
        RECT 135.615 191.380 136.585 191.630 ;
        RECT 136.755 192.480 136.925 192.980 ;
        RECT 137.095 192.735 139.110 192.990 ;
        RECT 137.095 192.650 138.080 192.735 ;
        RECT 138.735 192.630 139.110 192.735 ;
        RECT 138.235 192.480 138.565 192.565 ;
        RECT 136.755 192.070 137.355 192.480 ;
        RECT 137.525 192.215 138.565 192.480 ;
        RECT 139.475 192.365 139.645 193.160 ;
        RECT 139.925 192.535 140.095 193.150 ;
        RECT 140.265 193.025 140.595 193.170 ;
        RECT 140.265 192.705 141.555 193.025 ;
        RECT 141.725 192.535 141.895 193.250 ;
        RECT 139.925 192.365 141.895 192.535 ;
        RECT 142.195 193.160 143.530 193.450 ;
        RECT 144.190 193.160 145.810 193.450 ;
        RECT 146.470 193.160 147.805 193.450 ;
        RECT 142.195 192.375 142.365 193.160 ;
        RECT 142.535 192.680 144.735 192.990 ;
        RECT 142.535 192.550 143.165 192.680 ;
        RECT 144.175 192.550 144.735 192.680 ;
        RECT 135.615 191.030 135.785 191.380 ;
        RECT 136.755 191.325 136.925 192.070 ;
        RECT 136.755 191.200 137.345 191.325 ;
        RECT 134.375 190.860 135.785 191.030 ;
        RECT 135.955 190.995 137.345 191.200 ;
        RECT 137.525 191.205 137.695 192.215 ;
        RECT 138.735 192.195 139.645 192.365 ;
        RECT 139.475 192.090 139.645 192.195 ;
        RECT 137.865 191.545 138.035 192.000 ;
        RECT 138.235 191.715 138.565 192.045 ;
        RECT 138.735 191.745 139.110 191.915 ;
        RECT 139.475 191.880 140.175 192.090 ;
        RECT 138.735 191.545 138.905 191.745 ;
        RECT 137.865 191.375 138.905 191.545 ;
        RECT 137.525 191.035 139.305 191.205 ;
        RECT 139.475 191.120 139.645 191.880 ;
        RECT 140.555 191.660 140.885 192.365 ;
        RECT 141.090 191.640 141.465 192.195 ;
        RECT 142.195 192.185 143.215 192.375 ;
        RECT 141.695 192.060 143.215 192.185 ;
        RECT 143.385 192.340 144.005 192.510 ;
        RECT 144.915 192.380 145.085 193.160 ;
        RECT 141.695 191.870 142.365 192.060 ;
        RECT 143.385 191.890 143.555 192.340 ;
        RECT 139.860 191.490 140.385 191.620 ;
        RECT 141.090 191.490 142.025 191.640 ;
        RECT 139.860 191.300 142.025 191.490 ;
        RECT 139.860 191.290 140.885 191.300 ;
        RECT 135.955 190.870 136.925 190.995 ;
        RECT 130.175 190.410 132.575 190.690 ;
        RECT 128.935 189.970 129.485 190.140 ;
        RECT 128.595 189.460 129.145 189.790 ;
        RECT 129.315 189.645 129.485 189.970 ;
        RECT 129.665 189.870 130.035 190.210 ;
        RECT 130.215 189.970 131.145 190.150 ;
        RECT 130.215 189.645 130.385 189.970 ;
        RECT 131.315 189.790 132.575 190.410 ;
        RECT 129.315 189.475 130.385 189.645 ;
        RECT 121.535 188.095 122.605 188.265 ;
        RECT 117.255 187.765 117.885 187.880 ;
        RECT 118.795 187.880 119.125 187.965 ;
        RECT 120.435 187.880 120.605 188.080 ;
        RECT 121.850 187.980 122.180 188.095 ;
        RECT 122.775 188.080 123.325 188.410 ;
        RECT 117.255 187.710 118.625 187.765 ;
        RECT 117.715 187.595 118.625 187.710 ;
        RECT 118.795 187.615 119.835 187.880 ;
        RECT 113.665 186.695 113.835 186.710 ;
        RECT 112.775 186.525 113.835 186.695 ;
        RECT 112.275 185.770 112.940 186.165 ;
        RECT 113.305 186.135 113.835 186.525 ;
        RECT 11.950 185.465 90.610 185.635 ;
        RECT 12.035 184.375 13.245 185.465 ;
        RECT 13.415 184.375 16.005 185.465 ;
        RECT 12.035 183.665 12.555 184.205 ;
        RECT 12.725 183.835 13.245 184.375 ;
        RECT 13.415 183.685 14.625 184.205 ;
        RECT 14.795 183.855 16.005 184.375 ;
        RECT 16.175 184.325 16.455 185.465 ;
        RECT 16.625 184.315 16.955 185.295 ;
        RECT 17.125 184.325 17.385 185.465 ;
        RECT 17.615 184.405 17.945 185.250 ;
        RECT 18.115 184.455 18.285 185.465 ;
        RECT 18.455 184.735 18.795 185.295 ;
        RECT 19.025 184.965 19.340 185.465 ;
        RECT 19.520 184.995 20.405 185.165 ;
        RECT 17.555 184.325 17.945 184.405 ;
        RECT 18.455 184.360 19.350 184.735 ;
        RECT 16.185 183.885 16.520 184.155 ;
        RECT 16.690 183.715 16.860 184.315 ;
        RECT 17.555 184.275 17.770 184.325 ;
        RECT 17.030 183.905 17.365 184.155 ;
        RECT 12.035 182.915 13.245 183.665 ;
        RECT 13.415 182.915 16.005 183.685 ;
        RECT 16.175 182.915 16.485 183.715 ;
        RECT 16.690 183.085 17.385 183.715 ;
        RECT 17.555 183.695 17.725 184.275 ;
        RECT 18.455 184.155 18.645 184.360 ;
        RECT 19.520 184.155 19.690 184.995 ;
        RECT 20.630 184.965 20.880 185.295 ;
        RECT 17.895 183.825 18.645 184.155 ;
        RECT 18.815 183.825 19.690 184.155 ;
        RECT 17.555 183.655 17.780 183.695 ;
        RECT 18.445 183.655 18.645 183.825 ;
        RECT 17.555 183.570 17.935 183.655 ;
        RECT 17.605 183.135 17.935 183.570 ;
        RECT 18.105 182.915 18.275 183.525 ;
        RECT 18.445 183.130 18.775 183.655 ;
        RECT 19.035 182.915 19.245 183.445 ;
        RECT 19.520 183.365 19.690 183.825 ;
        RECT 19.860 183.865 20.180 184.825 ;
        RECT 20.350 184.075 20.540 184.795 ;
        RECT 20.710 183.895 20.880 184.965 ;
        RECT 21.050 184.665 21.220 185.465 ;
        RECT 21.390 185.020 22.495 185.190 ;
        RECT 21.390 184.405 21.560 185.020 ;
        RECT 22.705 184.870 22.955 185.295 ;
        RECT 23.125 185.005 23.390 185.465 ;
        RECT 21.730 184.485 22.260 184.850 ;
        RECT 22.705 184.740 23.010 184.870 ;
        RECT 21.050 184.315 21.560 184.405 ;
        RECT 21.050 184.145 21.920 184.315 ;
        RECT 21.050 184.075 21.220 184.145 ;
        RECT 21.340 183.895 21.540 183.925 ;
        RECT 19.860 183.535 20.325 183.865 ;
        RECT 20.710 183.595 21.540 183.895 ;
        RECT 20.710 183.365 20.880 183.595 ;
        RECT 19.520 183.195 20.305 183.365 ;
        RECT 20.475 183.195 20.880 183.365 ;
        RECT 21.060 182.915 21.430 183.415 ;
        RECT 21.750 183.365 21.920 184.145 ;
        RECT 22.090 183.785 22.260 184.485 ;
        RECT 22.430 183.955 22.670 184.550 ;
        RECT 22.090 183.565 22.615 183.785 ;
        RECT 22.840 183.635 23.010 184.740 ;
        RECT 22.785 183.505 23.010 183.635 ;
        RECT 23.180 183.545 23.460 184.495 ;
        RECT 22.785 183.365 22.955 183.505 ;
        RECT 21.750 183.195 22.425 183.365 ;
        RECT 22.620 183.195 22.955 183.365 ;
        RECT 23.125 182.915 23.375 183.375 ;
        RECT 23.630 183.175 23.815 185.295 ;
        RECT 23.985 184.965 24.315 185.465 ;
        RECT 24.485 184.795 24.655 185.295 ;
        RECT 23.990 184.625 24.655 184.795 ;
        RECT 23.990 183.635 24.220 184.625 ;
        RECT 24.390 183.805 24.740 184.455 ;
        RECT 24.915 184.300 25.205 185.465 ;
        RECT 26.295 184.595 26.570 185.295 ;
        RECT 26.740 184.920 26.995 185.465 ;
        RECT 27.165 184.955 27.645 185.295 ;
        RECT 27.820 184.910 28.425 185.465 ;
        RECT 27.810 184.810 28.425 184.910 ;
        RECT 27.810 184.785 27.995 184.810 ;
        RECT 23.990 183.465 24.655 183.635 ;
        RECT 23.985 182.915 24.315 183.295 ;
        RECT 24.485 183.175 24.655 183.465 ;
        RECT 24.915 182.915 25.205 183.640 ;
        RECT 26.295 183.565 26.465 184.595 ;
        RECT 26.740 184.465 27.495 184.715 ;
        RECT 27.665 184.540 27.995 184.785 ;
        RECT 26.740 184.430 27.510 184.465 ;
        RECT 26.740 184.420 27.525 184.430 ;
        RECT 26.635 184.405 27.530 184.420 ;
        RECT 26.635 184.390 27.550 184.405 ;
        RECT 26.635 184.380 27.570 184.390 ;
        RECT 26.635 184.370 27.595 184.380 ;
        RECT 26.635 184.340 27.665 184.370 ;
        RECT 26.635 184.310 27.685 184.340 ;
        RECT 26.635 184.280 27.705 184.310 ;
        RECT 26.635 184.255 27.735 184.280 ;
        RECT 26.635 184.220 27.770 184.255 ;
        RECT 26.635 184.215 27.800 184.220 ;
        RECT 26.635 183.820 26.865 184.215 ;
        RECT 27.410 184.210 27.800 184.215 ;
        RECT 27.435 184.200 27.800 184.210 ;
        RECT 27.450 184.195 27.800 184.200 ;
        RECT 27.465 184.190 27.800 184.195 ;
        RECT 28.165 184.190 28.425 184.640 ;
        RECT 27.465 184.185 28.425 184.190 ;
        RECT 27.475 184.175 28.425 184.185 ;
        RECT 27.485 184.170 28.425 184.175 ;
        RECT 27.495 184.160 28.425 184.170 ;
        RECT 27.500 184.150 28.425 184.160 ;
        RECT 27.505 184.145 28.425 184.150 ;
        RECT 27.515 184.130 28.425 184.145 ;
        RECT 27.520 184.115 28.425 184.130 ;
        RECT 27.530 184.090 28.425 184.115 ;
        RECT 27.035 183.620 27.365 184.045 ;
        RECT 26.295 183.085 26.555 183.565 ;
        RECT 26.725 182.915 26.975 183.455 ;
        RECT 27.145 183.135 27.365 183.620 ;
        RECT 27.535 184.020 28.425 184.090 ;
        RECT 28.605 184.405 28.935 185.255 ;
        RECT 27.535 183.295 27.705 184.020 ;
        RECT 27.875 183.465 28.425 183.850 ;
        RECT 28.605 183.640 28.795 184.405 ;
        RECT 29.105 184.325 29.355 185.465 ;
        RECT 29.545 184.825 29.795 185.245 ;
        RECT 30.025 184.995 30.355 185.465 ;
        RECT 30.585 184.825 30.835 185.245 ;
        RECT 29.545 184.655 30.835 184.825 ;
        RECT 31.015 184.825 31.345 185.255 ;
        RECT 31.015 184.655 31.470 184.825 ;
        RECT 29.535 184.155 29.750 184.485 ;
        RECT 28.965 183.825 29.275 184.155 ;
        RECT 29.445 183.825 29.750 184.155 ;
        RECT 29.925 183.825 30.210 184.485 ;
        RECT 30.405 183.825 30.670 184.485 ;
        RECT 30.885 183.825 31.130 184.485 ;
        RECT 29.105 183.655 29.275 183.825 ;
        RECT 31.300 183.655 31.470 184.655 ;
        RECT 27.535 183.125 28.425 183.295 ;
        RECT 28.605 183.130 28.935 183.640 ;
        RECT 29.105 183.485 31.470 183.655 ;
        RECT 29.105 182.915 29.435 183.315 ;
        RECT 30.485 183.145 30.815 183.485 ;
        RECT 30.985 182.915 31.315 183.315 ;
        RECT 31.825 183.095 32.085 185.285 ;
        RECT 32.255 184.735 32.595 185.465 ;
        RECT 32.775 184.555 33.045 185.285 ;
        RECT 32.275 184.335 33.045 184.555 ;
        RECT 33.225 184.575 33.455 185.285 ;
        RECT 33.625 184.755 33.955 185.465 ;
        RECT 34.125 184.575 34.385 185.285 ;
        RECT 33.225 184.335 34.385 184.575 ;
        RECT 34.575 184.745 35.035 185.295 ;
        RECT 35.225 184.745 35.555 185.465 ;
        RECT 32.275 183.665 32.565 184.335 ;
        RECT 32.745 183.845 33.210 184.155 ;
        RECT 33.390 183.845 33.915 184.155 ;
        RECT 32.275 183.465 33.505 183.665 ;
        RECT 32.345 182.915 33.015 183.285 ;
        RECT 33.195 183.095 33.505 183.465 ;
        RECT 33.685 183.205 33.915 183.845 ;
        RECT 34.095 183.825 34.395 184.155 ;
        RECT 34.095 182.915 34.385 183.645 ;
        RECT 34.575 183.375 34.825 184.745 ;
        RECT 35.755 184.575 36.055 185.125 ;
        RECT 36.225 184.795 36.505 185.465 ;
        RECT 35.115 184.405 36.055 184.575 ;
        RECT 35.115 184.155 35.285 184.405 ;
        RECT 36.425 184.155 36.690 184.515 ;
        RECT 36.885 184.495 37.215 185.295 ;
        RECT 37.385 184.665 37.615 185.465 ;
        RECT 37.785 184.495 38.115 185.295 ;
        RECT 36.885 184.325 38.115 184.495 ;
        RECT 38.285 184.325 38.540 185.465 ;
        RECT 38.715 184.615 39.095 185.295 ;
        RECT 39.685 184.615 39.855 185.465 ;
        RECT 40.025 184.785 40.355 185.295 ;
        RECT 40.525 184.955 40.695 185.465 ;
        RECT 40.865 184.785 41.265 185.295 ;
        RECT 40.025 184.615 41.265 184.785 ;
        RECT 34.995 183.825 35.285 184.155 ;
        RECT 35.455 183.905 35.795 184.155 ;
        RECT 36.015 183.905 36.690 184.155 ;
        RECT 36.875 183.825 37.185 184.155 ;
        RECT 35.115 183.735 35.285 183.825 ;
        RECT 35.115 183.545 36.505 183.735 ;
        RECT 34.575 183.085 35.135 183.375 ;
        RECT 35.305 182.915 35.555 183.375 ;
        RECT 36.175 183.185 36.505 183.545 ;
        RECT 36.885 183.425 37.215 183.655 ;
        RECT 37.390 183.595 37.765 184.155 ;
        RECT 37.935 183.425 38.115 184.325 ;
        RECT 38.300 183.575 38.520 184.155 ;
        RECT 38.715 183.655 38.885 184.615 ;
        RECT 39.055 184.275 40.360 184.445 ;
        RECT 41.445 184.365 41.765 185.295 ;
        RECT 41.935 184.375 45.445 185.465 ;
        RECT 45.620 185.040 45.955 185.465 ;
        RECT 46.125 184.860 46.310 185.265 ;
        RECT 39.055 183.825 39.300 184.275 ;
        RECT 39.470 183.905 40.020 184.105 ;
        RECT 40.190 184.075 40.360 184.275 ;
        RECT 41.135 184.195 41.765 184.365 ;
        RECT 40.190 183.905 40.565 184.075 ;
        RECT 40.735 183.655 40.965 184.155 ;
        RECT 38.715 183.485 40.965 183.655 ;
        RECT 36.885 183.085 38.115 183.425 ;
        RECT 38.285 182.915 38.540 183.405 ;
        RECT 38.765 182.915 39.095 183.305 ;
        RECT 39.265 183.165 39.435 183.485 ;
        RECT 41.135 183.315 41.305 184.195 ;
        RECT 39.605 182.915 39.935 183.305 ;
        RECT 40.350 183.145 41.305 183.315 ;
        RECT 41.475 182.915 41.765 183.750 ;
        RECT 41.935 183.685 43.585 184.205 ;
        RECT 43.755 183.855 45.445 184.375 ;
        RECT 45.645 184.685 46.310 184.860 ;
        RECT 46.515 184.685 46.845 185.465 ;
        RECT 41.935 182.915 45.445 183.685 ;
        RECT 45.645 183.655 45.985 184.685 ;
        RECT 47.015 184.495 47.285 185.265 ;
        RECT 46.155 184.325 47.285 184.495 ;
        RECT 47.455 184.375 50.045 185.465 ;
        RECT 46.155 183.825 46.405 184.325 ;
        RECT 45.645 183.485 46.330 183.655 ;
        RECT 46.585 183.575 46.945 184.155 ;
        RECT 45.620 182.915 45.955 183.315 ;
        RECT 46.125 183.085 46.330 183.485 ;
        RECT 47.115 183.415 47.285 184.325 ;
        RECT 46.540 182.915 46.815 183.395 ;
        RECT 47.025 183.085 47.285 183.415 ;
        RECT 47.455 183.685 48.665 184.205 ;
        RECT 48.835 183.855 50.045 184.375 ;
        RECT 50.675 184.300 50.965 185.465 ;
        RECT 47.455 182.915 50.045 183.685 ;
        RECT 50.675 182.915 50.965 183.640 ;
        RECT 51.145 183.095 51.405 185.285 ;
        RECT 51.575 184.735 51.915 185.465 ;
        RECT 52.095 184.555 52.365 185.285 ;
        RECT 51.595 184.335 52.365 184.555 ;
        RECT 52.545 184.575 52.775 185.285 ;
        RECT 52.945 184.755 53.275 185.465 ;
        RECT 53.445 184.575 53.705 185.285 ;
        RECT 52.545 184.335 53.705 184.575 ;
        RECT 53.895 184.375 57.405 185.465 ;
        RECT 51.595 183.665 51.885 184.335 ;
        RECT 52.065 183.845 52.530 184.155 ;
        RECT 52.710 183.845 53.235 184.155 ;
        RECT 51.595 183.465 52.825 183.665 ;
        RECT 51.665 182.915 52.335 183.285 ;
        RECT 52.515 183.095 52.825 183.465 ;
        RECT 53.005 183.205 53.235 183.845 ;
        RECT 53.415 183.825 53.715 184.155 ;
        RECT 53.895 183.685 55.545 184.205 ;
        RECT 55.715 183.855 57.405 184.375 ;
        RECT 58.035 184.495 58.325 185.295 ;
        RECT 58.495 184.665 58.730 185.465 ;
        RECT 58.915 185.125 60.450 185.295 ;
        RECT 58.915 184.495 59.245 185.125 ;
        RECT 58.035 184.325 59.245 184.495 ;
        RECT 58.035 183.825 58.280 184.155 ;
        RECT 53.415 182.915 53.705 183.645 ;
        RECT 53.895 182.915 57.405 183.685 ;
        RECT 58.450 183.655 58.620 184.325 ;
        RECT 59.415 184.155 59.650 184.900 ;
        RECT 58.790 183.825 59.190 184.155 ;
        RECT 59.360 183.825 59.650 184.155 ;
        RECT 59.840 184.155 60.110 184.900 ;
        RECT 60.280 184.495 60.450 185.125 ;
        RECT 60.620 184.665 61.025 185.465 ;
        RECT 60.280 184.325 61.025 184.495 ;
        RECT 59.840 183.825 60.180 184.155 ;
        RECT 60.350 183.825 60.685 184.155 ;
        RECT 60.855 183.825 61.025 184.325 ;
        RECT 61.195 183.900 61.545 185.295 ;
        RECT 58.035 183.085 58.620 183.655 ;
        RECT 58.870 183.485 60.265 183.655 ;
        RECT 58.870 183.140 59.200 183.485 ;
        RECT 59.415 182.915 59.790 183.315 ;
        RECT 59.970 183.140 60.265 183.485 ;
        RECT 60.435 182.915 61.105 183.655 ;
        RECT 61.275 183.085 61.545 183.900 ;
        RECT 61.715 184.745 62.175 185.295 ;
        RECT 62.365 184.745 62.695 185.465 ;
        RECT 61.715 183.375 61.965 184.745 ;
        RECT 62.895 184.575 63.195 185.125 ;
        RECT 63.365 184.795 63.645 185.465 ;
        RECT 62.255 184.405 63.195 184.575 ;
        RECT 62.255 184.155 62.425 184.405 ;
        RECT 63.565 184.155 63.830 184.515 ;
        RECT 64.055 184.325 64.285 185.465 ;
        RECT 64.455 184.315 64.785 185.295 ;
        RECT 64.955 184.325 65.165 185.465 ;
        RECT 65.855 184.955 66.115 185.465 ;
        RECT 62.135 183.825 62.425 184.155 ;
        RECT 62.595 183.905 62.935 184.155 ;
        RECT 63.155 183.905 63.830 184.155 ;
        RECT 64.035 183.905 64.365 184.155 ;
        RECT 62.255 183.735 62.425 183.825 ;
        RECT 62.255 183.545 63.645 183.735 ;
        RECT 61.715 183.085 62.275 183.375 ;
        RECT 62.445 182.915 62.695 183.375 ;
        RECT 63.315 183.185 63.645 183.545 ;
        RECT 64.055 182.915 64.285 183.735 ;
        RECT 64.535 183.715 64.785 184.315 ;
        RECT 65.855 183.905 66.195 184.785 ;
        RECT 66.365 184.075 66.535 185.295 ;
        RECT 66.775 184.960 67.390 185.465 ;
        RECT 66.775 184.425 67.025 184.790 ;
        RECT 67.195 184.785 67.390 184.960 ;
        RECT 67.560 184.955 68.035 185.295 ;
        RECT 68.205 184.920 68.420 185.465 ;
        RECT 67.195 184.595 67.525 184.785 ;
        RECT 67.745 184.425 68.460 184.720 ;
        RECT 68.630 184.595 68.905 185.295 ;
        RECT 66.775 184.255 68.565 184.425 ;
        RECT 66.365 183.825 67.160 184.075 ;
        RECT 66.365 183.735 66.615 183.825 ;
        RECT 64.455 183.085 64.785 183.715 ;
        RECT 64.955 182.915 65.165 183.735 ;
        RECT 65.855 182.915 66.115 183.735 ;
        RECT 66.285 183.315 66.615 183.735 ;
        RECT 67.330 183.400 67.585 184.255 ;
        RECT 66.795 183.135 67.585 183.400 ;
        RECT 67.755 183.555 68.165 184.075 ;
        RECT 68.335 183.825 68.565 184.255 ;
        RECT 68.735 183.565 68.905 184.595 ;
        RECT 69.135 184.405 69.465 185.250 ;
        RECT 69.635 184.455 69.805 185.465 ;
        RECT 69.975 184.735 70.315 185.295 ;
        RECT 70.545 184.965 70.860 185.465 ;
        RECT 71.040 184.995 71.925 185.165 ;
        RECT 69.075 184.325 69.465 184.405 ;
        RECT 69.975 184.360 70.870 184.735 ;
        RECT 69.075 184.275 69.290 184.325 ;
        RECT 69.075 183.695 69.245 184.275 ;
        RECT 69.975 184.155 70.165 184.360 ;
        RECT 71.040 184.155 71.210 184.995 ;
        RECT 72.150 184.965 72.400 185.295 ;
        RECT 69.415 183.825 70.165 184.155 ;
        RECT 70.335 183.825 71.210 184.155 ;
        RECT 69.075 183.655 69.300 183.695 ;
        RECT 69.965 183.655 70.165 183.825 ;
        RECT 69.075 183.570 69.455 183.655 ;
        RECT 67.755 183.135 67.955 183.555 ;
        RECT 68.145 182.915 68.475 183.375 ;
        RECT 68.645 183.085 68.905 183.565 ;
        RECT 69.125 183.135 69.455 183.570 ;
        RECT 69.625 182.915 69.795 183.525 ;
        RECT 69.965 183.130 70.295 183.655 ;
        RECT 70.555 182.915 70.765 183.445 ;
        RECT 71.040 183.365 71.210 183.825 ;
        RECT 71.380 183.865 71.700 184.825 ;
        RECT 71.870 184.075 72.060 184.795 ;
        RECT 72.230 183.895 72.400 184.965 ;
        RECT 72.570 184.665 72.740 185.465 ;
        RECT 72.910 185.020 74.015 185.190 ;
        RECT 72.910 184.405 73.080 185.020 ;
        RECT 74.225 184.870 74.475 185.295 ;
        RECT 74.645 185.005 74.910 185.465 ;
        RECT 73.250 184.485 73.780 184.850 ;
        RECT 74.225 184.740 74.530 184.870 ;
        RECT 72.570 184.315 73.080 184.405 ;
        RECT 72.570 184.145 73.440 184.315 ;
        RECT 72.570 184.075 72.740 184.145 ;
        RECT 72.860 183.895 73.060 183.925 ;
        RECT 71.380 183.535 71.845 183.865 ;
        RECT 72.230 183.595 73.060 183.895 ;
        RECT 72.230 183.365 72.400 183.595 ;
        RECT 71.040 183.195 71.825 183.365 ;
        RECT 71.995 183.195 72.400 183.365 ;
        RECT 72.580 182.915 72.950 183.415 ;
        RECT 73.270 183.365 73.440 184.145 ;
        RECT 73.610 183.785 73.780 184.485 ;
        RECT 73.950 183.955 74.190 184.550 ;
        RECT 73.610 183.565 74.135 183.785 ;
        RECT 74.360 183.635 74.530 184.740 ;
        RECT 74.305 183.505 74.530 183.635 ;
        RECT 74.700 183.545 74.980 184.495 ;
        RECT 74.305 183.365 74.475 183.505 ;
        RECT 73.270 183.195 73.945 183.365 ;
        RECT 74.140 183.195 74.475 183.365 ;
        RECT 74.645 182.915 74.895 183.375 ;
        RECT 75.150 183.175 75.335 185.295 ;
        RECT 75.505 184.965 75.835 185.465 ;
        RECT 76.005 184.795 76.175 185.295 ;
        RECT 75.510 184.625 76.175 184.795 ;
        RECT 75.510 183.635 75.740 184.625 ;
        RECT 75.910 183.805 76.260 184.455 ;
        RECT 76.435 184.300 76.725 185.465 ;
        RECT 76.895 185.030 82.240 185.465 ;
        RECT 82.415 185.030 87.760 185.465 ;
        RECT 75.510 183.465 76.175 183.635 ;
        RECT 75.505 182.915 75.835 183.295 ;
        RECT 76.005 183.175 76.175 183.465 ;
        RECT 76.435 182.915 76.725 183.640 ;
        RECT 78.480 183.460 78.820 184.290 ;
        RECT 80.300 183.780 80.650 185.030 ;
        RECT 84.000 183.460 84.340 184.290 ;
        RECT 85.820 183.780 86.170 185.030 ;
        RECT 87.935 184.375 89.145 185.465 ;
        RECT 87.935 183.665 88.455 184.205 ;
        RECT 88.625 183.835 89.145 184.375 ;
        RECT 89.315 184.375 90.525 185.465 ;
        RECT 112.275 184.710 112.445 185.770 ;
        RECT 113.305 185.710 113.685 186.135 ;
        RECT 114.005 185.840 114.315 186.535 ;
        RECT 114.995 186.530 115.940 186.960 ;
        RECT 114.525 186.250 115.940 186.530 ;
        RECT 116.110 186.595 116.325 187.130 ;
        RECT 116.495 186.780 116.725 187.250 ;
        RECT 116.895 187.210 117.165 187.540 ;
        RECT 117.280 187.075 117.545 187.080 ;
        RECT 117.275 187.070 117.545 187.075 ;
        RECT 117.265 187.065 117.545 187.070 ;
        RECT 117.260 187.060 117.545 187.065 ;
        RECT 117.250 187.055 117.545 187.060 ;
        RECT 117.245 187.045 117.545 187.055 ;
        RECT 117.235 187.035 117.545 187.045 ;
        RECT 117.225 187.020 117.545 187.035 ;
        RECT 116.895 186.720 117.545 187.020 ;
        RECT 116.895 186.595 117.085 186.720 ;
        RECT 116.110 186.310 117.085 186.595 ;
        RECT 117.715 186.480 117.885 187.595 ;
        RECT 118.250 187.145 118.625 187.315 ;
        RECT 118.455 186.945 118.625 187.145 ;
        RECT 118.795 187.115 119.125 187.445 ;
        RECT 119.325 186.945 119.495 187.400 ;
        RECT 118.455 186.775 119.495 186.945 ;
        RECT 119.665 186.605 119.835 187.615 ;
        RECT 120.005 187.470 120.605 187.880 ;
        RECT 120.775 187.810 121.680 187.910 ;
        RECT 122.480 187.810 122.985 187.900 ;
        RECT 120.775 187.640 122.985 187.810 ;
        RECT 123.155 187.780 123.325 188.080 ;
        RECT 123.505 188.080 125.705 188.390 ;
        RECT 123.505 187.950 124.065 188.080 ;
        RECT 125.075 187.950 125.705 188.080 ;
        RECT 125.875 188.305 127.145 188.635 ;
        RECT 120.435 186.990 120.605 187.470 ;
        RECT 120.775 187.300 122.825 187.470 ;
        RECT 120.775 187.200 121.745 187.300 ;
        RECT 122.480 187.200 122.825 187.300 ;
        RECT 123.155 187.330 124.065 187.780 ;
        RECT 124.235 187.740 124.855 187.910 ;
        RECT 125.875 187.775 126.045 188.305 ;
        RECT 127.395 188.205 127.605 188.850 ;
        RECT 127.775 188.365 128.410 188.695 ;
        RECT 121.915 187.030 122.245 187.130 ;
        RECT 120.435 186.725 121.405 186.990 ;
        RECT 117.255 186.310 117.885 186.480 ;
        RECT 118.055 186.435 119.835 186.605 ;
        RECT 114.525 185.845 115.165 186.250 ;
        RECT 116.770 186.080 117.545 186.140 ;
        RECT 112.615 185.535 113.135 185.600 ;
        RECT 113.940 185.535 114.725 185.665 ;
        RECT 112.615 185.360 114.725 185.535 ;
        RECT 114.995 184.710 115.165 185.845 ;
        RECT 115.335 185.800 117.545 186.080 ;
        RECT 117.715 185.705 117.885 186.310 ;
        RECT 118.055 185.875 118.705 186.205 ;
        RECT 117.715 185.535 118.355 185.705 ;
        RECT 117.715 184.710 117.885 185.535 ;
        RECT 118.535 185.365 118.705 185.875 ;
        RECT 118.875 185.695 119.085 186.265 ;
        RECT 119.255 186.225 119.835 186.435 ;
        RECT 120.015 186.710 121.405 186.725 ;
        RECT 121.575 186.860 122.585 187.030 ;
        RECT 123.155 187.010 123.325 187.330 ;
        RECT 124.235 187.180 124.515 187.570 ;
        RECT 124.685 187.290 124.855 187.740 ;
        RECT 125.025 187.460 126.045 187.775 ;
        RECT 126.215 187.505 127.225 187.830 ;
        RECT 125.875 187.335 126.045 187.460 ;
        RECT 120.015 186.395 120.605 186.710 ;
        RECT 119.255 185.900 120.265 186.225 ;
        RECT 118.070 185.035 118.705 185.365 ;
        RECT 118.875 184.880 119.085 185.525 ;
        RECT 120.435 185.425 120.605 186.395 ;
        RECT 119.335 185.095 120.605 185.425 ;
        RECT 120.435 184.710 120.605 185.095 ;
        RECT 120.825 184.885 121.115 186.540 ;
        RECT 121.575 186.475 121.745 186.860 ;
        RECT 121.285 186.305 121.745 186.475 ;
        RECT 121.285 185.205 121.455 186.305 ;
        RECT 121.915 186.285 122.245 186.690 ;
        RECT 122.415 186.460 122.585 186.860 ;
        RECT 122.755 186.820 123.325 187.010 ;
        RECT 123.495 186.990 124.065 187.160 ;
        RECT 124.685 187.120 125.705 187.290 ;
        RECT 122.755 186.630 123.725 186.820 ;
        RECT 122.415 186.290 122.935 186.460 ;
        RECT 123.155 186.400 123.725 186.630 ;
        RECT 121.625 185.405 122.245 186.115 ;
        RECT 122.415 185.590 122.585 186.290 ;
        RECT 123.155 186.120 123.325 186.400 ;
        RECT 123.895 186.230 124.065 186.990 ;
        RECT 124.235 186.950 124.565 186.995 ;
        RECT 124.235 186.750 125.365 186.950 ;
        RECT 124.235 186.300 125.365 186.550 ;
        RECT 122.755 185.790 123.325 186.120 ;
        RECT 123.495 186.000 124.065 186.230 ;
        RECT 125.535 186.110 125.705 187.120 ;
        RECT 122.415 185.420 122.935 185.590 ;
        RECT 121.285 184.885 121.745 185.205 ;
        RECT 121.915 184.885 122.485 185.235 ;
        RECT 123.155 185.220 123.325 185.790 ;
        RECT 123.495 185.510 124.065 185.830 ;
        RECT 124.235 185.680 124.565 186.085 ;
        RECT 124.735 185.860 125.705 186.110 ;
        RECT 125.875 187.005 126.465 187.335 ;
        RECT 126.645 187.295 127.225 187.505 ;
        RECT 127.395 187.465 127.605 188.035 ;
        RECT 127.775 187.855 127.945 188.365 ;
        RECT 128.595 188.195 128.765 189.460 ;
        RECT 129.740 189.370 130.070 189.475 ;
        RECT 130.555 189.460 132.575 189.790 ;
        RECT 132.745 190.670 134.205 190.690 ;
        RECT 132.745 190.430 135.015 190.670 ;
        RECT 132.745 189.760 134.205 190.430 ;
        RECT 135.195 190.340 135.445 190.690 ;
        RECT 135.615 190.350 136.570 190.680 ;
        RECT 134.375 190.170 135.015 190.260 ;
        RECT 135.615 190.170 135.785 190.350 ;
        RECT 134.375 190.000 135.785 190.170 ;
        RECT 136.755 190.025 136.925 190.870 ;
        RECT 137.525 190.825 138.105 191.035 ;
        RECT 139.475 190.950 140.255 191.120 ;
        RECT 137.095 190.500 138.105 190.825 ;
        RECT 138.275 190.295 138.485 190.865 ;
        RECT 138.655 190.475 139.305 190.805 ;
        RECT 134.375 189.930 135.015 190.000 ;
        RECT 132.745 189.490 135.015 189.760 ;
        RECT 132.745 189.480 134.205 189.490 ;
        RECT 135.195 189.480 135.445 189.830 ;
        RECT 136.755 189.820 138.025 190.025 ;
        RECT 135.615 189.695 138.025 189.820 ;
        RECT 135.615 189.490 136.925 189.695 ;
        RECT 131.315 189.310 132.575 189.460 ;
        RECT 128.935 189.200 129.440 189.280 ;
        RECT 130.240 189.200 131.145 189.290 ;
        RECT 128.935 189.020 131.145 189.200 ;
        RECT 128.950 188.365 129.585 188.695 ;
        RECT 128.125 188.025 129.235 188.195 ;
        RECT 127.775 187.525 128.425 187.855 ;
        RECT 126.645 187.125 128.425 187.295 ;
        RECT 125.875 186.260 126.045 187.005 ;
        RECT 124.735 185.510 124.905 185.860 ;
        RECT 125.875 185.850 126.475 186.260 ;
        RECT 126.645 186.115 126.815 187.125 ;
        RECT 126.985 186.785 128.025 186.955 ;
        RECT 126.985 186.330 127.155 186.785 ;
        RECT 127.355 186.285 127.685 186.615 ;
        RECT 127.855 186.585 128.025 186.785 ;
        RECT 127.855 186.415 128.230 186.585 ;
        RECT 128.595 186.135 128.765 188.025 ;
        RECT 129.415 187.855 129.585 188.365 ;
        RECT 129.755 188.205 129.965 188.850 ;
        RECT 131.315 188.635 133.095 189.310 ;
        RECT 130.215 188.305 133.095 188.635 ;
        RECT 131.315 188.100 133.095 188.305 ;
        RECT 133.265 188.225 134.205 189.480 ;
        RECT 134.570 188.595 136.585 188.850 ;
        RECT 134.570 188.490 134.945 188.595 ;
        RECT 135.600 188.510 136.585 188.595 ;
        RECT 136.755 188.800 136.925 189.490 ;
        RECT 138.275 189.480 138.485 190.125 ;
        RECT 138.655 189.965 138.825 190.475 ;
        RECT 139.475 190.305 139.645 190.950 ;
        RECT 139.865 190.625 140.385 190.780 ;
        RECT 140.555 190.740 140.885 191.290 ;
        RECT 142.195 191.130 142.365 191.870 ;
        RECT 141.185 190.960 142.365 191.130 ;
        RECT 139.865 190.570 140.425 190.625 ;
        RECT 141.055 190.615 141.980 190.790 ;
        RECT 141.005 190.570 141.980 190.615 ;
        RECT 139.865 190.460 141.980 190.570 ;
        RECT 139.865 190.450 141.135 190.460 ;
        RECT 140.300 190.400 141.135 190.450 ;
        RECT 139.005 190.135 139.645 190.305 ;
        RECT 138.655 189.635 139.290 189.965 ;
        RECT 139.475 189.605 139.645 190.135 ;
        RECT 142.195 190.280 142.365 190.960 ;
        RECT 142.535 191.720 143.555 191.890 ;
        RECT 143.725 191.780 144.005 192.170 ;
        RECT 144.175 192.065 145.085 192.380 ;
        RECT 147.635 192.065 147.805 193.160 ;
        RECT 144.175 191.930 145.925 192.065 ;
        RECT 144.915 191.805 145.925 191.930 ;
        RECT 146.485 191.805 147.805 192.065 ;
        RECT 142.535 190.710 142.705 191.720 ;
        RECT 143.675 191.550 144.005 191.595 ;
        RECT 142.875 191.350 144.005 191.550 ;
        RECT 144.175 191.590 144.745 191.760 ;
        RECT 142.875 190.900 144.005 191.150 ;
        RECT 144.175 190.830 144.345 191.590 ;
        RECT 144.915 191.420 145.085 191.805 ;
        RECT 144.515 191.205 145.085 191.420 ;
        RECT 145.255 191.460 147.465 191.630 ;
        RECT 145.255 191.375 145.830 191.460 ;
        RECT 146.560 191.375 147.465 191.460 ;
        RECT 145.995 191.205 146.325 191.290 ;
        RECT 147.635 191.205 147.805 191.805 ;
        RECT 144.515 191.000 145.465 191.205 ;
        RECT 144.915 190.875 145.465 191.000 ;
        RECT 145.635 191.035 146.705 191.205 ;
        RECT 142.535 190.460 143.505 190.710 ;
        RECT 142.195 189.950 143.165 190.280 ;
        RECT 143.335 190.110 143.505 190.460 ;
        RECT 143.675 190.280 144.005 190.685 ;
        RECT 144.175 190.600 144.745 190.830 ;
        RECT 144.175 190.110 144.745 190.430 ;
        RECT 139.475 189.365 140.155 189.605 ;
        RECT 137.095 189.055 139.110 189.310 ;
        RECT 137.095 188.970 138.080 189.055 ;
        RECT 138.735 188.950 139.110 189.055 ;
        RECT 138.235 188.800 138.565 188.885 ;
        RECT 135.115 188.340 135.445 188.425 ;
        RECT 136.755 188.390 137.355 188.800 ;
        RECT 137.525 188.535 138.565 188.800 ;
        RECT 139.475 188.685 139.645 189.365 ;
        RECT 140.325 189.355 140.885 189.710 ;
        RECT 141.055 189.195 141.400 189.585 ;
        RECT 142.195 189.200 142.365 189.950 ;
        RECT 143.335 189.940 144.745 190.110 ;
        RECT 144.915 190.230 145.085 190.875 ;
        RECT 145.635 190.660 145.805 191.035 ;
        RECT 145.255 190.490 145.805 190.660 ;
        RECT 145.985 190.400 146.355 190.755 ;
        RECT 146.535 190.660 146.705 191.035 ;
        RECT 146.875 190.875 147.805 191.205 ;
        RECT 146.535 190.490 147.465 190.660 ;
        RECT 147.635 190.230 147.805 190.875 ;
        RECT 142.535 189.370 143.215 189.655 ;
        RECT 141.055 189.185 141.225 189.195 ;
        RECT 139.825 189.015 141.225 189.185 ;
        RECT 139.825 188.905 140.155 189.015 ;
        RECT 138.735 188.675 139.645 188.685 ;
        RECT 136.755 188.340 136.925 188.390 ;
        RECT 133.265 188.100 134.945 188.225 ;
        RECT 128.935 187.525 129.585 187.855 ;
        RECT 129.755 187.465 129.965 188.035 ;
        RECT 130.135 187.505 131.145 187.830 ;
        RECT 130.135 187.295 130.715 187.505 ;
        RECT 131.315 187.460 131.485 188.100 ;
        RECT 134.035 188.055 134.945 188.100 ;
        RECT 135.115 188.075 136.155 188.340 ;
        RECT 131.315 187.335 132.625 187.460 ;
        RECT 128.935 187.125 130.715 187.295 ;
        RECT 129.335 186.785 130.375 186.955 ;
        RECT 129.335 186.585 129.505 186.785 ;
        RECT 129.130 186.415 129.505 186.585 ;
        RECT 129.675 186.285 130.005 186.615 ;
        RECT 130.205 186.330 130.375 186.785 ;
        RECT 126.645 185.850 127.685 186.115 ;
        RECT 127.855 185.965 129.505 186.135 ;
        RECT 130.545 186.115 130.715 187.125 ;
        RECT 130.895 187.130 132.625 187.335 ;
        RECT 130.895 187.005 131.485 187.130 ;
        RECT 132.795 187.120 133.045 187.470 ;
        RECT 134.035 187.460 134.205 188.055 ;
        RECT 134.570 187.605 134.945 187.775 ;
        RECT 133.225 187.190 134.205 187.460 ;
        RECT 134.775 187.405 134.945 187.605 ;
        RECT 135.115 187.575 135.445 187.905 ;
        RECT 135.645 187.405 135.815 187.860 ;
        RECT 134.775 187.235 135.815 187.405 ;
        RECT 131.315 186.260 131.485 187.005 ;
        RECT 133.225 186.950 133.865 187.020 ;
        RECT 132.455 186.780 133.865 186.950 ;
        RECT 132.455 186.600 132.625 186.780 ;
        RECT 133.225 186.690 133.865 186.780 ;
        RECT 131.670 186.270 132.625 186.600 ;
        RECT 132.795 186.260 133.045 186.610 ;
        RECT 134.035 186.520 134.205 187.190 ;
        RECT 135.985 187.065 136.155 188.075 ;
        RECT 136.325 187.930 136.925 188.340 ;
        RECT 136.755 187.645 136.925 187.930 ;
        RECT 136.755 187.315 137.345 187.645 ;
        RECT 137.525 187.525 137.695 188.535 ;
        RECT 138.735 188.515 140.155 188.675 ;
        RECT 140.325 188.580 140.885 188.845 ;
        RECT 139.475 188.460 140.155 188.515 ;
        RECT 137.865 187.865 138.035 188.320 ;
        RECT 138.235 188.035 138.565 188.365 ;
        RECT 138.735 188.065 139.110 188.235 ;
        RECT 138.735 187.865 138.905 188.065 ;
        RECT 137.865 187.695 138.905 187.865 ;
        RECT 137.525 187.355 139.305 187.525 ;
        RECT 136.755 187.185 136.925 187.315 ;
        RECT 134.375 186.895 136.155 187.065 ;
        RECT 133.225 186.280 134.205 186.520 ;
        RECT 134.375 186.335 135.025 186.665 ;
        RECT 125.875 185.680 126.045 185.850 ;
        RECT 127.355 185.765 127.685 185.850 ;
        RECT 123.495 185.340 124.905 185.510 ;
        RECT 125.075 185.350 126.045 185.680 ;
        RECT 122.655 184.890 123.325 185.220 ;
        RECT 123.155 184.710 123.325 184.890 ;
        RECT 125.875 184.710 126.045 185.350 ;
        RECT 126.215 185.595 127.200 185.680 ;
        RECT 127.855 185.595 128.230 185.700 ;
        RECT 126.215 185.570 128.230 185.595 ;
        RECT 126.215 185.400 128.255 185.570 ;
        RECT 126.215 185.340 128.230 185.400 ;
        RECT 128.595 184.710 128.765 185.965 ;
        RECT 129.675 185.850 130.715 186.115 ;
        RECT 130.885 185.850 131.485 186.260 ;
        RECT 134.035 186.165 134.205 186.280 ;
        RECT 129.675 185.765 130.005 185.850 ;
        RECT 129.130 185.595 129.505 185.700 ;
        RECT 130.160 185.595 131.145 185.680 ;
        RECT 129.130 185.340 131.145 185.595 ;
        RECT 131.315 185.650 131.485 185.850 ;
        RECT 131.655 185.920 133.865 186.090 ;
        RECT 131.655 185.820 132.560 185.920 ;
        RECT 133.360 185.830 133.865 185.920 ;
        RECT 134.035 185.995 134.675 186.165 ;
        RECT 131.315 185.320 132.245 185.650 ;
        RECT 132.730 185.635 133.060 185.750 ;
        RECT 134.035 185.650 134.205 185.995 ;
        RECT 134.855 185.825 135.025 186.335 ;
        RECT 135.195 186.155 135.405 186.725 ;
        RECT 135.575 186.685 136.155 186.895 ;
        RECT 136.335 186.855 136.925 187.185 ;
        RECT 137.525 187.145 138.105 187.355 ;
        RECT 135.575 186.360 136.585 186.685 ;
        RECT 136.755 186.345 136.925 186.855 ;
        RECT 137.095 186.820 138.105 187.145 ;
        RECT 138.275 186.615 138.485 187.185 ;
        RECT 138.655 186.795 139.305 187.125 ;
        RECT 139.475 187.030 139.645 188.460 ;
        RECT 141.055 188.330 141.225 189.015 ;
        RECT 142.195 188.930 142.825 189.200 ;
        RECT 142.195 188.710 142.365 188.930 ;
        RECT 141.395 188.380 142.365 188.710 ;
        RECT 142.995 188.910 143.215 189.370 ;
        RECT 143.385 189.080 143.945 189.770 ;
        RECT 144.915 189.710 146.375 190.230 ;
        RECT 144.115 189.370 144.745 189.655 ;
        RECT 144.115 188.910 144.285 189.370 ;
        RECT 144.915 189.200 145.835 189.710 ;
        RECT 146.545 189.540 147.805 190.230 ;
        RECT 144.455 189.020 145.835 189.200 ;
        RECT 146.005 189.020 147.805 189.540 ;
        RECT 144.455 188.930 145.085 189.020 ;
        RECT 142.995 188.700 144.285 188.910 ;
        RECT 139.815 187.990 140.385 188.290 ;
        RECT 140.555 188.160 141.225 188.330 ;
        RECT 141.405 187.990 142.025 188.210 ;
        RECT 139.815 187.675 142.025 187.990 ;
        RECT 139.815 187.210 140.365 187.380 ;
        RECT 136.755 186.015 138.025 186.345 ;
        RECT 132.415 185.465 133.485 185.635 ;
        RECT 131.315 184.710 131.485 185.320 ;
        RECT 132.415 185.140 132.585 185.465 ;
        RECT 131.655 184.970 132.585 185.140 ;
        RECT 132.765 184.900 133.135 185.230 ;
        RECT 133.315 185.140 133.485 185.465 ;
        RECT 133.655 185.320 134.205 185.650 ;
        RECT 134.390 185.495 135.025 185.825 ;
        RECT 135.195 185.340 135.405 185.985 ;
        RECT 136.755 185.885 136.925 186.015 ;
        RECT 135.655 185.555 136.925 185.885 ;
        RECT 138.275 185.800 138.485 186.445 ;
        RECT 138.655 186.285 138.825 186.795 ;
        RECT 139.475 186.700 140.025 187.030 ;
        RECT 140.195 186.885 140.365 187.210 ;
        RECT 140.545 187.120 140.915 187.450 ;
        RECT 141.095 187.210 142.025 187.380 ;
        RECT 141.095 186.885 141.265 187.210 ;
        RECT 142.195 187.140 142.365 188.380 ;
        RECT 142.535 188.130 144.745 188.530 ;
        RECT 144.915 188.410 145.085 188.930 ;
        RECT 145.255 188.680 147.465 188.850 ;
        RECT 145.255 188.590 145.760 188.680 ;
        RECT 146.560 188.580 147.465 188.680 ;
        RECT 142.535 187.660 143.215 187.940 ;
        RECT 142.995 187.265 143.215 187.660 ;
        RECT 143.385 187.435 143.945 188.130 ;
        RECT 144.915 188.080 145.465 188.410 ;
        RECT 146.060 188.395 146.390 188.510 ;
        RECT 147.635 188.410 147.805 189.020 ;
        RECT 145.635 188.225 146.705 188.395 ;
        RECT 144.115 187.660 144.745 187.940 ;
        RECT 144.115 187.265 144.285 187.660 ;
        RECT 142.195 187.030 142.825 187.140 ;
        RECT 140.195 186.715 141.265 186.885 ;
        RECT 141.435 186.815 142.825 187.030 ;
        RECT 142.995 186.815 144.285 187.265 ;
        RECT 144.915 187.140 145.085 188.080 ;
        RECT 145.635 187.900 145.805 188.225 ;
        RECT 145.255 187.730 145.805 187.900 ;
        RECT 145.985 187.660 146.355 187.990 ;
        RECT 146.535 187.900 146.705 188.225 ;
        RECT 146.875 188.080 147.805 188.410 ;
        RECT 146.535 187.730 147.465 187.900 ;
        RECT 145.255 187.300 147.465 187.470 ;
        RECT 145.255 187.210 145.760 187.300 ;
        RECT 146.560 187.200 147.465 187.300 ;
        RECT 144.455 187.030 145.085 187.140 ;
        RECT 144.455 186.815 145.465 187.030 ;
        RECT 146.060 187.015 146.390 187.130 ;
        RECT 147.635 187.030 147.805 188.080 ;
        RECT 139.475 186.625 139.645 186.700 ;
        RECT 139.005 186.455 139.645 186.625 ;
        RECT 140.620 186.600 140.950 186.715 ;
        RECT 141.435 186.700 142.365 186.815 ;
        RECT 143.675 186.710 144.005 186.815 ;
        RECT 138.655 185.955 139.290 186.285 ;
        RECT 133.315 184.970 133.865 185.140 ;
        RECT 134.035 184.710 134.205 185.320 ;
        RECT 136.755 184.710 136.925 185.555 ;
        RECT 139.475 185.650 139.645 186.455 ;
        RECT 139.815 186.430 140.320 186.520 ;
        RECT 141.120 186.430 142.025 186.530 ;
        RECT 139.815 186.260 142.025 186.430 ;
        RECT 139.815 185.910 142.025 186.090 ;
        RECT 139.815 185.830 140.320 185.910 ;
        RECT 141.120 185.820 142.025 185.910 ;
        RECT 139.475 185.320 140.025 185.650 ;
        RECT 140.620 185.635 140.950 185.740 ;
        RECT 142.195 185.650 142.365 186.700 ;
        RECT 144.915 186.700 145.465 186.815 ;
        RECT 145.635 186.845 146.705 187.015 ;
        RECT 142.535 186.540 143.505 186.645 ;
        RECT 144.175 186.540 144.745 186.645 ;
        RECT 142.535 186.260 144.745 186.540 ;
        RECT 142.535 185.910 144.745 186.090 ;
        RECT 142.535 185.820 143.440 185.910 ;
        RECT 144.240 185.830 144.745 185.910 ;
        RECT 140.195 185.465 141.265 185.635 ;
        RECT 139.475 184.710 139.645 185.320 ;
        RECT 140.195 185.140 140.365 185.465 ;
        RECT 139.815 184.970 140.365 185.140 ;
        RECT 140.545 184.900 140.915 185.240 ;
        RECT 141.095 185.140 141.265 185.465 ;
        RECT 141.435 185.320 143.125 185.650 ;
        RECT 143.610 185.635 143.940 185.740 ;
        RECT 144.915 185.650 145.085 186.700 ;
        RECT 145.635 186.520 145.805 186.845 ;
        RECT 145.255 186.350 145.805 186.520 ;
        RECT 145.985 186.280 146.355 186.610 ;
        RECT 146.535 186.520 146.705 186.845 ;
        RECT 146.875 186.700 147.805 187.030 ;
        RECT 146.535 186.350 147.465 186.520 ;
        RECT 145.255 185.910 147.465 186.090 ;
        RECT 145.255 185.830 145.760 185.910 ;
        RECT 146.560 185.820 147.465 185.910 ;
        RECT 143.295 185.465 144.365 185.635 ;
        RECT 141.095 184.960 142.025 185.140 ;
        RECT 142.195 184.710 142.365 185.320 ;
        RECT 143.295 185.140 143.465 185.465 ;
        RECT 142.535 184.960 143.465 185.140 ;
        RECT 143.645 184.900 144.015 185.240 ;
        RECT 144.195 185.140 144.365 185.465 ;
        RECT 144.535 185.320 145.465 185.650 ;
        RECT 146.060 185.635 146.390 185.740 ;
        RECT 147.635 185.650 147.805 186.700 ;
        RECT 145.635 185.465 146.705 185.635 ;
        RECT 144.195 184.970 144.745 185.140 ;
        RECT 144.915 184.710 145.085 185.320 ;
        RECT 145.635 185.140 145.805 185.465 ;
        RECT 145.255 184.970 145.805 185.140 ;
        RECT 145.985 184.900 146.355 185.240 ;
        RECT 146.535 185.140 146.705 185.465 ;
        RECT 146.875 185.320 147.805 185.650 ;
        RECT 146.535 184.960 147.465 185.140 ;
        RECT 147.635 184.710 147.805 185.320 ;
        RECT 89.315 183.835 89.835 184.375 ;
        RECT 90.005 183.665 90.525 184.205 ;
        RECT 76.895 182.915 82.240 183.460 ;
        RECT 82.415 182.915 87.760 183.460 ;
        RECT 87.935 182.915 89.145 183.665 ;
        RECT 89.315 182.915 90.525 183.665 ;
        RECT 112.275 184.020 113.195 184.710 ;
        RECT 113.365 184.190 116.795 184.710 ;
        RECT 112.275 183.500 113.735 184.020 ;
        RECT 113.905 183.500 116.255 184.190 ;
        RECT 116.965 184.020 118.635 184.710 ;
        RECT 118.805 184.190 122.235 184.710 ;
        RECT 116.425 183.500 119.175 184.020 ;
        RECT 119.345 183.500 121.695 184.190 ;
        RECT 122.405 184.020 124.075 184.710 ;
        RECT 124.245 184.190 127.675 184.710 ;
        RECT 121.865 183.500 124.615 184.020 ;
        RECT 124.785 183.500 127.135 184.190 ;
        RECT 127.845 184.020 129.515 184.710 ;
        RECT 129.685 184.190 133.115 184.710 ;
        RECT 127.305 183.500 130.055 184.020 ;
        RECT 130.225 183.500 132.575 184.190 ;
        RECT 133.285 184.020 134.955 184.710 ;
        RECT 135.125 184.190 138.555 184.710 ;
        RECT 132.745 183.500 135.495 184.020 ;
        RECT 135.665 183.500 138.015 184.190 ;
        RECT 138.725 184.020 140.395 184.710 ;
        RECT 140.565 184.190 143.995 184.710 ;
        RECT 138.185 183.500 140.935 184.020 ;
        RECT 141.105 183.500 143.455 184.190 ;
        RECT 144.165 184.020 145.835 184.710 ;
        RECT 146.005 184.190 147.805 184.710 ;
        RECT 143.625 183.500 146.375 184.020 ;
        RECT 146.545 183.500 147.805 184.190 ;
        RECT 112.275 183.415 112.445 183.500 ;
        RECT 114.995 183.415 115.165 183.500 ;
        RECT 117.715 183.415 117.885 183.500 ;
        RECT 120.435 183.415 120.605 183.500 ;
        RECT 123.155 183.415 123.325 183.500 ;
        RECT 125.875 183.415 126.045 183.500 ;
        RECT 128.595 183.415 128.765 183.500 ;
        RECT 131.315 183.415 131.485 183.500 ;
        RECT 134.035 183.415 134.205 183.500 ;
        RECT 136.755 183.415 136.925 183.500 ;
        RECT 139.475 183.415 139.645 183.500 ;
        RECT 142.195 183.415 142.365 183.500 ;
        RECT 144.915 183.415 145.085 183.500 ;
        RECT 147.635 183.415 147.805 183.500 ;
        RECT 11.950 182.745 90.610 182.915 ;
        RECT 12.035 181.995 13.245 182.745 ;
        RECT 13.415 182.200 18.760 182.745 ;
        RECT 12.035 181.455 12.555 181.995 ;
        RECT 12.725 181.285 13.245 181.825 ;
        RECT 15.000 181.370 15.340 182.200 ;
        RECT 18.935 181.975 20.605 182.745 ;
        RECT 20.810 182.005 21.425 182.575 ;
        RECT 21.595 182.235 21.810 182.745 ;
        RECT 22.040 182.235 22.320 182.565 ;
        RECT 22.500 182.235 22.740 182.745 ;
        RECT 12.035 180.195 13.245 181.285 ;
        RECT 16.820 180.630 17.170 181.880 ;
        RECT 18.935 181.455 19.685 181.975 ;
        RECT 19.855 181.285 20.605 181.805 ;
        RECT 13.415 180.195 18.760 180.630 ;
        RECT 18.935 180.195 20.605 181.285 ;
        RECT 20.810 180.985 21.125 182.005 ;
        RECT 21.295 181.335 21.465 181.835 ;
        RECT 21.715 181.505 21.980 182.065 ;
        RECT 22.150 181.335 22.320 182.235 ;
        RECT 23.075 182.200 28.420 182.745 ;
        RECT 22.490 181.505 22.845 182.065 ;
        RECT 24.660 181.370 25.000 182.200 ;
        RECT 29.055 182.025 29.395 182.535 ;
        RECT 21.295 181.165 22.720 181.335 ;
        RECT 20.810 180.365 21.345 180.985 ;
        RECT 21.515 180.195 21.845 180.995 ;
        RECT 22.330 180.990 22.720 181.165 ;
        RECT 26.480 180.630 26.830 181.880 ;
        RECT 23.075 180.195 28.420 180.630 ;
        RECT 29.055 180.625 29.315 182.025 ;
        RECT 29.565 181.945 29.835 182.745 ;
        RECT 29.490 181.505 29.820 181.755 ;
        RECT 30.015 181.505 30.295 182.475 ;
        RECT 30.475 181.505 30.775 182.475 ;
        RECT 30.955 181.505 31.305 182.470 ;
        RECT 31.525 182.245 32.020 182.575 ;
        RECT 29.505 181.335 29.820 181.505 ;
        RECT 31.525 181.335 31.695 182.245 ;
        RECT 29.505 181.165 31.695 181.335 ;
        RECT 29.055 180.365 29.395 180.625 ;
        RECT 29.565 180.195 29.895 180.995 ;
        RECT 30.360 180.365 30.610 181.165 ;
        RECT 30.795 180.195 31.125 180.915 ;
        RECT 31.345 180.365 31.595 181.165 ;
        RECT 31.865 180.755 32.105 182.065 ;
        RECT 32.735 182.005 33.175 182.565 ;
        RECT 33.345 182.005 33.795 182.745 ;
        RECT 33.965 182.175 34.135 182.575 ;
        RECT 34.305 182.345 34.725 182.745 ;
        RECT 34.895 182.175 35.125 182.575 ;
        RECT 33.965 182.005 35.125 182.175 ;
        RECT 35.295 182.005 35.785 182.575 ;
        RECT 32.735 180.995 33.045 182.005 ;
        RECT 33.215 181.385 33.385 181.835 ;
        RECT 33.555 181.555 33.945 181.835 ;
        RECT 34.130 181.505 34.375 181.835 ;
        RECT 33.215 181.215 34.005 181.385 ;
        RECT 31.765 180.195 32.100 180.575 ;
        RECT 32.735 180.365 33.175 180.995 ;
        RECT 33.350 180.195 33.665 181.045 ;
        RECT 33.835 180.535 34.005 181.215 ;
        RECT 34.175 180.705 34.375 181.505 ;
        RECT 34.575 180.705 34.825 181.835 ;
        RECT 35.040 181.505 35.445 181.835 ;
        RECT 35.615 181.335 35.785 182.005 ;
        RECT 35.955 181.975 37.625 182.745 ;
        RECT 37.795 182.020 38.085 182.745 ;
        RECT 39.175 182.005 39.640 182.550 ;
        RECT 35.955 181.455 36.705 181.975 ;
        RECT 35.015 181.165 35.785 181.335 ;
        RECT 36.875 181.285 37.625 181.805 ;
        RECT 35.015 180.535 35.265 181.165 ;
        RECT 33.835 180.365 35.265 180.535 ;
        RECT 35.445 180.195 35.775 180.995 ;
        RECT 35.955 180.195 37.625 181.285 ;
        RECT 37.795 180.195 38.085 181.360 ;
        RECT 39.175 181.045 39.345 182.005 ;
        RECT 40.145 181.925 40.315 182.745 ;
        RECT 40.485 182.095 40.815 182.575 ;
        RECT 40.985 182.355 41.335 182.745 ;
        RECT 41.505 182.175 41.735 182.575 ;
        RECT 41.225 182.095 41.735 182.175 ;
        RECT 40.485 182.005 41.735 182.095 ;
        RECT 41.905 182.005 42.225 182.485 ;
        RECT 40.485 181.925 41.395 182.005 ;
        RECT 39.515 181.385 39.760 181.835 ;
        RECT 40.020 181.555 40.715 181.755 ;
        RECT 40.885 181.585 41.485 181.755 ;
        RECT 40.885 181.385 41.055 181.585 ;
        RECT 41.715 181.415 41.885 181.835 ;
        RECT 39.515 181.215 41.055 181.385 ;
        RECT 41.225 181.245 41.885 181.415 ;
        RECT 41.225 181.045 41.395 181.245 ;
        RECT 42.055 181.075 42.225 182.005 ;
        RECT 42.395 181.945 43.090 182.575 ;
        RECT 43.295 181.945 43.605 182.745 ;
        RECT 43.940 182.235 44.180 182.745 ;
        RECT 44.360 182.235 44.640 182.565 ;
        RECT 44.870 182.235 45.085 182.745 ;
        RECT 42.915 181.895 43.090 181.945 ;
        RECT 42.415 181.505 42.750 181.755 ;
        RECT 42.920 181.345 43.090 181.895 ;
        RECT 43.260 181.505 43.595 181.775 ;
        RECT 43.835 181.505 44.190 182.065 ;
        RECT 39.175 180.875 41.395 181.045 ;
        RECT 41.565 180.875 42.225 181.075 ;
        RECT 39.175 180.195 39.475 180.705 ;
        RECT 39.645 180.365 39.975 180.875 ;
        RECT 41.565 180.705 41.735 180.875 ;
        RECT 40.145 180.195 40.775 180.705 ;
        RECT 41.355 180.535 41.735 180.705 ;
        RECT 41.905 180.195 42.205 180.705 ;
        RECT 42.395 180.195 42.655 181.335 ;
        RECT 42.825 180.365 43.155 181.345 ;
        RECT 44.360 181.335 44.530 182.235 ;
        RECT 44.700 181.505 44.965 182.065 ;
        RECT 45.255 182.005 45.870 182.575 ;
        RECT 46.160 182.175 46.335 182.575 ;
        RECT 46.505 182.365 46.835 182.745 ;
        RECT 47.080 182.245 47.310 182.575 ;
        RECT 46.160 182.005 46.790 182.175 ;
        RECT 45.215 181.335 45.385 181.835 ;
        RECT 43.325 180.195 43.605 181.335 ;
        RECT 43.960 181.165 45.385 181.335 ;
        RECT 43.960 180.990 44.350 181.165 ;
        RECT 44.835 180.195 45.165 180.995 ;
        RECT 45.555 180.985 45.870 182.005 ;
        RECT 46.620 181.835 46.790 182.005 ;
        RECT 46.075 181.155 46.440 181.835 ;
        RECT 46.620 181.505 46.970 181.835 ;
        RECT 46.620 180.985 46.790 181.505 ;
        RECT 45.335 180.365 45.870 180.985 ;
        RECT 46.160 180.815 46.790 180.985 ;
        RECT 47.140 180.955 47.310 182.245 ;
        RECT 47.510 181.135 47.790 182.410 ;
        RECT 48.015 182.405 48.285 182.410 ;
        RECT 47.975 182.235 48.285 182.405 ;
        RECT 48.745 182.365 49.075 182.745 ;
        RECT 49.245 182.490 49.580 182.535 ;
        RECT 48.015 181.135 48.285 182.235 ;
        RECT 48.475 181.135 48.815 182.165 ;
        RECT 49.245 182.025 49.585 182.490 ;
        RECT 49.760 182.215 50.050 182.565 ;
        RECT 50.245 182.385 50.575 182.745 ;
        RECT 50.745 182.215 50.975 182.520 ;
        RECT 49.760 182.045 50.975 182.215 ;
        RECT 51.165 182.405 51.335 182.440 ;
        RECT 51.165 182.235 51.365 182.405 ;
        RECT 48.985 181.505 49.245 181.835 ;
        RECT 48.985 180.955 49.155 181.505 ;
        RECT 49.415 181.335 49.585 182.025 ;
        RECT 51.165 181.875 51.335 182.235 ;
        RECT 51.735 182.150 52.055 182.575 ;
        RECT 52.225 182.320 52.555 182.745 ;
        RECT 52.725 182.325 53.815 182.575 ;
        RECT 54.005 182.325 55.095 182.575 ;
        RECT 52.725 182.150 52.895 182.325 ;
        RECT 51.735 181.980 52.895 182.150 ;
        RECT 53.065 181.985 54.755 182.155 ;
        RECT 54.925 182.150 55.095 182.325 ;
        RECT 55.265 182.320 55.595 182.745 ;
        RECT 55.765 182.150 56.015 182.575 ;
        RECT 49.820 181.725 50.080 181.835 ;
        RECT 49.815 181.555 50.080 181.725 ;
        RECT 49.820 181.505 50.080 181.555 ;
        RECT 50.260 181.505 50.645 181.835 ;
        RECT 50.815 181.705 51.335 181.875 ;
        RECT 51.610 181.725 52.720 181.755 ;
        RECT 46.160 180.365 46.335 180.815 ;
        RECT 47.140 180.785 49.155 180.955 ;
        RECT 46.505 180.195 46.835 180.635 ;
        RECT 47.140 180.365 47.310 180.785 ;
        RECT 47.545 180.195 48.215 180.605 ;
        RECT 48.430 180.365 48.600 180.785 ;
        RECT 48.800 180.195 49.130 180.605 ;
        RECT 49.325 180.365 49.585 181.335 ;
        RECT 49.760 180.195 50.080 181.335 ;
        RECT 50.260 180.455 50.455 181.505 ;
        RECT 50.815 181.325 50.985 181.705 ;
        RECT 51.610 181.555 52.745 181.725 ;
        RECT 53.010 181.555 53.665 181.755 ;
        RECT 50.635 181.045 50.985 181.325 ;
        RECT 51.175 181.175 51.420 181.535 ;
        RECT 53.950 181.345 54.240 181.985 ;
        RECT 54.925 181.980 56.015 182.150 ;
        RECT 56.195 182.160 56.505 182.575 ;
        RECT 56.700 182.365 57.030 182.745 ;
        RECT 57.200 182.405 58.605 182.575 ;
        RECT 57.200 182.175 57.370 182.405 ;
        RECT 54.410 181.555 55.040 181.755 ;
        RECT 55.330 181.725 55.960 181.755 ;
        RECT 55.330 181.555 55.965 181.725 ;
        RECT 51.805 181.175 53.735 181.345 ;
        RECT 50.635 180.365 50.965 181.045 ;
        RECT 51.165 180.195 51.420 180.995 ;
        RECT 51.805 180.365 52.135 181.175 ;
        RECT 52.305 180.195 52.475 181.005 ;
        RECT 52.645 180.365 52.975 181.175 ;
        RECT 53.145 180.195 53.315 181.005 ;
        RECT 53.485 180.535 53.735 181.175 ;
        RECT 53.950 181.175 56.015 181.345 ;
        RECT 53.950 180.705 54.335 181.175 ;
        RECT 54.505 180.535 54.675 181.005 ;
        RECT 54.845 180.705 55.175 181.175 ;
        RECT 55.345 180.535 55.595 181.005 ;
        RECT 53.485 180.365 55.595 180.535 ;
        RECT 55.765 180.365 56.015 181.175 ;
        RECT 56.195 181.045 56.365 182.160 ;
        RECT 56.675 182.005 57.370 182.175 ;
        RECT 58.435 182.175 58.605 182.405 ;
        RECT 58.875 182.345 59.205 182.745 ;
        RECT 59.445 182.175 59.615 182.575 ;
        RECT 56.675 181.835 56.845 182.005 ;
        RECT 56.535 181.505 56.845 181.835 ;
        RECT 57.015 181.505 57.350 181.835 ;
        RECT 57.620 181.505 57.815 182.080 ;
        RECT 58.075 181.835 58.265 182.065 ;
        RECT 58.435 182.005 59.615 182.175 ;
        RECT 60.335 181.925 60.595 182.745 ;
        RECT 60.765 181.925 61.095 182.345 ;
        RECT 61.275 182.175 61.535 182.575 ;
        RECT 61.705 182.345 62.035 182.745 ;
        RECT 62.205 182.175 62.375 182.525 ;
        RECT 62.545 182.345 62.920 182.745 ;
        RECT 61.275 182.005 62.940 182.175 ;
        RECT 63.110 182.070 63.385 182.415 ;
        RECT 60.845 181.835 61.095 181.925 ;
        RECT 62.770 181.835 62.940 182.005 ;
        RECT 58.075 181.505 58.420 181.835 ;
        RECT 58.730 181.505 59.205 181.835 ;
        RECT 59.460 181.505 59.645 181.835 ;
        RECT 60.340 181.505 60.675 181.755 ;
        RECT 60.845 181.505 61.560 181.835 ;
        RECT 61.775 181.505 62.600 181.835 ;
        RECT 62.770 181.505 63.045 181.835 ;
        RECT 56.675 181.335 56.845 181.505 ;
        RECT 56.675 181.165 59.615 181.335 ;
        RECT 56.195 180.405 56.535 181.045 ;
        RECT 57.125 180.825 58.685 180.995 ;
        RECT 56.705 180.195 56.950 180.655 ;
        RECT 57.125 180.365 57.375 180.825 ;
        RECT 57.565 180.195 58.235 180.575 ;
        RECT 58.435 180.365 58.685 180.825 ;
        RECT 59.445 180.365 59.615 181.165 ;
        RECT 60.335 180.195 60.595 181.335 ;
        RECT 60.845 180.945 61.015 181.505 ;
        RECT 61.275 181.045 61.605 181.335 ;
        RECT 61.775 181.215 62.020 181.505 ;
        RECT 62.770 181.335 62.940 181.505 ;
        RECT 63.215 181.335 63.385 182.070 ;
        RECT 63.555 182.020 63.845 182.745 ;
        RECT 64.015 182.095 64.275 182.575 ;
        RECT 64.445 182.285 64.775 182.745 ;
        RECT 64.965 182.105 65.165 182.525 ;
        RECT 62.280 181.165 62.940 181.335 ;
        RECT 62.280 181.045 62.450 181.165 ;
        RECT 61.275 180.875 62.450 181.045 ;
        RECT 60.835 180.375 62.450 180.705 ;
        RECT 62.620 180.195 62.900 180.995 ;
        RECT 63.110 180.365 63.385 181.335 ;
        RECT 63.555 180.195 63.845 181.360 ;
        RECT 64.015 181.065 64.185 182.095 ;
        RECT 64.355 181.405 64.585 181.835 ;
        RECT 64.755 181.585 65.165 182.105 ;
        RECT 65.335 182.260 66.125 182.525 ;
        RECT 65.335 181.405 65.590 182.260 ;
        RECT 66.305 181.925 66.635 182.345 ;
        RECT 66.805 181.925 67.065 182.745 ;
        RECT 67.235 182.365 68.125 182.535 ;
        RECT 66.305 181.835 66.555 181.925 ;
        RECT 65.760 181.585 66.555 181.835 ;
        RECT 67.235 181.810 67.785 182.195 ;
        RECT 64.355 181.235 66.145 181.405 ;
        RECT 64.015 180.365 64.290 181.065 ;
        RECT 64.460 180.940 65.175 181.235 ;
        RECT 65.395 180.875 65.725 181.065 ;
        RECT 64.500 180.195 64.715 180.740 ;
        RECT 64.885 180.365 65.360 180.705 ;
        RECT 65.530 180.700 65.725 180.875 ;
        RECT 65.895 180.870 66.145 181.235 ;
        RECT 65.530 180.195 66.145 180.700 ;
        RECT 66.385 180.365 66.555 181.585 ;
        RECT 66.725 180.875 67.065 181.755 ;
        RECT 67.955 181.640 68.125 182.365 ;
        RECT 67.235 181.570 68.125 181.640 ;
        RECT 68.295 182.040 68.515 182.525 ;
        RECT 68.685 182.205 68.935 182.745 ;
        RECT 69.105 182.095 69.365 182.575 ;
        RECT 68.295 181.615 68.625 182.040 ;
        RECT 67.235 181.545 68.130 181.570 ;
        RECT 67.235 181.530 68.140 181.545 ;
        RECT 67.235 181.515 68.145 181.530 ;
        RECT 67.235 181.510 68.155 181.515 ;
        RECT 67.235 181.500 68.160 181.510 ;
        RECT 67.235 181.490 68.165 181.500 ;
        RECT 67.235 181.485 68.175 181.490 ;
        RECT 67.235 181.475 68.185 181.485 ;
        RECT 67.235 181.470 68.195 181.475 ;
        RECT 67.235 181.020 67.495 181.470 ;
        RECT 67.860 181.465 68.195 181.470 ;
        RECT 67.860 181.460 68.210 181.465 ;
        RECT 67.860 181.450 68.225 181.460 ;
        RECT 67.860 181.445 68.250 181.450 ;
        RECT 68.795 181.445 69.025 181.840 ;
        RECT 67.860 181.440 69.025 181.445 ;
        RECT 67.890 181.405 69.025 181.440 ;
        RECT 67.925 181.380 69.025 181.405 ;
        RECT 67.955 181.350 69.025 181.380 ;
        RECT 67.975 181.320 69.025 181.350 ;
        RECT 67.995 181.290 69.025 181.320 ;
        RECT 68.065 181.280 69.025 181.290 ;
        RECT 68.090 181.270 69.025 181.280 ;
        RECT 68.110 181.255 69.025 181.270 ;
        RECT 68.130 181.240 69.025 181.255 ;
        RECT 68.135 181.230 68.920 181.240 ;
        RECT 68.150 181.195 68.920 181.230 ;
        RECT 67.665 180.875 67.995 181.120 ;
        RECT 68.165 180.945 68.920 181.195 ;
        RECT 69.195 181.065 69.365 182.095 ;
        RECT 69.625 182.195 69.795 182.485 ;
        RECT 69.965 182.365 70.295 182.745 ;
        RECT 69.625 182.025 70.290 182.195 ;
        RECT 69.540 181.205 69.890 181.855 ;
        RECT 67.665 180.850 67.850 180.875 ;
        RECT 67.235 180.750 67.850 180.850 ;
        RECT 66.805 180.195 67.065 180.705 ;
        RECT 67.235 180.195 67.840 180.750 ;
        RECT 68.015 180.365 68.495 180.705 ;
        RECT 68.665 180.195 68.920 180.740 ;
        RECT 69.090 180.365 69.365 181.065 ;
        RECT 70.060 181.035 70.290 182.025 ;
        RECT 69.625 180.865 70.290 181.035 ;
        RECT 69.625 180.365 69.795 180.865 ;
        RECT 69.965 180.195 70.295 180.695 ;
        RECT 70.465 180.365 70.650 182.485 ;
        RECT 70.905 182.285 71.155 182.745 ;
        RECT 71.325 182.295 71.660 182.465 ;
        RECT 71.855 182.295 72.530 182.465 ;
        RECT 71.325 182.155 71.495 182.295 ;
        RECT 70.820 181.165 71.100 182.115 ;
        RECT 71.270 182.025 71.495 182.155 ;
        RECT 71.270 180.920 71.440 182.025 ;
        RECT 71.665 181.875 72.190 182.095 ;
        RECT 71.610 181.110 71.850 181.705 ;
        RECT 72.020 181.175 72.190 181.875 ;
        RECT 72.360 181.515 72.530 182.295 ;
        RECT 72.850 182.245 73.220 182.745 ;
        RECT 73.400 182.295 73.805 182.465 ;
        RECT 73.975 182.295 74.760 182.465 ;
        RECT 73.400 182.065 73.570 182.295 ;
        RECT 72.740 181.765 73.570 182.065 ;
        RECT 73.955 181.795 74.420 182.125 ;
        RECT 72.740 181.735 72.940 181.765 ;
        RECT 73.060 181.515 73.230 181.585 ;
        RECT 72.360 181.345 73.230 181.515 ;
        RECT 72.720 181.255 73.230 181.345 ;
        RECT 71.270 180.790 71.575 180.920 ;
        RECT 72.020 180.810 72.550 181.175 ;
        RECT 70.890 180.195 71.155 180.655 ;
        RECT 71.325 180.365 71.575 180.790 ;
        RECT 72.720 180.640 72.890 181.255 ;
        RECT 71.785 180.470 72.890 180.640 ;
        RECT 73.060 180.195 73.230 180.995 ;
        RECT 73.400 180.695 73.570 181.765 ;
        RECT 73.740 180.865 73.930 181.585 ;
        RECT 74.100 180.835 74.420 181.795 ;
        RECT 74.590 181.835 74.760 182.295 ;
        RECT 75.035 182.215 75.245 182.745 ;
        RECT 75.505 182.005 75.835 182.530 ;
        RECT 76.005 182.135 76.175 182.745 ;
        RECT 76.345 182.090 76.675 182.525 ;
        RECT 76.895 182.200 82.240 182.745 ;
        RECT 82.415 182.200 87.760 182.745 ;
        RECT 76.345 182.005 76.725 182.090 ;
        RECT 75.635 181.835 75.835 182.005 ;
        RECT 76.500 181.965 76.725 182.005 ;
        RECT 74.590 181.505 75.465 181.835 ;
        RECT 75.635 181.505 76.385 181.835 ;
        RECT 73.400 180.365 73.650 180.695 ;
        RECT 74.590 180.665 74.760 181.505 ;
        RECT 75.635 181.300 75.825 181.505 ;
        RECT 76.555 181.385 76.725 181.965 ;
        RECT 76.510 181.335 76.725 181.385 ;
        RECT 78.480 181.370 78.820 182.200 ;
        RECT 74.930 180.925 75.825 181.300 ;
        RECT 76.335 181.255 76.725 181.335 ;
        RECT 73.875 180.495 74.760 180.665 ;
        RECT 74.940 180.195 75.255 180.695 ;
        RECT 75.485 180.365 75.825 180.925 ;
        RECT 75.995 180.195 76.165 181.205 ;
        RECT 76.335 180.410 76.665 181.255 ;
        RECT 80.300 180.630 80.650 181.880 ;
        RECT 84.000 181.370 84.340 182.200 ;
        RECT 87.935 181.995 89.145 182.745 ;
        RECT 89.315 181.995 90.525 182.745 ;
        RECT 85.820 180.630 86.170 181.880 ;
        RECT 87.935 181.455 88.455 181.995 ;
        RECT 88.625 181.285 89.145 181.825 ;
        RECT 76.895 180.195 82.240 180.630 ;
        RECT 82.415 180.195 87.760 180.630 ;
        RECT 87.935 180.195 89.145 181.285 ;
        RECT 89.315 181.285 89.835 181.825 ;
        RECT 90.005 181.455 90.525 181.995 ;
        RECT 89.315 180.195 90.525 181.285 ;
        RECT 11.950 180.025 90.610 180.195 ;
        RECT 12.035 178.935 13.245 180.025 ;
        RECT 13.415 178.935 16.925 180.025 ;
        RECT 17.615 178.965 17.945 179.810 ;
        RECT 18.115 179.015 18.285 180.025 ;
        RECT 18.455 179.295 18.795 179.855 ;
        RECT 19.025 179.525 19.340 180.025 ;
        RECT 19.520 179.555 20.405 179.725 ;
        RECT 12.035 178.225 12.555 178.765 ;
        RECT 12.725 178.395 13.245 178.935 ;
        RECT 13.415 178.245 15.065 178.765 ;
        RECT 15.235 178.415 16.925 178.935 ;
        RECT 17.555 178.885 17.945 178.965 ;
        RECT 18.455 178.920 19.350 179.295 ;
        RECT 17.555 178.835 17.770 178.885 ;
        RECT 17.555 178.255 17.725 178.835 ;
        RECT 18.455 178.715 18.645 178.920 ;
        RECT 19.520 178.715 19.690 179.555 ;
        RECT 20.630 179.525 20.880 179.855 ;
        RECT 17.895 178.385 18.645 178.715 ;
        RECT 18.815 178.385 19.690 178.715 ;
        RECT 12.035 177.475 13.245 178.225 ;
        RECT 13.415 177.475 16.925 178.245 ;
        RECT 17.555 178.215 17.780 178.255 ;
        RECT 18.445 178.215 18.645 178.385 ;
        RECT 17.555 178.130 17.935 178.215 ;
        RECT 17.605 177.695 17.935 178.130 ;
        RECT 18.105 177.475 18.275 178.085 ;
        RECT 18.445 177.690 18.775 178.215 ;
        RECT 19.035 177.475 19.245 178.005 ;
        RECT 19.520 177.925 19.690 178.385 ;
        RECT 19.860 178.425 20.180 179.385 ;
        RECT 20.350 178.635 20.540 179.355 ;
        RECT 20.710 178.455 20.880 179.525 ;
        RECT 21.050 179.225 21.220 180.025 ;
        RECT 21.390 179.580 22.495 179.750 ;
        RECT 21.390 178.965 21.560 179.580 ;
        RECT 22.705 179.430 22.955 179.855 ;
        RECT 23.125 179.565 23.390 180.025 ;
        RECT 21.730 179.045 22.260 179.410 ;
        RECT 22.705 179.300 23.010 179.430 ;
        RECT 21.050 178.875 21.560 178.965 ;
        RECT 21.050 178.705 21.920 178.875 ;
        RECT 21.050 178.635 21.220 178.705 ;
        RECT 21.340 178.455 21.540 178.485 ;
        RECT 19.860 178.095 20.325 178.425 ;
        RECT 20.710 178.155 21.540 178.455 ;
        RECT 20.710 177.925 20.880 178.155 ;
        RECT 19.520 177.755 20.305 177.925 ;
        RECT 20.475 177.755 20.880 177.925 ;
        RECT 21.060 177.475 21.430 177.975 ;
        RECT 21.750 177.925 21.920 178.705 ;
        RECT 22.090 178.345 22.260 179.045 ;
        RECT 22.430 178.515 22.670 179.110 ;
        RECT 22.090 178.125 22.615 178.345 ;
        RECT 22.840 178.195 23.010 179.300 ;
        RECT 22.785 178.065 23.010 178.195 ;
        RECT 23.180 178.105 23.460 179.055 ;
        RECT 22.785 177.925 22.955 178.065 ;
        RECT 21.750 177.755 22.425 177.925 ;
        RECT 22.620 177.755 22.955 177.925 ;
        RECT 23.125 177.475 23.375 177.935 ;
        RECT 23.630 177.735 23.815 179.855 ;
        RECT 23.985 179.525 24.315 180.025 ;
        RECT 24.485 179.355 24.655 179.855 ;
        RECT 23.990 179.185 24.655 179.355 ;
        RECT 23.990 178.195 24.220 179.185 ;
        RECT 24.390 178.365 24.740 179.015 ;
        RECT 24.915 178.860 25.205 180.025 ;
        RECT 25.375 179.515 25.635 180.025 ;
        RECT 25.375 178.465 25.715 179.345 ;
        RECT 25.885 178.635 26.055 179.855 ;
        RECT 26.295 179.520 26.910 180.025 ;
        RECT 26.295 178.985 26.545 179.350 ;
        RECT 26.715 179.345 26.910 179.520 ;
        RECT 27.080 179.515 27.555 179.855 ;
        RECT 27.725 179.480 27.940 180.025 ;
        RECT 26.715 179.155 27.045 179.345 ;
        RECT 27.265 178.985 27.980 179.280 ;
        RECT 28.150 179.155 28.425 179.855 ;
        RECT 28.685 179.355 28.855 179.855 ;
        RECT 29.025 179.525 29.355 180.025 ;
        RECT 28.685 179.185 29.350 179.355 ;
        RECT 26.295 178.815 28.085 178.985 ;
        RECT 25.885 178.385 26.680 178.635 ;
        RECT 25.885 178.295 26.135 178.385 ;
        RECT 23.990 178.025 24.655 178.195 ;
        RECT 23.985 177.475 24.315 177.855 ;
        RECT 24.485 177.735 24.655 178.025 ;
        RECT 24.915 177.475 25.205 178.200 ;
        RECT 25.375 177.475 25.635 178.295 ;
        RECT 25.805 177.875 26.135 178.295 ;
        RECT 26.850 177.960 27.105 178.815 ;
        RECT 26.315 177.695 27.105 177.960 ;
        RECT 27.275 178.115 27.685 178.635 ;
        RECT 27.855 178.385 28.085 178.815 ;
        RECT 28.255 178.125 28.425 179.155 ;
        RECT 28.600 178.365 28.950 179.015 ;
        RECT 29.120 178.195 29.350 179.185 ;
        RECT 27.275 177.695 27.475 178.115 ;
        RECT 27.665 177.475 27.995 177.935 ;
        RECT 28.165 177.645 28.425 178.125 ;
        RECT 28.685 178.025 29.350 178.195 ;
        RECT 28.685 177.735 28.855 178.025 ;
        RECT 29.025 177.475 29.355 177.855 ;
        RECT 29.525 177.735 29.710 179.855 ;
        RECT 29.950 179.565 30.215 180.025 ;
        RECT 30.385 179.430 30.635 179.855 ;
        RECT 30.845 179.580 31.950 179.750 ;
        RECT 30.330 179.300 30.635 179.430 ;
        RECT 29.880 178.105 30.160 179.055 ;
        RECT 30.330 178.195 30.500 179.300 ;
        RECT 30.670 178.515 30.910 179.110 ;
        RECT 31.080 179.045 31.610 179.410 ;
        RECT 31.080 178.345 31.250 179.045 ;
        RECT 31.780 178.965 31.950 179.580 ;
        RECT 32.120 179.225 32.290 180.025 ;
        RECT 32.460 179.525 32.710 179.855 ;
        RECT 32.935 179.555 33.820 179.725 ;
        RECT 31.780 178.875 32.290 178.965 ;
        RECT 30.330 178.065 30.555 178.195 ;
        RECT 30.725 178.125 31.250 178.345 ;
        RECT 31.420 178.705 32.290 178.875 ;
        RECT 29.965 177.475 30.215 177.935 ;
        RECT 30.385 177.925 30.555 178.065 ;
        RECT 31.420 177.925 31.590 178.705 ;
        RECT 32.120 178.635 32.290 178.705 ;
        RECT 31.800 178.455 32.000 178.485 ;
        RECT 32.460 178.455 32.630 179.525 ;
        RECT 32.800 178.635 32.990 179.355 ;
        RECT 31.800 178.155 32.630 178.455 ;
        RECT 33.160 178.425 33.480 179.385 ;
        RECT 30.385 177.755 30.720 177.925 ;
        RECT 30.915 177.755 31.590 177.925 ;
        RECT 31.910 177.475 32.280 177.975 ;
        RECT 32.460 177.925 32.630 178.155 ;
        RECT 33.015 178.095 33.480 178.425 ;
        RECT 33.650 178.715 33.820 179.555 ;
        RECT 34.000 179.525 34.315 180.025 ;
        RECT 34.545 179.295 34.885 179.855 ;
        RECT 33.990 178.920 34.885 179.295 ;
        RECT 35.055 179.015 35.225 180.025 ;
        RECT 34.695 178.715 34.885 178.920 ;
        RECT 35.395 178.965 35.725 179.810 ;
        RECT 36.435 178.970 36.740 179.755 ;
        RECT 36.920 179.555 37.605 180.025 ;
        RECT 36.915 179.035 37.610 179.345 ;
        RECT 35.395 178.885 35.785 178.965 ;
        RECT 35.570 178.835 35.785 178.885 ;
        RECT 33.650 178.385 34.525 178.715 ;
        RECT 34.695 178.385 35.445 178.715 ;
        RECT 33.650 177.925 33.820 178.385 ;
        RECT 34.695 178.215 34.895 178.385 ;
        RECT 35.615 178.255 35.785 178.835 ;
        RECT 35.560 178.215 35.785 178.255 ;
        RECT 32.460 177.755 32.865 177.925 ;
        RECT 33.035 177.755 33.820 177.925 ;
        RECT 34.095 177.475 34.305 178.005 ;
        RECT 34.565 177.690 34.895 178.215 ;
        RECT 35.405 178.130 35.785 178.215 ;
        RECT 36.435 178.165 36.610 178.970 ;
        RECT 37.785 178.865 38.070 179.810 ;
        RECT 38.245 179.575 38.575 180.025 ;
        RECT 38.745 179.405 38.915 179.835 ;
        RECT 39.175 179.590 44.520 180.025 ;
        RECT 37.210 178.715 38.070 178.865 ;
        RECT 36.785 178.695 38.070 178.715 ;
        RECT 38.240 179.175 38.915 179.405 ;
        RECT 36.785 178.335 37.770 178.695 ;
        RECT 38.240 178.525 38.475 179.175 ;
        RECT 35.065 177.475 35.235 178.085 ;
        RECT 35.405 177.695 35.735 178.130 ;
        RECT 36.435 177.645 36.675 178.165 ;
        RECT 37.600 178.000 37.770 178.335 ;
        RECT 37.940 178.195 38.475 178.525 ;
        RECT 38.255 178.045 38.475 178.195 ;
        RECT 38.645 178.155 38.945 179.005 ;
        RECT 36.845 177.475 37.240 177.970 ;
        RECT 37.600 177.805 37.975 178.000 ;
        RECT 37.805 177.660 37.975 177.805 ;
        RECT 38.255 177.670 38.495 178.045 ;
        RECT 40.760 178.020 41.100 178.850 ;
        RECT 42.580 178.340 42.930 179.590 ;
        RECT 44.880 179.055 45.270 179.230 ;
        RECT 45.755 179.225 46.085 180.025 ;
        RECT 46.255 179.235 46.790 179.855 ;
        RECT 47.460 179.515 49.115 179.805 ;
        RECT 44.880 178.885 46.305 179.055 ;
        RECT 44.755 178.155 45.110 178.715 ;
        RECT 38.665 177.475 39.000 177.980 ;
        RECT 39.175 177.475 44.520 178.020 ;
        RECT 45.280 177.985 45.450 178.885 ;
        RECT 45.620 178.155 45.885 178.715 ;
        RECT 46.135 178.385 46.305 178.885 ;
        RECT 46.475 178.215 46.790 179.235 ;
        RECT 47.460 179.175 49.050 179.345 ;
        RECT 49.285 179.225 49.565 180.025 ;
        RECT 47.460 178.885 47.780 179.175 ;
        RECT 48.880 179.055 49.050 179.175 ;
        RECT 47.975 178.835 48.690 179.005 ;
        RECT 48.880 178.885 49.605 179.055 ;
        RECT 49.775 178.885 50.045 179.855 ;
        RECT 44.860 177.475 45.100 177.985 ;
        RECT 45.280 177.655 45.560 177.985 ;
        RECT 45.790 177.475 46.005 177.985 ;
        RECT 46.175 177.645 46.790 178.215 ;
        RECT 47.460 178.145 47.810 178.715 ;
        RECT 47.980 178.385 48.690 178.835 ;
        RECT 49.435 178.715 49.605 178.885 ;
        RECT 48.860 178.385 49.265 178.715 ;
        RECT 49.435 178.385 49.705 178.715 ;
        RECT 49.435 178.215 49.605 178.385 ;
        RECT 47.995 178.045 49.605 178.215 ;
        RECT 49.875 178.150 50.045 178.885 ;
        RECT 50.675 178.860 50.965 180.025 ;
        RECT 47.465 177.475 47.795 177.975 ;
        RECT 47.995 177.695 48.165 178.045 ;
        RECT 48.365 177.475 48.695 177.875 ;
        RECT 48.865 177.695 49.035 178.045 ;
        RECT 49.205 177.475 49.585 177.875 ;
        RECT 49.775 177.805 50.045 178.150 ;
        RECT 50.675 177.475 50.965 178.200 ;
        RECT 51.135 177.755 51.415 179.855 ;
        RECT 51.605 179.265 52.390 180.025 ;
        RECT 52.785 179.195 53.170 179.855 ;
        RECT 52.785 179.095 53.195 179.195 ;
        RECT 51.585 178.885 53.195 179.095 ;
        RECT 53.495 179.005 53.695 179.795 ;
        RECT 51.585 178.285 51.860 178.885 ;
        RECT 53.365 178.835 53.695 179.005 ;
        RECT 53.865 178.845 54.185 180.025 ;
        RECT 54.815 178.885 55.075 180.025 ;
        RECT 55.245 178.875 55.575 179.855 ;
        RECT 55.745 178.885 56.025 180.025 ;
        RECT 56.195 179.155 56.470 179.855 ;
        RECT 56.640 179.480 56.895 180.025 ;
        RECT 57.065 179.515 57.545 179.855 ;
        RECT 57.720 179.470 58.325 180.025 ;
        RECT 57.710 179.370 58.325 179.470 ;
        RECT 57.710 179.345 57.895 179.370 ;
        RECT 53.365 178.715 53.545 178.835 ;
        RECT 52.030 178.465 52.385 178.715 ;
        RECT 52.580 178.665 53.045 178.715 ;
        RECT 52.575 178.495 53.045 178.665 ;
        RECT 52.580 178.465 53.045 178.495 ;
        RECT 53.215 178.465 53.545 178.715 ;
        RECT 53.720 178.465 54.185 178.665 ;
        RECT 54.835 178.465 55.170 178.715 ;
        RECT 51.585 178.105 52.835 178.285 ;
        RECT 55.340 178.275 55.510 178.875 ;
        RECT 55.680 178.445 56.015 178.715 ;
        RECT 52.470 178.035 52.835 178.105 ;
        RECT 53.005 178.085 54.185 178.255 ;
        RECT 51.645 177.475 51.815 177.935 ;
        RECT 53.005 177.865 53.335 178.085 ;
        RECT 52.085 177.685 53.335 177.865 ;
        RECT 53.505 177.475 53.675 177.915 ;
        RECT 53.845 177.670 54.185 178.085 ;
        RECT 54.815 177.645 55.510 178.275 ;
        RECT 55.715 177.475 56.025 178.275 ;
        RECT 56.195 178.125 56.365 179.155 ;
        RECT 56.640 179.025 57.395 179.275 ;
        RECT 57.565 179.100 57.895 179.345 ;
        RECT 58.500 179.225 58.815 180.025 ;
        RECT 59.080 179.670 60.160 179.840 ;
        RECT 56.640 178.990 57.410 179.025 ;
        RECT 56.640 178.980 57.425 178.990 ;
        RECT 56.535 178.965 57.430 178.980 ;
        RECT 56.535 178.950 57.450 178.965 ;
        RECT 56.535 178.940 57.470 178.950 ;
        RECT 56.535 178.930 57.495 178.940 ;
        RECT 56.535 178.900 57.565 178.930 ;
        RECT 56.535 178.870 57.585 178.900 ;
        RECT 56.535 178.840 57.605 178.870 ;
        RECT 56.535 178.815 57.635 178.840 ;
        RECT 56.535 178.780 57.670 178.815 ;
        RECT 56.535 178.775 57.700 178.780 ;
        RECT 56.535 178.380 56.765 178.775 ;
        RECT 57.310 178.770 57.700 178.775 ;
        RECT 57.335 178.760 57.700 178.770 ;
        RECT 57.350 178.755 57.700 178.760 ;
        RECT 57.365 178.750 57.700 178.755 ;
        RECT 58.065 178.750 58.325 179.200 ;
        RECT 59.080 179.055 59.250 179.670 ;
        RECT 57.365 178.745 58.325 178.750 ;
        RECT 57.375 178.735 58.325 178.745 ;
        RECT 57.385 178.730 58.325 178.735 ;
        RECT 57.395 178.720 58.325 178.730 ;
        RECT 57.400 178.710 58.325 178.720 ;
        RECT 57.405 178.705 58.325 178.710 ;
        RECT 57.415 178.690 58.325 178.705 ;
        RECT 57.420 178.675 58.325 178.690 ;
        RECT 57.430 178.650 58.325 178.675 ;
        RECT 56.935 178.180 57.265 178.605 ;
        RECT 56.195 177.645 56.455 178.125 ;
        RECT 56.625 177.475 56.875 178.015 ;
        RECT 57.045 177.695 57.265 178.180 ;
        RECT 57.435 178.580 58.325 178.650 ;
        RECT 57.435 177.855 57.605 178.580 ;
        RECT 57.775 178.025 58.325 178.410 ;
        RECT 58.495 178.045 58.765 179.055 ;
        RECT 58.935 178.885 59.250 179.055 ;
        RECT 58.935 178.215 59.105 178.885 ;
        RECT 59.420 178.715 59.655 179.395 ;
        RECT 59.825 178.885 60.160 179.670 ;
        RECT 61.255 178.885 61.595 179.855 ;
        RECT 61.765 178.885 61.935 180.025 ;
        RECT 62.205 179.225 62.455 180.025 ;
        RECT 63.100 179.055 63.430 179.855 ;
        RECT 63.730 179.225 64.060 180.025 ;
        RECT 64.230 179.055 64.560 179.855 ;
        RECT 62.125 178.885 64.560 179.055 ;
        RECT 64.935 178.935 68.445 180.025 ;
        RECT 59.275 178.385 59.655 178.715 ;
        RECT 59.825 178.385 60.160 178.715 ;
        RECT 61.255 178.275 61.430 178.885 ;
        RECT 62.125 178.635 62.295 178.885 ;
        RECT 61.600 178.465 62.295 178.635 ;
        RECT 62.470 178.465 62.890 178.665 ;
        RECT 63.060 178.465 63.390 178.665 ;
        RECT 63.560 178.465 63.890 178.665 ;
        RECT 58.935 178.045 60.160 178.215 ;
        RECT 57.435 177.685 58.325 177.855 ;
        RECT 58.565 177.475 58.895 177.875 ;
        RECT 59.065 177.775 59.235 178.045 ;
        RECT 59.405 177.475 59.735 177.875 ;
        RECT 59.905 177.775 60.160 178.045 ;
        RECT 61.255 177.645 61.595 178.275 ;
        RECT 61.765 177.475 62.015 178.275 ;
        RECT 62.205 178.125 63.430 178.295 ;
        RECT 62.205 177.645 62.535 178.125 ;
        RECT 62.705 177.475 62.930 177.935 ;
        RECT 63.100 177.645 63.430 178.125 ;
        RECT 64.060 178.255 64.230 178.885 ;
        RECT 64.415 178.465 64.765 178.715 ;
        RECT 64.060 177.645 64.560 178.255 ;
        RECT 64.935 178.245 66.585 178.765 ;
        RECT 66.755 178.415 68.445 178.935 ;
        RECT 68.625 178.885 68.955 180.025 ;
        RECT 69.485 179.055 69.815 179.840 ;
        RECT 69.135 178.885 69.815 179.055 ;
        RECT 70.005 179.055 70.335 179.840 ;
        RECT 70.005 178.885 70.685 179.055 ;
        RECT 70.865 178.885 71.195 180.025 ;
        RECT 71.375 178.935 74.885 180.025 ;
        RECT 75.055 178.935 76.265 180.025 ;
        RECT 68.615 178.465 68.965 178.715 ;
        RECT 69.135 178.285 69.305 178.885 ;
        RECT 69.475 178.465 69.825 178.715 ;
        RECT 69.995 178.465 70.345 178.715 ;
        RECT 70.515 178.285 70.685 178.885 ;
        RECT 70.855 178.465 71.205 178.715 ;
        RECT 64.935 177.475 68.445 178.245 ;
        RECT 68.625 177.475 68.895 178.285 ;
        RECT 69.065 177.645 69.395 178.285 ;
        RECT 69.565 177.475 69.805 178.285 ;
        RECT 70.015 177.475 70.255 178.285 ;
        RECT 70.425 177.645 70.755 178.285 ;
        RECT 70.925 177.475 71.195 178.285 ;
        RECT 71.375 178.245 73.025 178.765 ;
        RECT 73.195 178.415 74.885 178.935 ;
        RECT 71.375 177.475 74.885 178.245 ;
        RECT 75.055 178.225 75.575 178.765 ;
        RECT 75.745 178.395 76.265 178.935 ;
        RECT 76.435 178.860 76.725 180.025 ;
        RECT 76.895 179.590 82.240 180.025 ;
        RECT 82.415 179.590 87.760 180.025 ;
        RECT 75.055 177.475 76.265 178.225 ;
        RECT 76.435 177.475 76.725 178.200 ;
        RECT 78.480 178.020 78.820 178.850 ;
        RECT 80.300 178.340 80.650 179.590 ;
        RECT 84.000 178.020 84.340 178.850 ;
        RECT 85.820 178.340 86.170 179.590 ;
        RECT 87.935 178.935 89.145 180.025 ;
        RECT 87.935 178.225 88.455 178.765 ;
        RECT 88.625 178.395 89.145 178.935 ;
        RECT 89.315 178.935 90.525 180.025 ;
        RECT 89.315 178.395 89.835 178.935 ;
        RECT 90.005 178.225 90.525 178.765 ;
        RECT 76.895 177.475 82.240 178.020 ;
        RECT 82.415 177.475 87.760 178.020 ;
        RECT 87.935 177.475 89.145 178.225 ;
        RECT 89.315 177.475 90.525 178.225 ;
        RECT 11.950 177.305 90.610 177.475 ;
        RECT 12.035 176.555 13.245 177.305 ;
        RECT 13.415 176.760 18.760 177.305 ;
        RECT 19.400 176.800 19.735 177.305 ;
        RECT 12.035 176.015 12.555 176.555 ;
        RECT 12.725 175.845 13.245 176.385 ;
        RECT 15.000 175.930 15.340 176.760 ;
        RECT 19.905 176.735 20.145 177.110 ;
        RECT 20.425 176.975 20.595 177.120 ;
        RECT 20.425 176.780 20.800 176.975 ;
        RECT 21.160 176.810 21.555 177.305 ;
        RECT 12.035 174.755 13.245 175.845 ;
        RECT 16.820 175.190 17.170 176.440 ;
        RECT 19.455 175.775 19.755 176.625 ;
        RECT 19.925 176.585 20.145 176.735 ;
        RECT 19.925 176.255 20.460 176.585 ;
        RECT 20.630 176.445 20.800 176.780 ;
        RECT 21.725 176.615 21.965 177.135 ;
        RECT 22.155 176.760 27.500 177.305 ;
        RECT 27.675 176.760 33.020 177.305 ;
        RECT 19.925 175.605 20.160 176.255 ;
        RECT 20.630 176.085 21.615 176.445 ;
        RECT 19.485 175.375 20.160 175.605 ;
        RECT 20.330 176.065 21.615 176.085 ;
        RECT 20.330 175.915 21.190 176.065 ;
        RECT 13.415 174.755 18.760 175.190 ;
        RECT 19.485 174.945 19.655 175.375 ;
        RECT 19.825 174.755 20.155 175.205 ;
        RECT 20.330 174.970 20.615 175.915 ;
        RECT 21.790 175.810 21.965 176.615 ;
        RECT 23.740 175.930 24.080 176.760 ;
        RECT 20.790 175.435 21.485 175.745 ;
        RECT 20.795 174.755 21.480 175.225 ;
        RECT 21.660 175.025 21.965 175.810 ;
        RECT 25.560 175.190 25.910 176.440 ;
        RECT 29.260 175.930 29.600 176.760 ;
        RECT 33.195 176.535 36.705 177.305 ;
        RECT 37.795 176.580 38.085 177.305 ;
        RECT 38.255 176.535 41.765 177.305 ;
        RECT 41.935 176.555 43.145 177.305 ;
        RECT 31.080 175.190 31.430 176.440 ;
        RECT 33.195 176.015 34.845 176.535 ;
        RECT 35.015 175.845 36.705 176.365 ;
        RECT 38.255 176.015 39.905 176.535 ;
        RECT 22.155 174.755 27.500 175.190 ;
        RECT 27.675 174.755 33.020 175.190 ;
        RECT 33.195 174.755 36.705 175.845 ;
        RECT 37.795 174.755 38.085 175.920 ;
        RECT 40.075 175.845 41.765 176.365 ;
        RECT 41.935 176.015 42.455 176.555 ;
        RECT 43.335 176.495 43.575 177.305 ;
        RECT 43.745 176.495 44.075 177.135 ;
        RECT 44.245 176.495 44.515 177.305 ;
        RECT 44.695 176.760 50.040 177.305 ;
        RECT 50.215 176.760 55.560 177.305 ;
        RECT 55.735 176.760 61.080 177.305 ;
        RECT 42.625 175.845 43.145 176.385 ;
        RECT 43.315 176.065 43.665 176.315 ;
        RECT 43.835 175.895 44.005 176.495 ;
        RECT 44.175 176.065 44.525 176.315 ;
        RECT 46.280 175.930 46.620 176.760 ;
        RECT 38.255 174.755 41.765 175.845 ;
        RECT 41.935 174.755 43.145 175.845 ;
        RECT 43.325 175.725 44.005 175.895 ;
        RECT 43.325 174.940 43.655 175.725 ;
        RECT 44.185 174.755 44.515 175.895 ;
        RECT 48.100 175.190 48.450 176.440 ;
        RECT 51.800 175.930 52.140 176.760 ;
        RECT 53.620 175.190 53.970 176.440 ;
        RECT 57.320 175.930 57.660 176.760 ;
        RECT 61.255 176.535 62.925 177.305 ;
        RECT 63.555 176.580 63.845 177.305 ;
        RECT 64.015 176.535 66.605 177.305 ;
        RECT 59.140 175.190 59.490 176.440 ;
        RECT 61.255 176.015 62.005 176.535 ;
        RECT 62.175 175.845 62.925 176.365 ;
        RECT 64.015 176.015 65.225 176.535 ;
        RECT 66.835 176.485 67.045 177.305 ;
        RECT 67.215 176.505 67.545 177.135 ;
        RECT 44.695 174.755 50.040 175.190 ;
        RECT 50.215 174.755 55.560 175.190 ;
        RECT 55.735 174.755 61.080 175.190 ;
        RECT 61.255 174.755 62.925 175.845 ;
        RECT 63.555 174.755 63.845 175.920 ;
        RECT 65.395 175.845 66.605 176.365 ;
        RECT 67.215 175.905 67.465 176.505 ;
        RECT 67.715 176.485 67.945 177.305 ;
        RECT 69.095 176.495 69.335 177.305 ;
        RECT 69.505 176.495 69.835 177.135 ;
        RECT 70.005 176.495 70.275 177.305 ;
        RECT 70.465 176.495 70.735 177.305 ;
        RECT 70.905 176.495 71.235 177.135 ;
        RECT 71.405 176.495 71.645 177.305 ;
        RECT 71.835 176.505 72.530 177.135 ;
        RECT 72.735 176.505 73.045 177.305 ;
        RECT 73.215 176.760 78.560 177.305 ;
        RECT 78.735 176.760 84.080 177.305 ;
        RECT 67.635 176.065 67.965 176.315 ;
        RECT 69.075 176.065 69.425 176.315 ;
        RECT 64.015 174.755 66.605 175.845 ;
        RECT 66.835 174.755 67.045 175.895 ;
        RECT 67.215 174.925 67.545 175.905 ;
        RECT 69.595 175.895 69.765 176.495 ;
        RECT 69.935 176.065 70.285 176.315 ;
        RECT 70.455 176.065 70.805 176.315 ;
        RECT 70.975 175.895 71.145 176.495 ;
        RECT 72.355 176.455 72.530 176.505 ;
        RECT 71.315 176.065 71.665 176.315 ;
        RECT 71.855 176.065 72.190 176.315 ;
        RECT 72.360 175.905 72.530 176.455 ;
        RECT 72.700 176.065 73.035 176.335 ;
        RECT 74.800 175.930 75.140 176.760 ;
        RECT 67.715 174.755 67.945 175.895 ;
        RECT 69.085 175.725 69.765 175.895 ;
        RECT 69.085 174.940 69.415 175.725 ;
        RECT 69.945 174.755 70.275 175.895 ;
        RECT 70.465 174.755 70.795 175.895 ;
        RECT 70.975 175.725 71.655 175.895 ;
        RECT 71.325 174.940 71.655 175.725 ;
        RECT 71.835 174.755 72.095 175.895 ;
        RECT 72.265 174.925 72.595 175.905 ;
        RECT 72.765 174.755 73.045 175.895 ;
        RECT 76.620 175.190 76.970 176.440 ;
        RECT 80.320 175.930 80.660 176.760 ;
        RECT 84.255 176.535 87.765 177.305 ;
        RECT 87.935 176.555 89.145 177.305 ;
        RECT 89.315 176.555 90.525 177.305 ;
        RECT 100.630 176.790 106.370 176.800 ;
        RECT 82.140 175.190 82.490 176.440 ;
        RECT 84.255 176.015 85.905 176.535 ;
        RECT 86.075 175.845 87.765 176.365 ;
        RECT 87.935 176.015 88.455 176.555 ;
        RECT 88.625 175.845 89.145 176.385 ;
        RECT 73.215 174.755 78.560 175.190 ;
        RECT 78.735 174.755 84.080 175.190 ;
        RECT 84.255 174.755 87.765 175.845 ;
        RECT 87.935 174.755 89.145 175.845 ;
        RECT 89.315 175.845 89.835 176.385 ;
        RECT 90.005 176.015 90.525 176.555 ;
        RECT 100.140 176.630 106.370 176.790 ;
        RECT 89.315 174.755 90.525 175.845 ;
        RECT 11.950 174.585 90.610 174.755 ;
        RECT 12.035 173.495 13.245 174.585 ;
        RECT 13.415 174.150 18.760 174.585 ;
        RECT 18.935 174.150 24.280 174.585 ;
        RECT 12.035 172.785 12.555 173.325 ;
        RECT 12.725 172.955 13.245 173.495 ;
        RECT 12.035 172.035 13.245 172.785 ;
        RECT 15.000 172.580 15.340 173.410 ;
        RECT 16.820 172.900 17.170 174.150 ;
        RECT 20.520 172.580 20.860 173.410 ;
        RECT 22.340 172.900 22.690 174.150 ;
        RECT 24.915 173.420 25.205 174.585 ;
        RECT 25.375 173.495 27.965 174.585 ;
        RECT 28.595 174.030 29.200 174.585 ;
        RECT 29.375 174.075 29.855 174.415 ;
        RECT 30.025 174.040 30.280 174.585 ;
        RECT 28.595 173.930 29.210 174.030 ;
        RECT 29.025 173.905 29.210 173.930 ;
        RECT 25.375 172.805 26.585 173.325 ;
        RECT 26.755 172.975 27.965 173.495 ;
        RECT 28.595 173.310 28.855 173.760 ;
        RECT 29.025 173.660 29.355 173.905 ;
        RECT 29.525 173.585 30.280 173.835 ;
        RECT 30.450 173.715 30.725 174.415 ;
        RECT 29.510 173.550 30.280 173.585 ;
        RECT 29.495 173.540 30.280 173.550 ;
        RECT 29.490 173.525 30.385 173.540 ;
        RECT 29.470 173.510 30.385 173.525 ;
        RECT 29.450 173.500 30.385 173.510 ;
        RECT 29.425 173.490 30.385 173.500 ;
        RECT 29.355 173.460 30.385 173.490 ;
        RECT 29.335 173.430 30.385 173.460 ;
        RECT 29.315 173.400 30.385 173.430 ;
        RECT 29.285 173.375 30.385 173.400 ;
        RECT 29.250 173.340 30.385 173.375 ;
        RECT 29.220 173.335 30.385 173.340 ;
        RECT 29.220 173.330 29.610 173.335 ;
        RECT 29.220 173.320 29.585 173.330 ;
        RECT 29.220 173.315 29.570 173.320 ;
        RECT 29.220 173.310 29.555 173.315 ;
        RECT 28.595 173.305 29.555 173.310 ;
        RECT 28.595 173.295 29.545 173.305 ;
        RECT 28.595 173.290 29.535 173.295 ;
        RECT 28.595 173.280 29.525 173.290 ;
        RECT 28.595 173.270 29.520 173.280 ;
        RECT 28.595 173.265 29.515 173.270 ;
        RECT 28.595 173.250 29.505 173.265 ;
        RECT 28.595 173.235 29.500 173.250 ;
        RECT 28.595 173.210 29.490 173.235 ;
        RECT 28.595 173.140 29.485 173.210 ;
        RECT 13.415 172.035 18.760 172.580 ;
        RECT 18.935 172.035 24.280 172.580 ;
        RECT 24.915 172.035 25.205 172.760 ;
        RECT 25.375 172.035 27.965 172.805 ;
        RECT 28.595 172.585 29.145 172.970 ;
        RECT 29.315 172.415 29.485 173.140 ;
        RECT 28.595 172.245 29.485 172.415 ;
        RECT 29.655 172.740 29.985 173.165 ;
        RECT 30.155 172.940 30.385 173.335 ;
        RECT 29.655 172.255 29.875 172.740 ;
        RECT 30.555 172.685 30.725 173.715 ;
        RECT 30.045 172.035 30.295 172.575 ;
        RECT 30.465 172.205 30.725 172.685 ;
        RECT 30.895 173.715 31.170 174.415 ;
        RECT 31.340 174.040 31.595 174.585 ;
        RECT 31.765 174.075 32.245 174.415 ;
        RECT 32.420 174.030 33.025 174.585 ;
        RECT 32.410 173.930 33.025 174.030 ;
        RECT 32.410 173.905 32.595 173.930 ;
        RECT 30.895 172.685 31.065 173.715 ;
        RECT 31.340 173.585 32.095 173.835 ;
        RECT 32.265 173.660 32.595 173.905 ;
        RECT 31.340 173.550 32.110 173.585 ;
        RECT 31.340 173.540 32.125 173.550 ;
        RECT 31.235 173.525 32.130 173.540 ;
        RECT 31.235 173.510 32.150 173.525 ;
        RECT 31.235 173.500 32.170 173.510 ;
        RECT 31.235 173.490 32.195 173.500 ;
        RECT 31.235 173.460 32.265 173.490 ;
        RECT 31.235 173.430 32.285 173.460 ;
        RECT 31.235 173.400 32.305 173.430 ;
        RECT 31.235 173.375 32.335 173.400 ;
        RECT 31.235 173.340 32.370 173.375 ;
        RECT 31.235 173.335 32.400 173.340 ;
        RECT 31.235 172.940 31.465 173.335 ;
        RECT 32.010 173.330 32.400 173.335 ;
        RECT 32.035 173.320 32.400 173.330 ;
        RECT 32.050 173.315 32.400 173.320 ;
        RECT 32.065 173.310 32.400 173.315 ;
        RECT 32.765 173.310 33.025 173.760 ;
        RECT 33.195 173.495 35.785 174.585 ;
        RECT 36.665 173.855 36.960 174.585 ;
        RECT 37.130 173.685 37.390 174.410 ;
        RECT 37.560 173.855 37.820 174.585 ;
        RECT 37.990 173.685 38.250 174.410 ;
        RECT 38.420 173.855 38.680 174.585 ;
        RECT 38.850 173.685 39.110 174.410 ;
        RECT 39.280 173.855 39.540 174.585 ;
        RECT 39.710 173.685 39.970 174.410 ;
        RECT 32.065 173.305 33.025 173.310 ;
        RECT 32.075 173.295 33.025 173.305 ;
        RECT 32.085 173.290 33.025 173.295 ;
        RECT 32.095 173.280 33.025 173.290 ;
        RECT 32.100 173.270 33.025 173.280 ;
        RECT 32.105 173.265 33.025 173.270 ;
        RECT 32.115 173.250 33.025 173.265 ;
        RECT 32.120 173.235 33.025 173.250 ;
        RECT 32.130 173.210 33.025 173.235 ;
        RECT 31.635 172.740 31.965 173.165 ;
        RECT 31.715 172.715 31.965 172.740 ;
        RECT 30.895 172.205 31.155 172.685 ;
        RECT 31.325 172.035 31.575 172.575 ;
        RECT 31.745 172.255 31.965 172.715 ;
        RECT 32.135 173.140 33.025 173.210 ;
        RECT 32.135 172.415 32.305 173.140 ;
        RECT 32.475 172.585 33.025 172.970 ;
        RECT 33.195 172.805 34.405 173.325 ;
        RECT 34.575 172.975 35.785 173.495 ;
        RECT 36.660 173.445 39.970 173.685 ;
        RECT 40.140 173.475 40.400 174.585 ;
        RECT 36.660 172.855 37.630 173.445 ;
        RECT 40.570 173.275 40.820 174.410 ;
        RECT 41.000 173.475 41.295 174.585 ;
        RECT 41.475 173.715 41.750 174.415 ;
        RECT 41.920 174.040 42.175 174.585 ;
        RECT 42.345 174.075 42.825 174.415 ;
        RECT 43.000 174.030 43.605 174.585 ;
        RECT 42.990 173.930 43.605 174.030 ;
        RECT 42.990 173.905 43.175 173.930 ;
        RECT 37.800 173.025 40.820 173.275 ;
        RECT 32.135 172.245 33.025 172.415 ;
        RECT 33.195 172.035 35.785 172.805 ;
        RECT 36.660 172.685 39.970 172.855 ;
        RECT 36.660 172.035 36.960 172.515 ;
        RECT 37.130 172.230 37.390 172.685 ;
        RECT 37.560 172.035 37.820 172.515 ;
        RECT 37.990 172.230 38.250 172.685 ;
        RECT 38.420 172.035 38.680 172.515 ;
        RECT 38.850 172.230 39.110 172.685 ;
        RECT 39.280 172.035 39.540 172.515 ;
        RECT 39.710 172.230 39.970 172.685 ;
        RECT 40.140 172.035 40.400 172.560 ;
        RECT 40.570 172.215 40.820 173.025 ;
        RECT 40.990 172.665 41.305 173.275 ;
        RECT 41.475 172.685 41.645 173.715 ;
        RECT 41.920 173.585 42.675 173.835 ;
        RECT 42.845 173.660 43.175 173.905 ;
        RECT 41.920 173.550 42.690 173.585 ;
        RECT 41.920 173.540 42.705 173.550 ;
        RECT 41.815 173.525 42.710 173.540 ;
        RECT 41.815 173.510 42.730 173.525 ;
        RECT 41.815 173.500 42.750 173.510 ;
        RECT 41.815 173.490 42.775 173.500 ;
        RECT 41.815 173.460 42.845 173.490 ;
        RECT 41.815 173.430 42.865 173.460 ;
        RECT 41.815 173.400 42.885 173.430 ;
        RECT 41.815 173.375 42.915 173.400 ;
        RECT 41.815 173.340 42.950 173.375 ;
        RECT 41.815 173.335 42.980 173.340 ;
        RECT 41.815 172.940 42.045 173.335 ;
        RECT 42.590 173.330 42.980 173.335 ;
        RECT 42.615 173.320 42.980 173.330 ;
        RECT 42.630 173.315 42.980 173.320 ;
        RECT 42.645 173.310 42.980 173.315 ;
        RECT 43.345 173.310 43.605 173.760 ;
        RECT 42.645 173.305 43.605 173.310 ;
        RECT 42.655 173.295 43.605 173.305 ;
        RECT 42.665 173.290 43.605 173.295 ;
        RECT 42.675 173.280 43.605 173.290 ;
        RECT 42.680 173.270 43.605 173.280 ;
        RECT 42.685 173.265 43.605 173.270 ;
        RECT 42.695 173.250 43.605 173.265 ;
        RECT 42.700 173.235 43.605 173.250 ;
        RECT 42.710 173.210 43.605 173.235 ;
        RECT 42.215 172.740 42.545 173.165 ;
        RECT 41.000 172.035 41.245 172.495 ;
        RECT 41.475 172.205 41.735 172.685 ;
        RECT 41.905 172.035 42.155 172.575 ;
        RECT 42.325 172.255 42.545 172.740 ;
        RECT 42.715 173.140 43.605 173.210 ;
        RECT 43.775 173.715 44.050 174.415 ;
        RECT 44.220 174.040 44.475 174.585 ;
        RECT 44.645 174.075 45.125 174.415 ;
        RECT 45.300 174.030 45.905 174.585 ;
        RECT 45.290 173.930 45.905 174.030 ;
        RECT 46.085 173.975 46.415 174.405 ;
        RECT 46.595 174.145 46.790 174.585 ;
        RECT 46.960 173.975 47.290 174.405 ;
        RECT 45.290 173.905 45.475 173.930 ;
        RECT 42.715 172.415 42.885 173.140 ;
        RECT 43.055 172.585 43.605 172.970 ;
        RECT 43.775 172.685 43.945 173.715 ;
        RECT 44.220 173.585 44.975 173.835 ;
        RECT 45.145 173.660 45.475 173.905 ;
        RECT 46.085 173.805 47.290 173.975 ;
        RECT 44.220 173.550 44.990 173.585 ;
        RECT 44.220 173.540 45.005 173.550 ;
        RECT 44.115 173.525 45.010 173.540 ;
        RECT 44.115 173.510 45.030 173.525 ;
        RECT 44.115 173.500 45.050 173.510 ;
        RECT 44.115 173.490 45.075 173.500 ;
        RECT 44.115 173.460 45.145 173.490 ;
        RECT 44.115 173.430 45.165 173.460 ;
        RECT 44.115 173.400 45.185 173.430 ;
        RECT 44.115 173.375 45.215 173.400 ;
        RECT 44.115 173.340 45.250 173.375 ;
        RECT 44.115 173.335 45.280 173.340 ;
        RECT 44.115 172.940 44.345 173.335 ;
        RECT 44.890 173.330 45.280 173.335 ;
        RECT 44.915 173.320 45.280 173.330 ;
        RECT 44.930 173.315 45.280 173.320 ;
        RECT 44.945 173.310 45.280 173.315 ;
        RECT 45.645 173.310 45.905 173.760 ;
        RECT 46.085 173.475 46.980 173.805 ;
        RECT 47.460 173.635 47.735 174.405 ;
        RECT 44.945 173.305 45.905 173.310 ;
        RECT 44.955 173.295 45.905 173.305 ;
        RECT 44.965 173.290 45.905 173.295 ;
        RECT 44.975 173.280 45.905 173.290 ;
        RECT 44.980 173.270 45.905 173.280 ;
        RECT 47.150 173.445 47.735 173.635 ;
        RECT 47.915 173.495 50.505 174.585 ;
        RECT 44.985 173.265 45.905 173.270 ;
        RECT 44.995 173.250 45.905 173.265 ;
        RECT 45.000 173.235 45.905 173.250 ;
        RECT 45.010 173.210 45.905 173.235 ;
        RECT 44.515 172.740 44.845 173.165 ;
        RECT 42.715 172.245 43.605 172.415 ;
        RECT 43.775 172.205 44.035 172.685 ;
        RECT 44.205 172.035 44.455 172.575 ;
        RECT 44.625 172.255 44.845 172.740 ;
        RECT 45.015 173.140 45.905 173.210 ;
        RECT 45.015 172.415 45.185 173.140 ;
        RECT 45.355 172.585 45.905 172.970 ;
        RECT 46.090 172.945 46.385 173.275 ;
        RECT 46.565 172.945 46.980 173.275 ;
        RECT 45.015 172.245 45.905 172.415 ;
        RECT 46.085 172.035 46.385 172.765 ;
        RECT 46.565 172.325 46.795 172.945 ;
        RECT 47.150 172.775 47.325 173.445 ;
        RECT 46.995 172.595 47.325 172.775 ;
        RECT 47.495 172.625 47.735 173.275 ;
        RECT 47.915 172.805 49.125 173.325 ;
        RECT 49.295 172.975 50.505 173.495 ;
        RECT 50.675 173.420 50.965 174.585 ;
        RECT 51.135 173.615 51.405 174.385 ;
        RECT 51.575 173.805 51.905 174.585 ;
        RECT 52.110 173.980 52.295 174.385 ;
        RECT 52.465 174.160 52.800 174.585 ;
        RECT 52.980 174.160 53.315 174.585 ;
        RECT 53.485 173.980 53.670 174.385 ;
        RECT 52.110 173.805 52.775 173.980 ;
        RECT 51.135 173.445 52.265 173.615 ;
        RECT 46.995 172.215 47.220 172.595 ;
        RECT 47.390 172.035 47.720 172.425 ;
        RECT 47.915 172.035 50.505 172.805 ;
        RECT 50.675 172.035 50.965 172.760 ;
        RECT 51.135 172.535 51.305 173.445 ;
        RECT 51.475 172.695 51.835 173.275 ;
        RECT 52.015 172.945 52.265 173.445 ;
        RECT 52.435 172.775 52.775 173.805 ;
        RECT 52.090 172.605 52.775 172.775 ;
        RECT 53.005 173.805 53.670 173.980 ;
        RECT 53.875 173.805 54.205 174.585 ;
        RECT 53.005 172.775 53.345 173.805 ;
        RECT 54.375 173.615 54.645 174.385 ;
        RECT 53.515 173.445 54.645 173.615 ;
        RECT 54.815 173.495 56.025 174.585 ;
        RECT 53.515 172.945 53.765 173.445 ;
        RECT 53.005 172.605 53.690 172.775 ;
        RECT 53.945 172.695 54.305 173.275 ;
        RECT 51.135 172.205 51.395 172.535 ;
        RECT 51.605 172.035 51.880 172.515 ;
        RECT 52.090 172.205 52.295 172.605 ;
        RECT 52.465 172.035 52.800 172.435 ;
        RECT 52.980 172.035 53.315 172.435 ;
        RECT 53.485 172.205 53.690 172.605 ;
        RECT 54.475 172.535 54.645 173.445 ;
        RECT 53.900 172.035 54.175 172.515 ;
        RECT 54.385 172.205 54.645 172.535 ;
        RECT 54.815 172.785 55.335 173.325 ;
        RECT 55.505 172.955 56.025 173.495 ;
        RECT 56.205 173.445 56.535 174.585 ;
        RECT 57.065 173.615 57.395 174.400 ;
        RECT 56.715 173.445 57.395 173.615 ;
        RECT 57.575 173.735 57.835 174.415 ;
        RECT 58.005 173.805 58.255 174.585 ;
        RECT 58.505 174.035 58.755 174.415 ;
        RECT 58.925 174.205 59.280 174.585 ;
        RECT 60.285 174.195 60.620 174.415 ;
        RECT 59.885 174.035 60.115 174.075 ;
        RECT 58.505 173.835 60.115 174.035 ;
        RECT 58.505 173.825 59.340 173.835 ;
        RECT 59.930 173.745 60.115 173.835 ;
        RECT 56.195 173.025 56.545 173.275 ;
        RECT 56.715 172.845 56.885 173.445 ;
        RECT 57.055 173.025 57.405 173.275 ;
        RECT 54.815 172.035 56.025 172.785 ;
        RECT 56.205 172.035 56.475 172.845 ;
        RECT 56.645 172.205 56.975 172.845 ;
        RECT 57.145 172.035 57.385 172.845 ;
        RECT 57.575 172.535 57.745 173.735 ;
        RECT 59.445 173.635 59.775 173.665 ;
        RECT 57.975 173.575 59.775 173.635 ;
        RECT 60.365 173.575 60.620 174.195 ;
        RECT 61.295 174.125 61.510 174.585 ;
        RECT 61.680 173.955 62.010 174.415 ;
        RECT 57.915 173.465 60.620 173.575 ;
        RECT 57.915 173.430 58.115 173.465 ;
        RECT 57.915 172.855 58.085 173.430 ;
        RECT 59.445 173.405 60.620 173.465 ;
        RECT 60.840 173.785 62.010 173.955 ;
        RECT 62.180 173.785 62.430 174.585 ;
        RECT 58.315 172.990 58.725 173.295 ;
        RECT 58.895 173.025 59.225 173.235 ;
        RECT 57.915 172.735 58.185 172.855 ;
        RECT 57.915 172.690 58.760 172.735 ;
        RECT 58.005 172.565 58.760 172.690 ;
        RECT 59.015 172.625 59.225 173.025 ;
        RECT 59.470 173.025 59.945 173.235 ;
        RECT 60.135 173.025 60.625 173.225 ;
        RECT 59.470 172.625 59.690 173.025 ;
        RECT 57.575 172.205 57.835 172.535 ;
        RECT 58.590 172.415 58.760 172.565 ;
        RECT 58.005 172.035 58.335 172.395 ;
        RECT 58.590 172.205 59.890 172.415 ;
        RECT 60.165 172.035 60.620 172.800 ;
        RECT 60.840 172.495 61.210 173.785 ;
        RECT 62.640 173.615 62.920 173.775 ;
        RECT 61.585 173.445 62.920 173.615 ;
        RECT 63.095 173.495 64.765 174.585 ;
        RECT 61.585 173.275 61.755 173.445 ;
        RECT 61.380 173.025 61.755 173.275 ;
        RECT 61.925 173.025 62.400 173.265 ;
        RECT 62.570 173.025 62.920 173.265 ;
        RECT 61.585 172.855 61.755 173.025 ;
        RECT 61.585 172.685 62.920 172.855 ;
        RECT 60.840 172.205 61.590 172.495 ;
        RECT 62.100 172.035 62.430 172.495 ;
        RECT 62.650 172.475 62.920 172.685 ;
        RECT 63.095 172.805 63.845 173.325 ;
        RECT 64.015 172.975 64.765 173.495 ;
        RECT 65.395 174.155 65.735 174.415 ;
        RECT 63.095 172.035 64.765 172.805 ;
        RECT 65.395 172.755 65.655 174.155 ;
        RECT 65.905 173.785 66.235 174.585 ;
        RECT 66.700 173.615 66.950 174.415 ;
        RECT 67.135 173.865 67.465 174.585 ;
        RECT 67.685 173.615 67.935 174.415 ;
        RECT 68.105 174.205 68.440 174.585 ;
        RECT 65.845 173.445 68.035 173.615 ;
        RECT 65.845 173.275 66.160 173.445 ;
        RECT 65.830 173.025 66.160 173.275 ;
        RECT 65.395 172.245 65.735 172.755 ;
        RECT 65.905 172.035 66.175 172.835 ;
        RECT 66.355 172.305 66.635 173.275 ;
        RECT 66.815 172.305 67.115 173.275 ;
        RECT 67.295 172.310 67.645 173.275 ;
        RECT 67.865 172.535 68.035 173.445 ;
        RECT 68.205 172.715 68.445 174.025 ;
        RECT 68.615 173.865 69.075 174.415 ;
        RECT 69.265 173.865 69.595 174.585 ;
        RECT 67.865 172.205 68.360 172.535 ;
        RECT 68.615 172.495 68.865 173.865 ;
        RECT 69.795 173.695 70.095 174.245 ;
        RECT 70.265 173.915 70.545 174.585 ;
        RECT 70.920 174.205 71.255 174.585 ;
        RECT 69.155 173.525 70.095 173.695 ;
        RECT 69.155 173.275 69.325 173.525 ;
        RECT 70.465 173.275 70.730 173.635 ;
        RECT 69.035 172.945 69.325 173.275 ;
        RECT 69.495 173.025 69.835 173.275 ;
        RECT 70.055 173.025 70.730 173.275 ;
        RECT 69.155 172.855 69.325 172.945 ;
        RECT 69.155 172.665 70.545 172.855 ;
        RECT 70.915 172.715 71.155 174.025 ;
        RECT 71.425 173.615 71.675 174.415 ;
        RECT 71.895 173.865 72.225 174.585 ;
        RECT 72.410 173.615 72.660 174.415 ;
        RECT 73.125 173.785 73.455 174.585 ;
        RECT 73.625 174.155 73.965 174.415 ;
        RECT 71.325 173.445 73.515 173.615 ;
        RECT 68.615 172.205 69.175 172.495 ;
        RECT 69.345 172.035 69.595 172.495 ;
        RECT 70.215 172.305 70.545 172.665 ;
        RECT 71.325 172.535 71.495 173.445 ;
        RECT 73.200 173.275 73.515 173.445 ;
        RECT 71.000 172.205 71.495 172.535 ;
        RECT 71.715 172.310 72.065 173.275 ;
        RECT 72.245 172.305 72.545 173.275 ;
        RECT 72.725 172.305 73.005 173.275 ;
        RECT 73.200 173.025 73.530 173.275 ;
        RECT 73.185 172.035 73.455 172.835 ;
        RECT 73.705 172.755 73.965 174.155 ;
        RECT 73.625 172.245 73.965 172.755 ;
        RECT 74.170 173.795 74.705 174.415 ;
        RECT 74.170 172.775 74.485 173.795 ;
        RECT 74.875 173.785 75.205 174.585 ;
        RECT 75.690 173.615 76.080 173.790 ;
        RECT 74.655 173.445 76.080 173.615 ;
        RECT 74.655 172.945 74.825 173.445 ;
        RECT 74.170 172.205 74.785 172.775 ;
        RECT 75.075 172.715 75.340 173.275 ;
        RECT 75.510 172.545 75.680 173.445 ;
        RECT 76.435 173.420 76.725 174.585 ;
        RECT 76.985 173.915 77.155 174.415 ;
        RECT 77.325 174.085 77.655 174.585 ;
        RECT 76.985 173.745 77.650 173.915 ;
        RECT 75.850 172.715 76.205 173.275 ;
        RECT 76.900 172.925 77.250 173.575 ;
        RECT 74.955 172.035 75.170 172.545 ;
        RECT 75.400 172.215 75.680 172.545 ;
        RECT 75.860 172.035 76.100 172.545 ;
        RECT 76.435 172.035 76.725 172.760 ;
        RECT 77.420 172.755 77.650 173.745 ;
        RECT 76.985 172.585 77.650 172.755 ;
        RECT 76.985 172.295 77.155 172.585 ;
        RECT 77.325 172.035 77.655 172.415 ;
        RECT 77.825 172.295 78.010 174.415 ;
        RECT 78.250 174.125 78.515 174.585 ;
        RECT 78.685 173.990 78.935 174.415 ;
        RECT 79.145 174.140 80.250 174.310 ;
        RECT 78.630 173.860 78.935 173.990 ;
        RECT 78.180 172.665 78.460 173.615 ;
        RECT 78.630 172.755 78.800 173.860 ;
        RECT 78.970 173.075 79.210 173.670 ;
        RECT 79.380 173.605 79.910 173.970 ;
        RECT 79.380 172.905 79.550 173.605 ;
        RECT 80.080 173.525 80.250 174.140 ;
        RECT 80.420 173.785 80.590 174.585 ;
        RECT 80.760 174.085 81.010 174.415 ;
        RECT 81.235 174.115 82.120 174.285 ;
        RECT 80.080 173.435 80.590 173.525 ;
        RECT 78.630 172.625 78.855 172.755 ;
        RECT 79.025 172.685 79.550 172.905 ;
        RECT 79.720 173.265 80.590 173.435 ;
        RECT 78.265 172.035 78.515 172.495 ;
        RECT 78.685 172.485 78.855 172.625 ;
        RECT 79.720 172.485 79.890 173.265 ;
        RECT 80.420 173.195 80.590 173.265 ;
        RECT 80.100 173.015 80.300 173.045 ;
        RECT 80.760 173.015 80.930 174.085 ;
        RECT 81.100 173.195 81.290 173.915 ;
        RECT 80.100 172.715 80.930 173.015 ;
        RECT 81.460 172.985 81.780 173.945 ;
        RECT 78.685 172.315 79.020 172.485 ;
        RECT 79.215 172.315 79.890 172.485 ;
        RECT 80.210 172.035 80.580 172.535 ;
        RECT 80.760 172.485 80.930 172.715 ;
        RECT 81.315 172.655 81.780 172.985 ;
        RECT 81.950 173.275 82.120 174.115 ;
        RECT 82.300 174.085 82.615 174.585 ;
        RECT 82.845 173.855 83.185 174.415 ;
        RECT 82.290 173.480 83.185 173.855 ;
        RECT 83.355 173.575 83.525 174.585 ;
        RECT 82.995 173.275 83.185 173.480 ;
        RECT 83.695 173.525 84.025 174.370 ;
        RECT 83.695 173.445 84.085 173.525 ;
        RECT 84.255 173.495 87.765 174.585 ;
        RECT 87.935 173.495 89.145 174.585 ;
        RECT 83.870 173.395 84.085 173.445 ;
        RECT 81.950 172.945 82.825 173.275 ;
        RECT 82.995 172.945 83.745 173.275 ;
        RECT 81.950 172.485 82.120 172.945 ;
        RECT 82.995 172.775 83.195 172.945 ;
        RECT 83.915 172.815 84.085 173.395 ;
        RECT 83.860 172.775 84.085 172.815 ;
        RECT 80.760 172.315 81.165 172.485 ;
        RECT 81.335 172.315 82.120 172.485 ;
        RECT 82.395 172.035 82.605 172.565 ;
        RECT 82.865 172.250 83.195 172.775 ;
        RECT 83.705 172.690 84.085 172.775 ;
        RECT 84.255 172.805 85.905 173.325 ;
        RECT 86.075 172.975 87.765 173.495 ;
        RECT 83.365 172.035 83.535 172.645 ;
        RECT 83.705 172.255 84.035 172.690 ;
        RECT 84.255 172.035 87.765 172.805 ;
        RECT 87.935 172.785 88.455 173.325 ;
        RECT 88.625 172.955 89.145 173.495 ;
        RECT 89.315 173.495 90.525 174.585 ;
        RECT 100.140 174.370 100.810 176.630 ;
        RECT 101.480 176.060 105.520 176.230 ;
        RECT 101.140 175.000 101.310 176.000 ;
        RECT 105.690 175.000 105.860 176.000 ;
        RECT 101.480 174.770 105.520 174.940 ;
        RECT 106.200 174.370 106.370 176.630 ;
        RECT 100.140 174.200 106.370 174.370 ;
        RECT 89.315 172.955 89.835 173.495 ;
        RECT 90.005 172.785 90.525 173.325 ;
        RECT 87.935 172.035 89.145 172.785 ;
        RECT 89.315 172.035 90.525 172.785 ;
        RECT 11.950 171.865 90.610 172.035 ;
        RECT 12.035 171.115 13.245 171.865 ;
        RECT 13.415 171.320 18.760 171.865 ;
        RECT 12.035 170.575 12.555 171.115 ;
        RECT 12.725 170.405 13.245 170.945 ;
        RECT 15.000 170.490 15.340 171.320 ;
        RECT 18.935 171.095 20.605 171.865 ;
        RECT 20.865 171.315 21.035 171.605 ;
        RECT 21.205 171.485 21.535 171.865 ;
        RECT 20.865 171.145 21.530 171.315 ;
        RECT 12.035 169.315 13.245 170.405 ;
        RECT 16.820 169.750 17.170 171.000 ;
        RECT 18.935 170.575 19.685 171.095 ;
        RECT 19.855 170.405 20.605 170.925 ;
        RECT 13.415 169.315 18.760 169.750 ;
        RECT 18.935 169.315 20.605 170.405 ;
        RECT 20.780 170.325 21.130 170.975 ;
        RECT 21.300 170.155 21.530 171.145 ;
        RECT 20.865 169.985 21.530 170.155 ;
        RECT 20.865 169.485 21.035 169.985 ;
        RECT 21.205 169.315 21.535 169.815 ;
        RECT 21.705 169.485 21.890 171.605 ;
        RECT 22.145 171.405 22.395 171.865 ;
        RECT 22.565 171.415 22.900 171.585 ;
        RECT 23.095 171.415 23.770 171.585 ;
        RECT 22.565 171.275 22.735 171.415 ;
        RECT 22.060 170.285 22.340 171.235 ;
        RECT 22.510 171.145 22.735 171.275 ;
        RECT 22.510 170.040 22.680 171.145 ;
        RECT 22.905 170.995 23.430 171.215 ;
        RECT 22.850 170.230 23.090 170.825 ;
        RECT 23.260 170.295 23.430 170.995 ;
        RECT 23.600 170.635 23.770 171.415 ;
        RECT 24.090 171.365 24.460 171.865 ;
        RECT 24.640 171.415 25.045 171.585 ;
        RECT 25.215 171.415 26.000 171.585 ;
        RECT 24.640 171.185 24.810 171.415 ;
        RECT 23.980 170.885 24.810 171.185 ;
        RECT 25.195 170.915 25.660 171.245 ;
        RECT 23.980 170.855 24.180 170.885 ;
        RECT 24.300 170.635 24.470 170.705 ;
        RECT 23.600 170.465 24.470 170.635 ;
        RECT 23.960 170.375 24.470 170.465 ;
        RECT 22.510 169.910 22.815 170.040 ;
        RECT 23.260 169.930 23.790 170.295 ;
        RECT 22.130 169.315 22.395 169.775 ;
        RECT 22.565 169.485 22.815 169.910 ;
        RECT 23.960 169.760 24.130 170.375 ;
        RECT 23.025 169.590 24.130 169.760 ;
        RECT 24.300 169.315 24.470 170.115 ;
        RECT 24.640 169.815 24.810 170.885 ;
        RECT 24.980 169.985 25.170 170.705 ;
        RECT 25.340 169.955 25.660 170.915 ;
        RECT 25.830 170.955 26.000 171.415 ;
        RECT 26.275 171.335 26.485 171.865 ;
        RECT 26.745 171.125 27.075 171.650 ;
        RECT 27.245 171.255 27.415 171.865 ;
        RECT 27.585 171.210 27.915 171.645 ;
        RECT 27.585 171.125 27.965 171.210 ;
        RECT 26.875 170.955 27.075 171.125 ;
        RECT 27.740 171.085 27.965 171.125 ;
        RECT 25.830 170.625 26.705 170.955 ;
        RECT 26.875 170.625 27.625 170.955 ;
        RECT 24.640 169.485 24.890 169.815 ;
        RECT 25.830 169.785 26.000 170.625 ;
        RECT 26.875 170.420 27.065 170.625 ;
        RECT 27.795 170.505 27.965 171.085 ;
        RECT 28.135 171.065 28.445 171.865 ;
        RECT 28.650 171.065 29.345 171.695 ;
        RECT 29.605 171.315 29.775 171.605 ;
        RECT 29.945 171.485 30.275 171.865 ;
        RECT 29.605 171.145 30.270 171.315 ;
        RECT 28.145 170.625 28.480 170.895 ;
        RECT 27.750 170.455 27.965 170.505 ;
        RECT 28.650 170.465 28.820 171.065 ;
        RECT 28.990 170.625 29.325 170.875 ;
        RECT 26.170 170.045 27.065 170.420 ;
        RECT 27.575 170.375 27.965 170.455 ;
        RECT 25.115 169.615 26.000 169.785 ;
        RECT 26.180 169.315 26.495 169.815 ;
        RECT 26.725 169.485 27.065 170.045 ;
        RECT 27.235 169.315 27.405 170.325 ;
        RECT 27.575 169.530 27.905 170.375 ;
        RECT 28.135 169.315 28.415 170.455 ;
        RECT 28.585 169.485 28.915 170.465 ;
        RECT 29.085 169.315 29.345 170.455 ;
        RECT 29.520 170.325 29.870 170.975 ;
        RECT 30.040 170.155 30.270 171.145 ;
        RECT 29.605 169.985 30.270 170.155 ;
        RECT 29.605 169.485 29.775 169.985 ;
        RECT 29.945 169.315 30.275 169.815 ;
        RECT 30.445 169.485 30.630 171.605 ;
        RECT 30.885 171.405 31.135 171.865 ;
        RECT 31.305 171.415 31.640 171.585 ;
        RECT 31.835 171.415 32.510 171.585 ;
        RECT 31.305 171.275 31.475 171.415 ;
        RECT 30.800 170.285 31.080 171.235 ;
        RECT 31.250 171.145 31.475 171.275 ;
        RECT 31.250 170.040 31.420 171.145 ;
        RECT 31.645 170.995 32.170 171.215 ;
        RECT 31.590 170.230 31.830 170.825 ;
        RECT 32.000 170.295 32.170 170.995 ;
        RECT 32.340 170.635 32.510 171.415 ;
        RECT 32.830 171.365 33.200 171.865 ;
        RECT 33.380 171.415 33.785 171.585 ;
        RECT 33.955 171.415 34.740 171.585 ;
        RECT 33.380 171.185 33.550 171.415 ;
        RECT 32.720 170.885 33.550 171.185 ;
        RECT 33.935 170.915 34.400 171.245 ;
        RECT 32.720 170.855 32.920 170.885 ;
        RECT 33.040 170.635 33.210 170.705 ;
        RECT 32.340 170.465 33.210 170.635 ;
        RECT 32.700 170.375 33.210 170.465 ;
        RECT 31.250 169.910 31.555 170.040 ;
        RECT 32.000 169.930 32.530 170.295 ;
        RECT 30.870 169.315 31.135 169.775 ;
        RECT 31.305 169.485 31.555 169.910 ;
        RECT 32.700 169.760 32.870 170.375 ;
        RECT 31.765 169.590 32.870 169.760 ;
        RECT 33.040 169.315 33.210 170.115 ;
        RECT 33.380 169.815 33.550 170.885 ;
        RECT 33.720 169.985 33.910 170.705 ;
        RECT 34.080 169.955 34.400 170.915 ;
        RECT 34.570 170.955 34.740 171.415 ;
        RECT 35.015 171.335 35.225 171.865 ;
        RECT 35.485 171.125 35.815 171.650 ;
        RECT 35.985 171.255 36.155 171.865 ;
        RECT 36.325 171.210 36.655 171.645 ;
        RECT 36.325 171.125 36.705 171.210 ;
        RECT 37.795 171.140 38.085 171.865 ;
        RECT 38.340 171.475 40.350 171.695 ;
        RECT 35.615 170.955 35.815 171.125 ;
        RECT 36.480 171.085 36.705 171.125 ;
        RECT 34.570 170.625 35.445 170.955 ;
        RECT 35.615 170.625 36.365 170.955 ;
        RECT 33.380 169.485 33.630 169.815 ;
        RECT 34.570 169.785 34.740 170.625 ;
        RECT 35.615 170.420 35.805 170.625 ;
        RECT 36.535 170.505 36.705 171.085 ;
        RECT 36.490 170.455 36.705 170.505 ;
        RECT 38.255 171.045 39.930 171.305 ;
        RECT 40.100 171.225 40.350 171.475 ;
        RECT 40.520 171.395 40.690 171.865 ;
        RECT 40.860 171.225 41.190 171.695 ;
        RECT 41.360 171.395 41.530 171.865 ;
        RECT 41.700 171.225 42.030 171.695 ;
        RECT 40.100 171.045 42.030 171.225 ;
        RECT 42.205 171.045 42.480 171.865 ;
        RECT 42.650 171.225 42.980 171.695 ;
        RECT 43.150 171.395 43.320 171.865 ;
        RECT 43.490 171.225 43.820 171.695 ;
        RECT 43.990 171.395 44.160 171.865 ;
        RECT 44.330 171.225 44.660 171.695 ;
        RECT 44.830 171.395 45.000 171.865 ;
        RECT 45.170 171.225 45.500 171.695 ;
        RECT 45.670 171.395 45.940 171.865 ;
        RECT 46.130 171.475 48.140 171.645 ;
        RECT 42.650 171.215 45.600 171.225 ;
        RECT 46.130 171.215 46.380 171.475 ;
        RECT 48.465 171.315 48.635 171.605 ;
        RECT 48.805 171.485 49.135 171.865 ;
        RECT 42.650 171.045 46.380 171.215 ;
        RECT 46.550 171.045 48.205 171.305 ;
        RECT 48.465 171.145 49.130 171.315 ;
        RECT 38.255 170.505 38.490 171.045 ;
        RECT 38.660 170.675 40.025 170.875 ;
        RECT 40.345 170.675 43.560 170.875 ;
        RECT 43.730 170.675 45.600 170.875 ;
        RECT 45.770 170.675 47.815 170.875 ;
        RECT 39.855 170.505 40.025 170.675 ;
        RECT 43.730 170.505 43.900 170.675 ;
        RECT 45.770 170.505 45.940 170.675 ;
        RECT 47.985 170.505 48.205 171.045 ;
        RECT 34.910 170.045 35.805 170.420 ;
        RECT 36.315 170.375 36.705 170.455 ;
        RECT 33.855 169.615 34.740 169.785 ;
        RECT 34.920 169.315 35.235 169.815 ;
        RECT 35.465 169.485 35.805 170.045 ;
        RECT 35.975 169.315 36.145 170.325 ;
        RECT 36.315 169.530 36.645 170.375 ;
        RECT 37.795 169.315 38.085 170.480 ;
        RECT 38.255 170.335 39.470 170.505 ;
        RECT 39.855 170.335 43.900 170.505 ;
        RECT 44.070 170.335 45.940 170.505 ;
        RECT 38.255 169.485 38.630 170.335 ;
        RECT 39.220 170.165 39.470 170.335 ;
        RECT 46.130 170.285 48.205 170.505 ;
        RECT 48.380 170.325 48.730 170.975 ;
        RECT 46.130 170.165 46.420 170.285 ;
        RECT 38.800 169.315 39.050 170.115 ;
        RECT 39.220 169.945 41.990 170.165 ;
        RECT 39.220 169.485 39.470 169.945 ;
        RECT 39.640 169.315 39.890 169.775 ;
        RECT 40.060 169.485 40.310 169.945 ;
        RECT 40.480 169.315 40.730 169.775 ;
        RECT 40.900 169.485 41.150 169.945 ;
        RECT 41.320 169.315 41.570 169.775 ;
        RECT 41.740 169.485 41.990 169.945 ;
        RECT 42.205 169.945 44.160 170.165 ;
        RECT 42.205 169.485 42.520 169.945 ;
        RECT 42.690 169.315 42.940 169.775 ;
        RECT 43.110 169.485 43.360 169.945 ;
        RECT 43.530 169.315 43.780 169.775 ;
        RECT 43.950 169.735 44.160 169.945 ;
        RECT 44.330 169.905 46.420 170.165 ;
        RECT 43.950 169.485 45.920 169.735 ;
        RECT 46.130 169.485 46.420 169.905 ;
        RECT 46.590 169.315 46.840 170.115 ;
        RECT 47.010 169.485 47.260 170.285 ;
        RECT 47.430 169.315 47.680 170.115 ;
        RECT 47.850 169.485 48.205 170.285 ;
        RECT 48.900 170.155 49.130 171.145 ;
        RECT 48.465 169.985 49.130 170.155 ;
        RECT 48.465 169.485 48.635 169.985 ;
        RECT 48.805 169.315 49.135 169.815 ;
        RECT 49.305 169.485 49.490 171.605 ;
        RECT 49.745 171.405 49.995 171.865 ;
        RECT 50.165 171.415 50.500 171.585 ;
        RECT 50.695 171.415 51.370 171.585 ;
        RECT 50.165 171.275 50.335 171.415 ;
        RECT 49.660 170.285 49.940 171.235 ;
        RECT 50.110 171.145 50.335 171.275 ;
        RECT 50.110 170.040 50.280 171.145 ;
        RECT 50.505 170.995 51.030 171.215 ;
        RECT 50.450 170.230 50.690 170.825 ;
        RECT 50.860 170.295 51.030 170.995 ;
        RECT 51.200 170.635 51.370 171.415 ;
        RECT 51.690 171.365 52.060 171.865 ;
        RECT 52.240 171.415 52.645 171.585 ;
        RECT 52.815 171.415 53.600 171.585 ;
        RECT 52.240 171.185 52.410 171.415 ;
        RECT 51.580 170.885 52.410 171.185 ;
        RECT 52.795 170.915 53.260 171.245 ;
        RECT 51.580 170.855 51.780 170.885 ;
        RECT 51.900 170.635 52.070 170.705 ;
        RECT 51.200 170.465 52.070 170.635 ;
        RECT 51.560 170.375 52.070 170.465 ;
        RECT 50.110 169.910 50.415 170.040 ;
        RECT 50.860 169.930 51.390 170.295 ;
        RECT 49.730 169.315 49.995 169.775 ;
        RECT 50.165 169.485 50.415 169.910 ;
        RECT 51.560 169.760 51.730 170.375 ;
        RECT 50.625 169.590 51.730 169.760 ;
        RECT 51.900 169.315 52.070 170.115 ;
        RECT 52.240 169.815 52.410 170.885 ;
        RECT 52.580 169.985 52.770 170.705 ;
        RECT 52.940 169.955 53.260 170.915 ;
        RECT 53.430 170.955 53.600 171.415 ;
        RECT 53.875 171.335 54.085 171.865 ;
        RECT 54.345 171.125 54.675 171.650 ;
        RECT 54.845 171.255 55.015 171.865 ;
        RECT 55.185 171.210 55.515 171.645 ;
        RECT 55.735 171.255 56.075 171.670 ;
        RECT 56.245 171.425 56.415 171.865 ;
        RECT 56.605 171.475 57.865 171.655 ;
        RECT 56.605 171.255 56.935 171.475 ;
        RECT 55.185 171.125 55.565 171.210 ;
        RECT 54.475 170.955 54.675 171.125 ;
        RECT 55.340 171.085 55.565 171.125 ;
        RECT 55.735 171.125 56.935 171.255 ;
        RECT 57.105 171.125 57.455 171.305 ;
        RECT 55.735 171.085 56.765 171.125 ;
        RECT 53.430 170.625 54.305 170.955 ;
        RECT 54.475 170.625 55.225 170.955 ;
        RECT 52.240 169.485 52.490 169.815 ;
        RECT 53.430 169.785 53.600 170.625 ;
        RECT 54.475 170.420 54.665 170.625 ;
        RECT 55.395 170.505 55.565 171.085 ;
        RECT 55.735 170.675 56.195 170.875 ;
        RECT 56.365 170.705 56.730 170.875 ;
        RECT 56.365 170.505 56.545 170.705 ;
        RECT 56.945 170.535 57.115 170.955 ;
        RECT 55.350 170.455 55.565 170.505 ;
        RECT 53.770 170.045 54.665 170.420 ;
        RECT 55.175 170.375 55.565 170.455 ;
        RECT 52.715 169.615 53.600 169.785 ;
        RECT 53.780 169.315 54.095 169.815 ;
        RECT 54.325 169.485 54.665 170.045 ;
        RECT 54.835 169.315 55.005 170.325 ;
        RECT 55.175 169.530 55.505 170.375 ;
        RECT 55.735 169.315 56.055 170.495 ;
        RECT 56.225 170.335 56.545 170.505 ;
        RECT 56.225 169.545 56.425 170.335 ;
        RECT 56.715 170.285 57.115 170.535 ;
        RECT 57.285 170.115 57.455 171.125 ;
        RECT 56.615 169.905 57.455 170.115 ;
        RECT 57.625 169.960 57.865 171.285 ;
        RECT 58.960 171.025 59.220 171.865 ;
        RECT 59.395 171.120 59.650 171.695 ;
        RECT 59.820 171.485 60.150 171.865 ;
        RECT 60.365 171.315 60.535 171.695 ;
        RECT 59.820 171.145 60.535 171.315 ;
        RECT 56.615 169.485 57.115 169.905 ;
        RECT 57.605 169.315 57.815 169.775 ;
        RECT 58.960 169.315 59.220 170.465 ;
        RECT 59.395 170.390 59.565 171.120 ;
        RECT 59.820 170.955 59.990 171.145 ;
        RECT 60.795 171.095 63.385 171.865 ;
        RECT 63.555 171.140 63.845 171.865 ;
        RECT 64.015 171.125 64.355 171.695 ;
        RECT 64.550 171.200 64.720 171.865 ;
        RECT 65.000 171.525 65.220 171.570 ;
        RECT 64.995 171.355 65.220 171.525 ;
        RECT 65.390 171.385 65.835 171.555 ;
        RECT 65.000 171.215 65.220 171.355 ;
        RECT 59.735 170.625 59.990 170.955 ;
        RECT 59.820 170.415 59.990 170.625 ;
        RECT 60.270 170.595 60.625 170.965 ;
        RECT 60.795 170.575 62.005 171.095 ;
        RECT 59.395 169.485 59.650 170.390 ;
        RECT 59.820 170.245 60.535 170.415 ;
        RECT 62.175 170.405 63.385 170.925 ;
        RECT 59.820 169.315 60.150 170.075 ;
        RECT 60.365 169.485 60.535 170.245 ;
        RECT 60.795 169.315 63.385 170.405 ;
        RECT 63.555 169.315 63.845 170.480 ;
        RECT 64.015 170.155 64.190 171.125 ;
        RECT 65.000 171.045 65.495 171.215 ;
        RECT 64.360 170.505 64.530 170.955 ;
        RECT 64.700 170.675 65.150 170.875 ;
        RECT 65.320 170.850 65.495 171.045 ;
        RECT 65.665 170.595 65.835 171.385 ;
        RECT 66.005 171.260 66.255 171.630 ;
        RECT 66.085 170.875 66.255 171.260 ;
        RECT 66.425 171.225 66.675 171.630 ;
        RECT 66.845 171.395 67.015 171.865 ;
        RECT 67.185 171.225 67.525 171.630 ;
        RECT 66.425 171.045 67.525 171.225 ;
        RECT 67.695 171.095 69.365 171.865 ;
        RECT 69.585 171.210 69.915 171.645 ;
        RECT 70.085 171.255 70.255 171.865 ;
        RECT 69.535 171.125 69.915 171.210 ;
        RECT 70.425 171.125 70.755 171.650 ;
        RECT 71.015 171.335 71.225 171.865 ;
        RECT 71.500 171.415 72.285 171.585 ;
        RECT 72.455 171.415 72.860 171.585 ;
        RECT 66.085 170.705 66.280 170.875 ;
        RECT 64.360 170.335 64.755 170.505 ;
        RECT 65.665 170.455 65.940 170.595 ;
        RECT 64.015 169.485 64.275 170.155 ;
        RECT 64.585 170.065 64.755 170.335 ;
        RECT 64.925 170.235 65.940 170.455 ;
        RECT 66.110 170.455 66.280 170.705 ;
        RECT 66.450 170.625 67.010 170.875 ;
        RECT 66.110 170.065 66.665 170.455 ;
        RECT 64.585 169.895 66.665 170.065 ;
        RECT 64.445 169.315 64.775 169.715 ;
        RECT 65.645 169.315 66.045 169.715 ;
        RECT 66.335 169.660 66.665 169.895 ;
        RECT 66.835 169.525 67.010 170.625 ;
        RECT 67.180 170.305 67.525 170.875 ;
        RECT 67.695 170.575 68.445 171.095 ;
        RECT 69.535 171.085 69.760 171.125 ;
        RECT 68.615 170.405 69.365 170.925 ;
        RECT 67.180 169.315 67.525 170.135 ;
        RECT 67.695 169.315 69.365 170.405 ;
        RECT 69.535 170.505 69.705 171.085 ;
        RECT 70.425 170.955 70.625 171.125 ;
        RECT 71.500 170.955 71.670 171.415 ;
        RECT 69.875 170.625 70.625 170.955 ;
        RECT 70.795 170.625 71.670 170.955 ;
        RECT 69.535 170.455 69.750 170.505 ;
        RECT 69.535 170.375 69.925 170.455 ;
        RECT 69.595 169.530 69.925 170.375 ;
        RECT 70.435 170.420 70.625 170.625 ;
        RECT 70.095 169.315 70.265 170.325 ;
        RECT 70.435 170.045 71.330 170.420 ;
        RECT 70.435 169.485 70.775 170.045 ;
        RECT 71.005 169.315 71.320 169.815 ;
        RECT 71.500 169.785 71.670 170.625 ;
        RECT 71.840 170.915 72.305 171.245 ;
        RECT 72.690 171.185 72.860 171.415 ;
        RECT 73.040 171.365 73.410 171.865 ;
        RECT 73.730 171.415 74.405 171.585 ;
        RECT 74.600 171.415 74.935 171.585 ;
        RECT 71.840 169.955 72.160 170.915 ;
        RECT 72.690 170.885 73.520 171.185 ;
        RECT 72.330 169.985 72.520 170.705 ;
        RECT 72.690 169.815 72.860 170.885 ;
        RECT 73.320 170.855 73.520 170.885 ;
        RECT 73.030 170.635 73.200 170.705 ;
        RECT 73.730 170.635 73.900 171.415 ;
        RECT 74.765 171.275 74.935 171.415 ;
        RECT 75.105 171.405 75.355 171.865 ;
        RECT 73.030 170.465 73.900 170.635 ;
        RECT 74.070 170.995 74.595 171.215 ;
        RECT 74.765 171.145 74.990 171.275 ;
        RECT 73.030 170.375 73.540 170.465 ;
        RECT 71.500 169.615 72.385 169.785 ;
        RECT 72.610 169.485 72.860 169.815 ;
        RECT 73.030 169.315 73.200 170.115 ;
        RECT 73.370 169.760 73.540 170.375 ;
        RECT 74.070 170.295 74.240 170.995 ;
        RECT 73.710 169.930 74.240 170.295 ;
        RECT 74.410 170.230 74.650 170.825 ;
        RECT 74.820 170.040 74.990 171.145 ;
        RECT 75.160 170.285 75.440 171.235 ;
        RECT 74.685 169.910 74.990 170.040 ;
        RECT 73.370 169.590 74.475 169.760 ;
        RECT 74.685 169.485 74.935 169.910 ;
        RECT 75.105 169.315 75.370 169.775 ;
        RECT 75.610 169.485 75.795 171.605 ;
        RECT 75.965 171.485 76.295 171.865 ;
        RECT 76.465 171.315 76.635 171.605 ;
        RECT 76.895 171.320 82.240 171.865 ;
        RECT 82.415 171.320 87.760 171.865 ;
        RECT 75.970 171.145 76.635 171.315 ;
        RECT 75.970 170.155 76.200 171.145 ;
        RECT 76.370 170.325 76.720 170.975 ;
        RECT 78.480 170.490 78.820 171.320 ;
        RECT 75.970 169.985 76.635 170.155 ;
        RECT 75.965 169.315 76.295 169.815 ;
        RECT 76.465 169.485 76.635 169.985 ;
        RECT 80.300 169.750 80.650 171.000 ;
        RECT 84.000 170.490 84.340 171.320 ;
        RECT 87.935 171.115 89.145 171.865 ;
        RECT 89.315 171.115 90.525 171.865 ;
        RECT 85.820 169.750 86.170 171.000 ;
        RECT 87.935 170.575 88.455 171.115 ;
        RECT 88.625 170.405 89.145 170.945 ;
        RECT 76.895 169.315 82.240 169.750 ;
        RECT 82.415 169.315 87.760 169.750 ;
        RECT 87.935 169.315 89.145 170.405 ;
        RECT 89.315 170.405 89.835 170.945 ;
        RECT 90.005 170.575 90.525 171.115 ;
        RECT 100.140 170.940 100.810 174.200 ;
        RECT 101.480 173.630 105.520 173.800 ;
        RECT 101.140 171.570 101.310 173.570 ;
        RECT 105.690 171.570 105.860 173.570 ;
        RECT 101.480 171.340 105.520 171.510 ;
        RECT 106.200 170.940 106.370 174.200 ;
        RECT 100.140 170.770 106.370 170.940 ;
        RECT 89.315 169.315 90.525 170.405 ;
        RECT 11.950 169.145 90.610 169.315 ;
        RECT 12.035 168.055 13.245 169.145 ;
        RECT 13.415 168.710 18.760 169.145 ;
        RECT 12.035 167.345 12.555 167.885 ;
        RECT 12.725 167.515 13.245 168.055 ;
        RECT 12.035 166.595 13.245 167.345 ;
        RECT 15.000 167.140 15.340 167.970 ;
        RECT 16.820 167.460 17.170 168.710 ;
        RECT 18.935 168.055 20.605 169.145 ;
        RECT 18.935 167.365 19.685 167.885 ;
        RECT 19.855 167.535 20.605 168.055 ;
        RECT 21.235 168.275 21.510 168.975 ;
        RECT 21.720 168.600 21.935 169.145 ;
        RECT 22.105 168.635 22.580 168.975 ;
        RECT 22.750 168.640 23.365 169.145 ;
        RECT 22.750 168.465 22.945 168.640 ;
        RECT 13.415 166.595 18.760 167.140 ;
        RECT 18.935 166.595 20.605 167.365 ;
        RECT 21.235 167.245 21.405 168.275 ;
        RECT 21.680 168.105 22.395 168.400 ;
        RECT 22.615 168.275 22.945 168.465 ;
        RECT 23.115 168.105 23.365 168.470 ;
        RECT 21.575 167.935 23.365 168.105 ;
        RECT 21.575 167.505 21.805 167.935 ;
        RECT 21.235 166.765 21.495 167.245 ;
        RECT 21.975 167.235 22.385 167.755 ;
        RECT 21.665 166.595 21.995 167.055 ;
        RECT 22.185 166.815 22.385 167.235 ;
        RECT 22.555 167.080 22.810 167.935 ;
        RECT 23.605 167.755 23.775 168.975 ;
        RECT 24.025 168.635 24.285 169.145 ;
        RECT 22.980 167.505 23.775 167.755 ;
        RECT 23.945 167.585 24.285 168.465 ;
        RECT 24.915 167.980 25.205 169.145 ;
        RECT 23.525 167.415 23.775 167.505 ;
        RECT 22.555 166.815 23.345 167.080 ;
        RECT 23.525 166.995 23.855 167.415 ;
        RECT 24.025 166.595 24.285 167.415 ;
        RECT 24.915 166.595 25.205 167.320 ;
        RECT 25.385 166.775 25.645 168.965 ;
        RECT 25.815 168.415 26.155 169.145 ;
        RECT 26.335 168.235 26.605 168.965 ;
        RECT 25.835 168.015 26.605 168.235 ;
        RECT 26.785 168.255 27.015 168.965 ;
        RECT 27.185 168.435 27.515 169.145 ;
        RECT 27.685 168.255 27.945 168.965 ;
        RECT 28.305 168.345 28.560 169.145 ;
        RECT 26.785 168.015 27.945 168.255 ;
        RECT 28.730 168.175 29.060 168.975 ;
        RECT 29.230 168.345 29.400 169.145 ;
        RECT 29.570 168.175 29.900 168.975 ;
        RECT 30.070 168.345 30.240 169.145 ;
        RECT 30.410 168.175 30.740 168.975 ;
        RECT 30.910 168.345 31.080 169.145 ;
        RECT 31.250 168.175 31.580 168.975 ;
        RECT 31.750 168.345 32.050 169.145 ;
        RECT 25.835 167.345 26.125 168.015 ;
        RECT 28.135 168.005 32.105 168.175 ;
        RECT 32.275 168.055 33.945 169.145 ;
        RECT 26.305 167.525 26.770 167.835 ;
        RECT 26.950 167.525 27.475 167.835 ;
        RECT 25.835 167.145 27.065 167.345 ;
        RECT 25.905 166.595 26.575 166.965 ;
        RECT 26.755 166.775 27.065 167.145 ;
        RECT 27.245 166.885 27.475 167.525 ;
        RECT 27.655 167.505 27.955 167.835 ;
        RECT 28.135 167.415 28.480 168.005 ;
        RECT 28.730 167.585 31.585 167.835 ;
        RECT 31.785 167.415 32.105 168.005 ;
        RECT 27.655 166.595 27.945 167.325 ;
        RECT 28.135 167.225 32.105 167.415 ;
        RECT 32.275 167.365 33.025 167.885 ;
        RECT 33.195 167.535 33.945 168.055 ;
        RECT 34.300 168.175 34.690 168.350 ;
        RECT 35.175 168.345 35.505 169.145 ;
        RECT 35.675 168.355 36.210 168.975 ;
        RECT 34.300 168.005 35.725 168.175 ;
        RECT 28.305 166.595 28.560 167.055 ;
        RECT 28.730 166.765 29.060 167.225 ;
        RECT 29.230 166.595 29.400 167.055 ;
        RECT 29.570 166.765 29.900 167.225 ;
        RECT 30.070 166.595 30.240 167.055 ;
        RECT 30.410 166.765 30.740 167.225 ;
        RECT 30.910 166.595 31.080 167.055 ;
        RECT 31.250 166.765 31.580 167.225 ;
        RECT 31.750 166.595 32.055 167.055 ;
        RECT 32.275 166.595 33.945 167.365 ;
        RECT 34.175 167.275 34.530 167.835 ;
        RECT 34.700 167.105 34.870 168.005 ;
        RECT 35.040 167.275 35.305 167.835 ;
        RECT 35.555 167.505 35.725 168.005 ;
        RECT 35.895 167.335 36.210 168.355 ;
        RECT 36.460 168.005 36.755 169.145 ;
        RECT 37.015 168.175 37.345 168.975 ;
        RECT 37.515 168.345 37.685 169.145 ;
        RECT 37.855 168.175 38.185 168.975 ;
        RECT 38.355 168.345 38.525 169.145 ;
        RECT 38.695 168.195 39.025 168.975 ;
        RECT 39.195 168.685 39.365 169.145 ;
        RECT 39.725 168.475 39.895 168.975 ;
        RECT 40.065 168.645 40.395 169.145 ;
        RECT 39.725 168.305 40.390 168.475 ;
        RECT 38.695 168.175 39.465 168.195 ;
        RECT 37.015 168.005 39.465 168.175 ;
        RECT 36.435 167.585 38.945 167.835 ;
        RECT 39.115 167.415 39.465 168.005 ;
        RECT 39.640 167.485 39.990 168.135 ;
        RECT 34.280 166.595 34.520 167.105 ;
        RECT 34.700 166.775 34.980 167.105 ;
        RECT 35.210 166.595 35.425 167.105 ;
        RECT 35.595 166.765 36.210 167.335 ;
        RECT 37.095 167.235 39.465 167.415 ;
        RECT 40.160 167.315 40.390 168.305 ;
        RECT 36.460 166.595 36.725 167.055 ;
        RECT 37.095 166.765 37.265 167.235 ;
        RECT 37.515 166.595 37.685 167.055 ;
        RECT 37.935 166.765 38.105 167.235 ;
        RECT 38.355 166.595 38.525 167.055 ;
        RECT 38.775 166.765 38.945 167.235 ;
        RECT 39.725 167.145 40.390 167.315 ;
        RECT 39.115 166.595 39.365 167.060 ;
        RECT 39.725 166.855 39.895 167.145 ;
        RECT 40.065 166.595 40.395 166.975 ;
        RECT 40.565 166.855 40.750 168.975 ;
        RECT 40.990 168.685 41.255 169.145 ;
        RECT 41.425 168.550 41.675 168.975 ;
        RECT 41.885 168.700 42.990 168.870 ;
        RECT 41.370 168.420 41.675 168.550 ;
        RECT 40.920 167.225 41.200 168.175 ;
        RECT 41.370 167.315 41.540 168.420 ;
        RECT 41.710 167.635 41.950 168.230 ;
        RECT 42.120 168.165 42.650 168.530 ;
        RECT 42.120 167.465 42.290 168.165 ;
        RECT 42.820 168.085 42.990 168.700 ;
        RECT 43.160 168.345 43.330 169.145 ;
        RECT 43.500 168.645 43.750 168.975 ;
        RECT 43.975 168.675 44.860 168.845 ;
        RECT 42.820 167.995 43.330 168.085 ;
        RECT 41.370 167.185 41.595 167.315 ;
        RECT 41.765 167.245 42.290 167.465 ;
        RECT 42.460 167.825 43.330 167.995 ;
        RECT 41.005 166.595 41.255 167.055 ;
        RECT 41.425 167.045 41.595 167.185 ;
        RECT 42.460 167.045 42.630 167.825 ;
        RECT 43.160 167.755 43.330 167.825 ;
        RECT 42.840 167.575 43.040 167.605 ;
        RECT 43.500 167.575 43.670 168.645 ;
        RECT 43.840 167.755 44.030 168.475 ;
        RECT 42.840 167.275 43.670 167.575 ;
        RECT 44.200 167.545 44.520 168.505 ;
        RECT 41.425 166.875 41.760 167.045 ;
        RECT 41.955 166.875 42.630 167.045 ;
        RECT 42.950 166.595 43.320 167.095 ;
        RECT 43.500 167.045 43.670 167.275 ;
        RECT 44.055 167.215 44.520 167.545 ;
        RECT 44.690 167.835 44.860 168.675 ;
        RECT 45.040 168.645 45.355 169.145 ;
        RECT 45.585 168.415 45.925 168.975 ;
        RECT 45.030 168.040 45.925 168.415 ;
        RECT 46.095 168.135 46.265 169.145 ;
        RECT 45.735 167.835 45.925 168.040 ;
        RECT 46.435 168.085 46.765 168.930 ;
        RECT 47.200 168.175 47.530 168.975 ;
        RECT 47.700 168.345 48.030 169.145 ;
        RECT 48.330 168.175 48.660 168.975 ;
        RECT 49.305 168.345 49.555 169.145 ;
        RECT 46.435 168.005 46.825 168.085 ;
        RECT 47.200 168.005 49.635 168.175 ;
        RECT 49.825 168.005 49.995 169.145 ;
        RECT 50.165 168.005 50.505 168.975 ;
        RECT 46.610 167.955 46.825 168.005 ;
        RECT 44.690 167.505 45.565 167.835 ;
        RECT 45.735 167.505 46.485 167.835 ;
        RECT 44.690 167.045 44.860 167.505 ;
        RECT 45.735 167.335 45.935 167.505 ;
        RECT 46.655 167.375 46.825 167.955 ;
        RECT 46.995 167.585 47.345 167.835 ;
        RECT 47.530 167.375 47.700 168.005 ;
        RECT 47.870 167.585 48.200 167.785 ;
        RECT 48.370 167.585 48.700 167.785 ;
        RECT 48.870 167.585 49.290 167.785 ;
        RECT 49.465 167.755 49.635 168.005 ;
        RECT 49.465 167.585 50.160 167.755 ;
        RECT 46.600 167.335 46.825 167.375 ;
        RECT 43.500 166.875 43.905 167.045 ;
        RECT 44.075 166.875 44.860 167.045 ;
        RECT 45.135 166.595 45.345 167.125 ;
        RECT 45.605 166.810 45.935 167.335 ;
        RECT 46.445 167.250 46.825 167.335 ;
        RECT 46.105 166.595 46.275 167.205 ;
        RECT 46.445 166.815 46.775 167.250 ;
        RECT 47.200 166.765 47.700 167.375 ;
        RECT 48.330 167.245 49.555 167.415 ;
        RECT 50.330 167.395 50.505 168.005 ;
        RECT 50.675 167.980 50.965 169.145 ;
        RECT 51.135 168.005 51.415 169.145 ;
        RECT 51.585 167.995 51.915 168.975 ;
        RECT 52.085 168.005 52.345 169.145 ;
        RECT 52.555 168.005 52.785 169.145 ;
        RECT 52.955 167.995 53.285 168.975 ;
        RECT 53.455 168.005 53.665 169.145 ;
        RECT 53.985 168.525 54.155 168.955 ;
        RECT 54.325 168.695 54.655 169.145 ;
        RECT 53.985 168.295 54.660 168.525 ;
        RECT 51.145 167.565 51.480 167.835 ;
        RECT 51.650 167.395 51.820 167.995 ;
        RECT 51.990 167.585 52.325 167.835 ;
        RECT 52.535 167.585 52.865 167.835 ;
        RECT 48.330 166.765 48.660 167.245 ;
        RECT 48.830 166.595 49.055 167.055 ;
        RECT 49.225 166.765 49.555 167.245 ;
        RECT 49.745 166.595 49.995 167.395 ;
        RECT 50.165 166.765 50.505 167.395 ;
        RECT 50.675 166.595 50.965 167.320 ;
        RECT 51.135 166.595 51.445 167.395 ;
        RECT 51.650 166.765 52.345 167.395 ;
        RECT 52.555 166.595 52.785 167.415 ;
        RECT 53.035 167.395 53.285 167.995 ;
        RECT 52.955 166.765 53.285 167.395 ;
        RECT 53.455 166.595 53.665 167.415 ;
        RECT 53.955 167.275 54.255 168.125 ;
        RECT 54.425 167.645 54.660 168.295 ;
        RECT 54.830 167.985 55.115 168.930 ;
        RECT 55.295 168.675 55.980 169.145 ;
        RECT 55.290 168.155 55.985 168.465 ;
        RECT 56.160 168.090 56.465 168.875 ;
        RECT 54.830 167.835 55.690 167.985 ;
        RECT 56.255 167.955 56.465 168.090 ;
        RECT 56.665 168.035 56.960 169.145 ;
        RECT 54.830 167.815 56.115 167.835 ;
        RECT 54.425 167.315 54.960 167.645 ;
        RECT 55.130 167.455 56.115 167.815 ;
        RECT 54.425 167.165 54.645 167.315 ;
        RECT 53.900 166.595 54.235 167.100 ;
        RECT 54.405 166.790 54.645 167.165 ;
        RECT 55.130 167.120 55.300 167.455 ;
        RECT 56.290 167.285 56.465 167.955 ;
        RECT 57.140 167.835 57.390 168.970 ;
        RECT 57.560 168.035 57.820 169.145 ;
        RECT 57.990 168.245 58.250 168.970 ;
        RECT 58.420 168.415 58.680 169.145 ;
        RECT 58.850 168.245 59.110 168.970 ;
        RECT 59.280 168.415 59.540 169.145 ;
        RECT 59.710 168.245 59.970 168.970 ;
        RECT 60.140 168.415 60.400 169.145 ;
        RECT 60.570 168.245 60.830 168.970 ;
        RECT 61.000 168.415 61.295 169.145 ;
        RECT 61.715 168.295 62.095 168.975 ;
        RECT 62.685 168.295 62.855 169.145 ;
        RECT 63.025 168.465 63.355 168.975 ;
        RECT 63.525 168.635 63.695 169.145 ;
        RECT 63.865 168.465 64.265 168.975 ;
        RECT 63.025 168.295 64.265 168.465 ;
        RECT 57.990 168.005 61.300 168.245 ;
        RECT 54.925 166.925 55.300 167.120 ;
        RECT 54.925 166.780 55.095 166.925 ;
        RECT 55.660 166.595 56.055 167.090 ;
        RECT 56.225 166.765 56.465 167.285 ;
        RECT 56.655 167.225 56.970 167.835 ;
        RECT 57.140 167.585 60.160 167.835 ;
        RECT 56.715 166.595 56.960 167.055 ;
        RECT 57.140 166.775 57.390 167.585 ;
        RECT 60.330 167.415 61.300 168.005 ;
        RECT 57.990 167.245 61.300 167.415 ;
        RECT 61.715 167.335 61.885 168.295 ;
        RECT 62.055 167.955 63.360 168.125 ;
        RECT 64.445 168.045 64.765 168.975 ;
        RECT 64.935 168.055 66.605 169.145 ;
        RECT 62.055 167.505 62.300 167.955 ;
        RECT 62.470 167.585 63.020 167.785 ;
        RECT 63.190 167.755 63.360 167.955 ;
        RECT 64.135 167.875 64.765 168.045 ;
        RECT 63.190 167.585 63.565 167.755 ;
        RECT 63.735 167.335 63.965 167.835 ;
        RECT 57.560 166.595 57.820 167.120 ;
        RECT 57.990 166.790 58.250 167.245 ;
        RECT 58.420 166.595 58.680 167.075 ;
        RECT 58.850 166.790 59.110 167.245 ;
        RECT 59.280 166.595 59.540 167.075 ;
        RECT 59.710 166.790 59.970 167.245 ;
        RECT 60.140 166.595 60.400 167.075 ;
        RECT 60.570 166.790 60.830 167.245 ;
        RECT 61.715 167.165 63.965 167.335 ;
        RECT 61.000 166.595 61.300 167.075 ;
        RECT 61.765 166.595 62.095 166.985 ;
        RECT 62.265 166.845 62.435 167.165 ;
        RECT 64.135 166.995 64.305 167.875 ;
        RECT 62.605 166.595 62.935 166.985 ;
        RECT 63.350 166.825 64.305 166.995 ;
        RECT 64.475 166.595 64.765 167.430 ;
        RECT 64.935 167.365 65.685 167.885 ;
        RECT 65.855 167.535 66.605 168.055 ;
        RECT 67.280 168.005 67.575 169.145 ;
        RECT 67.835 168.175 68.165 168.975 ;
        RECT 68.335 168.345 68.505 169.145 ;
        RECT 68.675 168.175 69.005 168.975 ;
        RECT 69.175 168.345 69.345 169.145 ;
        RECT 69.515 168.195 69.845 168.975 ;
        RECT 70.015 168.685 70.185 169.145 ;
        RECT 70.455 168.275 70.730 168.975 ;
        RECT 70.900 168.600 71.155 169.145 ;
        RECT 71.325 168.635 71.805 168.975 ;
        RECT 71.980 168.590 72.585 169.145 ;
        RECT 71.970 168.490 72.585 168.590 ;
        RECT 71.970 168.465 72.155 168.490 ;
        RECT 69.515 168.175 70.285 168.195 ;
        RECT 67.835 168.005 70.285 168.175 ;
        RECT 67.255 167.585 69.765 167.835 ;
        RECT 69.935 167.415 70.285 168.005 ;
        RECT 64.935 166.595 66.605 167.365 ;
        RECT 67.915 167.235 70.285 167.415 ;
        RECT 70.455 167.245 70.625 168.275 ;
        RECT 70.900 168.145 71.655 168.395 ;
        RECT 71.825 168.220 72.155 168.465 ;
        RECT 70.900 168.110 71.670 168.145 ;
        RECT 70.900 168.100 71.685 168.110 ;
        RECT 70.795 168.085 71.690 168.100 ;
        RECT 70.795 168.070 71.710 168.085 ;
        RECT 70.795 168.060 71.730 168.070 ;
        RECT 70.795 168.050 71.755 168.060 ;
        RECT 70.795 168.020 71.825 168.050 ;
        RECT 70.795 167.990 71.845 168.020 ;
        RECT 70.795 167.960 71.865 167.990 ;
        RECT 70.795 167.935 71.895 167.960 ;
        RECT 70.795 167.900 71.930 167.935 ;
        RECT 70.795 167.895 71.960 167.900 ;
        RECT 70.795 167.500 71.025 167.895 ;
        RECT 71.570 167.890 71.960 167.895 ;
        RECT 71.595 167.880 71.960 167.890 ;
        RECT 71.610 167.875 71.960 167.880 ;
        RECT 71.625 167.870 71.960 167.875 ;
        RECT 72.325 167.870 72.585 168.320 ;
        RECT 72.755 168.055 76.265 169.145 ;
        RECT 71.625 167.865 72.585 167.870 ;
        RECT 71.635 167.855 72.585 167.865 ;
        RECT 71.645 167.850 72.585 167.855 ;
        RECT 71.655 167.840 72.585 167.850 ;
        RECT 71.660 167.830 72.585 167.840 ;
        RECT 71.665 167.825 72.585 167.830 ;
        RECT 71.675 167.810 72.585 167.825 ;
        RECT 71.680 167.795 72.585 167.810 ;
        RECT 71.690 167.770 72.585 167.795 ;
        RECT 71.195 167.300 71.525 167.725 ;
        RECT 71.275 167.275 71.525 167.300 ;
        RECT 67.280 166.595 67.545 167.055 ;
        RECT 67.915 166.765 68.085 167.235 ;
        RECT 68.335 166.595 68.505 167.055 ;
        RECT 68.755 166.765 68.925 167.235 ;
        RECT 69.175 166.595 69.345 167.055 ;
        RECT 69.595 166.765 69.765 167.235 ;
        RECT 69.935 166.595 70.185 167.060 ;
        RECT 70.455 166.765 70.715 167.245 ;
        RECT 70.885 166.595 71.135 167.135 ;
        RECT 71.305 166.815 71.525 167.275 ;
        RECT 71.695 167.700 72.585 167.770 ;
        RECT 71.695 166.975 71.865 167.700 ;
        RECT 72.035 167.145 72.585 167.530 ;
        RECT 72.755 167.365 74.405 167.885 ;
        RECT 74.575 167.535 76.265 168.055 ;
        RECT 76.435 167.980 76.725 169.145 ;
        RECT 76.895 168.710 82.240 169.145 ;
        RECT 82.415 168.710 87.760 169.145 ;
        RECT 71.695 166.805 72.585 166.975 ;
        RECT 72.755 166.595 76.265 167.365 ;
        RECT 76.435 166.595 76.725 167.320 ;
        RECT 78.480 167.140 78.820 167.970 ;
        RECT 80.300 167.460 80.650 168.710 ;
        RECT 84.000 167.140 84.340 167.970 ;
        RECT 85.820 167.460 86.170 168.710 ;
        RECT 87.935 168.055 89.145 169.145 ;
        RECT 87.935 167.345 88.455 167.885 ;
        RECT 88.625 167.515 89.145 168.055 ;
        RECT 89.315 168.055 90.525 169.145 ;
        RECT 89.315 167.515 89.835 168.055 ;
        RECT 90.005 167.345 90.525 167.885 ;
        RECT 100.140 167.510 100.810 170.770 ;
        RECT 101.480 170.200 105.520 170.370 ;
        RECT 101.140 168.140 101.310 170.140 ;
        RECT 105.690 168.140 105.860 170.140 ;
        RECT 101.480 167.910 105.520 168.080 ;
        RECT 106.200 167.510 106.370 170.770 ;
        RECT 100.140 167.500 106.370 167.510 ;
        RECT 107.960 176.770 117.790 176.810 ;
        RECT 140.540 176.790 146.280 176.800 ;
        RECT 107.960 176.640 118.590 176.770 ;
        RECT 120.510 176.740 126.250 176.750 ;
        RECT 107.960 174.380 108.130 176.640 ;
        RECT 108.855 176.070 116.895 176.240 ;
        RECT 108.470 175.010 108.640 176.010 ;
        RECT 117.110 175.010 117.280 176.010 ;
        RECT 108.855 174.780 116.895 174.950 ;
        RECT 117.620 174.380 118.590 176.640 ;
        RECT 107.960 174.210 118.590 174.380 ;
        RECT 107.960 170.950 108.130 174.210 ;
        RECT 108.855 173.640 116.895 173.810 ;
        RECT 108.470 171.580 108.640 173.580 ;
        RECT 117.110 171.580 117.280 173.580 ;
        RECT 108.855 171.350 116.895 171.520 ;
        RECT 117.620 170.950 118.590 174.210 ;
        RECT 107.960 170.780 118.590 170.950 ;
        RECT 107.960 167.520 108.130 170.780 ;
        RECT 108.855 170.210 116.895 170.380 ;
        RECT 108.470 168.150 108.640 170.150 ;
        RECT 117.110 168.150 117.280 170.150 ;
        RECT 108.855 167.920 116.895 168.090 ;
        RECT 117.620 167.520 118.590 170.780 ;
        RECT 100.140 167.400 106.380 167.500 ;
        RECT 76.895 166.595 82.240 167.140 ;
        RECT 82.415 166.595 87.760 167.140 ;
        RECT 87.935 166.595 89.145 167.345 ;
        RECT 89.315 166.595 90.525 167.345 ;
        RECT 100.130 166.840 106.380 167.400 ;
        RECT 100.130 166.820 105.300 166.840 ;
        RECT 100.130 166.750 104.120 166.820 ;
        RECT 11.950 166.425 90.610 166.595 ;
        RECT 12.035 165.675 13.245 166.425 ;
        RECT 13.415 165.880 18.760 166.425 ;
        RECT 12.035 165.135 12.555 165.675 ;
        RECT 12.725 164.965 13.245 165.505 ;
        RECT 15.000 165.050 15.340 165.880 ;
        RECT 18.935 165.655 22.445 166.425 ;
        RECT 22.780 165.915 23.020 166.425 ;
        RECT 23.200 165.915 23.480 166.245 ;
        RECT 23.710 165.915 23.925 166.425 ;
        RECT 12.035 163.875 13.245 164.965 ;
        RECT 16.820 164.310 17.170 165.560 ;
        RECT 18.935 165.135 20.585 165.655 ;
        RECT 20.755 164.965 22.445 165.485 ;
        RECT 22.675 165.185 23.030 165.745 ;
        RECT 23.200 165.015 23.370 165.915 ;
        RECT 23.540 165.185 23.805 165.745 ;
        RECT 24.095 165.685 24.710 166.255 ;
        RECT 24.055 165.015 24.225 165.515 ;
        RECT 13.415 163.875 18.760 164.310 ;
        RECT 18.935 163.875 22.445 164.965 ;
        RECT 22.800 164.845 24.225 165.015 ;
        RECT 22.800 164.670 23.190 164.845 ;
        RECT 23.675 163.875 24.005 164.675 ;
        RECT 24.395 164.665 24.710 165.685 ;
        RECT 24.175 164.045 24.710 164.665 ;
        RECT 24.915 165.705 25.255 166.215 ;
        RECT 24.915 164.305 25.175 165.705 ;
        RECT 25.425 165.625 25.695 166.425 ;
        RECT 25.350 165.185 25.680 165.435 ;
        RECT 25.875 165.185 26.155 166.155 ;
        RECT 26.335 165.185 26.635 166.155 ;
        RECT 26.815 165.185 27.165 166.150 ;
        RECT 27.385 165.925 27.880 166.255 ;
        RECT 28.380 165.945 28.680 166.425 ;
        RECT 25.365 165.015 25.680 165.185 ;
        RECT 27.385 165.015 27.555 165.925 ;
        RECT 28.850 165.775 29.110 166.230 ;
        RECT 29.280 165.945 29.540 166.425 ;
        RECT 29.710 165.775 29.970 166.230 ;
        RECT 30.140 165.945 30.400 166.425 ;
        RECT 30.570 165.775 30.830 166.230 ;
        RECT 31.000 165.945 31.260 166.425 ;
        RECT 31.430 165.775 31.690 166.230 ;
        RECT 31.860 165.900 32.120 166.425 ;
        RECT 25.365 164.845 27.555 165.015 ;
        RECT 24.915 164.045 25.255 164.305 ;
        RECT 25.425 163.875 25.755 164.675 ;
        RECT 26.220 164.045 26.470 164.845 ;
        RECT 26.655 163.875 26.985 164.595 ;
        RECT 27.205 164.045 27.455 164.845 ;
        RECT 27.725 164.435 27.965 165.745 ;
        RECT 28.380 165.605 31.690 165.775 ;
        RECT 28.380 165.015 29.350 165.605 ;
        RECT 32.290 165.435 32.540 166.245 ;
        RECT 32.720 165.965 32.965 166.425 ;
        RECT 29.520 165.185 32.540 165.435 ;
        RECT 32.710 165.185 33.025 165.795 ;
        RECT 28.380 164.775 31.690 165.015 ;
        RECT 27.625 163.875 27.960 164.255 ;
        RECT 28.385 163.875 28.680 164.605 ;
        RECT 28.850 164.050 29.110 164.775 ;
        RECT 29.280 163.875 29.540 164.605 ;
        RECT 29.710 164.050 29.970 164.775 ;
        RECT 30.140 163.875 30.400 164.605 ;
        RECT 30.570 164.050 30.830 164.775 ;
        RECT 31.000 163.875 31.260 164.605 ;
        RECT 31.430 164.050 31.690 164.775 ;
        RECT 31.860 163.875 32.120 164.985 ;
        RECT 32.290 164.050 32.540 165.185 ;
        RECT 32.720 163.875 33.015 164.985 ;
        RECT 33.205 164.055 33.465 166.245 ;
        RECT 33.725 166.055 34.395 166.425 ;
        RECT 34.575 165.875 34.885 166.245 ;
        RECT 33.655 165.675 34.885 165.875 ;
        RECT 33.655 165.005 33.945 165.675 ;
        RECT 35.065 165.495 35.295 166.135 ;
        RECT 35.475 165.695 35.765 166.425 ;
        RECT 35.955 165.655 37.625 166.425 ;
        RECT 37.795 165.700 38.085 166.425 ;
        RECT 38.255 165.880 43.600 166.425 ;
        RECT 43.775 165.880 49.120 166.425 ;
        RECT 49.295 165.880 54.640 166.425 ;
        RECT 34.125 165.185 34.590 165.495 ;
        RECT 34.770 165.185 35.295 165.495 ;
        RECT 35.475 165.185 35.775 165.515 ;
        RECT 35.955 165.135 36.705 165.655 ;
        RECT 33.655 164.785 34.425 165.005 ;
        RECT 33.635 163.875 33.975 164.605 ;
        RECT 34.155 164.055 34.425 164.785 ;
        RECT 34.605 164.765 35.765 165.005 ;
        RECT 36.875 164.965 37.625 165.485 ;
        RECT 39.840 165.050 40.180 165.880 ;
        RECT 34.605 164.055 34.835 164.765 ;
        RECT 35.005 163.875 35.335 164.585 ;
        RECT 35.505 164.055 35.765 164.765 ;
        RECT 35.955 163.875 37.625 164.965 ;
        RECT 37.795 163.875 38.085 165.040 ;
        RECT 41.660 164.310 42.010 165.560 ;
        RECT 45.360 165.050 45.700 165.880 ;
        RECT 47.180 164.310 47.530 165.560 ;
        RECT 50.880 165.050 51.220 165.880 ;
        RECT 54.815 165.655 56.485 166.425 ;
        RECT 56.825 165.965 57.080 166.425 ;
        RECT 57.250 165.795 57.580 166.255 ;
        RECT 57.750 165.965 57.920 166.425 ;
        RECT 58.090 165.795 58.420 166.255 ;
        RECT 58.590 165.965 58.760 166.425 ;
        RECT 58.930 165.795 59.260 166.255 ;
        RECT 59.430 165.965 59.600 166.425 ;
        RECT 59.770 165.795 60.100 166.255 ;
        RECT 60.270 165.965 60.575 166.425 ;
        RECT 52.700 164.310 53.050 165.560 ;
        RECT 54.815 165.135 55.565 165.655 ;
        RECT 56.655 165.605 60.625 165.795 ;
        RECT 61.260 165.775 61.530 165.985 ;
        RECT 61.750 165.965 62.080 166.425 ;
        RECT 62.590 165.965 63.340 166.255 ;
        RECT 61.260 165.605 62.595 165.775 ;
        RECT 55.735 164.965 56.485 165.485 ;
        RECT 38.255 163.875 43.600 164.310 ;
        RECT 43.775 163.875 49.120 164.310 ;
        RECT 49.295 163.875 54.640 164.310 ;
        RECT 54.815 163.875 56.485 164.965 ;
        RECT 56.655 165.015 57.000 165.605 ;
        RECT 57.250 165.405 60.105 165.435 ;
        RECT 57.175 165.235 60.105 165.405 ;
        RECT 57.250 165.185 60.105 165.235 ;
        RECT 60.305 165.015 60.625 165.605 ;
        RECT 62.425 165.435 62.595 165.605 ;
        RECT 61.260 165.195 61.610 165.435 ;
        RECT 61.780 165.195 62.255 165.435 ;
        RECT 62.425 165.185 62.800 165.435 ;
        RECT 62.425 165.015 62.595 165.185 ;
        RECT 56.655 164.845 60.625 165.015 ;
        RECT 61.260 164.845 62.595 165.015 ;
        RECT 56.825 163.875 57.080 164.675 ;
        RECT 57.250 164.045 57.580 164.845 ;
        RECT 57.750 163.875 57.920 164.675 ;
        RECT 58.090 164.045 58.420 164.845 ;
        RECT 58.590 163.875 58.760 164.675 ;
        RECT 58.930 164.045 59.260 164.845 ;
        RECT 59.430 163.875 59.600 164.675 ;
        RECT 59.770 164.045 60.100 164.845 ;
        RECT 61.260 164.685 61.540 164.845 ;
        RECT 62.970 164.675 63.340 165.965 ;
        RECT 63.555 165.700 63.845 166.425 ;
        RECT 64.015 165.925 64.315 166.255 ;
        RECT 64.485 165.945 64.760 166.425 ;
        RECT 60.270 163.875 60.570 164.675 ;
        RECT 61.750 163.875 62.000 164.675 ;
        RECT 62.170 164.505 63.340 164.675 ;
        RECT 62.170 164.045 62.500 164.505 ;
        RECT 62.670 163.875 62.885 164.335 ;
        RECT 63.555 163.875 63.845 165.040 ;
        RECT 64.015 165.015 64.185 165.925 ;
        RECT 64.940 165.775 65.235 166.165 ;
        RECT 65.405 165.945 65.660 166.425 ;
        RECT 65.835 165.775 66.095 166.165 ;
        RECT 66.265 165.945 66.545 166.425 ;
        RECT 67.295 165.965 67.540 166.425 ;
        RECT 64.355 165.185 64.705 165.755 ;
        RECT 64.940 165.605 66.590 165.775 ;
        RECT 64.875 165.265 66.015 165.435 ;
        RECT 64.875 165.015 65.045 165.265 ;
        RECT 66.185 165.095 66.590 165.605 ;
        RECT 67.235 165.185 67.550 165.795 ;
        RECT 67.720 165.435 67.970 166.245 ;
        RECT 68.140 165.900 68.400 166.425 ;
        RECT 68.570 165.775 68.830 166.230 ;
        RECT 69.000 165.945 69.260 166.425 ;
        RECT 69.430 165.775 69.690 166.230 ;
        RECT 69.860 165.945 70.120 166.425 ;
        RECT 70.290 165.775 70.550 166.230 ;
        RECT 70.720 165.945 70.980 166.425 ;
        RECT 71.150 165.775 71.410 166.230 ;
        RECT 71.580 165.945 71.880 166.425 ;
        RECT 72.295 165.880 77.640 166.425 ;
        RECT 77.815 165.880 83.160 166.425 ;
        RECT 83.335 165.880 88.680 166.425 ;
        RECT 68.570 165.605 71.880 165.775 ;
        RECT 67.720 165.185 70.740 165.435 ;
        RECT 64.015 164.845 65.045 165.015 ;
        RECT 65.835 164.925 66.590 165.095 ;
        RECT 64.015 164.045 64.325 164.845 ;
        RECT 65.835 164.675 66.095 164.925 ;
        RECT 64.495 163.875 64.805 164.675 ;
        RECT 64.975 164.505 66.095 164.675 ;
        RECT 64.975 164.045 65.235 164.505 ;
        RECT 65.405 163.875 65.660 164.335 ;
        RECT 65.835 164.045 66.095 164.505 ;
        RECT 66.265 163.875 66.550 164.745 ;
        RECT 67.245 163.875 67.540 164.985 ;
        RECT 67.720 164.050 67.970 165.185 ;
        RECT 70.910 165.015 71.880 165.605 ;
        RECT 73.880 165.050 74.220 165.880 ;
        RECT 68.140 163.875 68.400 164.985 ;
        RECT 68.570 164.775 71.880 165.015 ;
        RECT 68.570 164.050 68.830 164.775 ;
        RECT 69.000 163.875 69.260 164.605 ;
        RECT 69.430 164.050 69.690 164.775 ;
        RECT 69.860 163.875 70.120 164.605 ;
        RECT 70.290 164.050 70.550 164.775 ;
        RECT 70.720 163.875 70.980 164.605 ;
        RECT 71.150 164.050 71.410 164.775 ;
        RECT 71.580 163.875 71.875 164.605 ;
        RECT 75.700 164.310 76.050 165.560 ;
        RECT 79.400 165.050 79.740 165.880 ;
        RECT 81.220 164.310 81.570 165.560 ;
        RECT 84.920 165.050 85.260 165.880 ;
        RECT 89.315 165.675 90.525 166.425 ;
        RECT 86.740 164.310 87.090 165.560 ;
        RECT 89.315 164.965 89.835 165.505 ;
        RECT 90.005 165.135 90.525 165.675 ;
        RECT 100.130 165.480 102.050 166.750 ;
        RECT 103.560 166.740 104.120 166.750 ;
        RECT 103.790 165.650 104.120 166.740 ;
        RECT 104.490 166.270 105.530 166.440 ;
        RECT 104.490 165.830 105.530 166.000 ;
        RECT 105.700 165.970 105.870 166.300 ;
        RECT 103.950 165.430 104.120 165.650 ;
        RECT 106.210 165.430 106.380 166.840 ;
        RECT 103.950 165.260 106.380 165.430 ;
        RECT 107.960 167.350 118.590 167.520 ;
        RECT 120.020 176.580 126.250 176.740 ;
        RECT 120.020 174.320 120.690 176.580 ;
        RECT 121.360 176.010 125.400 176.180 ;
        RECT 121.020 174.950 121.190 175.950 ;
        RECT 125.570 174.950 125.740 175.950 ;
        RECT 121.360 174.720 125.400 174.890 ;
        RECT 126.080 174.320 126.250 176.580 ;
        RECT 120.020 174.150 126.250 174.320 ;
        RECT 120.020 170.890 120.690 174.150 ;
        RECT 121.360 173.580 125.400 173.750 ;
        RECT 121.020 171.520 121.190 173.520 ;
        RECT 125.570 171.520 125.740 173.520 ;
        RECT 121.360 171.290 125.400 171.460 ;
        RECT 126.080 170.890 126.250 174.150 ;
        RECT 120.020 170.720 126.250 170.890 ;
        RECT 120.020 167.460 120.690 170.720 ;
        RECT 121.360 170.150 125.400 170.320 ;
        RECT 121.020 168.090 121.190 170.090 ;
        RECT 125.570 168.090 125.740 170.090 ;
        RECT 121.360 167.860 125.400 168.030 ;
        RECT 126.080 167.460 126.250 170.720 ;
        RECT 120.020 167.450 126.250 167.460 ;
        RECT 127.840 176.720 137.670 176.760 ;
        RECT 127.840 176.590 138.470 176.720 ;
        RECT 127.840 174.330 128.010 176.590 ;
        RECT 128.735 176.020 136.775 176.190 ;
        RECT 128.350 174.960 128.520 175.960 ;
        RECT 136.990 174.960 137.160 175.960 ;
        RECT 128.735 174.730 136.775 174.900 ;
        RECT 137.500 174.330 138.470 176.590 ;
        RECT 127.840 174.160 138.470 174.330 ;
        RECT 127.840 170.900 128.010 174.160 ;
        RECT 128.735 173.590 136.775 173.760 ;
        RECT 128.350 171.530 128.520 173.530 ;
        RECT 136.990 171.530 137.160 173.530 ;
        RECT 128.735 171.300 136.775 171.470 ;
        RECT 137.500 170.900 138.470 174.160 ;
        RECT 127.840 170.730 138.470 170.900 ;
        RECT 127.840 167.470 128.010 170.730 ;
        RECT 128.735 170.160 136.775 170.330 ;
        RECT 128.350 168.100 128.520 170.100 ;
        RECT 136.990 168.100 137.160 170.100 ;
        RECT 128.735 167.870 136.775 168.040 ;
        RECT 137.500 167.470 138.470 170.730 ;
        RECT 120.020 167.350 126.260 167.450 ;
        RECT 107.960 165.090 108.130 167.350 ;
        RECT 108.855 166.780 116.895 166.950 ;
        RECT 108.470 165.720 108.640 166.720 ;
        RECT 117.110 165.720 117.280 166.720 ;
        RECT 108.855 165.490 116.895 165.660 ;
        RECT 117.620 165.090 118.590 167.350 ;
        RECT 120.010 166.790 126.260 167.350 ;
        RECT 120.010 166.770 125.180 166.790 ;
        RECT 120.010 166.700 124.000 166.770 ;
        RECT 120.010 165.430 121.930 166.700 ;
        RECT 123.440 166.690 124.000 166.700 ;
        RECT 123.670 165.600 124.000 166.690 ;
        RECT 124.370 166.220 125.410 166.390 ;
        RECT 124.370 165.780 125.410 165.950 ;
        RECT 125.580 165.920 125.750 166.250 ;
        RECT 123.830 165.380 124.000 165.600 ;
        RECT 126.090 165.380 126.260 166.790 ;
        RECT 123.830 165.210 126.260 165.380 ;
        RECT 127.840 167.300 138.470 167.470 ;
        RECT 140.050 176.630 146.280 176.790 ;
        RECT 140.050 174.370 140.720 176.630 ;
        RECT 141.390 176.060 145.430 176.230 ;
        RECT 141.050 175.000 141.220 176.000 ;
        RECT 145.600 175.000 145.770 176.000 ;
        RECT 141.390 174.770 145.430 174.940 ;
        RECT 146.110 174.370 146.280 176.630 ;
        RECT 140.050 174.200 146.280 174.370 ;
        RECT 140.050 170.940 140.720 174.200 ;
        RECT 141.390 173.630 145.430 173.800 ;
        RECT 141.050 171.570 141.220 173.570 ;
        RECT 145.600 171.570 145.770 173.570 ;
        RECT 141.390 171.340 145.430 171.510 ;
        RECT 146.110 170.940 146.280 174.200 ;
        RECT 140.050 170.770 146.280 170.940 ;
        RECT 140.050 167.510 140.720 170.770 ;
        RECT 141.390 170.200 145.430 170.370 ;
        RECT 141.050 168.140 141.220 170.140 ;
        RECT 145.600 168.140 145.770 170.140 ;
        RECT 141.390 167.910 145.430 168.080 ;
        RECT 146.110 167.510 146.280 170.770 ;
        RECT 140.050 167.500 146.280 167.510 ;
        RECT 147.870 176.770 157.700 176.810 ;
        RECT 147.870 176.640 158.500 176.770 ;
        RECT 147.870 174.380 148.040 176.640 ;
        RECT 148.765 176.070 156.805 176.240 ;
        RECT 148.380 175.010 148.550 176.010 ;
        RECT 157.020 175.010 157.190 176.010 ;
        RECT 148.765 174.780 156.805 174.950 ;
        RECT 157.530 174.380 158.500 176.640 ;
        RECT 147.870 174.210 158.500 174.380 ;
        RECT 147.870 170.950 148.040 174.210 ;
        RECT 148.765 173.640 156.805 173.810 ;
        RECT 148.380 171.580 148.550 173.580 ;
        RECT 157.020 171.580 157.190 173.580 ;
        RECT 148.765 171.350 156.805 171.520 ;
        RECT 157.530 170.950 158.500 174.210 ;
        RECT 147.870 170.780 158.500 170.950 ;
        RECT 147.870 167.520 148.040 170.780 ;
        RECT 148.765 170.210 156.805 170.380 ;
        RECT 148.380 168.150 148.550 170.150 ;
        RECT 157.020 168.150 157.190 170.150 ;
        RECT 148.765 167.920 156.805 168.090 ;
        RECT 157.530 167.520 158.500 170.780 ;
        RECT 140.050 167.400 146.290 167.500 ;
        RECT 107.960 165.060 118.590 165.090 ;
        RECT 72.295 163.875 77.640 164.310 ;
        RECT 77.815 163.875 83.160 164.310 ;
        RECT 83.335 163.875 88.680 164.310 ;
        RECT 89.315 163.875 90.525 164.965 ;
        RECT 107.930 164.950 118.590 165.060 ;
        RECT 127.840 165.040 128.010 167.300 ;
        RECT 128.735 166.730 136.775 166.900 ;
        RECT 128.350 165.670 128.520 166.670 ;
        RECT 136.990 165.670 137.160 166.670 ;
        RECT 128.735 165.440 136.775 165.610 ;
        RECT 137.500 165.040 138.470 167.300 ;
        RECT 140.040 166.840 146.290 167.400 ;
        RECT 140.040 166.820 145.210 166.840 ;
        RECT 140.040 166.750 144.030 166.820 ;
        RECT 140.040 165.480 141.960 166.750 ;
        RECT 143.470 166.740 144.030 166.750 ;
        RECT 143.700 165.650 144.030 166.740 ;
        RECT 144.400 166.270 145.440 166.440 ;
        RECT 144.400 165.830 145.440 166.000 ;
        RECT 145.610 165.970 145.780 166.300 ;
        RECT 143.860 165.430 144.030 165.650 ;
        RECT 146.120 165.430 146.290 166.840 ;
        RECT 143.860 165.260 146.290 165.430 ;
        RECT 147.870 167.350 158.500 167.520 ;
        RECT 147.870 165.090 148.040 167.350 ;
        RECT 148.765 166.780 156.805 166.950 ;
        RECT 148.380 165.720 148.550 166.720 ;
        RECT 157.020 165.720 157.190 166.720 ;
        RECT 148.765 165.490 156.805 165.660 ;
        RECT 157.530 165.090 158.500 167.350 ;
        RECT 147.870 165.060 158.500 165.090 ;
        RECT 127.840 165.010 138.470 165.040 ;
        RECT 106.180 164.900 118.590 164.950 ;
        RECT 127.810 164.900 138.470 165.010 ;
        RECT 147.840 164.950 158.500 165.060 ;
        RECT 146.090 164.900 158.500 164.950 ;
        RECT 101.840 164.730 118.590 164.900 ;
        RECT 126.060 164.850 138.470 164.900 ;
        RECT 11.950 163.705 90.610 163.875 ;
        RECT 12.035 162.615 13.245 163.705 ;
        RECT 13.415 163.270 18.760 163.705 ;
        RECT 18.935 163.270 24.280 163.705 ;
        RECT 12.035 161.905 12.555 162.445 ;
        RECT 12.725 162.075 13.245 162.615 ;
        RECT 12.035 161.155 13.245 161.905 ;
        RECT 15.000 161.700 15.340 162.530 ;
        RECT 16.820 162.020 17.170 163.270 ;
        RECT 20.520 161.700 20.860 162.530 ;
        RECT 22.340 162.020 22.690 163.270 ;
        RECT 24.915 162.540 25.205 163.705 ;
        RECT 25.375 163.195 25.635 163.705 ;
        RECT 25.375 162.145 25.715 163.025 ;
        RECT 25.885 162.315 26.055 163.535 ;
        RECT 26.295 163.200 26.910 163.705 ;
        RECT 26.295 162.665 26.545 163.030 ;
        RECT 26.715 163.025 26.910 163.200 ;
        RECT 27.080 163.195 27.555 163.535 ;
        RECT 27.725 163.160 27.940 163.705 ;
        RECT 26.715 162.835 27.045 163.025 ;
        RECT 27.265 162.665 27.980 162.960 ;
        RECT 28.150 162.835 28.425 163.535 ;
        RECT 26.295 162.495 28.085 162.665 ;
        RECT 25.885 162.065 26.680 162.315 ;
        RECT 25.885 161.975 26.135 162.065 ;
        RECT 13.415 161.155 18.760 161.700 ;
        RECT 18.935 161.155 24.280 161.700 ;
        RECT 24.915 161.155 25.205 161.880 ;
        RECT 25.375 161.155 25.635 161.975 ;
        RECT 25.805 161.555 26.135 161.975 ;
        RECT 26.850 161.640 27.105 162.495 ;
        RECT 26.315 161.375 27.105 161.640 ;
        RECT 27.275 161.795 27.685 162.315 ;
        RECT 27.855 162.065 28.085 162.495 ;
        RECT 28.255 161.805 28.425 162.835 ;
        RECT 28.780 162.735 29.170 162.910 ;
        RECT 29.655 162.905 29.985 163.705 ;
        RECT 30.155 162.915 30.690 163.535 ;
        RECT 28.780 162.565 30.205 162.735 ;
        RECT 28.655 161.835 29.010 162.395 ;
        RECT 27.275 161.375 27.475 161.795 ;
        RECT 27.665 161.155 27.995 161.615 ;
        RECT 28.165 161.325 28.425 161.805 ;
        RECT 29.180 161.665 29.350 162.565 ;
        RECT 29.520 161.835 29.785 162.395 ;
        RECT 30.035 162.065 30.205 162.565 ;
        RECT 30.375 161.895 30.690 162.915 ;
        RECT 31.510 162.695 31.810 163.535 ;
        RECT 32.005 162.865 32.255 163.705 ;
        RECT 32.845 163.115 33.650 163.535 ;
        RECT 32.425 162.945 33.990 163.115 ;
        RECT 32.425 162.695 32.595 162.945 ;
        RECT 31.510 162.525 32.595 162.695 ;
        RECT 31.355 162.065 31.685 162.355 ;
        RECT 31.855 161.895 32.025 162.525 ;
        RECT 32.765 162.395 33.085 162.775 ;
        RECT 33.275 162.685 33.650 162.775 ;
        RECT 33.255 162.515 33.650 162.685 ;
        RECT 33.820 162.695 33.990 162.945 ;
        RECT 34.160 162.865 34.490 163.705 ;
        RECT 34.660 162.945 35.325 163.535 ;
        RECT 33.820 162.525 34.740 162.695 ;
        RECT 32.195 162.145 32.525 162.355 ;
        RECT 32.705 162.145 33.085 162.395 ;
        RECT 33.275 162.355 33.650 162.515 ;
        RECT 34.570 162.355 34.740 162.525 ;
        RECT 33.275 162.145 33.760 162.355 ;
        RECT 33.950 162.145 34.400 162.355 ;
        RECT 34.570 162.145 34.905 162.355 ;
        RECT 35.075 161.975 35.325 162.945 ;
        RECT 28.760 161.155 29.000 161.665 ;
        RECT 29.180 161.335 29.460 161.665 ;
        RECT 29.690 161.155 29.905 161.665 ;
        RECT 30.075 161.325 30.690 161.895 ;
        RECT 31.515 161.715 32.025 161.895 ;
        RECT 32.430 161.805 34.130 161.975 ;
        RECT 32.430 161.715 32.815 161.805 ;
        RECT 31.515 161.325 31.845 161.715 ;
        RECT 32.015 161.375 33.200 161.545 ;
        RECT 33.460 161.155 33.630 161.625 ;
        RECT 33.800 161.340 34.130 161.805 ;
        RECT 34.300 161.155 34.470 161.975 ;
        RECT 34.640 161.335 35.325 161.975 ;
        RECT 35.495 162.100 35.775 163.535 ;
        RECT 35.945 162.930 36.655 163.705 ;
        RECT 36.825 162.760 37.155 163.535 ;
        RECT 36.005 162.545 37.155 162.760 ;
        RECT 35.495 161.325 35.835 162.100 ;
        RECT 36.005 161.975 36.290 162.545 ;
        RECT 36.475 162.145 36.945 162.375 ;
        RECT 37.350 162.345 37.565 163.460 ;
        RECT 37.745 162.985 38.075 163.705 ;
        RECT 39.195 163.195 39.495 163.705 ;
        RECT 39.665 163.195 40.045 163.365 ;
        RECT 40.625 163.195 41.255 163.705 ;
        RECT 39.665 163.025 39.835 163.195 ;
        RECT 41.425 163.025 41.755 163.535 ;
        RECT 41.925 163.195 42.225 163.705 ;
        RECT 39.175 162.825 39.835 163.025 ;
        RECT 40.005 162.855 42.225 163.025 ;
        RECT 37.855 162.345 38.085 162.685 ;
        RECT 37.115 162.165 37.565 162.345 ;
        RECT 37.115 162.145 37.445 162.165 ;
        RECT 37.755 162.145 38.085 162.345 ;
        RECT 36.005 161.785 36.715 161.975 ;
        RECT 36.415 161.645 36.715 161.785 ;
        RECT 36.905 161.785 38.085 161.975 ;
        RECT 36.905 161.705 37.235 161.785 ;
        RECT 36.415 161.635 36.730 161.645 ;
        RECT 36.415 161.625 36.740 161.635 ;
        RECT 36.415 161.620 36.750 161.625 ;
        RECT 36.005 161.155 36.175 161.615 ;
        RECT 36.415 161.610 36.755 161.620 ;
        RECT 36.415 161.605 36.760 161.610 ;
        RECT 36.415 161.595 36.765 161.605 ;
        RECT 36.415 161.590 36.770 161.595 ;
        RECT 36.415 161.325 36.775 161.590 ;
        RECT 37.405 161.155 37.575 161.615 ;
        RECT 37.745 161.325 38.085 161.785 ;
        RECT 39.175 161.895 39.345 162.825 ;
        RECT 40.005 162.655 40.175 162.855 ;
        RECT 39.515 162.485 40.175 162.655 ;
        RECT 40.345 162.515 41.885 162.685 ;
        RECT 39.515 162.065 39.685 162.485 ;
        RECT 40.345 162.315 40.515 162.515 ;
        RECT 39.915 162.145 40.515 162.315 ;
        RECT 40.685 162.145 41.380 162.345 ;
        RECT 41.640 162.065 41.885 162.515 ;
        RECT 40.005 161.895 40.915 161.975 ;
        RECT 39.175 161.415 39.495 161.895 ;
        RECT 39.665 161.805 40.915 161.895 ;
        RECT 39.665 161.725 40.175 161.805 ;
        RECT 39.665 161.325 39.895 161.725 ;
        RECT 40.065 161.155 40.415 161.545 ;
        RECT 40.585 161.325 40.915 161.805 ;
        RECT 41.085 161.155 41.255 161.975 ;
        RECT 42.055 161.895 42.225 162.855 ;
        RECT 42.395 162.615 44.985 163.705 ;
        RECT 45.620 163.280 45.955 163.705 ;
        RECT 46.125 163.100 46.310 163.505 ;
        RECT 41.760 161.350 42.225 161.895 ;
        RECT 42.395 161.925 43.605 162.445 ;
        RECT 43.775 162.095 44.985 162.615 ;
        RECT 45.645 162.925 46.310 163.100 ;
        RECT 46.515 162.925 46.845 163.705 ;
        RECT 42.395 161.155 44.985 161.925 ;
        RECT 45.645 161.895 45.985 162.925 ;
        RECT 47.015 162.735 47.285 163.505 ;
        RECT 46.155 162.565 47.285 162.735 ;
        RECT 46.155 162.065 46.405 162.565 ;
        RECT 45.645 161.725 46.330 161.895 ;
        RECT 46.585 161.815 46.945 162.395 ;
        RECT 45.620 161.155 45.955 161.555 ;
        RECT 46.125 161.325 46.330 161.725 ;
        RECT 47.115 161.655 47.285 162.565 ;
        RECT 46.540 161.155 46.815 161.635 ;
        RECT 47.025 161.325 47.285 161.655 ;
        RECT 47.465 162.645 47.795 163.495 ;
        RECT 47.465 161.880 47.655 162.645 ;
        RECT 47.965 162.565 48.215 163.705 ;
        RECT 48.405 163.065 48.655 163.485 ;
        RECT 48.885 163.235 49.215 163.705 ;
        RECT 49.445 163.065 49.695 163.485 ;
        RECT 48.405 162.895 49.695 163.065 ;
        RECT 49.875 163.065 50.205 163.495 ;
        RECT 49.875 162.895 50.330 163.065 ;
        RECT 48.395 162.395 48.610 162.725 ;
        RECT 47.825 162.065 48.135 162.395 ;
        RECT 48.305 162.065 48.610 162.395 ;
        RECT 48.785 162.065 49.070 162.725 ;
        RECT 49.265 162.065 49.530 162.725 ;
        RECT 49.745 162.065 49.990 162.725 ;
        RECT 47.965 161.895 48.135 162.065 ;
        RECT 50.160 161.895 50.330 162.895 ;
        RECT 50.675 162.540 50.965 163.705 ;
        RECT 51.135 162.615 52.345 163.705 ;
        RECT 47.465 161.370 47.795 161.880 ;
        RECT 47.965 161.725 50.330 161.895 ;
        RECT 51.135 161.905 51.655 162.445 ;
        RECT 51.825 162.075 52.345 162.615 ;
        RECT 52.550 162.915 53.085 163.535 ;
        RECT 47.965 161.155 48.295 161.555 ;
        RECT 49.345 161.385 49.675 161.725 ;
        RECT 49.845 161.155 50.175 161.555 ;
        RECT 50.675 161.155 50.965 161.880 ;
        RECT 51.135 161.155 52.345 161.905 ;
        RECT 52.550 161.895 52.865 162.915 ;
        RECT 53.255 162.905 53.585 163.705 ;
        RECT 54.070 162.735 54.460 162.910 ;
        RECT 53.035 162.565 54.460 162.735 ;
        RECT 54.905 162.775 55.075 163.535 ;
        RECT 55.290 162.945 55.620 163.705 ;
        RECT 54.905 162.605 55.620 162.775 ;
        RECT 55.790 162.630 56.045 163.535 ;
        RECT 53.035 162.065 53.205 162.565 ;
        RECT 52.550 161.325 53.165 161.895 ;
        RECT 53.455 161.835 53.720 162.395 ;
        RECT 53.890 161.665 54.060 162.565 ;
        RECT 54.230 161.835 54.585 162.395 ;
        RECT 54.815 162.055 55.170 162.425 ;
        RECT 55.450 162.395 55.620 162.605 ;
        RECT 55.450 162.065 55.705 162.395 ;
        RECT 55.450 161.875 55.620 162.065 ;
        RECT 55.875 161.900 56.045 162.630 ;
        RECT 56.220 162.555 56.480 163.705 ;
        RECT 57.585 162.565 57.915 163.705 ;
        RECT 58.445 162.735 58.775 163.520 ;
        RECT 58.095 162.565 58.775 162.735 ;
        RECT 58.960 163.315 59.295 163.535 ;
        RECT 60.300 163.325 60.655 163.705 ;
        RECT 58.960 162.695 59.215 163.315 ;
        RECT 59.465 163.155 59.695 163.195 ;
        RECT 60.825 163.155 61.075 163.535 ;
        RECT 59.465 162.955 61.075 163.155 ;
        RECT 59.465 162.865 59.650 162.955 ;
        RECT 60.240 162.945 61.075 162.955 ;
        RECT 61.325 162.925 61.575 163.705 ;
        RECT 61.745 162.855 62.005 163.535 ;
        RECT 62.675 163.245 62.890 163.705 ;
        RECT 63.060 163.075 63.390 163.535 ;
        RECT 59.805 162.755 60.135 162.785 ;
        RECT 59.805 162.695 61.605 162.755 ;
        RECT 58.960 162.585 61.665 162.695 ;
        RECT 57.575 162.145 57.925 162.395 ;
        RECT 54.905 161.705 55.620 161.875 ;
        RECT 53.335 161.155 53.550 161.665 ;
        RECT 53.780 161.335 54.060 161.665 ;
        RECT 54.240 161.155 54.480 161.665 ;
        RECT 54.905 161.325 55.075 161.705 ;
        RECT 55.290 161.155 55.620 161.535 ;
        RECT 55.790 161.325 56.045 161.900 ;
        RECT 56.220 161.155 56.480 161.995 ;
        RECT 58.095 161.965 58.265 162.565 ;
        RECT 58.960 162.525 60.135 162.585 ;
        RECT 61.465 162.550 61.665 162.585 ;
        RECT 58.435 162.145 58.785 162.395 ;
        RECT 58.955 162.145 59.445 162.345 ;
        RECT 59.635 162.145 60.110 162.355 ;
        RECT 57.585 161.155 57.855 161.965 ;
        RECT 58.025 161.325 58.355 161.965 ;
        RECT 58.525 161.155 58.765 161.965 ;
        RECT 58.960 161.155 59.415 161.920 ;
        RECT 59.890 161.745 60.110 162.145 ;
        RECT 60.355 162.145 60.685 162.355 ;
        RECT 60.355 161.745 60.565 162.145 ;
        RECT 60.855 162.110 61.265 162.415 ;
        RECT 61.495 161.975 61.665 162.550 ;
        RECT 61.395 161.855 61.665 161.975 ;
        RECT 60.820 161.810 61.665 161.855 ;
        RECT 60.820 161.685 61.575 161.810 ;
        RECT 60.820 161.535 60.990 161.685 ;
        RECT 61.835 161.665 62.005 162.855 ;
        RECT 61.775 161.655 62.005 161.665 ;
        RECT 59.690 161.325 60.990 161.535 ;
        RECT 61.245 161.155 61.575 161.515 ;
        RECT 61.745 161.325 62.005 161.655 ;
        RECT 62.220 162.905 63.390 163.075 ;
        RECT 63.560 162.905 63.810 163.705 ;
        RECT 62.220 161.615 62.590 162.905 ;
        RECT 64.020 162.735 64.300 162.895 ;
        RECT 62.965 162.565 64.300 162.735 ;
        RECT 64.475 162.615 66.145 163.705 ;
        RECT 62.965 162.395 63.135 162.565 ;
        RECT 62.760 162.145 63.135 162.395 ;
        RECT 63.305 162.145 63.780 162.385 ;
        RECT 63.950 162.145 64.300 162.385 ;
        RECT 62.965 161.975 63.135 162.145 ;
        RECT 62.965 161.805 64.300 161.975 ;
        RECT 62.220 161.325 62.970 161.615 ;
        RECT 63.480 161.155 63.810 161.615 ;
        RECT 64.030 161.595 64.300 161.805 ;
        RECT 64.475 161.925 65.225 162.445 ;
        RECT 65.395 162.095 66.145 162.615 ;
        RECT 66.315 162.855 66.695 163.535 ;
        RECT 67.285 162.855 67.455 163.705 ;
        RECT 67.625 163.025 67.955 163.535 ;
        RECT 68.125 163.195 68.295 163.705 ;
        RECT 68.465 163.025 68.865 163.535 ;
        RECT 67.625 162.855 68.865 163.025 ;
        RECT 64.475 161.155 66.145 161.925 ;
        RECT 66.315 161.895 66.485 162.855 ;
        RECT 66.655 162.515 67.960 162.685 ;
        RECT 69.045 162.605 69.365 163.535 ;
        RECT 69.620 163.085 69.795 163.535 ;
        RECT 69.965 163.265 70.295 163.705 ;
        RECT 70.600 163.115 70.770 163.535 ;
        RECT 71.005 163.295 71.675 163.705 ;
        RECT 71.890 163.115 72.060 163.535 ;
        RECT 72.260 163.295 72.590 163.705 ;
        RECT 69.620 162.915 70.250 163.085 ;
        RECT 66.655 162.065 66.900 162.515 ;
        RECT 67.070 162.145 67.620 162.345 ;
        RECT 67.790 162.315 67.960 162.515 ;
        RECT 68.735 162.435 69.365 162.605 ;
        RECT 67.790 162.145 68.165 162.315 ;
        RECT 68.335 161.895 68.565 162.395 ;
        RECT 66.315 161.725 68.565 161.895 ;
        RECT 66.365 161.155 66.695 161.545 ;
        RECT 66.865 161.405 67.035 161.725 ;
        RECT 68.735 161.555 68.905 162.435 ;
        RECT 69.535 162.065 69.900 162.745 ;
        RECT 70.080 162.395 70.250 162.915 ;
        RECT 70.600 162.945 72.615 163.115 ;
        RECT 70.080 162.065 70.430 162.395 ;
        RECT 67.205 161.155 67.535 161.545 ;
        RECT 67.950 161.385 68.905 161.555 ;
        RECT 69.075 161.155 69.365 161.990 ;
        RECT 70.080 161.895 70.250 162.065 ;
        RECT 69.620 161.725 70.250 161.895 ;
        RECT 69.620 161.325 69.795 161.725 ;
        RECT 70.600 161.655 70.770 162.945 ;
        RECT 69.965 161.155 70.295 161.535 ;
        RECT 70.540 161.325 70.770 161.655 ;
        RECT 70.970 161.490 71.250 162.765 ;
        RECT 71.475 162.345 71.745 162.765 ;
        RECT 71.435 162.175 71.745 162.345 ;
        RECT 71.475 161.490 71.745 162.175 ;
        RECT 71.935 161.735 72.275 162.765 ;
        RECT 72.445 162.395 72.615 162.945 ;
        RECT 72.785 162.565 73.045 163.535 ;
        RECT 73.215 162.615 75.805 163.705 ;
        RECT 72.445 162.065 72.705 162.395 ;
        RECT 72.875 161.875 73.045 162.565 ;
        RECT 72.205 161.155 72.535 161.535 ;
        RECT 72.705 161.410 73.045 161.875 ;
        RECT 73.215 161.925 74.425 162.445 ;
        RECT 74.595 162.095 75.805 162.615 ;
        RECT 76.435 162.540 76.725 163.705 ;
        RECT 76.895 163.270 82.240 163.705 ;
        RECT 82.415 163.270 87.760 163.705 ;
        RECT 72.705 161.365 73.040 161.410 ;
        RECT 73.215 161.155 75.805 161.925 ;
        RECT 76.435 161.155 76.725 161.880 ;
        RECT 78.480 161.700 78.820 162.530 ;
        RECT 80.300 162.020 80.650 163.270 ;
        RECT 84.000 161.700 84.340 162.530 ;
        RECT 85.820 162.020 86.170 163.270 ;
        RECT 87.935 162.615 89.145 163.705 ;
        RECT 87.935 161.905 88.455 162.445 ;
        RECT 88.625 162.075 89.145 162.615 ;
        RECT 89.315 162.615 90.525 163.705 ;
        RECT 101.840 163.320 102.010 164.730 ;
        RECT 102.380 164.160 105.420 164.330 ;
        RECT 102.380 163.720 105.420 163.890 ;
        RECT 105.635 163.860 105.805 164.190 ;
        RECT 106.140 163.970 118.590 164.730 ;
        RECT 121.720 164.680 138.470 164.850 ;
        RECT 106.140 163.960 118.480 163.970 ;
        RECT 106.140 163.950 112.020 163.960 ;
        RECT 106.140 163.930 106.710 163.950 ;
        RECT 107.930 163.940 112.020 163.950 ;
        RECT 106.150 163.320 106.320 163.930 ;
        RECT 101.840 163.150 106.320 163.320 ;
        RECT 121.720 163.270 121.890 164.680 ;
        RECT 122.260 164.110 125.300 164.280 ;
        RECT 122.260 163.670 125.300 163.840 ;
        RECT 125.515 163.810 125.685 164.140 ;
        RECT 126.020 163.920 138.470 164.680 ;
        RECT 141.750 164.730 158.500 164.900 ;
        RECT 126.020 163.910 138.360 163.920 ;
        RECT 126.020 163.900 131.900 163.910 ;
        RECT 126.020 163.880 126.590 163.900 ;
        RECT 127.810 163.890 131.900 163.900 ;
        RECT 126.030 163.270 126.200 163.880 ;
        RECT 121.720 163.100 126.200 163.270 ;
        RECT 141.750 163.320 141.920 164.730 ;
        RECT 142.290 164.160 145.330 164.330 ;
        RECT 142.290 163.720 145.330 163.890 ;
        RECT 145.545 163.860 145.715 164.190 ;
        RECT 146.050 163.970 158.500 164.730 ;
        RECT 146.050 163.960 158.390 163.970 ;
        RECT 146.050 163.950 151.930 163.960 ;
        RECT 146.050 163.930 146.620 163.950 ;
        RECT 147.840 163.940 151.930 163.950 ;
        RECT 146.060 163.320 146.230 163.930 ;
        RECT 141.750 163.150 146.230 163.320 ;
        RECT 89.315 162.075 89.835 162.615 ;
        RECT 90.005 161.905 90.525 162.445 ;
        RECT 76.895 161.155 82.240 161.700 ;
        RECT 82.415 161.155 87.760 161.700 ;
        RECT 87.935 161.155 89.145 161.905 ;
        RECT 89.315 161.155 90.525 161.905 ;
        RECT 100.630 161.790 106.370 161.800 ;
        RECT 100.140 161.630 106.370 161.790 ;
        RECT 11.950 160.985 90.610 161.155 ;
        RECT 12.035 160.235 13.245 160.985 ;
        RECT 13.415 160.440 18.760 160.985 ;
        RECT 12.035 159.695 12.555 160.235 ;
        RECT 12.725 159.525 13.245 160.065 ;
        RECT 15.000 159.610 15.340 160.440 ;
        RECT 18.935 160.215 22.445 160.985 ;
        RECT 23.125 160.330 23.455 160.765 ;
        RECT 23.625 160.375 23.795 160.985 ;
        RECT 23.075 160.245 23.455 160.330 ;
        RECT 23.965 160.245 24.295 160.770 ;
        RECT 24.555 160.455 24.765 160.985 ;
        RECT 25.040 160.535 25.825 160.705 ;
        RECT 25.995 160.535 26.400 160.705 ;
        RECT 12.035 158.435 13.245 159.525 ;
        RECT 16.820 158.870 17.170 160.120 ;
        RECT 18.935 159.695 20.585 160.215 ;
        RECT 23.075 160.205 23.300 160.245 ;
        RECT 20.755 159.525 22.445 160.045 ;
        RECT 13.415 158.435 18.760 158.870 ;
        RECT 18.935 158.435 22.445 159.525 ;
        RECT 23.075 159.625 23.245 160.205 ;
        RECT 23.965 160.075 24.165 160.245 ;
        RECT 25.040 160.075 25.210 160.535 ;
        RECT 23.415 159.745 24.165 160.075 ;
        RECT 24.335 159.745 25.210 160.075 ;
        RECT 23.075 159.575 23.290 159.625 ;
        RECT 23.075 159.495 23.465 159.575 ;
        RECT 23.135 158.650 23.465 159.495 ;
        RECT 23.975 159.540 24.165 159.745 ;
        RECT 23.635 158.435 23.805 159.445 ;
        RECT 23.975 159.165 24.870 159.540 ;
        RECT 23.975 158.605 24.315 159.165 ;
        RECT 24.545 158.435 24.860 158.935 ;
        RECT 25.040 158.905 25.210 159.745 ;
        RECT 25.380 160.035 25.845 160.365 ;
        RECT 26.230 160.305 26.400 160.535 ;
        RECT 26.580 160.485 26.950 160.985 ;
        RECT 27.270 160.535 27.945 160.705 ;
        RECT 28.140 160.535 28.475 160.705 ;
        RECT 25.380 159.075 25.700 160.035 ;
        RECT 26.230 160.005 27.060 160.305 ;
        RECT 25.870 159.105 26.060 159.825 ;
        RECT 26.230 158.935 26.400 160.005 ;
        RECT 26.860 159.975 27.060 160.005 ;
        RECT 26.570 159.755 26.740 159.825 ;
        RECT 27.270 159.755 27.440 160.535 ;
        RECT 28.305 160.395 28.475 160.535 ;
        RECT 28.645 160.525 28.895 160.985 ;
        RECT 26.570 159.585 27.440 159.755 ;
        RECT 27.610 160.115 28.135 160.335 ;
        RECT 28.305 160.265 28.530 160.395 ;
        RECT 26.570 159.495 27.080 159.585 ;
        RECT 25.040 158.735 25.925 158.905 ;
        RECT 26.150 158.605 26.400 158.935 ;
        RECT 26.570 158.435 26.740 159.235 ;
        RECT 26.910 158.880 27.080 159.495 ;
        RECT 27.610 159.415 27.780 160.115 ;
        RECT 27.250 159.050 27.780 159.415 ;
        RECT 27.950 159.350 28.190 159.945 ;
        RECT 28.360 159.160 28.530 160.265 ;
        RECT 28.700 159.405 28.980 160.355 ;
        RECT 28.225 159.030 28.530 159.160 ;
        RECT 26.910 158.710 28.015 158.880 ;
        RECT 28.225 158.605 28.475 159.030 ;
        RECT 28.645 158.435 28.910 158.895 ;
        RECT 29.150 158.605 29.335 160.725 ;
        RECT 29.505 160.605 29.835 160.985 ;
        RECT 30.005 160.435 30.175 160.725 ;
        RECT 29.510 160.265 30.175 160.435 ;
        RECT 29.510 159.275 29.740 160.265 ;
        RECT 29.910 159.445 30.260 160.095 ;
        RECT 31.355 160.040 31.695 160.815 ;
        RECT 31.865 160.525 32.035 160.985 ;
        RECT 32.275 160.550 32.635 160.815 ;
        RECT 32.275 160.545 32.630 160.550 ;
        RECT 32.275 160.535 32.625 160.545 ;
        RECT 32.275 160.530 32.620 160.535 ;
        RECT 32.275 160.520 32.615 160.530 ;
        RECT 33.265 160.525 33.435 160.985 ;
        RECT 32.275 160.515 32.610 160.520 ;
        RECT 32.275 160.505 32.600 160.515 ;
        RECT 32.275 160.495 32.590 160.505 ;
        RECT 32.275 160.355 32.575 160.495 ;
        RECT 31.865 160.165 32.575 160.355 ;
        RECT 32.765 160.355 33.095 160.435 ;
        RECT 33.605 160.355 33.945 160.815 ;
        RECT 32.765 160.165 33.945 160.355 ;
        RECT 34.115 160.215 35.785 160.985 ;
        RECT 29.510 159.105 30.175 159.275 ;
        RECT 29.505 158.435 29.835 158.935 ;
        RECT 30.005 158.605 30.175 159.105 ;
        RECT 31.355 158.605 31.635 160.040 ;
        RECT 31.865 159.595 32.150 160.165 ;
        RECT 32.335 159.765 32.805 159.995 ;
        RECT 32.975 159.975 33.305 159.995 ;
        RECT 32.975 159.795 33.425 159.975 ;
        RECT 33.615 159.795 33.945 159.995 ;
        RECT 31.865 159.380 33.015 159.595 ;
        RECT 31.805 158.435 32.515 159.210 ;
        RECT 32.685 158.605 33.015 159.380 ;
        RECT 33.210 158.680 33.425 159.795 ;
        RECT 33.715 159.455 33.945 159.795 ;
        RECT 34.115 159.695 34.865 160.215 ;
        RECT 36.415 160.185 36.725 160.985 ;
        RECT 36.930 160.185 37.625 160.815 ;
        RECT 37.795 160.260 38.085 160.985 ;
        RECT 38.805 160.435 38.975 160.725 ;
        RECT 39.145 160.605 39.475 160.985 ;
        RECT 38.805 160.265 39.470 160.435 ;
        RECT 35.035 159.525 35.785 160.045 ;
        RECT 36.425 159.745 36.760 160.015 ;
        RECT 36.930 159.585 37.100 160.185 ;
        RECT 37.270 159.745 37.605 159.995 ;
        RECT 33.605 158.435 33.935 159.155 ;
        RECT 34.115 158.435 35.785 159.525 ;
        RECT 36.415 158.435 36.695 159.575 ;
        RECT 36.865 158.605 37.195 159.585 ;
        RECT 37.365 158.435 37.625 159.575 ;
        RECT 37.795 158.435 38.085 159.600 ;
        RECT 38.720 159.445 39.070 160.095 ;
        RECT 39.240 159.275 39.470 160.265 ;
        RECT 38.805 159.105 39.470 159.275 ;
        RECT 38.805 158.605 38.975 159.105 ;
        RECT 39.145 158.435 39.475 158.935 ;
        RECT 39.645 158.605 39.830 160.725 ;
        RECT 40.085 160.525 40.335 160.985 ;
        RECT 40.505 160.535 40.840 160.705 ;
        RECT 41.035 160.535 41.710 160.705 ;
        RECT 40.505 160.395 40.675 160.535 ;
        RECT 40.000 159.405 40.280 160.355 ;
        RECT 40.450 160.265 40.675 160.395 ;
        RECT 40.450 159.160 40.620 160.265 ;
        RECT 40.845 160.115 41.370 160.335 ;
        RECT 40.790 159.350 41.030 159.945 ;
        RECT 41.200 159.415 41.370 160.115 ;
        RECT 41.540 159.755 41.710 160.535 ;
        RECT 42.030 160.485 42.400 160.985 ;
        RECT 42.580 160.535 42.985 160.705 ;
        RECT 43.155 160.535 43.940 160.705 ;
        RECT 42.580 160.305 42.750 160.535 ;
        RECT 41.920 160.005 42.750 160.305 ;
        RECT 43.135 160.035 43.600 160.365 ;
        RECT 41.920 159.975 42.120 160.005 ;
        RECT 42.240 159.755 42.410 159.825 ;
        RECT 41.540 159.585 42.410 159.755 ;
        RECT 41.900 159.495 42.410 159.585 ;
        RECT 40.450 159.030 40.755 159.160 ;
        RECT 41.200 159.050 41.730 159.415 ;
        RECT 40.070 158.435 40.335 158.895 ;
        RECT 40.505 158.605 40.755 159.030 ;
        RECT 41.900 158.880 42.070 159.495 ;
        RECT 40.965 158.710 42.070 158.880 ;
        RECT 42.240 158.435 42.410 159.235 ;
        RECT 42.580 158.935 42.750 160.005 ;
        RECT 42.920 159.105 43.110 159.825 ;
        RECT 43.280 159.075 43.600 160.035 ;
        RECT 43.770 160.075 43.940 160.535 ;
        RECT 44.215 160.455 44.425 160.985 ;
        RECT 44.685 160.245 45.015 160.770 ;
        RECT 45.185 160.375 45.355 160.985 ;
        RECT 45.525 160.330 45.855 160.765 ;
        RECT 46.165 160.435 46.335 160.725 ;
        RECT 46.505 160.605 46.835 160.985 ;
        RECT 45.525 160.245 45.905 160.330 ;
        RECT 46.165 160.265 46.830 160.435 ;
        RECT 44.815 160.075 45.015 160.245 ;
        RECT 45.680 160.205 45.905 160.245 ;
        RECT 43.770 159.745 44.645 160.075 ;
        RECT 44.815 159.745 45.565 160.075 ;
        RECT 42.580 158.605 42.830 158.935 ;
        RECT 43.770 158.905 43.940 159.745 ;
        RECT 44.815 159.540 45.005 159.745 ;
        RECT 45.735 159.625 45.905 160.205 ;
        RECT 45.690 159.575 45.905 159.625 ;
        RECT 44.110 159.165 45.005 159.540 ;
        RECT 45.515 159.495 45.905 159.575 ;
        RECT 43.055 158.735 43.940 158.905 ;
        RECT 44.120 158.435 44.435 158.935 ;
        RECT 44.665 158.605 45.005 159.165 ;
        RECT 45.175 158.435 45.345 159.445 ;
        RECT 45.515 158.650 45.845 159.495 ;
        RECT 46.080 159.445 46.430 160.095 ;
        RECT 46.600 159.275 46.830 160.265 ;
        RECT 46.165 159.105 46.830 159.275 ;
        RECT 46.165 158.605 46.335 159.105 ;
        RECT 46.505 158.435 46.835 158.935 ;
        RECT 47.005 158.605 47.190 160.725 ;
        RECT 47.445 160.525 47.695 160.985 ;
        RECT 47.865 160.535 48.200 160.705 ;
        RECT 48.395 160.535 49.070 160.705 ;
        RECT 47.865 160.395 48.035 160.535 ;
        RECT 47.360 159.405 47.640 160.355 ;
        RECT 47.810 160.265 48.035 160.395 ;
        RECT 47.810 159.160 47.980 160.265 ;
        RECT 48.205 160.115 48.730 160.335 ;
        RECT 48.150 159.350 48.390 159.945 ;
        RECT 48.560 159.415 48.730 160.115 ;
        RECT 48.900 159.755 49.070 160.535 ;
        RECT 49.390 160.485 49.760 160.985 ;
        RECT 49.940 160.535 50.345 160.705 ;
        RECT 50.515 160.535 51.300 160.705 ;
        RECT 49.940 160.305 50.110 160.535 ;
        RECT 49.280 160.005 50.110 160.305 ;
        RECT 50.495 160.035 50.960 160.365 ;
        RECT 49.280 159.975 49.480 160.005 ;
        RECT 49.600 159.755 49.770 159.825 ;
        RECT 48.900 159.585 49.770 159.755 ;
        RECT 49.260 159.495 49.770 159.585 ;
        RECT 47.810 159.030 48.115 159.160 ;
        RECT 48.560 159.050 49.090 159.415 ;
        RECT 47.430 158.435 47.695 158.895 ;
        RECT 47.865 158.605 48.115 159.030 ;
        RECT 49.260 158.880 49.430 159.495 ;
        RECT 48.325 158.710 49.430 158.880 ;
        RECT 49.600 158.435 49.770 159.235 ;
        RECT 49.940 158.935 50.110 160.005 ;
        RECT 50.280 159.105 50.470 159.825 ;
        RECT 50.640 159.075 50.960 160.035 ;
        RECT 51.130 160.075 51.300 160.535 ;
        RECT 51.575 160.455 51.785 160.985 ;
        RECT 52.045 160.245 52.375 160.770 ;
        RECT 52.545 160.375 52.715 160.985 ;
        RECT 52.885 160.330 53.215 160.765 ;
        RECT 52.885 160.245 53.265 160.330 ;
        RECT 52.175 160.075 52.375 160.245 ;
        RECT 53.040 160.205 53.265 160.245 ;
        RECT 51.130 159.745 52.005 160.075 ;
        RECT 52.175 159.745 52.925 160.075 ;
        RECT 49.940 158.605 50.190 158.935 ;
        RECT 51.130 158.905 51.300 159.745 ;
        RECT 52.175 159.540 52.365 159.745 ;
        RECT 53.095 159.625 53.265 160.205 ;
        RECT 53.435 160.235 54.645 160.985 ;
        RECT 53.435 159.695 53.955 160.235 ;
        RECT 53.050 159.575 53.265 159.625 ;
        RECT 51.470 159.165 52.365 159.540 ;
        RECT 52.875 159.495 53.265 159.575 ;
        RECT 54.125 159.525 54.645 160.065 ;
        RECT 50.415 158.735 51.300 158.905 ;
        RECT 51.480 158.435 51.795 158.935 ;
        RECT 52.025 158.605 52.365 159.165 ;
        RECT 52.535 158.435 52.705 159.445 ;
        RECT 52.875 158.650 53.205 159.495 ;
        RECT 53.435 158.435 54.645 159.525 ;
        RECT 54.815 160.040 55.155 160.815 ;
        RECT 55.325 160.525 55.495 160.985 ;
        RECT 55.735 160.550 56.095 160.815 ;
        RECT 55.735 160.545 56.090 160.550 ;
        RECT 55.735 160.535 56.085 160.545 ;
        RECT 55.735 160.530 56.080 160.535 ;
        RECT 55.735 160.520 56.075 160.530 ;
        RECT 56.725 160.525 56.895 160.985 ;
        RECT 55.735 160.515 56.070 160.520 ;
        RECT 55.735 160.505 56.060 160.515 ;
        RECT 55.735 160.495 56.050 160.505 ;
        RECT 55.735 160.355 56.035 160.495 ;
        RECT 55.325 160.165 56.035 160.355 ;
        RECT 56.225 160.355 56.555 160.435 ;
        RECT 57.065 160.355 57.405 160.815 ;
        RECT 57.575 160.440 62.920 160.985 ;
        RECT 56.225 160.165 57.405 160.355 ;
        RECT 54.815 158.605 55.095 160.040 ;
        RECT 55.325 159.595 55.610 160.165 ;
        RECT 55.795 159.765 56.265 159.995 ;
        RECT 56.435 159.975 56.765 159.995 ;
        RECT 56.435 159.795 56.885 159.975 ;
        RECT 57.075 159.795 57.405 159.995 ;
        RECT 55.325 159.380 56.475 159.595 ;
        RECT 55.265 158.435 55.975 159.210 ;
        RECT 56.145 158.605 56.475 159.380 ;
        RECT 56.670 158.680 56.885 159.795 ;
        RECT 57.175 159.455 57.405 159.795 ;
        RECT 59.160 159.610 59.500 160.440 ;
        RECT 63.555 160.260 63.845 160.985 ;
        RECT 64.015 160.440 69.360 160.985 ;
        RECT 57.065 158.435 57.395 159.155 ;
        RECT 60.980 158.870 61.330 160.120 ;
        RECT 65.600 159.610 65.940 160.440 ;
        RECT 69.535 160.215 71.205 160.985 ;
        RECT 71.925 160.435 72.095 160.725 ;
        RECT 72.265 160.605 72.595 160.985 ;
        RECT 71.925 160.265 72.590 160.435 ;
        RECT 57.575 158.435 62.920 158.870 ;
        RECT 63.555 158.435 63.845 159.600 ;
        RECT 67.420 158.870 67.770 160.120 ;
        RECT 69.535 159.695 70.285 160.215 ;
        RECT 70.455 159.525 71.205 160.045 ;
        RECT 64.015 158.435 69.360 158.870 ;
        RECT 69.535 158.435 71.205 159.525 ;
        RECT 71.840 159.445 72.190 160.095 ;
        RECT 72.360 159.275 72.590 160.265 ;
        RECT 71.925 159.105 72.590 159.275 ;
        RECT 71.925 158.605 72.095 159.105 ;
        RECT 72.265 158.435 72.595 158.935 ;
        RECT 72.765 158.605 72.950 160.725 ;
        RECT 73.205 160.525 73.455 160.985 ;
        RECT 73.625 160.535 73.960 160.705 ;
        RECT 74.155 160.535 74.830 160.705 ;
        RECT 73.625 160.395 73.795 160.535 ;
        RECT 73.120 159.405 73.400 160.355 ;
        RECT 73.570 160.265 73.795 160.395 ;
        RECT 73.570 159.160 73.740 160.265 ;
        RECT 73.965 160.115 74.490 160.335 ;
        RECT 73.910 159.350 74.150 159.945 ;
        RECT 74.320 159.415 74.490 160.115 ;
        RECT 74.660 159.755 74.830 160.535 ;
        RECT 75.150 160.485 75.520 160.985 ;
        RECT 75.700 160.535 76.105 160.705 ;
        RECT 76.275 160.535 77.060 160.705 ;
        RECT 75.700 160.305 75.870 160.535 ;
        RECT 75.040 160.005 75.870 160.305 ;
        RECT 76.255 160.035 76.720 160.365 ;
        RECT 75.040 159.975 75.240 160.005 ;
        RECT 75.360 159.755 75.530 159.825 ;
        RECT 74.660 159.585 75.530 159.755 ;
        RECT 75.020 159.495 75.530 159.585 ;
        RECT 73.570 159.030 73.875 159.160 ;
        RECT 74.320 159.050 74.850 159.415 ;
        RECT 73.190 158.435 73.455 158.895 ;
        RECT 73.625 158.605 73.875 159.030 ;
        RECT 75.020 158.880 75.190 159.495 ;
        RECT 74.085 158.710 75.190 158.880 ;
        RECT 75.360 158.435 75.530 159.235 ;
        RECT 75.700 158.935 75.870 160.005 ;
        RECT 76.040 159.105 76.230 159.825 ;
        RECT 76.400 159.075 76.720 160.035 ;
        RECT 76.890 160.075 77.060 160.535 ;
        RECT 77.335 160.455 77.545 160.985 ;
        RECT 77.805 160.245 78.135 160.770 ;
        RECT 78.305 160.375 78.475 160.985 ;
        RECT 78.645 160.330 78.975 160.765 ;
        RECT 79.195 160.440 84.540 160.985 ;
        RECT 78.645 160.245 79.025 160.330 ;
        RECT 77.935 160.075 78.135 160.245 ;
        RECT 78.800 160.205 79.025 160.245 ;
        RECT 76.890 159.745 77.765 160.075 ;
        RECT 77.935 159.745 78.685 160.075 ;
        RECT 75.700 158.605 75.950 158.935 ;
        RECT 76.890 158.905 77.060 159.745 ;
        RECT 77.935 159.540 78.125 159.745 ;
        RECT 78.855 159.625 79.025 160.205 ;
        RECT 78.810 159.575 79.025 159.625 ;
        RECT 80.780 159.610 81.120 160.440 ;
        RECT 84.715 160.215 88.225 160.985 ;
        RECT 89.315 160.235 90.525 160.985 ;
        RECT 77.230 159.165 78.125 159.540 ;
        RECT 78.635 159.495 79.025 159.575 ;
        RECT 76.175 158.735 77.060 158.905 ;
        RECT 77.240 158.435 77.555 158.935 ;
        RECT 77.785 158.605 78.125 159.165 ;
        RECT 78.295 158.435 78.465 159.445 ;
        RECT 78.635 158.650 78.965 159.495 ;
        RECT 82.600 158.870 82.950 160.120 ;
        RECT 84.715 159.695 86.365 160.215 ;
        RECT 86.535 159.525 88.225 160.045 ;
        RECT 79.195 158.435 84.540 158.870 ;
        RECT 84.715 158.435 88.225 159.525 ;
        RECT 89.315 159.525 89.835 160.065 ;
        RECT 90.005 159.695 90.525 160.235 ;
        RECT 89.315 158.435 90.525 159.525 ;
        RECT 100.140 159.370 100.810 161.630 ;
        RECT 101.480 161.060 105.520 161.230 ;
        RECT 101.140 160.000 101.310 161.000 ;
        RECT 105.690 160.000 105.860 161.000 ;
        RECT 101.480 159.770 105.520 159.940 ;
        RECT 106.200 159.370 106.370 161.630 ;
        RECT 100.140 159.200 106.370 159.370 ;
        RECT 11.950 158.265 90.610 158.435 ;
        RECT 12.035 157.175 13.245 158.265 ;
        RECT 13.415 157.830 18.760 158.265 ;
        RECT 18.935 157.830 24.280 158.265 ;
        RECT 12.035 156.465 12.555 157.005 ;
        RECT 12.725 156.635 13.245 157.175 ;
        RECT 12.035 155.715 13.245 156.465 ;
        RECT 15.000 156.260 15.340 157.090 ;
        RECT 16.820 156.580 17.170 157.830 ;
        RECT 20.520 156.260 20.860 157.090 ;
        RECT 22.340 156.580 22.690 157.830 ;
        RECT 24.915 157.100 25.205 158.265 ;
        RECT 25.375 157.125 25.635 158.265 ;
        RECT 25.805 157.115 26.135 158.095 ;
        RECT 26.305 157.125 26.585 158.265 ;
        RECT 26.755 157.175 30.265 158.265 ;
        RECT 30.435 157.175 31.645 158.265 ;
        RECT 25.395 156.705 25.730 156.955 ;
        RECT 25.900 156.515 26.070 157.115 ;
        RECT 26.240 156.685 26.575 156.955 ;
        RECT 13.415 155.715 18.760 156.260 ;
        RECT 18.935 155.715 24.280 156.260 ;
        RECT 24.915 155.715 25.205 156.440 ;
        RECT 25.375 155.885 26.070 156.515 ;
        RECT 26.275 155.715 26.585 156.515 ;
        RECT 26.755 156.485 28.405 157.005 ;
        RECT 28.575 156.655 30.265 157.175 ;
        RECT 26.755 155.715 30.265 156.485 ;
        RECT 30.435 156.465 30.955 157.005 ;
        RECT 31.125 156.635 31.645 157.175 ;
        RECT 31.815 157.545 32.275 158.095 ;
        RECT 32.465 157.545 32.795 158.265 ;
        RECT 30.435 155.715 31.645 156.465 ;
        RECT 31.815 156.175 32.065 157.545 ;
        RECT 32.995 157.375 33.295 157.925 ;
        RECT 33.465 157.595 33.745 158.265 ;
        RECT 32.355 157.205 33.295 157.375 ;
        RECT 32.355 156.955 32.525 157.205 ;
        RECT 33.665 156.955 33.930 157.315 ;
        RECT 34.115 157.175 37.625 158.265 ;
        RECT 37.795 157.175 39.005 158.265 ;
        RECT 32.235 156.625 32.525 156.955 ;
        RECT 32.695 156.705 33.035 156.955 ;
        RECT 33.255 156.705 33.930 156.955 ;
        RECT 32.355 156.535 32.525 156.625 ;
        RECT 32.355 156.345 33.745 156.535 ;
        RECT 31.815 155.885 32.375 156.175 ;
        RECT 32.545 155.715 32.795 156.175 ;
        RECT 33.415 155.985 33.745 156.345 ;
        RECT 34.115 156.485 35.765 157.005 ;
        RECT 35.935 156.655 37.625 157.175 ;
        RECT 34.115 155.715 37.625 156.485 ;
        RECT 37.795 156.465 38.315 157.005 ;
        RECT 38.485 156.635 39.005 157.175 ;
        RECT 39.175 157.125 39.435 158.095 ;
        RECT 39.630 157.855 39.960 158.265 ;
        RECT 40.160 157.675 40.330 158.095 ;
        RECT 40.545 157.855 41.215 158.265 ;
        RECT 41.450 157.675 41.620 158.095 ;
        RECT 41.925 157.825 42.255 158.265 ;
        RECT 39.605 157.505 41.620 157.675 ;
        RECT 42.425 157.645 42.600 158.095 ;
        RECT 37.795 155.715 39.005 156.465 ;
        RECT 39.175 156.435 39.345 157.125 ;
        RECT 39.605 156.955 39.775 157.505 ;
        RECT 39.515 156.625 39.775 156.955 ;
        RECT 39.175 155.970 39.515 156.435 ;
        RECT 39.945 156.295 40.285 157.325 ;
        RECT 40.475 156.225 40.745 157.325 ;
        RECT 39.180 155.925 39.515 155.970 ;
        RECT 39.685 155.715 40.015 156.095 ;
        RECT 40.475 156.055 40.785 156.225 ;
        RECT 40.475 156.050 40.745 156.055 ;
        RECT 40.970 156.050 41.250 157.325 ;
        RECT 41.450 156.215 41.620 157.505 ;
        RECT 41.970 157.475 42.600 157.645 ;
        RECT 41.970 156.955 42.140 157.475 ;
        RECT 41.790 156.625 42.140 156.955 ;
        RECT 42.320 156.625 42.685 157.305 ;
        RECT 42.855 157.175 44.065 158.265 ;
        RECT 44.320 157.645 44.495 158.095 ;
        RECT 44.665 157.825 44.995 158.265 ;
        RECT 45.300 157.675 45.470 158.095 ;
        RECT 45.705 157.855 46.375 158.265 ;
        RECT 46.590 157.675 46.760 158.095 ;
        RECT 46.960 157.855 47.290 158.265 ;
        RECT 44.320 157.475 44.950 157.645 ;
        RECT 41.970 156.455 42.140 156.625 ;
        RECT 42.855 156.465 43.375 157.005 ;
        RECT 43.545 156.635 44.065 157.175 ;
        RECT 44.235 156.625 44.600 157.305 ;
        RECT 44.780 156.955 44.950 157.475 ;
        RECT 45.300 157.505 47.315 157.675 ;
        RECT 44.780 156.625 45.130 156.955 ;
        RECT 41.970 156.285 42.600 156.455 ;
        RECT 41.450 155.885 41.680 156.215 ;
        RECT 41.925 155.715 42.255 156.095 ;
        RECT 42.425 155.885 42.600 156.285 ;
        RECT 42.855 155.715 44.065 156.465 ;
        RECT 44.780 156.455 44.950 156.625 ;
        RECT 44.320 156.285 44.950 156.455 ;
        RECT 44.320 155.885 44.495 156.285 ;
        RECT 45.300 156.215 45.470 157.505 ;
        RECT 44.665 155.715 44.995 156.095 ;
        RECT 45.240 155.885 45.470 156.215 ;
        RECT 45.670 156.050 45.950 157.325 ;
        RECT 46.175 156.225 46.445 157.325 ;
        RECT 46.635 156.295 46.975 157.325 ;
        RECT 47.145 156.955 47.315 157.505 ;
        RECT 47.485 157.125 47.745 158.095 ;
        RECT 47.915 157.175 50.505 158.265 ;
        RECT 47.145 156.625 47.405 156.955 ;
        RECT 47.575 156.435 47.745 157.125 ;
        RECT 46.135 156.055 46.445 156.225 ;
        RECT 46.175 156.050 46.445 156.055 ;
        RECT 46.905 155.715 47.235 156.095 ;
        RECT 47.405 155.970 47.745 156.435 ;
        RECT 47.915 156.485 49.125 157.005 ;
        RECT 49.295 156.655 50.505 157.175 ;
        RECT 50.675 157.100 50.965 158.265 ;
        RECT 51.135 157.175 52.805 158.265 ;
        RECT 51.135 156.485 51.885 157.005 ;
        RECT 52.055 156.655 52.805 157.175 ;
        RECT 52.975 157.425 53.235 158.095 ;
        RECT 53.405 157.865 53.735 158.265 ;
        RECT 54.605 157.865 55.005 158.265 ;
        RECT 55.295 157.685 55.625 157.920 ;
        RECT 53.545 157.515 55.625 157.685 ;
        RECT 47.405 155.925 47.740 155.970 ;
        RECT 47.915 155.715 50.505 156.485 ;
        RECT 50.675 155.715 50.965 156.440 ;
        RECT 51.135 155.715 52.805 156.485 ;
        RECT 52.975 156.455 53.150 157.425 ;
        RECT 53.545 157.245 53.715 157.515 ;
        RECT 53.320 157.075 53.715 157.245 ;
        RECT 53.885 157.125 54.900 157.345 ;
        RECT 53.320 156.625 53.490 157.075 ;
        RECT 54.625 156.985 54.900 157.125 ;
        RECT 55.070 157.125 55.625 157.515 ;
        RECT 53.660 156.705 54.110 156.905 ;
        RECT 54.280 156.535 54.455 156.730 ;
        RECT 52.975 155.885 53.315 156.455 ;
        RECT 53.510 155.715 53.680 156.380 ;
        RECT 53.960 156.365 54.455 156.535 ;
        RECT 53.960 156.225 54.180 156.365 ;
        RECT 53.955 156.055 54.180 156.225 ;
        RECT 54.625 156.195 54.795 156.985 ;
        RECT 55.070 156.875 55.240 157.125 ;
        RECT 55.795 156.955 55.970 158.055 ;
        RECT 56.140 157.445 56.485 158.265 ;
        RECT 55.045 156.705 55.240 156.875 ;
        RECT 55.410 156.705 55.970 156.955 ;
        RECT 56.140 156.705 56.485 157.275 ;
        RECT 56.655 157.125 56.930 158.095 ;
        RECT 57.140 157.465 57.420 158.265 ;
        RECT 57.590 157.925 59.640 158.045 ;
        RECT 57.590 157.755 59.645 157.925 ;
        RECT 57.590 157.415 59.220 157.585 ;
        RECT 57.590 157.295 57.760 157.415 ;
        RECT 57.100 157.125 57.760 157.295 ;
        RECT 55.045 156.320 55.215 156.705 ;
        RECT 53.960 156.010 54.180 156.055 ;
        RECT 54.350 156.025 54.795 156.195 ;
        RECT 54.965 155.950 55.215 156.320 ;
        RECT 55.385 156.355 56.485 156.535 ;
        RECT 55.385 155.950 55.635 156.355 ;
        RECT 55.805 155.715 55.975 156.185 ;
        RECT 56.145 155.950 56.485 156.355 ;
        RECT 56.655 156.390 56.825 157.125 ;
        RECT 57.100 156.955 57.270 157.125 ;
        RECT 56.995 156.625 57.270 156.955 ;
        RECT 57.440 156.625 57.820 156.955 ;
        RECT 57.990 156.625 58.730 157.245 ;
        RECT 58.900 157.125 59.220 157.415 ;
        RECT 59.415 156.955 59.655 157.550 ;
        RECT 59.825 157.190 60.165 158.265 ;
        RECT 60.340 157.315 60.605 158.085 ;
        RECT 60.775 157.545 61.105 158.265 ;
        RECT 61.295 157.725 61.555 158.085 ;
        RECT 61.725 157.895 62.055 158.265 ;
        RECT 62.225 157.725 62.485 158.085 ;
        RECT 61.295 157.495 62.485 157.725 ;
        RECT 63.055 157.315 63.345 158.085 ;
        RECT 63.575 157.755 63.875 158.265 ;
        RECT 64.045 157.755 64.425 157.925 ;
        RECT 65.005 157.755 65.635 158.265 ;
        RECT 64.045 157.585 64.215 157.755 ;
        RECT 65.805 157.585 66.135 158.095 ;
        RECT 66.305 157.755 66.605 158.265 ;
        RECT 66.795 157.755 67.095 158.265 ;
        RECT 67.265 157.755 67.645 157.925 ;
        RECT 68.225 157.755 68.855 158.265 ;
        RECT 67.265 157.585 67.435 157.755 ;
        RECT 69.025 157.585 69.355 158.095 ;
        RECT 69.525 157.755 69.825 158.265 ;
        RECT 59.000 156.625 59.655 156.955 ;
        RECT 57.100 156.455 57.270 156.625 ;
        RECT 56.655 156.045 56.930 156.390 ;
        RECT 57.100 156.285 58.685 156.455 ;
        RECT 57.120 155.715 57.500 156.115 ;
        RECT 57.670 155.935 57.840 156.285 ;
        RECT 58.010 155.715 58.340 156.115 ;
        RECT 58.515 155.935 58.685 156.285 ;
        RECT 58.885 155.715 59.215 156.215 ;
        RECT 59.410 155.935 59.655 156.625 ;
        RECT 59.825 156.385 60.165 156.955 ;
        RECT 59.825 155.715 60.165 156.215 ;
        RECT 60.340 155.895 60.675 157.315 ;
        RECT 60.850 157.135 63.345 157.315 ;
        RECT 63.555 157.385 64.215 157.585 ;
        RECT 64.385 157.415 66.605 157.585 ;
        RECT 60.850 156.445 61.075 157.135 ;
        RECT 61.275 156.625 61.555 156.955 ;
        RECT 61.735 156.625 62.310 156.955 ;
        RECT 62.490 156.625 62.925 156.955 ;
        RECT 63.105 156.625 63.375 156.955 ;
        RECT 63.555 156.455 63.725 157.385 ;
        RECT 64.385 157.215 64.555 157.415 ;
        RECT 63.895 157.045 64.555 157.215 ;
        RECT 64.725 157.075 66.265 157.245 ;
        RECT 63.895 156.625 64.065 157.045 ;
        RECT 64.725 156.875 64.895 157.075 ;
        RECT 64.295 156.705 64.895 156.875 ;
        RECT 65.065 156.705 65.760 156.905 ;
        RECT 66.020 156.625 66.265 157.075 ;
        RECT 64.385 156.455 65.295 156.535 ;
        RECT 60.850 156.255 63.335 156.445 ;
        RECT 60.855 155.715 61.600 156.085 ;
        RECT 62.165 155.895 62.420 156.255 ;
        RECT 62.600 155.715 62.930 156.085 ;
        RECT 63.110 155.895 63.335 156.255 ;
        RECT 63.555 155.975 63.875 156.455 ;
        RECT 64.045 156.365 65.295 156.455 ;
        RECT 64.045 156.285 64.555 156.365 ;
        RECT 64.045 155.885 64.275 156.285 ;
        RECT 64.445 155.715 64.795 156.105 ;
        RECT 64.965 155.885 65.295 156.365 ;
        RECT 65.465 155.715 65.635 156.535 ;
        RECT 66.435 156.455 66.605 157.415 ;
        RECT 66.140 155.910 66.605 156.455 ;
        RECT 66.775 157.385 67.435 157.585 ;
        RECT 67.605 157.415 69.825 157.585 ;
        RECT 66.775 156.455 66.945 157.385 ;
        RECT 67.605 157.215 67.775 157.415 ;
        RECT 67.115 157.045 67.775 157.215 ;
        RECT 67.945 157.075 69.485 157.245 ;
        RECT 67.115 156.625 67.285 157.045 ;
        RECT 67.945 156.875 68.115 157.075 ;
        RECT 67.515 156.705 68.115 156.875 ;
        RECT 68.285 156.705 68.980 156.905 ;
        RECT 69.240 156.625 69.485 157.075 ;
        RECT 67.605 156.455 68.515 156.535 ;
        RECT 66.775 155.975 67.095 156.455 ;
        RECT 67.265 156.365 68.515 156.455 ;
        RECT 67.265 156.285 67.775 156.365 ;
        RECT 67.265 155.885 67.495 156.285 ;
        RECT 67.665 155.715 68.015 156.105 ;
        RECT 68.185 155.885 68.515 156.365 ;
        RECT 68.685 155.715 68.855 156.535 ;
        RECT 69.655 156.455 69.825 157.415 ;
        RECT 70.465 157.125 70.795 158.265 ;
        RECT 71.325 157.295 71.655 158.080 ;
        RECT 71.920 157.645 72.095 158.095 ;
        RECT 72.265 157.825 72.595 158.265 ;
        RECT 72.900 157.675 73.070 158.095 ;
        RECT 73.305 157.855 73.975 158.265 ;
        RECT 74.190 157.675 74.360 158.095 ;
        RECT 74.560 157.855 74.890 158.265 ;
        RECT 71.920 157.475 72.550 157.645 ;
        RECT 70.975 157.125 71.655 157.295 ;
        RECT 70.455 156.705 70.805 156.955 ;
        RECT 70.975 156.525 71.145 157.125 ;
        RECT 71.315 156.705 71.665 156.955 ;
        RECT 71.835 156.625 72.200 157.305 ;
        RECT 72.380 156.955 72.550 157.475 ;
        RECT 72.900 157.505 74.915 157.675 ;
        RECT 72.380 156.625 72.730 156.955 ;
        RECT 69.360 155.910 69.825 156.455 ;
        RECT 70.465 155.715 70.735 156.525 ;
        RECT 70.905 155.885 71.235 156.525 ;
        RECT 71.405 155.715 71.645 156.525 ;
        RECT 72.380 156.455 72.550 156.625 ;
        RECT 71.920 156.285 72.550 156.455 ;
        RECT 71.920 155.885 72.095 156.285 ;
        RECT 72.900 156.215 73.070 157.505 ;
        RECT 72.265 155.715 72.595 156.095 ;
        RECT 72.840 155.885 73.070 156.215 ;
        RECT 73.270 156.050 73.550 157.325 ;
        RECT 73.775 156.905 74.045 157.325 ;
        RECT 73.735 156.735 74.045 156.905 ;
        RECT 73.775 156.050 74.045 156.735 ;
        RECT 74.235 156.295 74.575 157.325 ;
        RECT 74.745 156.955 74.915 157.505 ;
        RECT 75.085 157.125 75.345 158.095 ;
        RECT 74.745 156.625 75.005 156.955 ;
        RECT 75.175 156.435 75.345 157.125 ;
        RECT 76.435 157.100 76.725 158.265 ;
        RECT 76.985 157.595 77.155 158.095 ;
        RECT 77.325 157.765 77.655 158.265 ;
        RECT 76.985 157.425 77.650 157.595 ;
        RECT 76.900 156.605 77.250 157.255 ;
        RECT 74.505 155.715 74.835 156.095 ;
        RECT 75.005 155.970 75.345 156.435 ;
        RECT 75.005 155.925 75.340 155.970 ;
        RECT 76.435 155.715 76.725 156.440 ;
        RECT 77.420 156.435 77.650 157.425 ;
        RECT 76.985 156.265 77.650 156.435 ;
        RECT 76.985 155.975 77.155 156.265 ;
        RECT 77.325 155.715 77.655 156.095 ;
        RECT 77.825 155.975 78.010 158.095 ;
        RECT 78.250 157.805 78.515 158.265 ;
        RECT 78.685 157.670 78.935 158.095 ;
        RECT 79.145 157.820 80.250 157.990 ;
        RECT 78.630 157.540 78.935 157.670 ;
        RECT 78.180 156.345 78.460 157.295 ;
        RECT 78.630 156.435 78.800 157.540 ;
        RECT 78.970 156.755 79.210 157.350 ;
        RECT 79.380 157.285 79.910 157.650 ;
        RECT 79.380 156.585 79.550 157.285 ;
        RECT 80.080 157.205 80.250 157.820 ;
        RECT 80.420 157.465 80.590 158.265 ;
        RECT 80.760 157.765 81.010 158.095 ;
        RECT 81.235 157.795 82.120 157.965 ;
        RECT 80.080 157.115 80.590 157.205 ;
        RECT 78.630 156.305 78.855 156.435 ;
        RECT 79.025 156.365 79.550 156.585 ;
        RECT 79.720 156.945 80.590 157.115 ;
        RECT 78.265 155.715 78.515 156.175 ;
        RECT 78.685 156.165 78.855 156.305 ;
        RECT 79.720 156.165 79.890 156.945 ;
        RECT 80.420 156.875 80.590 156.945 ;
        RECT 80.100 156.695 80.300 156.725 ;
        RECT 80.760 156.695 80.930 157.765 ;
        RECT 81.100 156.875 81.290 157.595 ;
        RECT 80.100 156.395 80.930 156.695 ;
        RECT 81.460 156.665 81.780 157.625 ;
        RECT 78.685 155.995 79.020 156.165 ;
        RECT 79.215 155.995 79.890 156.165 ;
        RECT 80.210 155.715 80.580 156.215 ;
        RECT 80.760 156.165 80.930 156.395 ;
        RECT 81.315 156.335 81.780 156.665 ;
        RECT 81.950 156.955 82.120 157.795 ;
        RECT 82.300 157.765 82.615 158.265 ;
        RECT 82.845 157.535 83.185 158.095 ;
        RECT 82.290 157.160 83.185 157.535 ;
        RECT 83.355 157.255 83.525 158.265 ;
        RECT 82.995 156.955 83.185 157.160 ;
        RECT 83.695 157.205 84.025 158.050 ;
        RECT 83.695 157.125 84.085 157.205 ;
        RECT 84.255 157.175 87.765 158.265 ;
        RECT 87.935 157.175 89.145 158.265 ;
        RECT 83.870 157.075 84.085 157.125 ;
        RECT 81.950 156.625 82.825 156.955 ;
        RECT 82.995 156.625 83.745 156.955 ;
        RECT 81.950 156.165 82.120 156.625 ;
        RECT 82.995 156.455 83.195 156.625 ;
        RECT 83.915 156.495 84.085 157.075 ;
        RECT 83.860 156.455 84.085 156.495 ;
        RECT 80.760 155.995 81.165 156.165 ;
        RECT 81.335 155.995 82.120 156.165 ;
        RECT 82.395 155.715 82.605 156.245 ;
        RECT 82.865 155.930 83.195 156.455 ;
        RECT 83.705 156.370 84.085 156.455 ;
        RECT 84.255 156.485 85.905 157.005 ;
        RECT 86.075 156.655 87.765 157.175 ;
        RECT 83.365 155.715 83.535 156.325 ;
        RECT 83.705 155.935 84.035 156.370 ;
        RECT 84.255 155.715 87.765 156.485 ;
        RECT 87.935 156.465 88.455 157.005 ;
        RECT 88.625 156.635 89.145 157.175 ;
        RECT 89.315 157.175 90.525 158.265 ;
        RECT 89.315 156.635 89.835 157.175 ;
        RECT 90.005 156.465 90.525 157.005 ;
        RECT 87.935 155.715 89.145 156.465 ;
        RECT 89.315 155.715 90.525 156.465 ;
        RECT 100.140 155.940 100.810 159.200 ;
        RECT 101.480 158.630 105.520 158.800 ;
        RECT 101.140 156.570 101.310 158.570 ;
        RECT 105.690 156.570 105.860 158.570 ;
        RECT 101.480 156.340 105.520 156.510 ;
        RECT 106.200 155.940 106.370 159.200 ;
        RECT 100.140 155.770 106.370 155.940 ;
        RECT 11.950 155.545 90.610 155.715 ;
        RECT 12.035 154.795 13.245 155.545 ;
        RECT 13.415 155.000 18.760 155.545 ;
        RECT 12.035 154.255 12.555 154.795 ;
        RECT 12.725 154.085 13.245 154.625 ;
        RECT 15.000 154.170 15.340 155.000 ;
        RECT 18.935 154.775 20.605 155.545 ;
        RECT 21.235 155.165 22.125 155.335 ;
        RECT 12.035 152.995 13.245 154.085 ;
        RECT 16.820 153.430 17.170 154.680 ;
        RECT 18.935 154.255 19.685 154.775 ;
        RECT 21.235 154.610 21.785 154.995 ;
        RECT 19.855 154.085 20.605 154.605 ;
        RECT 21.955 154.440 22.125 155.165 ;
        RECT 13.415 152.995 18.760 153.430 ;
        RECT 18.935 152.995 20.605 154.085 ;
        RECT 21.235 154.370 22.125 154.440 ;
        RECT 22.295 154.865 22.515 155.325 ;
        RECT 22.685 155.005 22.935 155.545 ;
        RECT 23.105 154.895 23.365 155.375 ;
        RECT 22.295 154.840 22.545 154.865 ;
        RECT 22.295 154.415 22.625 154.840 ;
        RECT 21.235 154.345 22.130 154.370 ;
        RECT 21.235 154.330 22.140 154.345 ;
        RECT 21.235 154.315 22.145 154.330 ;
        RECT 21.235 154.310 22.155 154.315 ;
        RECT 21.235 154.300 22.160 154.310 ;
        RECT 21.235 154.290 22.165 154.300 ;
        RECT 21.235 154.285 22.175 154.290 ;
        RECT 21.235 154.275 22.185 154.285 ;
        RECT 21.235 154.270 22.195 154.275 ;
        RECT 21.235 153.820 21.495 154.270 ;
        RECT 21.860 154.265 22.195 154.270 ;
        RECT 21.860 154.260 22.210 154.265 ;
        RECT 21.860 154.250 22.225 154.260 ;
        RECT 21.860 154.245 22.250 154.250 ;
        RECT 22.795 154.245 23.025 154.640 ;
        RECT 21.860 154.240 23.025 154.245 ;
        RECT 21.890 154.205 23.025 154.240 ;
        RECT 21.925 154.180 23.025 154.205 ;
        RECT 21.955 154.150 23.025 154.180 ;
        RECT 21.975 154.120 23.025 154.150 ;
        RECT 21.995 154.090 23.025 154.120 ;
        RECT 22.065 154.080 23.025 154.090 ;
        RECT 22.090 154.070 23.025 154.080 ;
        RECT 22.110 154.055 23.025 154.070 ;
        RECT 22.130 154.040 23.025 154.055 ;
        RECT 22.135 154.030 22.920 154.040 ;
        RECT 22.150 153.995 22.920 154.030 ;
        RECT 21.665 153.675 21.995 153.920 ;
        RECT 22.165 153.745 22.920 153.995 ;
        RECT 23.195 153.865 23.365 154.895 ;
        RECT 21.665 153.650 21.850 153.675 ;
        RECT 21.235 153.550 21.850 153.650 ;
        RECT 21.235 152.995 21.840 153.550 ;
        RECT 22.015 153.165 22.495 153.505 ;
        RECT 22.665 152.995 22.920 153.540 ;
        RECT 23.090 153.165 23.365 153.865 ;
        RECT 23.570 154.805 24.185 155.375 ;
        RECT 24.355 155.035 24.570 155.545 ;
        RECT 24.800 155.035 25.080 155.365 ;
        RECT 25.260 155.035 25.500 155.545 ;
        RECT 23.570 153.785 23.885 154.805 ;
        RECT 24.055 154.135 24.225 154.635 ;
        RECT 24.475 154.305 24.740 154.865 ;
        RECT 24.910 154.135 25.080 155.035 ;
        RECT 25.925 154.995 26.095 155.285 ;
        RECT 26.265 155.165 26.595 155.545 ;
        RECT 25.250 154.305 25.605 154.865 ;
        RECT 25.925 154.825 26.590 154.995 ;
        RECT 24.055 153.965 25.480 154.135 ;
        RECT 25.840 154.005 26.190 154.655 ;
        RECT 23.570 153.165 24.105 153.785 ;
        RECT 24.275 152.995 24.605 153.795 ;
        RECT 25.090 153.790 25.480 153.965 ;
        RECT 26.360 153.835 26.590 154.825 ;
        RECT 25.925 153.665 26.590 153.835 ;
        RECT 25.925 153.165 26.095 153.665 ;
        RECT 26.265 152.995 26.595 153.495 ;
        RECT 26.765 153.165 26.950 155.285 ;
        RECT 27.205 155.085 27.455 155.545 ;
        RECT 27.625 155.095 27.960 155.265 ;
        RECT 28.155 155.095 28.830 155.265 ;
        RECT 27.625 154.955 27.795 155.095 ;
        RECT 27.120 153.965 27.400 154.915 ;
        RECT 27.570 154.825 27.795 154.955 ;
        RECT 27.570 153.720 27.740 154.825 ;
        RECT 27.965 154.675 28.490 154.895 ;
        RECT 27.910 153.910 28.150 154.505 ;
        RECT 28.320 153.975 28.490 154.675 ;
        RECT 28.660 154.315 28.830 155.095 ;
        RECT 29.150 155.045 29.520 155.545 ;
        RECT 29.700 155.095 30.105 155.265 ;
        RECT 30.275 155.095 31.060 155.265 ;
        RECT 29.700 154.865 29.870 155.095 ;
        RECT 29.040 154.565 29.870 154.865 ;
        RECT 30.255 154.595 30.720 154.925 ;
        RECT 29.040 154.535 29.240 154.565 ;
        RECT 29.360 154.315 29.530 154.385 ;
        RECT 28.660 154.145 29.530 154.315 ;
        RECT 29.020 154.055 29.530 154.145 ;
        RECT 27.570 153.590 27.875 153.720 ;
        RECT 28.320 153.610 28.850 153.975 ;
        RECT 27.190 152.995 27.455 153.455 ;
        RECT 27.625 153.165 27.875 153.590 ;
        RECT 29.020 153.440 29.190 154.055 ;
        RECT 28.085 153.270 29.190 153.440 ;
        RECT 29.360 152.995 29.530 153.795 ;
        RECT 29.700 153.495 29.870 154.565 ;
        RECT 30.040 153.665 30.230 154.385 ;
        RECT 30.400 153.635 30.720 154.595 ;
        RECT 30.890 154.635 31.060 155.095 ;
        RECT 31.335 155.015 31.545 155.545 ;
        RECT 31.805 154.805 32.135 155.330 ;
        RECT 32.305 154.935 32.475 155.545 ;
        RECT 32.645 154.890 32.975 155.325 ;
        RECT 32.645 154.805 33.025 154.890 ;
        RECT 31.935 154.635 32.135 154.805 ;
        RECT 32.800 154.765 33.025 154.805 ;
        RECT 30.890 154.305 31.765 154.635 ;
        RECT 31.935 154.305 32.685 154.635 ;
        RECT 29.700 153.165 29.950 153.495 ;
        RECT 30.890 153.465 31.060 154.305 ;
        RECT 31.935 154.100 32.125 154.305 ;
        RECT 32.855 154.185 33.025 154.765 ;
        RECT 33.195 154.775 36.705 155.545 ;
        RECT 37.795 154.820 38.085 155.545 ;
        RECT 38.255 155.000 43.600 155.545 ;
        RECT 33.195 154.255 34.845 154.775 ;
        RECT 32.810 154.135 33.025 154.185 ;
        RECT 31.230 153.725 32.125 154.100 ;
        RECT 32.635 154.055 33.025 154.135 ;
        RECT 35.015 154.085 36.705 154.605 ;
        RECT 39.840 154.170 40.180 155.000 ;
        RECT 43.775 154.775 47.285 155.545 ;
        RECT 47.455 154.795 48.665 155.545 ;
        RECT 30.175 153.295 31.060 153.465 ;
        RECT 31.240 152.995 31.555 153.495 ;
        RECT 31.785 153.165 32.125 153.725 ;
        RECT 32.295 152.995 32.465 154.005 ;
        RECT 32.635 153.210 32.965 154.055 ;
        RECT 33.195 152.995 36.705 154.085 ;
        RECT 37.795 152.995 38.085 154.160 ;
        RECT 41.660 153.430 42.010 154.680 ;
        RECT 43.775 154.255 45.425 154.775 ;
        RECT 45.595 154.085 47.285 154.605 ;
        RECT 47.455 154.255 47.975 154.795 ;
        RECT 48.855 154.735 49.095 155.545 ;
        RECT 49.265 154.735 49.595 155.375 ;
        RECT 49.765 154.735 50.035 155.545 ;
        RECT 50.215 154.805 50.655 155.365 ;
        RECT 50.825 154.805 51.275 155.545 ;
        RECT 51.445 154.975 51.615 155.375 ;
        RECT 51.785 155.145 52.205 155.545 ;
        RECT 52.375 154.975 52.605 155.375 ;
        RECT 51.445 154.805 52.605 154.975 ;
        RECT 52.775 154.805 53.265 155.375 ;
        RECT 53.445 155.045 53.775 155.545 ;
        RECT 53.975 154.975 54.145 155.325 ;
        RECT 54.345 155.145 54.675 155.545 ;
        RECT 54.845 154.975 55.015 155.325 ;
        RECT 55.185 155.145 55.565 155.545 ;
        RECT 48.145 154.085 48.665 154.625 ;
        RECT 48.835 154.305 49.185 154.555 ;
        RECT 49.355 154.135 49.525 154.735 ;
        RECT 49.695 154.305 50.045 154.555 ;
        RECT 38.255 152.995 43.600 153.430 ;
        RECT 43.775 152.995 47.285 154.085 ;
        RECT 47.455 152.995 48.665 154.085 ;
        RECT 48.845 153.965 49.525 154.135 ;
        RECT 48.845 153.180 49.175 153.965 ;
        RECT 49.705 152.995 50.035 154.135 ;
        RECT 50.215 153.795 50.525 154.805 ;
        RECT 50.695 154.185 50.865 154.635 ;
        RECT 51.035 154.355 51.425 154.635 ;
        RECT 51.610 154.305 51.855 154.635 ;
        RECT 50.695 154.015 51.485 154.185 ;
        RECT 50.215 153.165 50.655 153.795 ;
        RECT 50.830 152.995 51.145 153.845 ;
        RECT 51.315 153.335 51.485 154.015 ;
        RECT 51.655 153.505 51.855 154.305 ;
        RECT 52.055 153.505 52.305 154.635 ;
        RECT 52.520 154.305 52.925 154.635 ;
        RECT 53.095 154.135 53.265 154.805 ;
        RECT 53.440 154.305 53.790 154.875 ;
        RECT 53.975 154.805 55.585 154.975 ;
        RECT 55.755 154.870 56.025 155.215 ;
        RECT 55.415 154.635 55.585 154.805 ;
        RECT 53.960 154.185 54.670 154.635 ;
        RECT 54.840 154.305 55.245 154.635 ;
        RECT 55.415 154.305 55.685 154.635 ;
        RECT 52.495 153.965 53.265 154.135 ;
        RECT 52.495 153.335 52.745 153.965 ;
        RECT 53.440 153.845 53.760 154.135 ;
        RECT 53.955 154.015 54.670 154.185 ;
        RECT 55.415 154.135 55.585 154.305 ;
        RECT 55.855 154.135 56.025 154.870 ;
        RECT 56.195 154.775 59.705 155.545 ;
        RECT 60.800 154.870 61.075 155.215 ;
        RECT 61.265 155.145 61.645 155.545 ;
        RECT 61.815 154.975 61.985 155.325 ;
        RECT 62.155 155.145 62.485 155.545 ;
        RECT 62.655 154.975 62.910 155.325 ;
        RECT 56.195 154.255 57.845 154.775 ;
        RECT 54.860 153.965 55.585 154.135 ;
        RECT 54.860 153.845 55.030 153.965 ;
        RECT 51.315 153.165 52.745 153.335 ;
        RECT 52.925 152.995 53.255 153.795 ;
        RECT 53.440 153.675 55.030 153.845 ;
        RECT 53.440 153.215 55.095 153.505 ;
        RECT 55.265 152.995 55.545 153.795 ;
        RECT 55.755 153.165 56.025 154.135 ;
        RECT 58.015 154.085 59.705 154.605 ;
        RECT 56.195 152.995 59.705 154.085 ;
        RECT 60.800 154.135 60.970 154.870 ;
        RECT 61.245 154.805 62.910 154.975 ;
        RECT 63.555 154.820 63.845 155.545 ;
        RECT 64.940 154.870 65.215 155.215 ;
        RECT 65.405 155.145 65.785 155.545 ;
        RECT 65.955 154.975 66.125 155.325 ;
        RECT 66.295 155.145 66.625 155.545 ;
        RECT 66.795 154.975 67.050 155.325 ;
        RECT 61.245 154.635 61.415 154.805 ;
        RECT 61.140 154.305 61.415 154.635 ;
        RECT 61.585 154.305 62.410 154.635 ;
        RECT 62.580 154.305 62.925 154.635 ;
        RECT 61.245 154.135 61.415 154.305 ;
        RECT 60.800 153.165 61.075 154.135 ;
        RECT 61.245 153.965 61.905 154.135 ;
        RECT 62.215 154.015 62.410 154.305 ;
        RECT 61.735 153.845 61.905 153.965 ;
        RECT 62.580 153.845 62.905 154.135 ;
        RECT 61.285 152.995 61.565 153.795 ;
        RECT 61.735 153.675 62.905 153.845 ;
        RECT 61.735 153.215 62.925 153.505 ;
        RECT 63.555 152.995 63.845 154.160 ;
        RECT 64.940 154.135 65.110 154.870 ;
        RECT 65.385 154.805 67.050 154.975 ;
        RECT 68.155 154.825 68.495 155.335 ;
        RECT 65.385 154.635 65.555 154.805 ;
        RECT 65.280 154.305 65.555 154.635 ;
        RECT 65.725 154.305 66.550 154.635 ;
        RECT 66.720 154.305 67.065 154.635 ;
        RECT 65.385 154.135 65.555 154.305 ;
        RECT 64.940 153.165 65.215 154.135 ;
        RECT 65.385 153.965 66.045 154.135 ;
        RECT 66.355 154.015 66.550 154.305 ;
        RECT 65.875 153.845 66.045 153.965 ;
        RECT 66.720 153.845 67.045 154.135 ;
        RECT 65.425 152.995 65.705 153.795 ;
        RECT 65.875 153.675 67.045 153.845 ;
        RECT 65.875 153.215 67.065 153.505 ;
        RECT 68.155 153.425 68.415 154.825 ;
        RECT 68.665 154.745 68.935 155.545 ;
        RECT 68.590 154.305 68.920 154.555 ;
        RECT 69.115 154.305 69.395 155.275 ;
        RECT 69.575 154.305 69.875 155.275 ;
        RECT 70.055 154.305 70.405 155.270 ;
        RECT 70.625 155.045 71.120 155.375 ;
        RECT 68.605 154.135 68.920 154.305 ;
        RECT 70.625 154.135 70.795 155.045 ;
        RECT 68.605 153.965 70.795 154.135 ;
        RECT 68.155 153.165 68.495 153.425 ;
        RECT 68.665 152.995 68.995 153.795 ;
        RECT 69.460 153.165 69.710 153.965 ;
        RECT 69.895 152.995 70.225 153.715 ;
        RECT 70.445 153.165 70.695 153.965 ;
        RECT 70.965 153.555 71.205 154.865 ;
        RECT 71.375 154.775 73.045 155.545 ;
        RECT 73.215 154.895 73.475 155.375 ;
        RECT 73.645 155.005 73.895 155.545 ;
        RECT 71.375 154.255 72.125 154.775 ;
        RECT 72.295 154.085 73.045 154.605 ;
        RECT 70.865 152.995 71.200 153.375 ;
        RECT 71.375 152.995 73.045 154.085 ;
        RECT 73.215 153.865 73.385 154.895 ;
        RECT 74.065 154.865 74.285 155.325 ;
        RECT 74.035 154.840 74.285 154.865 ;
        RECT 73.555 154.245 73.785 154.640 ;
        RECT 73.955 154.415 74.285 154.840 ;
        RECT 74.455 155.165 75.345 155.335 ;
        RECT 74.455 154.440 74.625 155.165 ;
        RECT 74.795 154.610 75.345 154.995 ;
        RECT 75.525 154.815 75.825 155.545 ;
        RECT 76.005 154.635 76.235 155.255 ;
        RECT 76.435 154.985 76.660 155.365 ;
        RECT 76.830 155.155 77.160 155.545 ;
        RECT 77.355 155.000 82.700 155.545 ;
        RECT 82.875 155.000 88.220 155.545 ;
        RECT 76.435 154.805 76.765 154.985 ;
        RECT 74.455 154.370 75.345 154.440 ;
        RECT 74.450 154.345 75.345 154.370 ;
        RECT 74.440 154.330 75.345 154.345 ;
        RECT 74.435 154.315 75.345 154.330 ;
        RECT 74.425 154.310 75.345 154.315 ;
        RECT 74.420 154.300 75.345 154.310 ;
        RECT 75.530 154.305 75.825 154.635 ;
        RECT 76.005 154.305 76.420 154.635 ;
        RECT 74.415 154.290 75.345 154.300 ;
        RECT 74.405 154.285 75.345 154.290 ;
        RECT 74.395 154.275 75.345 154.285 ;
        RECT 74.385 154.270 75.345 154.275 ;
        RECT 74.385 154.265 74.720 154.270 ;
        RECT 74.370 154.260 74.720 154.265 ;
        RECT 74.355 154.250 74.720 154.260 ;
        RECT 74.330 154.245 74.720 154.250 ;
        RECT 73.555 154.240 74.720 154.245 ;
        RECT 73.555 154.205 74.690 154.240 ;
        RECT 73.555 154.180 74.655 154.205 ;
        RECT 73.555 154.150 74.625 154.180 ;
        RECT 73.555 154.120 74.605 154.150 ;
        RECT 73.555 154.090 74.585 154.120 ;
        RECT 73.555 154.080 74.515 154.090 ;
        RECT 73.555 154.070 74.490 154.080 ;
        RECT 73.555 154.055 74.470 154.070 ;
        RECT 73.555 154.040 74.450 154.055 ;
        RECT 73.660 154.030 74.445 154.040 ;
        RECT 73.660 153.995 74.430 154.030 ;
        RECT 73.215 153.165 73.490 153.865 ;
        RECT 73.660 153.745 74.415 153.995 ;
        RECT 74.585 153.675 74.915 153.920 ;
        RECT 75.085 153.820 75.345 154.270 ;
        RECT 76.590 154.135 76.765 154.805 ;
        RECT 76.935 154.305 77.175 154.955 ;
        RECT 78.940 154.170 79.280 155.000 ;
        RECT 74.730 153.650 74.915 153.675 ;
        RECT 75.525 153.775 76.420 154.105 ;
        RECT 76.590 153.945 77.175 154.135 ;
        RECT 74.730 153.550 75.345 153.650 ;
        RECT 73.660 152.995 73.915 153.540 ;
        RECT 74.085 153.165 74.565 153.505 ;
        RECT 74.740 152.995 75.345 153.550 ;
        RECT 75.525 153.605 76.730 153.775 ;
        RECT 75.525 153.175 75.855 153.605 ;
        RECT 76.035 152.995 76.230 153.435 ;
        RECT 76.400 153.175 76.730 153.605 ;
        RECT 76.900 153.175 77.175 153.945 ;
        RECT 80.760 153.430 81.110 154.680 ;
        RECT 84.460 154.170 84.800 155.000 ;
        RECT 89.315 154.795 90.525 155.545 ;
        RECT 86.280 153.430 86.630 154.680 ;
        RECT 89.315 154.085 89.835 154.625 ;
        RECT 90.005 154.255 90.525 154.795 ;
        RECT 77.355 152.995 82.700 153.430 ;
        RECT 82.875 152.995 88.220 153.430 ;
        RECT 89.315 152.995 90.525 154.085 ;
        RECT 11.950 152.825 90.610 152.995 ;
        RECT 12.035 151.735 13.245 152.825 ;
        RECT 13.415 151.735 16.925 152.825 ;
        RECT 17.645 152.155 17.815 152.655 ;
        RECT 17.985 152.325 18.315 152.825 ;
        RECT 17.645 151.985 18.310 152.155 ;
        RECT 12.035 151.025 12.555 151.565 ;
        RECT 12.725 151.195 13.245 151.735 ;
        RECT 13.415 151.045 15.065 151.565 ;
        RECT 15.235 151.215 16.925 151.735 ;
        RECT 17.560 151.165 17.910 151.815 ;
        RECT 12.035 150.275 13.245 151.025 ;
        RECT 13.415 150.275 16.925 151.045 ;
        RECT 18.080 150.995 18.310 151.985 ;
        RECT 17.645 150.825 18.310 150.995 ;
        RECT 17.645 150.535 17.815 150.825 ;
        RECT 17.985 150.275 18.315 150.655 ;
        RECT 18.485 150.535 18.670 152.655 ;
        RECT 18.910 152.365 19.175 152.825 ;
        RECT 19.345 152.230 19.595 152.655 ;
        RECT 19.805 152.380 20.910 152.550 ;
        RECT 19.290 152.100 19.595 152.230 ;
        RECT 18.840 150.905 19.120 151.855 ;
        RECT 19.290 150.995 19.460 152.100 ;
        RECT 19.630 151.315 19.870 151.910 ;
        RECT 20.040 151.845 20.570 152.210 ;
        RECT 20.040 151.145 20.210 151.845 ;
        RECT 20.740 151.765 20.910 152.380 ;
        RECT 21.080 152.025 21.250 152.825 ;
        RECT 21.420 152.325 21.670 152.655 ;
        RECT 21.895 152.355 22.780 152.525 ;
        RECT 20.740 151.675 21.250 151.765 ;
        RECT 19.290 150.865 19.515 150.995 ;
        RECT 19.685 150.925 20.210 151.145 ;
        RECT 20.380 151.505 21.250 151.675 ;
        RECT 18.925 150.275 19.175 150.735 ;
        RECT 19.345 150.725 19.515 150.865 ;
        RECT 20.380 150.725 20.550 151.505 ;
        RECT 21.080 151.435 21.250 151.505 ;
        RECT 20.760 151.255 20.960 151.285 ;
        RECT 21.420 151.255 21.590 152.325 ;
        RECT 21.760 151.435 21.950 152.155 ;
        RECT 20.760 150.955 21.590 151.255 ;
        RECT 22.120 151.225 22.440 152.185 ;
        RECT 19.345 150.555 19.680 150.725 ;
        RECT 19.875 150.555 20.550 150.725 ;
        RECT 20.870 150.275 21.240 150.775 ;
        RECT 21.420 150.725 21.590 150.955 ;
        RECT 21.975 150.895 22.440 151.225 ;
        RECT 22.610 151.515 22.780 152.355 ;
        RECT 22.960 152.325 23.275 152.825 ;
        RECT 23.505 152.095 23.845 152.655 ;
        RECT 22.950 151.720 23.845 152.095 ;
        RECT 24.015 151.815 24.185 152.825 ;
        RECT 23.655 151.515 23.845 151.720 ;
        RECT 24.355 151.765 24.685 152.610 ;
        RECT 24.355 151.685 24.745 151.765 ;
        RECT 24.530 151.635 24.745 151.685 ;
        RECT 24.915 151.660 25.205 152.825 ;
        RECT 22.610 151.185 23.485 151.515 ;
        RECT 23.655 151.185 24.405 151.515 ;
        RECT 22.610 150.725 22.780 151.185 ;
        RECT 23.655 151.015 23.855 151.185 ;
        RECT 24.575 151.055 24.745 151.635 ;
        RECT 24.520 151.015 24.745 151.055 ;
        RECT 21.420 150.555 21.825 150.725 ;
        RECT 21.995 150.555 22.780 150.725 ;
        RECT 23.055 150.275 23.265 150.805 ;
        RECT 23.525 150.490 23.855 151.015 ;
        RECT 24.365 150.930 24.745 151.015 ;
        RECT 24.025 150.275 24.195 150.885 ;
        RECT 24.365 150.495 24.695 150.930 ;
        RECT 24.915 150.275 25.205 151.000 ;
        RECT 25.385 150.455 25.645 152.645 ;
        RECT 25.815 152.095 26.155 152.825 ;
        RECT 26.335 151.915 26.605 152.645 ;
        RECT 25.835 151.695 26.605 151.915 ;
        RECT 26.785 151.935 27.015 152.645 ;
        RECT 27.185 152.115 27.515 152.825 ;
        RECT 27.685 151.935 27.945 152.645 ;
        RECT 26.785 151.695 27.945 151.935 ;
        RECT 28.135 151.735 30.725 152.825 ;
        RECT 25.835 151.025 26.125 151.695 ;
        RECT 26.305 151.205 26.770 151.515 ;
        RECT 26.950 151.205 27.475 151.515 ;
        RECT 25.835 150.825 27.065 151.025 ;
        RECT 25.905 150.275 26.575 150.645 ;
        RECT 26.755 150.455 27.065 150.825 ;
        RECT 27.245 150.565 27.475 151.205 ;
        RECT 27.655 151.185 27.955 151.515 ;
        RECT 28.135 151.045 29.345 151.565 ;
        RECT 29.515 151.215 30.725 151.735 ;
        RECT 30.985 151.815 31.155 152.655 ;
        RECT 31.325 152.485 32.495 152.655 ;
        RECT 31.325 151.985 31.655 152.485 ;
        RECT 32.165 152.445 32.495 152.485 ;
        RECT 32.685 152.405 33.040 152.825 ;
        RECT 31.825 152.225 32.055 152.315 ;
        RECT 33.210 152.225 33.460 152.655 ;
        RECT 31.825 151.985 33.460 152.225 ;
        RECT 33.630 152.065 33.960 152.825 ;
        RECT 34.130 151.985 34.385 152.655 ;
        RECT 30.985 151.645 34.045 151.815 ;
        RECT 30.900 151.265 31.250 151.475 ;
        RECT 31.420 151.265 31.865 151.465 ;
        RECT 32.035 151.265 32.510 151.465 ;
        RECT 27.655 150.275 27.945 151.005 ;
        RECT 28.135 150.275 30.725 151.045 ;
        RECT 30.985 150.925 32.050 151.095 ;
        RECT 30.985 150.445 31.155 150.925 ;
        RECT 31.325 150.275 31.655 150.755 ;
        RECT 31.880 150.695 32.050 150.925 ;
        RECT 32.230 150.865 32.510 151.265 ;
        RECT 32.780 151.265 33.110 151.465 ;
        RECT 33.280 151.295 33.655 151.465 ;
        RECT 33.280 151.265 33.645 151.295 ;
        RECT 32.780 150.865 33.065 151.265 ;
        RECT 33.875 151.095 34.045 151.645 ;
        RECT 33.245 150.925 34.045 151.095 ;
        RECT 33.245 150.695 33.415 150.925 ;
        RECT 34.215 150.855 34.385 151.985 ;
        RECT 34.575 151.735 35.785 152.825 ;
        RECT 36.455 152.365 36.670 152.825 ;
        RECT 36.840 152.195 37.170 152.655 ;
        RECT 34.200 150.785 34.385 150.855 ;
        RECT 34.175 150.775 34.385 150.785 ;
        RECT 31.880 150.445 33.415 150.695 ;
        RECT 33.585 150.275 33.915 150.755 ;
        RECT 34.130 150.445 34.385 150.775 ;
        RECT 34.575 151.025 35.095 151.565 ;
        RECT 35.265 151.195 35.785 151.735 ;
        RECT 36.000 152.025 37.170 152.195 ;
        RECT 37.340 152.025 37.590 152.825 ;
        RECT 34.575 150.275 35.785 151.025 ;
        RECT 36.000 150.735 36.370 152.025 ;
        RECT 37.800 151.855 38.080 152.015 ;
        RECT 36.745 151.685 38.080 151.855 ;
        RECT 38.715 151.975 39.095 152.655 ;
        RECT 39.685 151.975 39.855 152.825 ;
        RECT 40.025 152.145 40.355 152.655 ;
        RECT 40.525 152.315 40.695 152.825 ;
        RECT 40.865 152.145 41.265 152.655 ;
        RECT 40.025 151.975 41.265 152.145 ;
        RECT 36.745 151.515 36.915 151.685 ;
        RECT 36.540 151.265 36.915 151.515 ;
        RECT 37.085 151.265 37.560 151.505 ;
        RECT 37.730 151.265 38.080 151.505 ;
        RECT 36.745 151.095 36.915 151.265 ;
        RECT 36.745 150.925 38.080 151.095 ;
        RECT 36.000 150.445 36.750 150.735 ;
        RECT 37.260 150.275 37.590 150.735 ;
        RECT 37.810 150.715 38.080 150.925 ;
        RECT 38.715 151.015 38.885 151.975 ;
        RECT 39.055 151.635 40.360 151.805 ;
        RECT 41.445 151.725 41.765 152.655 ;
        RECT 41.935 151.735 43.145 152.825 ;
        RECT 43.315 152.315 43.615 152.825 ;
        RECT 43.785 152.145 44.115 152.655 ;
        RECT 44.285 152.315 44.915 152.825 ;
        RECT 45.495 152.315 45.875 152.485 ;
        RECT 46.045 152.315 46.345 152.825 ;
        RECT 45.705 152.145 45.875 152.315 ;
        RECT 39.055 151.185 39.300 151.635 ;
        RECT 39.470 151.265 40.020 151.465 ;
        RECT 40.190 151.435 40.360 151.635 ;
        RECT 41.135 151.555 41.765 151.725 ;
        RECT 40.190 151.265 40.565 151.435 ;
        RECT 40.735 151.015 40.965 151.515 ;
        RECT 38.715 150.845 40.965 151.015 ;
        RECT 38.765 150.275 39.095 150.665 ;
        RECT 39.265 150.525 39.435 150.845 ;
        RECT 41.135 150.675 41.305 151.555 ;
        RECT 39.605 150.275 39.935 150.665 ;
        RECT 40.350 150.505 41.305 150.675 ;
        RECT 41.475 150.275 41.765 151.110 ;
        RECT 41.935 151.025 42.455 151.565 ;
        RECT 42.625 151.195 43.145 151.735 ;
        RECT 43.315 151.975 45.535 152.145 ;
        RECT 41.935 150.275 43.145 151.025 ;
        RECT 43.315 151.015 43.485 151.975 ;
        RECT 43.655 151.635 45.195 151.805 ;
        RECT 43.655 151.185 43.900 151.635 ;
        RECT 44.160 151.265 44.855 151.465 ;
        RECT 45.025 151.435 45.195 151.635 ;
        RECT 45.365 151.775 45.535 151.975 ;
        RECT 45.705 151.945 46.365 152.145 ;
        RECT 45.365 151.605 46.025 151.775 ;
        RECT 45.025 151.265 45.625 151.435 ;
        RECT 45.855 151.185 46.025 151.605 ;
        RECT 43.315 150.470 43.780 151.015 ;
        RECT 44.285 150.275 44.455 151.095 ;
        RECT 44.625 151.015 45.535 151.095 ;
        RECT 46.195 151.015 46.365 151.945 ;
        RECT 46.535 151.735 47.745 152.825 ;
        RECT 47.920 152.315 49.575 152.605 ;
        RECT 44.625 150.925 45.875 151.015 ;
        RECT 44.625 150.445 44.955 150.925 ;
        RECT 45.365 150.845 45.875 150.925 ;
        RECT 45.125 150.275 45.475 150.665 ;
        RECT 45.645 150.445 45.875 150.845 ;
        RECT 46.045 150.535 46.365 151.015 ;
        RECT 46.535 151.025 47.055 151.565 ;
        RECT 47.225 151.195 47.745 151.735 ;
        RECT 47.920 151.975 49.510 152.145 ;
        RECT 49.745 152.025 50.025 152.825 ;
        RECT 47.920 151.685 48.240 151.975 ;
        RECT 49.340 151.855 49.510 151.975 ;
        RECT 46.535 150.275 47.745 151.025 ;
        RECT 47.920 150.945 48.270 151.515 ;
        RECT 48.440 151.185 49.150 151.805 ;
        RECT 49.340 151.685 50.065 151.855 ;
        RECT 50.235 151.685 50.505 152.655 ;
        RECT 49.895 151.515 50.065 151.685 ;
        RECT 49.320 151.185 49.725 151.515 ;
        RECT 49.895 151.185 50.165 151.515 ;
        RECT 49.895 151.015 50.065 151.185 ;
        RECT 48.455 150.845 50.065 151.015 ;
        RECT 50.335 150.950 50.505 151.685 ;
        RECT 50.675 151.660 50.965 152.825 ;
        RECT 51.140 151.855 51.435 152.825 ;
        RECT 52.005 152.465 52.335 152.825 ;
        RECT 52.505 152.465 54.485 152.655 ;
        RECT 51.605 152.295 51.825 152.380 ;
        RECT 52.505 152.295 52.685 152.465 ;
        RECT 54.665 152.385 54.935 152.825 ;
        RECT 55.485 152.465 55.815 152.825 ;
        RECT 56.330 152.465 56.660 152.825 ;
        RECT 57.170 152.465 57.505 152.825 ;
        RECT 58.405 152.465 58.735 152.825 ;
        RECT 51.605 152.125 52.685 152.295 ;
        RECT 52.855 152.215 54.520 152.295 ;
        RECT 55.095 152.215 58.730 152.295 ;
        RECT 51.605 152.050 51.825 152.125 ;
        RECT 52.855 152.045 58.730 152.215 ;
        RECT 52.015 151.705 54.680 151.875 ;
        RECT 52.015 151.520 52.460 151.705 ;
        RECT 51.450 151.265 52.460 151.520 ;
        RECT 52.755 151.265 54.230 151.535 ;
        RECT 54.400 151.185 54.680 151.705 ;
        RECT 55.310 151.705 58.050 151.875 ;
        RECT 55.310 151.600 56.025 151.705 ;
        RECT 54.850 151.185 56.025 151.600 ;
        RECT 56.420 151.265 57.490 151.535 ;
        RECT 57.880 151.185 58.050 151.705 ;
        RECT 58.220 151.530 58.730 152.045 ;
        RECT 59.045 151.815 59.215 152.655 ;
        RECT 59.385 152.485 60.555 152.655 ;
        RECT 59.385 151.985 59.715 152.485 ;
        RECT 60.225 152.445 60.555 152.485 ;
        RECT 60.745 152.405 61.100 152.825 ;
        RECT 59.885 152.225 60.115 152.315 ;
        RECT 61.270 152.225 61.520 152.655 ;
        RECT 59.885 151.985 61.520 152.225 ;
        RECT 61.690 152.065 62.020 152.825 ;
        RECT 62.190 151.985 62.445 152.655 ;
        RECT 59.045 151.645 62.105 151.815 ;
        RECT 51.205 151.055 52.845 151.095 ;
        RECT 47.925 150.275 48.255 150.775 ;
        RECT 48.455 150.495 48.625 150.845 ;
        RECT 48.825 150.275 49.155 150.675 ;
        RECT 49.325 150.495 49.495 150.845 ;
        RECT 49.665 150.275 50.045 150.675 ;
        RECT 50.235 150.605 50.505 150.950 ;
        RECT 50.675 150.275 50.965 151.000 ;
        RECT 51.205 150.985 54.180 151.055 ;
        RECT 58.220 151.015 58.400 151.530 ;
        RECT 58.960 151.265 59.310 151.475 ;
        RECT 59.480 151.265 59.925 151.465 ;
        RECT 60.095 151.265 60.570 151.465 ;
        RECT 51.205 150.885 54.885 150.985 ;
        RECT 51.205 150.815 52.290 150.885 ;
        RECT 52.825 150.815 54.885 150.885 ;
        RECT 55.055 150.825 57.220 151.005 ;
        RECT 57.615 150.845 58.400 151.015 ;
        RECT 59.045 150.925 60.110 151.095 ;
        RECT 51.205 150.725 51.405 150.815 ;
        RECT 51.575 150.275 51.905 150.635 ;
        RECT 52.075 150.615 52.290 150.815 ;
        RECT 52.515 150.275 52.685 150.715 ;
        RECT 54.655 150.645 54.885 150.815 ;
        RECT 53.295 150.275 53.625 150.635 ;
        RECT 54.155 150.275 54.485 150.635 ;
        RECT 54.655 150.445 55.970 150.645 ;
        RECT 57.615 150.640 57.785 150.845 ;
        RECT 58.560 150.670 58.730 150.785 ;
        RECT 56.330 150.460 57.785 150.640 ;
        RECT 58.030 150.500 58.730 150.670 ;
        RECT 59.045 150.445 59.215 150.925 ;
        RECT 59.385 150.275 59.715 150.755 ;
        RECT 59.940 150.695 60.110 150.925 ;
        RECT 60.290 150.865 60.570 151.265 ;
        RECT 60.840 151.265 61.170 151.465 ;
        RECT 61.340 151.265 61.705 151.465 ;
        RECT 60.840 150.865 61.125 151.265 ;
        RECT 61.935 151.095 62.105 151.645 ;
        RECT 61.305 150.925 62.105 151.095 ;
        RECT 61.305 150.695 61.475 150.925 ;
        RECT 62.275 150.855 62.445 151.985 ;
        RECT 62.635 151.685 62.895 152.825 ;
        RECT 63.065 151.675 63.395 152.655 ;
        RECT 63.565 151.685 63.845 152.825 ;
        RECT 64.015 152.390 69.360 152.825 ;
        RECT 62.655 151.265 62.990 151.515 ;
        RECT 63.160 151.075 63.330 151.675 ;
        RECT 63.500 151.245 63.835 151.515 ;
        RECT 62.260 150.785 62.445 150.855 ;
        RECT 62.235 150.775 62.445 150.785 ;
        RECT 59.940 150.445 61.475 150.695 ;
        RECT 61.645 150.275 61.975 150.755 ;
        RECT 62.190 150.445 62.445 150.775 ;
        RECT 62.635 150.445 63.330 151.075 ;
        RECT 63.535 150.275 63.845 151.075 ;
        RECT 65.600 150.820 65.940 151.650 ;
        RECT 67.420 151.140 67.770 152.390 ;
        RECT 69.535 151.735 72.125 152.825 ;
        RECT 69.535 151.045 70.745 151.565 ;
        RECT 70.915 151.215 72.125 151.735 ;
        RECT 72.305 151.685 72.635 152.825 ;
        RECT 73.165 151.855 73.495 152.640 ;
        RECT 72.815 151.685 73.495 151.855 ;
        RECT 73.685 151.855 74.015 152.640 ;
        RECT 73.685 151.685 74.365 151.855 ;
        RECT 74.545 151.685 74.875 152.825 ;
        RECT 75.055 151.735 76.265 152.825 ;
        RECT 72.295 151.265 72.645 151.515 ;
        RECT 72.815 151.085 72.985 151.685 ;
        RECT 73.155 151.265 73.505 151.515 ;
        RECT 73.675 151.265 74.025 151.515 ;
        RECT 74.195 151.085 74.365 151.685 ;
        RECT 74.535 151.265 74.885 151.515 ;
        RECT 64.015 150.275 69.360 150.820 ;
        RECT 69.535 150.275 72.125 151.045 ;
        RECT 72.305 150.275 72.575 151.085 ;
        RECT 72.745 150.445 73.075 151.085 ;
        RECT 73.245 150.275 73.485 151.085 ;
        RECT 73.695 150.275 73.935 151.085 ;
        RECT 74.105 150.445 74.435 151.085 ;
        RECT 74.605 150.275 74.875 151.085 ;
        RECT 75.055 151.025 75.575 151.565 ;
        RECT 75.745 151.195 76.265 151.735 ;
        RECT 76.435 151.660 76.725 152.825 ;
        RECT 76.895 152.390 82.240 152.825 ;
        RECT 82.415 152.390 87.760 152.825 ;
        RECT 75.055 150.275 76.265 151.025 ;
        RECT 76.435 150.275 76.725 151.000 ;
        RECT 78.480 150.820 78.820 151.650 ;
        RECT 80.300 151.140 80.650 152.390 ;
        RECT 84.000 150.820 84.340 151.650 ;
        RECT 85.820 151.140 86.170 152.390 ;
        RECT 87.935 151.735 89.145 152.825 ;
        RECT 87.935 151.025 88.455 151.565 ;
        RECT 88.625 151.195 89.145 151.735 ;
        RECT 89.315 151.735 90.525 152.825 ;
        RECT 100.140 152.510 100.810 155.770 ;
        RECT 101.480 155.200 105.520 155.370 ;
        RECT 101.140 153.140 101.310 155.140 ;
        RECT 105.690 153.140 105.860 155.140 ;
        RECT 101.480 152.910 105.520 153.080 ;
        RECT 106.200 152.510 106.370 155.770 ;
        RECT 100.140 152.500 106.370 152.510 ;
        RECT 107.960 161.770 117.790 161.810 ;
        RECT 120.510 161.790 126.250 161.800 ;
        RECT 107.960 161.640 118.590 161.770 ;
        RECT 107.960 159.380 108.130 161.640 ;
        RECT 108.855 161.070 116.895 161.240 ;
        RECT 108.470 160.010 108.640 161.010 ;
        RECT 117.110 160.010 117.280 161.010 ;
        RECT 108.855 159.780 116.895 159.950 ;
        RECT 117.620 159.380 118.590 161.640 ;
        RECT 107.960 159.210 118.590 159.380 ;
        RECT 107.960 155.950 108.130 159.210 ;
        RECT 108.855 158.640 116.895 158.810 ;
        RECT 108.470 156.580 108.640 158.580 ;
        RECT 117.110 156.580 117.280 158.580 ;
        RECT 108.855 156.350 116.895 156.520 ;
        RECT 117.620 155.950 118.590 159.210 ;
        RECT 107.960 155.780 118.590 155.950 ;
        RECT 107.960 152.520 108.130 155.780 ;
        RECT 108.855 155.210 116.895 155.380 ;
        RECT 108.470 153.150 108.640 155.150 ;
        RECT 117.110 153.150 117.280 155.150 ;
        RECT 108.855 152.920 116.895 153.090 ;
        RECT 117.620 152.520 118.590 155.780 ;
        RECT 100.140 152.400 106.380 152.500 ;
        RECT 100.130 151.840 106.380 152.400 ;
        RECT 100.130 151.820 105.300 151.840 ;
        RECT 100.130 151.750 104.120 151.820 ;
        RECT 89.315 151.195 89.835 151.735 ;
        RECT 90.005 151.025 90.525 151.565 ;
        RECT 76.895 150.275 82.240 150.820 ;
        RECT 82.415 150.275 87.760 150.820 ;
        RECT 87.935 150.275 89.145 151.025 ;
        RECT 89.315 150.275 90.525 151.025 ;
        RECT 100.130 150.480 102.050 151.750 ;
        RECT 103.560 151.740 104.120 151.750 ;
        RECT 103.790 150.650 104.120 151.740 ;
        RECT 104.490 151.270 105.530 151.440 ;
        RECT 104.490 150.830 105.530 151.000 ;
        RECT 105.700 150.970 105.870 151.300 ;
        RECT 103.950 150.430 104.120 150.650 ;
        RECT 106.210 150.430 106.380 151.840 ;
        RECT 11.950 150.105 90.610 150.275 ;
        RECT 103.950 150.260 106.380 150.430 ;
        RECT 107.960 152.350 118.590 152.520 ;
        RECT 120.020 161.630 126.250 161.790 ;
        RECT 120.020 159.370 120.690 161.630 ;
        RECT 121.360 161.060 125.400 161.230 ;
        RECT 121.020 160.000 121.190 161.000 ;
        RECT 125.570 160.000 125.740 161.000 ;
        RECT 121.360 159.770 125.400 159.940 ;
        RECT 126.080 159.370 126.250 161.630 ;
        RECT 120.020 159.200 126.250 159.370 ;
        RECT 120.020 155.940 120.690 159.200 ;
        RECT 121.360 158.630 125.400 158.800 ;
        RECT 121.020 156.570 121.190 158.570 ;
        RECT 125.570 156.570 125.740 158.570 ;
        RECT 121.360 156.340 125.400 156.510 ;
        RECT 126.080 155.940 126.250 159.200 ;
        RECT 120.020 155.770 126.250 155.940 ;
        RECT 120.020 152.510 120.690 155.770 ;
        RECT 121.360 155.200 125.400 155.370 ;
        RECT 121.020 153.140 121.190 155.140 ;
        RECT 125.570 153.140 125.740 155.140 ;
        RECT 121.360 152.910 125.400 153.080 ;
        RECT 126.080 152.510 126.250 155.770 ;
        RECT 120.020 152.500 126.250 152.510 ;
        RECT 127.840 161.770 137.670 161.810 ;
        RECT 127.840 161.640 138.470 161.770 ;
        RECT 140.590 161.740 146.330 161.750 ;
        RECT 127.840 159.380 128.010 161.640 ;
        RECT 128.735 161.070 136.775 161.240 ;
        RECT 128.350 160.010 128.520 161.010 ;
        RECT 136.990 160.010 137.160 161.010 ;
        RECT 128.735 159.780 136.775 159.950 ;
        RECT 137.500 159.380 138.470 161.640 ;
        RECT 127.840 159.210 138.470 159.380 ;
        RECT 127.840 155.950 128.010 159.210 ;
        RECT 128.735 158.640 136.775 158.810 ;
        RECT 128.350 156.580 128.520 158.580 ;
        RECT 136.990 156.580 137.160 158.580 ;
        RECT 128.735 156.350 136.775 156.520 ;
        RECT 137.500 155.950 138.470 159.210 ;
        RECT 127.840 155.780 138.470 155.950 ;
        RECT 127.840 152.520 128.010 155.780 ;
        RECT 128.735 155.210 136.775 155.380 ;
        RECT 128.350 153.150 128.520 155.150 ;
        RECT 136.990 153.150 137.160 155.150 ;
        RECT 128.735 152.920 136.775 153.090 ;
        RECT 137.500 152.520 138.470 155.780 ;
        RECT 120.020 152.400 126.260 152.500 ;
        RECT 12.035 149.355 13.245 150.105 ;
        RECT 13.415 149.560 18.760 150.105 ;
        RECT 12.035 148.815 12.555 149.355 ;
        RECT 12.725 148.645 13.245 149.185 ;
        RECT 15.000 148.730 15.340 149.560 ;
        RECT 18.935 149.455 19.195 149.935 ;
        RECT 19.365 149.645 19.695 150.105 ;
        RECT 19.885 149.465 20.085 149.885 ;
        RECT 12.035 147.555 13.245 148.645 ;
        RECT 16.820 147.990 17.170 149.240 ;
        RECT 18.935 148.425 19.105 149.455 ;
        RECT 19.275 148.765 19.505 149.195 ;
        RECT 19.675 148.945 20.085 149.465 ;
        RECT 20.255 149.620 21.045 149.885 ;
        RECT 20.255 148.765 20.510 149.620 ;
        RECT 21.225 149.285 21.555 149.705 ;
        RECT 21.725 149.285 21.985 150.105 ;
        RECT 22.615 149.455 22.875 149.935 ;
        RECT 23.045 149.565 23.295 150.105 ;
        RECT 21.225 149.195 21.475 149.285 ;
        RECT 20.680 148.945 21.475 149.195 ;
        RECT 19.275 148.595 21.065 148.765 ;
        RECT 13.415 147.555 18.760 147.990 ;
        RECT 18.935 147.725 19.210 148.425 ;
        RECT 19.380 148.300 20.095 148.595 ;
        RECT 20.315 148.235 20.645 148.425 ;
        RECT 19.420 147.555 19.635 148.100 ;
        RECT 19.805 147.725 20.280 148.065 ;
        RECT 20.450 148.060 20.645 148.235 ;
        RECT 20.815 148.230 21.065 148.595 ;
        RECT 20.450 147.555 21.065 148.060 ;
        RECT 21.305 147.725 21.475 148.945 ;
        RECT 21.645 148.235 21.985 149.115 ;
        RECT 22.615 148.425 22.785 149.455 ;
        RECT 23.465 149.400 23.685 149.885 ;
        RECT 22.955 148.805 23.185 149.200 ;
        RECT 23.355 148.975 23.685 149.400 ;
        RECT 23.855 149.725 24.745 149.895 ;
        RECT 23.855 149.000 24.025 149.725 ;
        RECT 24.915 149.560 30.260 150.105 ;
        RECT 24.195 149.170 24.745 149.555 ;
        RECT 23.855 148.930 24.745 149.000 ;
        RECT 23.850 148.905 24.745 148.930 ;
        RECT 23.840 148.890 24.745 148.905 ;
        RECT 23.835 148.875 24.745 148.890 ;
        RECT 23.825 148.870 24.745 148.875 ;
        RECT 23.820 148.860 24.745 148.870 ;
        RECT 23.815 148.850 24.745 148.860 ;
        RECT 23.805 148.845 24.745 148.850 ;
        RECT 23.795 148.835 24.745 148.845 ;
        RECT 23.785 148.830 24.745 148.835 ;
        RECT 23.785 148.825 24.120 148.830 ;
        RECT 23.770 148.820 24.120 148.825 ;
        RECT 23.755 148.810 24.120 148.820 ;
        RECT 23.730 148.805 24.120 148.810 ;
        RECT 22.955 148.800 24.120 148.805 ;
        RECT 22.955 148.765 24.090 148.800 ;
        RECT 22.955 148.740 24.055 148.765 ;
        RECT 22.955 148.710 24.025 148.740 ;
        RECT 22.955 148.680 24.005 148.710 ;
        RECT 22.955 148.650 23.985 148.680 ;
        RECT 22.955 148.640 23.915 148.650 ;
        RECT 22.955 148.630 23.890 148.640 ;
        RECT 22.955 148.615 23.870 148.630 ;
        RECT 22.955 148.600 23.850 148.615 ;
        RECT 23.060 148.590 23.845 148.600 ;
        RECT 23.060 148.555 23.830 148.590 ;
        RECT 21.725 147.555 21.985 148.065 ;
        RECT 22.615 147.725 22.890 148.425 ;
        RECT 23.060 148.305 23.815 148.555 ;
        RECT 23.985 148.235 24.315 148.480 ;
        RECT 24.485 148.380 24.745 148.830 ;
        RECT 26.500 148.730 26.840 149.560 ;
        RECT 30.435 149.455 30.775 149.935 ;
        RECT 31.140 149.625 31.470 149.935 ;
        RECT 31.640 149.625 31.890 150.105 ;
        RECT 31.300 149.455 31.470 149.625 ;
        RECT 32.060 149.455 32.390 149.935 ;
        RECT 32.560 149.625 32.810 150.105 ;
        RECT 32.980 149.455 33.310 149.935 ;
        RECT 30.435 149.285 31.130 149.455 ;
        RECT 31.300 149.285 33.310 149.455 ;
        RECT 33.655 149.335 37.165 150.105 ;
        RECT 37.795 149.380 38.085 150.105 ;
        RECT 38.305 149.450 38.635 149.885 ;
        RECT 38.805 149.495 38.975 150.105 ;
        RECT 38.255 149.365 38.635 149.450 ;
        RECT 39.145 149.365 39.475 149.890 ;
        RECT 39.735 149.575 39.945 150.105 ;
        RECT 40.220 149.655 41.005 149.825 ;
        RECT 41.175 149.655 41.580 149.825 ;
        RECT 24.130 148.210 24.315 148.235 ;
        RECT 24.130 148.110 24.745 148.210 ;
        RECT 23.060 147.555 23.315 148.100 ;
        RECT 23.485 147.725 23.965 148.065 ;
        RECT 24.140 147.555 24.745 148.110 ;
        RECT 28.320 147.990 28.670 149.240 ;
        RECT 30.455 148.915 30.790 149.115 ;
        RECT 24.915 147.555 30.260 147.990 ;
        RECT 30.435 147.555 30.695 148.745 ;
        RECT 30.960 148.705 31.130 149.285 ;
        RECT 31.340 148.945 31.670 149.115 ;
        RECT 30.865 147.725 31.195 148.705 ;
        RECT 31.365 147.835 31.670 148.945 ;
        RECT 31.850 148.945 32.180 149.115 ;
        RECT 31.850 147.835 32.170 148.945 ;
        RECT 32.350 148.775 32.680 149.115 ;
        RECT 32.850 148.865 33.430 149.115 ;
        RECT 33.655 148.815 35.305 149.335 ;
        RECT 38.255 149.325 38.480 149.365 ;
        RECT 32.340 147.835 32.680 148.775 ;
        RECT 32.980 147.555 33.310 148.695 ;
        RECT 35.475 148.645 37.165 149.165 ;
        RECT 38.255 148.745 38.425 149.325 ;
        RECT 39.145 149.195 39.345 149.365 ;
        RECT 40.220 149.195 40.390 149.655 ;
        RECT 38.595 148.865 39.345 149.195 ;
        RECT 39.515 148.865 40.390 149.195 ;
        RECT 33.655 147.555 37.165 148.645 ;
        RECT 37.795 147.555 38.085 148.720 ;
        RECT 38.255 148.695 38.470 148.745 ;
        RECT 38.255 148.615 38.645 148.695 ;
        RECT 38.315 147.770 38.645 148.615 ;
        RECT 39.155 148.660 39.345 148.865 ;
        RECT 38.815 147.555 38.985 148.565 ;
        RECT 39.155 148.285 40.050 148.660 ;
        RECT 39.155 147.725 39.495 148.285 ;
        RECT 39.725 147.555 40.040 148.055 ;
        RECT 40.220 148.025 40.390 148.865 ;
        RECT 40.560 149.155 41.025 149.485 ;
        RECT 41.410 149.425 41.580 149.655 ;
        RECT 41.760 149.605 42.130 150.105 ;
        RECT 42.450 149.655 43.125 149.825 ;
        RECT 43.320 149.655 43.655 149.825 ;
        RECT 40.560 148.195 40.880 149.155 ;
        RECT 41.410 149.125 42.240 149.425 ;
        RECT 41.050 148.225 41.240 148.945 ;
        RECT 41.410 148.055 41.580 149.125 ;
        RECT 42.040 149.095 42.240 149.125 ;
        RECT 41.750 148.875 41.920 148.945 ;
        RECT 42.450 148.875 42.620 149.655 ;
        RECT 43.485 149.515 43.655 149.655 ;
        RECT 43.825 149.645 44.075 150.105 ;
        RECT 41.750 148.705 42.620 148.875 ;
        RECT 42.790 149.235 43.315 149.455 ;
        RECT 43.485 149.385 43.710 149.515 ;
        RECT 41.750 148.615 42.260 148.705 ;
        RECT 40.220 147.855 41.105 148.025 ;
        RECT 41.330 147.725 41.580 148.055 ;
        RECT 41.750 147.555 41.920 148.355 ;
        RECT 42.090 148.000 42.260 148.615 ;
        RECT 42.790 148.535 42.960 149.235 ;
        RECT 42.430 148.170 42.960 148.535 ;
        RECT 43.130 148.470 43.370 149.065 ;
        RECT 43.540 148.280 43.710 149.385 ;
        RECT 43.880 148.525 44.160 149.475 ;
        RECT 43.405 148.150 43.710 148.280 ;
        RECT 42.090 147.830 43.195 148.000 ;
        RECT 43.405 147.725 43.655 148.150 ;
        RECT 43.825 147.555 44.090 148.015 ;
        RECT 44.330 147.725 44.515 149.845 ;
        RECT 44.685 149.725 45.015 150.105 ;
        RECT 45.185 149.555 45.355 149.845 ;
        RECT 44.690 149.385 45.355 149.555 ;
        RECT 44.690 148.395 44.920 149.385 ;
        RECT 45.615 149.335 47.285 150.105 ;
        RECT 47.935 149.375 48.225 150.105 ;
        RECT 45.090 148.565 45.440 149.215 ;
        RECT 45.615 148.815 46.365 149.335 ;
        RECT 46.535 148.645 47.285 149.165 ;
        RECT 47.925 148.865 48.225 149.195 ;
        RECT 48.405 149.175 48.635 149.815 ;
        RECT 48.815 149.555 49.125 149.925 ;
        RECT 49.305 149.735 49.975 150.105 ;
        RECT 48.815 149.355 50.045 149.555 ;
        RECT 48.405 148.865 48.930 149.175 ;
        RECT 49.110 148.865 49.575 149.175 ;
        RECT 49.755 148.685 50.045 149.355 ;
        RECT 44.690 148.225 45.355 148.395 ;
        RECT 44.685 147.555 45.015 148.055 ;
        RECT 45.185 147.725 45.355 148.225 ;
        RECT 45.615 147.555 47.285 148.645 ;
        RECT 47.935 148.445 49.095 148.685 ;
        RECT 47.935 147.735 48.195 148.445 ;
        RECT 48.365 147.555 48.695 148.265 ;
        RECT 48.865 147.735 49.095 148.445 ;
        RECT 49.275 148.465 50.045 148.685 ;
        RECT 49.275 147.735 49.545 148.465 ;
        RECT 49.725 147.555 50.065 148.285 ;
        RECT 50.235 147.735 50.495 149.925 ;
        RECT 50.675 149.560 56.020 150.105 ;
        RECT 52.260 148.730 52.600 149.560 ;
        RECT 56.195 149.355 57.405 150.105 ;
        RECT 57.740 149.595 57.980 150.105 ;
        RECT 58.160 149.595 58.440 149.925 ;
        RECT 58.670 149.595 58.885 150.105 ;
        RECT 54.080 147.990 54.430 149.240 ;
        RECT 56.195 148.815 56.715 149.355 ;
        RECT 56.885 148.645 57.405 149.185 ;
        RECT 57.635 148.865 57.990 149.425 ;
        RECT 58.160 148.695 58.330 149.595 ;
        RECT 58.500 148.865 58.765 149.425 ;
        RECT 59.055 149.365 59.670 149.935 ;
        RECT 59.015 148.695 59.185 149.195 ;
        RECT 50.675 147.555 56.020 147.990 ;
        RECT 56.195 147.555 57.405 148.645 ;
        RECT 57.760 148.525 59.185 148.695 ;
        RECT 57.760 148.350 58.150 148.525 ;
        RECT 58.635 147.555 58.965 148.355 ;
        RECT 59.355 148.345 59.670 149.365 ;
        RECT 59.135 147.725 59.670 148.345 ;
        RECT 59.875 149.305 60.215 149.935 ;
        RECT 60.385 149.305 60.635 150.105 ;
        RECT 60.825 149.455 61.155 149.935 ;
        RECT 61.325 149.645 61.550 150.105 ;
        RECT 61.720 149.455 62.050 149.935 ;
        RECT 59.875 148.695 60.050 149.305 ;
        RECT 60.825 149.285 62.050 149.455 ;
        RECT 62.680 149.325 63.180 149.935 ;
        RECT 63.555 149.380 63.845 150.105 ;
        RECT 60.220 148.945 60.915 149.115 ;
        RECT 60.745 148.695 60.915 148.945 ;
        RECT 61.090 148.915 61.510 149.115 ;
        RECT 61.680 148.915 62.010 149.115 ;
        RECT 62.180 148.915 62.510 149.115 ;
        RECT 62.680 148.695 62.850 149.325 ;
        RECT 64.015 149.305 64.355 149.935 ;
        RECT 64.525 149.305 64.775 150.105 ;
        RECT 64.965 149.455 65.295 149.935 ;
        RECT 65.465 149.645 65.690 150.105 ;
        RECT 65.860 149.455 66.190 149.935 ;
        RECT 64.015 149.255 64.245 149.305 ;
        RECT 64.965 149.285 66.190 149.455 ;
        RECT 66.820 149.325 67.320 149.935 ;
        RECT 67.740 149.645 68.490 149.935 ;
        RECT 69.000 149.645 69.330 150.105 ;
        RECT 63.035 148.865 63.385 149.115 ;
        RECT 59.875 147.725 60.215 148.695 ;
        RECT 60.385 147.555 60.555 148.695 ;
        RECT 60.745 148.525 63.180 148.695 ;
        RECT 60.825 147.555 61.075 148.355 ;
        RECT 61.720 147.725 62.050 148.525 ;
        RECT 62.350 147.555 62.680 148.355 ;
        RECT 62.850 147.725 63.180 148.525 ;
        RECT 63.555 147.555 63.845 148.720 ;
        RECT 64.015 148.695 64.190 149.255 ;
        RECT 64.360 148.945 65.055 149.115 ;
        RECT 64.885 148.695 65.055 148.945 ;
        RECT 65.230 148.915 65.650 149.115 ;
        RECT 65.820 148.915 66.150 149.115 ;
        RECT 66.320 148.915 66.650 149.115 ;
        RECT 66.820 148.695 66.990 149.325 ;
        RECT 67.175 148.865 67.525 149.115 ;
        RECT 64.015 147.725 64.355 148.695 ;
        RECT 64.525 147.555 64.695 148.695 ;
        RECT 64.885 148.525 67.320 148.695 ;
        RECT 64.965 147.555 65.215 148.355 ;
        RECT 65.860 147.725 66.190 148.525 ;
        RECT 66.490 147.555 66.820 148.355 ;
        RECT 66.990 147.725 67.320 148.525 ;
        RECT 67.740 148.355 68.110 149.645 ;
        RECT 69.550 149.455 69.820 149.665 ;
        RECT 68.485 149.285 69.820 149.455 ;
        RECT 70.080 149.535 70.255 149.935 ;
        RECT 70.425 149.725 70.755 150.105 ;
        RECT 71.000 149.605 71.230 149.935 ;
        RECT 70.080 149.365 70.710 149.535 ;
        RECT 68.485 149.115 68.655 149.285 ;
        RECT 70.540 149.195 70.710 149.365 ;
        RECT 68.280 148.865 68.655 149.115 ;
        RECT 68.825 148.875 69.300 149.115 ;
        RECT 69.470 148.875 69.820 149.115 ;
        RECT 68.485 148.695 68.655 148.865 ;
        RECT 68.485 148.525 69.820 148.695 ;
        RECT 69.540 148.365 69.820 148.525 ;
        RECT 69.995 148.515 70.360 149.195 ;
        RECT 70.540 148.865 70.890 149.195 ;
        RECT 67.740 148.185 68.910 148.355 ;
        RECT 68.195 147.555 68.410 148.015 ;
        RECT 68.580 147.725 68.910 148.185 ;
        RECT 69.080 147.555 69.330 148.355 ;
        RECT 70.540 148.345 70.710 148.865 ;
        RECT 70.080 148.175 70.710 148.345 ;
        RECT 71.060 148.315 71.230 149.605 ;
        RECT 71.430 148.495 71.710 149.770 ;
        RECT 71.935 149.765 72.205 149.770 ;
        RECT 71.895 149.595 72.205 149.765 ;
        RECT 72.665 149.725 72.995 150.105 ;
        RECT 73.165 149.850 73.500 149.895 ;
        RECT 71.935 148.495 72.205 149.595 ;
        RECT 72.395 148.495 72.735 149.525 ;
        RECT 73.165 149.385 73.505 149.850 ;
        RECT 73.765 149.555 73.935 149.845 ;
        RECT 74.105 149.725 74.435 150.105 ;
        RECT 73.765 149.385 74.430 149.555 ;
        RECT 72.905 148.865 73.165 149.195 ;
        RECT 72.905 148.315 73.075 148.865 ;
        RECT 73.335 148.695 73.505 149.385 ;
        RECT 70.080 147.725 70.255 148.175 ;
        RECT 71.060 148.145 73.075 148.315 ;
        RECT 70.425 147.555 70.755 147.995 ;
        RECT 71.060 147.725 71.230 148.145 ;
        RECT 71.465 147.555 72.135 147.965 ;
        RECT 72.350 147.725 72.520 148.145 ;
        RECT 72.720 147.555 73.050 147.965 ;
        RECT 73.245 147.725 73.505 148.695 ;
        RECT 73.680 148.565 74.030 149.215 ;
        RECT 74.200 148.395 74.430 149.385 ;
        RECT 73.765 148.225 74.430 148.395 ;
        RECT 73.765 147.725 73.935 148.225 ;
        RECT 74.105 147.555 74.435 148.055 ;
        RECT 74.605 147.725 74.790 149.845 ;
        RECT 75.045 149.645 75.295 150.105 ;
        RECT 75.465 149.655 75.800 149.825 ;
        RECT 75.995 149.655 76.670 149.825 ;
        RECT 75.465 149.515 75.635 149.655 ;
        RECT 74.960 148.525 75.240 149.475 ;
        RECT 75.410 149.385 75.635 149.515 ;
        RECT 75.410 148.280 75.580 149.385 ;
        RECT 75.805 149.235 76.330 149.455 ;
        RECT 75.750 148.470 75.990 149.065 ;
        RECT 76.160 148.535 76.330 149.235 ;
        RECT 76.500 148.875 76.670 149.655 ;
        RECT 76.990 149.605 77.360 150.105 ;
        RECT 77.540 149.655 77.945 149.825 ;
        RECT 78.115 149.655 78.900 149.825 ;
        RECT 77.540 149.425 77.710 149.655 ;
        RECT 76.880 149.125 77.710 149.425 ;
        RECT 78.095 149.155 78.560 149.485 ;
        RECT 76.880 149.095 77.080 149.125 ;
        RECT 77.200 148.875 77.370 148.945 ;
        RECT 76.500 148.705 77.370 148.875 ;
        RECT 76.860 148.615 77.370 148.705 ;
        RECT 75.410 148.150 75.715 148.280 ;
        RECT 76.160 148.170 76.690 148.535 ;
        RECT 75.030 147.555 75.295 148.015 ;
        RECT 75.465 147.725 75.715 148.150 ;
        RECT 76.860 148.000 77.030 148.615 ;
        RECT 75.925 147.830 77.030 148.000 ;
        RECT 77.200 147.555 77.370 148.355 ;
        RECT 77.540 148.055 77.710 149.125 ;
        RECT 77.880 148.225 78.070 148.945 ;
        RECT 78.240 148.195 78.560 149.155 ;
        RECT 78.730 149.195 78.900 149.655 ;
        RECT 79.175 149.575 79.385 150.105 ;
        RECT 79.645 149.365 79.975 149.890 ;
        RECT 80.145 149.495 80.315 150.105 ;
        RECT 80.485 149.450 80.815 149.885 ;
        RECT 81.035 149.560 86.380 150.105 ;
        RECT 80.485 149.365 80.865 149.450 ;
        RECT 79.775 149.195 79.975 149.365 ;
        RECT 80.640 149.325 80.865 149.365 ;
        RECT 78.730 148.865 79.605 149.195 ;
        RECT 79.775 148.865 80.525 149.195 ;
        RECT 77.540 147.725 77.790 148.055 ;
        RECT 78.730 148.025 78.900 148.865 ;
        RECT 79.775 148.660 79.965 148.865 ;
        RECT 80.695 148.745 80.865 149.325 ;
        RECT 80.650 148.695 80.865 148.745 ;
        RECT 82.620 148.730 82.960 149.560 ;
        RECT 86.555 149.335 89.145 150.105 ;
        RECT 89.315 149.355 90.525 150.105 ;
        RECT 107.960 150.090 108.130 152.350 ;
        RECT 108.855 151.780 116.895 151.950 ;
        RECT 108.470 150.720 108.640 151.720 ;
        RECT 117.110 150.720 117.280 151.720 ;
        RECT 108.855 150.490 116.895 150.660 ;
        RECT 117.620 150.090 118.590 152.350 ;
        RECT 120.010 151.840 126.260 152.400 ;
        RECT 120.010 151.820 125.180 151.840 ;
        RECT 120.010 151.750 124.000 151.820 ;
        RECT 120.010 150.480 121.930 151.750 ;
        RECT 123.440 151.740 124.000 151.750 ;
        RECT 123.670 150.650 124.000 151.740 ;
        RECT 124.370 151.270 125.410 151.440 ;
        RECT 124.370 150.830 125.410 151.000 ;
        RECT 125.580 150.970 125.750 151.300 ;
        RECT 123.830 150.430 124.000 150.650 ;
        RECT 126.090 150.430 126.260 151.840 ;
        RECT 123.830 150.260 126.260 150.430 ;
        RECT 127.840 152.350 138.470 152.520 ;
        RECT 140.100 161.580 146.330 161.740 ;
        RECT 140.100 159.320 140.770 161.580 ;
        RECT 141.440 161.010 145.480 161.180 ;
        RECT 141.100 159.950 141.270 160.950 ;
        RECT 145.650 159.950 145.820 160.950 ;
        RECT 141.440 159.720 145.480 159.890 ;
        RECT 146.160 159.320 146.330 161.580 ;
        RECT 140.100 159.150 146.330 159.320 ;
        RECT 140.100 155.890 140.770 159.150 ;
        RECT 141.440 158.580 145.480 158.750 ;
        RECT 141.100 156.520 141.270 158.520 ;
        RECT 145.650 156.520 145.820 158.520 ;
        RECT 141.440 156.290 145.480 156.460 ;
        RECT 146.160 155.890 146.330 159.150 ;
        RECT 140.100 155.720 146.330 155.890 ;
        RECT 140.100 152.460 140.770 155.720 ;
        RECT 141.440 155.150 145.480 155.320 ;
        RECT 141.100 153.090 141.270 155.090 ;
        RECT 145.650 153.090 145.820 155.090 ;
        RECT 141.440 152.860 145.480 153.030 ;
        RECT 146.160 152.460 146.330 155.720 ;
        RECT 140.100 152.450 146.330 152.460 ;
        RECT 147.920 161.720 157.750 161.760 ;
        RECT 147.920 161.590 158.550 161.720 ;
        RECT 147.920 159.330 148.090 161.590 ;
        RECT 148.815 161.020 156.855 161.190 ;
        RECT 148.430 159.960 148.600 160.960 ;
        RECT 157.070 159.960 157.240 160.960 ;
        RECT 148.815 159.730 156.855 159.900 ;
        RECT 157.580 159.330 158.550 161.590 ;
        RECT 147.920 159.160 158.550 159.330 ;
        RECT 147.920 155.900 148.090 159.160 ;
        RECT 148.815 158.590 156.855 158.760 ;
        RECT 148.430 156.530 148.600 158.530 ;
        RECT 157.070 156.530 157.240 158.530 ;
        RECT 148.815 156.300 156.855 156.470 ;
        RECT 157.580 155.900 158.550 159.160 ;
        RECT 147.920 155.730 158.550 155.900 ;
        RECT 147.920 152.470 148.090 155.730 ;
        RECT 148.815 155.160 156.855 155.330 ;
        RECT 148.430 153.100 148.600 155.100 ;
        RECT 157.070 153.100 157.240 155.100 ;
        RECT 148.815 152.870 156.855 153.040 ;
        RECT 157.580 152.470 158.550 155.730 ;
        RECT 140.100 152.350 146.340 152.450 ;
        RECT 107.960 150.060 118.590 150.090 ;
        RECT 127.840 150.090 128.010 152.350 ;
        RECT 128.735 151.780 136.775 151.950 ;
        RECT 128.350 150.720 128.520 151.720 ;
        RECT 136.990 150.720 137.160 151.720 ;
        RECT 128.735 150.490 136.775 150.660 ;
        RECT 137.500 150.090 138.470 152.350 ;
        RECT 140.090 151.790 146.340 152.350 ;
        RECT 140.090 151.770 145.260 151.790 ;
        RECT 140.090 151.700 144.080 151.770 ;
        RECT 140.090 150.430 142.010 151.700 ;
        RECT 143.520 151.690 144.080 151.700 ;
        RECT 143.750 150.600 144.080 151.690 ;
        RECT 144.450 151.220 145.490 151.390 ;
        RECT 144.450 150.780 145.490 150.950 ;
        RECT 145.660 150.920 145.830 151.250 ;
        RECT 143.910 150.380 144.080 150.600 ;
        RECT 146.170 150.380 146.340 151.790 ;
        RECT 143.910 150.210 146.340 150.380 ;
        RECT 147.920 152.300 158.550 152.470 ;
        RECT 127.840 150.060 138.470 150.090 ;
        RECT 107.930 149.950 118.590 150.060 ;
        RECT 127.810 149.950 138.470 150.060 ;
        RECT 147.920 150.040 148.090 152.300 ;
        RECT 148.815 151.730 156.855 151.900 ;
        RECT 148.430 150.670 148.600 151.670 ;
        RECT 157.070 150.670 157.240 151.670 ;
        RECT 148.815 150.440 156.855 150.610 ;
        RECT 157.580 150.040 158.550 152.300 ;
        RECT 147.920 150.010 158.550 150.040 ;
        RECT 106.180 149.900 118.590 149.950 ;
        RECT 126.060 149.900 138.470 149.950 ;
        RECT 147.890 149.900 158.550 150.010 ;
        RECT 79.070 148.285 79.965 148.660 ;
        RECT 80.475 148.615 80.865 148.695 ;
        RECT 78.015 147.855 78.900 148.025 ;
        RECT 79.080 147.555 79.395 148.055 ;
        RECT 79.625 147.725 79.965 148.285 ;
        RECT 80.135 147.555 80.305 148.565 ;
        RECT 80.475 147.770 80.805 148.615 ;
        RECT 84.440 147.990 84.790 149.240 ;
        RECT 86.555 148.815 87.765 149.335 ;
        RECT 87.935 148.645 89.145 149.165 ;
        RECT 81.035 147.555 86.380 147.990 ;
        RECT 86.555 147.555 89.145 148.645 ;
        RECT 89.315 148.645 89.835 149.185 ;
        RECT 90.005 148.815 90.525 149.355 ;
        RECT 101.840 149.730 118.590 149.900 ;
        RECT 89.315 147.555 90.525 148.645 ;
        RECT 101.840 148.320 102.010 149.730 ;
        RECT 102.380 149.160 105.420 149.330 ;
        RECT 102.380 148.720 105.420 148.890 ;
        RECT 105.635 148.860 105.805 149.190 ;
        RECT 106.140 148.970 118.590 149.730 ;
        RECT 121.720 149.730 138.470 149.900 ;
        RECT 146.140 149.850 158.550 149.900 ;
        RECT 106.140 148.960 118.480 148.970 ;
        RECT 106.140 148.950 112.020 148.960 ;
        RECT 106.140 148.930 106.710 148.950 ;
        RECT 107.930 148.940 112.020 148.950 ;
        RECT 106.150 148.320 106.320 148.930 ;
        RECT 101.840 148.150 106.320 148.320 ;
        RECT 121.720 148.320 121.890 149.730 ;
        RECT 122.260 149.160 125.300 149.330 ;
        RECT 122.260 148.720 125.300 148.890 ;
        RECT 125.515 148.860 125.685 149.190 ;
        RECT 126.020 148.970 138.470 149.730 ;
        RECT 141.800 149.680 158.550 149.850 ;
        RECT 126.020 148.960 138.360 148.970 ;
        RECT 126.020 148.950 131.900 148.960 ;
        RECT 126.020 148.930 126.590 148.950 ;
        RECT 127.810 148.940 131.900 148.950 ;
        RECT 126.030 148.320 126.200 148.930 ;
        RECT 121.720 148.150 126.200 148.320 ;
        RECT 141.800 148.270 141.970 149.680 ;
        RECT 142.340 149.110 145.380 149.280 ;
        RECT 142.340 148.670 145.380 148.840 ;
        RECT 145.595 148.810 145.765 149.140 ;
        RECT 146.100 148.920 158.550 149.680 ;
        RECT 146.100 148.910 158.440 148.920 ;
        RECT 146.100 148.900 151.980 148.910 ;
        RECT 146.100 148.880 146.670 148.900 ;
        RECT 147.890 148.890 151.980 148.900 ;
        RECT 146.110 148.270 146.280 148.880 ;
        RECT 141.800 148.100 146.280 148.270 ;
        RECT 11.950 147.385 90.610 147.555 ;
        RECT 12.035 146.295 13.245 147.385 ;
        RECT 13.415 146.950 18.760 147.385 ;
        RECT 18.935 146.950 24.280 147.385 ;
        RECT 12.035 145.585 12.555 146.125 ;
        RECT 12.725 145.755 13.245 146.295 ;
        RECT 12.035 144.835 13.245 145.585 ;
        RECT 15.000 145.380 15.340 146.210 ;
        RECT 16.820 145.700 17.170 146.950 ;
        RECT 20.520 145.380 20.860 146.210 ;
        RECT 22.340 145.700 22.690 146.950 ;
        RECT 24.915 146.220 25.205 147.385 ;
        RECT 25.375 146.295 26.585 147.385 ;
        RECT 25.375 145.585 25.895 146.125 ;
        RECT 26.065 145.755 26.585 146.295 ;
        RECT 26.755 146.245 27.035 147.385 ;
        RECT 27.205 146.235 27.535 147.215 ;
        RECT 27.705 146.245 27.965 147.385 ;
        RECT 26.765 145.805 27.100 146.075 ;
        RECT 27.270 145.635 27.440 146.235 ;
        RECT 27.610 145.825 27.945 146.075 ;
        RECT 13.415 144.835 18.760 145.380 ;
        RECT 18.935 144.835 24.280 145.380 ;
        RECT 24.915 144.835 25.205 145.560 ;
        RECT 25.375 144.835 26.585 145.585 ;
        RECT 26.755 144.835 27.065 145.635 ;
        RECT 27.270 145.005 27.965 145.635 ;
        RECT 29.065 145.015 29.325 147.205 ;
        RECT 29.495 146.655 29.835 147.385 ;
        RECT 30.015 146.475 30.285 147.205 ;
        RECT 29.515 146.255 30.285 146.475 ;
        RECT 30.465 146.495 30.695 147.205 ;
        RECT 30.865 146.675 31.195 147.385 ;
        RECT 31.365 146.495 31.625 147.205 ;
        RECT 31.930 146.755 32.215 147.215 ;
        RECT 32.385 146.925 32.655 147.385 ;
        RECT 31.930 146.535 32.885 146.755 ;
        RECT 30.465 146.255 31.625 146.495 ;
        RECT 29.515 145.585 29.805 146.255 ;
        RECT 29.985 145.765 30.450 146.075 ;
        RECT 30.630 145.765 31.155 146.075 ;
        RECT 29.515 145.385 30.745 145.585 ;
        RECT 29.585 144.835 30.255 145.205 ;
        RECT 30.435 145.015 30.745 145.385 ;
        RECT 30.925 145.125 31.155 145.765 ;
        RECT 31.335 145.745 31.635 146.075 ;
        RECT 31.815 145.805 32.505 146.365 ;
        RECT 32.675 145.635 32.885 146.535 ;
        RECT 31.335 144.835 31.625 145.565 ;
        RECT 31.930 145.465 32.885 145.635 ;
        RECT 33.055 146.365 33.455 147.215 ;
        RECT 33.645 146.755 33.925 147.215 ;
        RECT 34.445 146.925 34.770 147.385 ;
        RECT 33.645 146.535 34.770 146.755 ;
        RECT 33.055 145.805 34.150 146.365 ;
        RECT 34.320 146.075 34.770 146.535 ;
        RECT 34.940 146.245 35.325 147.215 ;
        RECT 35.680 146.415 36.070 146.590 ;
        RECT 36.555 146.585 36.885 147.385 ;
        RECT 37.055 146.595 37.590 147.215 ;
        RECT 35.680 146.245 37.105 146.415 ;
        RECT 31.930 145.005 32.215 145.465 ;
        RECT 32.385 144.835 32.655 145.295 ;
        RECT 33.055 145.005 33.455 145.805 ;
        RECT 34.320 145.745 34.875 146.075 ;
        RECT 34.320 145.635 34.770 145.745 ;
        RECT 33.645 145.465 34.770 145.635 ;
        RECT 35.045 145.575 35.325 146.245 ;
        RECT 33.645 145.005 33.925 145.465 ;
        RECT 34.445 144.835 34.770 145.295 ;
        RECT 34.940 145.005 35.325 145.575 ;
        RECT 35.555 145.515 35.910 146.075 ;
        RECT 36.080 145.345 36.250 146.245 ;
        RECT 36.420 145.515 36.685 146.075 ;
        RECT 36.935 145.745 37.105 146.245 ;
        RECT 37.275 145.575 37.590 146.595 ;
        RECT 37.835 146.245 38.065 147.385 ;
        RECT 38.235 146.235 38.565 147.215 ;
        RECT 38.735 146.245 38.945 147.385 ;
        RECT 39.260 146.765 39.435 147.215 ;
        RECT 39.605 146.945 39.935 147.385 ;
        RECT 40.240 146.795 40.410 147.215 ;
        RECT 40.645 146.975 41.315 147.385 ;
        RECT 41.530 146.795 41.700 147.215 ;
        RECT 41.900 146.975 42.230 147.385 ;
        RECT 39.260 146.595 39.890 146.765 ;
        RECT 37.815 145.825 38.145 146.075 ;
        RECT 35.660 144.835 35.900 145.345 ;
        RECT 36.080 145.015 36.360 145.345 ;
        RECT 36.590 144.835 36.805 145.345 ;
        RECT 36.975 145.005 37.590 145.575 ;
        RECT 37.835 144.835 38.065 145.655 ;
        RECT 38.315 145.635 38.565 146.235 ;
        RECT 39.175 145.745 39.540 146.425 ;
        RECT 39.720 146.075 39.890 146.595 ;
        RECT 40.240 146.625 42.255 146.795 ;
        RECT 39.720 145.745 40.070 146.075 ;
        RECT 38.235 145.005 38.565 145.635 ;
        RECT 38.735 144.835 38.945 145.655 ;
        RECT 39.720 145.575 39.890 145.745 ;
        RECT 39.260 145.405 39.890 145.575 ;
        RECT 39.260 145.005 39.435 145.405 ;
        RECT 40.240 145.335 40.410 146.625 ;
        RECT 39.605 144.835 39.935 145.215 ;
        RECT 40.180 145.005 40.410 145.335 ;
        RECT 40.610 145.170 40.890 146.445 ;
        RECT 41.115 146.365 41.385 146.445 ;
        RECT 41.075 146.195 41.385 146.365 ;
        RECT 41.115 145.170 41.385 146.195 ;
        RECT 41.575 145.415 41.915 146.445 ;
        RECT 42.085 146.075 42.255 146.625 ;
        RECT 42.425 146.245 42.685 147.215 ;
        RECT 42.855 146.950 48.200 147.385 ;
        RECT 42.085 145.745 42.345 146.075 ;
        RECT 42.515 145.555 42.685 146.245 ;
        RECT 41.845 144.835 42.175 145.215 ;
        RECT 42.345 145.090 42.685 145.555 ;
        RECT 44.440 145.380 44.780 146.210 ;
        RECT 46.260 145.700 46.610 146.950 ;
        RECT 48.375 146.295 50.045 147.385 ;
        RECT 48.375 145.605 49.125 146.125 ;
        RECT 49.295 145.775 50.045 146.295 ;
        RECT 50.675 146.220 50.965 147.385 ;
        RECT 51.135 146.950 56.480 147.385 ;
        RECT 42.345 145.045 42.680 145.090 ;
        RECT 42.855 144.835 48.200 145.380 ;
        RECT 48.375 144.835 50.045 145.605 ;
        RECT 50.675 144.835 50.965 145.560 ;
        RECT 52.720 145.380 53.060 146.210 ;
        RECT 54.540 145.700 54.890 146.950 ;
        RECT 57.315 146.715 57.595 147.385 ;
        RECT 57.765 146.495 58.065 147.045 ;
        RECT 58.265 146.665 58.595 147.385 ;
        RECT 58.785 146.665 59.245 147.215 ;
        RECT 57.130 146.075 57.395 146.435 ;
        RECT 57.765 146.325 58.705 146.495 ;
        RECT 58.535 146.075 58.705 146.325 ;
        RECT 57.130 145.825 57.805 146.075 ;
        RECT 58.025 145.825 58.365 146.075 ;
        RECT 58.535 145.745 58.825 146.075 ;
        RECT 58.535 145.655 58.705 145.745 ;
        RECT 57.315 145.465 58.705 145.655 ;
        RECT 51.135 144.835 56.480 145.380 ;
        RECT 57.315 145.105 57.645 145.465 ;
        RECT 58.995 145.295 59.245 146.665 ;
        RECT 59.415 146.245 59.675 147.385 ;
        RECT 59.915 146.875 61.530 147.205 ;
        RECT 59.925 146.075 60.095 146.635 ;
        RECT 60.355 146.535 61.530 146.705 ;
        RECT 61.700 146.585 61.980 147.385 ;
        RECT 60.355 146.245 60.685 146.535 ;
        RECT 61.360 146.415 61.530 146.535 ;
        RECT 60.855 146.075 61.100 146.365 ;
        RECT 61.360 146.245 62.020 146.415 ;
        RECT 62.190 146.245 62.465 147.215 ;
        RECT 62.735 146.925 62.905 147.385 ;
        RECT 63.075 146.435 63.405 147.215 ;
        RECT 63.575 146.585 63.745 147.385 ;
        RECT 61.850 146.075 62.020 146.245 ;
        RECT 59.420 145.825 59.755 146.075 ;
        RECT 59.925 145.745 60.640 146.075 ;
        RECT 60.855 145.745 61.680 146.075 ;
        RECT 61.850 145.745 62.125 146.075 ;
        RECT 59.925 145.655 60.175 145.745 ;
        RECT 58.265 144.835 58.515 145.295 ;
        RECT 58.685 145.005 59.245 145.295 ;
        RECT 59.415 144.835 59.675 145.655 ;
        RECT 59.845 145.235 60.175 145.655 ;
        RECT 61.850 145.575 62.020 145.745 ;
        RECT 60.355 145.405 62.020 145.575 ;
        RECT 62.295 145.510 62.465 146.245 ;
        RECT 60.355 145.005 60.615 145.405 ;
        RECT 60.785 144.835 61.115 145.235 ;
        RECT 61.285 145.055 61.455 145.405 ;
        RECT 61.625 144.835 62.000 145.235 ;
        RECT 62.190 145.165 62.465 145.510 ;
        RECT 62.635 146.415 63.405 146.435 ;
        RECT 63.915 146.415 64.245 147.215 ;
        RECT 64.415 146.585 64.585 147.385 ;
        RECT 64.755 146.415 65.085 147.215 ;
        RECT 62.635 146.245 65.085 146.415 ;
        RECT 65.345 146.245 65.640 147.385 ;
        RECT 65.865 146.275 66.160 147.385 ;
        RECT 62.635 145.655 62.985 146.245 ;
        RECT 66.340 146.075 66.590 147.210 ;
        RECT 66.760 146.275 67.020 147.385 ;
        RECT 67.190 146.485 67.450 147.210 ;
        RECT 67.620 146.655 67.880 147.385 ;
        RECT 68.050 146.485 68.310 147.210 ;
        RECT 68.480 146.655 68.740 147.385 ;
        RECT 68.910 146.485 69.170 147.210 ;
        RECT 69.340 146.655 69.600 147.385 ;
        RECT 69.770 146.485 70.030 147.210 ;
        RECT 70.200 146.655 70.495 147.385 ;
        RECT 67.190 146.245 70.500 146.485 ;
        RECT 63.155 145.825 65.665 146.075 ;
        RECT 62.635 145.475 65.005 145.655 ;
        RECT 62.735 144.835 62.985 145.300 ;
        RECT 63.155 145.005 63.325 145.475 ;
        RECT 63.575 144.835 63.745 145.295 ;
        RECT 63.995 145.005 64.165 145.475 ;
        RECT 64.415 144.835 64.585 145.295 ;
        RECT 64.835 145.005 65.005 145.475 ;
        RECT 65.855 145.465 66.170 146.075 ;
        RECT 66.340 145.825 69.360 146.075 ;
        RECT 65.375 144.835 65.640 145.295 ;
        RECT 65.915 144.835 66.160 145.295 ;
        RECT 66.340 145.015 66.590 145.825 ;
        RECT 69.530 145.655 70.500 146.245 ;
        RECT 67.190 145.485 70.500 145.655 ;
        RECT 66.760 144.835 67.020 145.360 ;
        RECT 67.190 145.030 67.450 145.485 ;
        RECT 67.620 144.835 67.880 145.315 ;
        RECT 68.050 145.030 68.310 145.485 ;
        RECT 68.480 144.835 68.740 145.315 ;
        RECT 68.910 145.030 69.170 145.485 ;
        RECT 69.340 144.835 69.600 145.315 ;
        RECT 69.770 145.030 70.030 145.485 ;
        RECT 70.200 144.835 70.500 145.315 ;
        RECT 70.915 145.005 71.175 147.215 ;
        RECT 71.345 147.005 71.675 147.385 ;
        RECT 72.100 146.835 72.270 147.215 ;
        RECT 72.530 147.005 72.860 147.385 ;
        RECT 73.055 146.835 73.225 147.215 ;
        RECT 73.435 147.005 73.765 147.385 ;
        RECT 74.015 146.835 74.205 147.215 ;
        RECT 74.445 147.005 74.775 147.385 ;
        RECT 75.085 146.885 75.345 147.215 ;
        RECT 71.345 146.665 73.295 146.835 ;
        RECT 71.345 145.745 71.515 146.665 ;
        RECT 71.885 146.075 72.080 146.385 ;
        RECT 72.350 146.075 72.535 146.385 ;
        RECT 71.825 145.745 72.080 146.075 ;
        RECT 72.305 145.745 72.535 146.075 ;
        RECT 71.345 144.835 71.675 145.215 ;
        RECT 71.885 145.170 72.080 145.745 ;
        RECT 72.350 145.165 72.535 145.745 ;
        RECT 72.785 145.175 72.955 146.075 ;
        RECT 73.125 145.675 73.295 146.665 ;
        RECT 73.465 146.665 74.205 146.835 ;
        RECT 73.465 146.155 73.635 146.665 ;
        RECT 73.805 146.325 74.385 146.495 ;
        RECT 74.655 146.375 75.005 146.705 ;
        RECT 74.215 146.205 74.385 146.325 ;
        RECT 75.175 146.205 75.345 146.885 ;
        RECT 76.435 146.220 76.725 147.385 ;
        RECT 76.895 146.310 77.165 147.215 ;
        RECT 77.335 146.625 77.665 147.385 ;
        RECT 77.845 146.455 78.015 147.215 ;
        RECT 78.275 146.950 83.620 147.385 ;
        RECT 83.795 146.950 89.140 147.385 ;
        RECT 73.465 145.985 74.035 146.155 ;
        RECT 74.215 146.035 75.345 146.205 ;
        RECT 73.125 145.345 73.675 145.675 ;
        RECT 73.865 145.505 74.035 145.985 ;
        RECT 74.205 145.695 74.825 145.865 ;
        RECT 74.615 145.515 74.825 145.695 ;
        RECT 73.865 145.175 74.265 145.505 ;
        RECT 75.175 145.335 75.345 146.035 ;
        RECT 72.785 145.005 74.265 145.175 ;
        RECT 74.445 144.835 74.775 145.215 ;
        RECT 75.085 145.005 75.345 145.335 ;
        RECT 76.435 144.835 76.725 145.560 ;
        RECT 76.895 145.510 77.065 146.310 ;
        RECT 77.350 146.285 78.015 146.455 ;
        RECT 77.350 146.140 77.520 146.285 ;
        RECT 77.235 145.810 77.520 146.140 ;
        RECT 77.350 145.555 77.520 145.810 ;
        RECT 77.755 145.735 78.085 146.105 ;
        RECT 76.895 145.005 77.155 145.510 ;
        RECT 77.350 145.385 78.015 145.555 ;
        RECT 77.335 144.835 77.665 145.215 ;
        RECT 77.845 145.005 78.015 145.385 ;
        RECT 79.860 145.380 80.200 146.210 ;
        RECT 81.680 145.700 82.030 146.950 ;
        RECT 85.380 145.380 85.720 146.210 ;
        RECT 87.200 145.700 87.550 146.950 ;
        RECT 89.315 146.295 90.525 147.385 ;
        RECT 100.630 146.740 106.370 146.750 ;
        RECT 100.140 146.580 106.370 146.740 ;
        RECT 89.315 145.755 89.835 146.295 ;
        RECT 90.005 145.585 90.525 146.125 ;
        RECT 78.275 144.835 83.620 145.380 ;
        RECT 83.795 144.835 89.140 145.380 ;
        RECT 89.315 144.835 90.525 145.585 ;
        RECT 11.950 144.665 90.610 144.835 ;
        RECT 12.035 143.915 13.245 144.665 ;
        RECT 13.415 144.120 18.760 144.665 ;
        RECT 12.035 143.375 12.555 143.915 ;
        RECT 12.725 143.205 13.245 143.745 ;
        RECT 15.000 143.290 15.340 144.120 ;
        RECT 18.935 143.895 21.525 144.665 ;
        RECT 21.695 144.205 22.255 144.495 ;
        RECT 22.425 144.205 22.675 144.665 ;
        RECT 12.035 142.115 13.245 143.205 ;
        RECT 16.820 142.550 17.170 143.800 ;
        RECT 18.935 143.375 20.145 143.895 ;
        RECT 20.315 143.205 21.525 143.725 ;
        RECT 13.415 142.115 18.760 142.550 ;
        RECT 18.935 142.115 21.525 143.205 ;
        RECT 21.695 142.835 21.945 144.205 ;
        RECT 23.295 144.035 23.625 144.395 ;
        RECT 24.160 144.155 24.400 144.665 ;
        RECT 24.580 144.155 24.860 144.485 ;
        RECT 25.090 144.155 25.305 144.665 ;
        RECT 22.235 143.845 23.625 144.035 ;
        RECT 22.235 143.755 22.405 143.845 ;
        RECT 22.115 143.425 22.405 143.755 ;
        RECT 22.575 143.425 22.915 143.675 ;
        RECT 23.135 143.425 23.810 143.675 ;
        RECT 24.055 143.425 24.410 143.985 ;
        RECT 22.235 143.175 22.405 143.425 ;
        RECT 22.235 143.005 23.175 143.175 ;
        RECT 23.545 143.065 23.810 143.425 ;
        RECT 24.580 143.255 24.750 144.155 ;
        RECT 24.920 143.425 25.185 143.985 ;
        RECT 25.475 143.925 26.090 144.495 ;
        RECT 26.295 144.165 26.635 144.665 ;
        RECT 25.435 143.255 25.605 143.755 ;
        RECT 24.180 143.085 25.605 143.255 ;
        RECT 21.695 142.285 22.155 142.835 ;
        RECT 22.345 142.115 22.675 142.835 ;
        RECT 22.875 142.455 23.175 143.005 ;
        RECT 24.180 142.910 24.570 143.085 ;
        RECT 23.345 142.115 23.625 142.785 ;
        RECT 25.055 142.115 25.385 142.915 ;
        RECT 25.775 142.905 26.090 143.925 ;
        RECT 26.295 143.425 26.635 143.995 ;
        RECT 26.805 143.755 27.050 144.445 ;
        RECT 27.245 144.165 27.575 144.665 ;
        RECT 27.775 144.095 27.945 144.445 ;
        RECT 28.120 144.265 28.450 144.665 ;
        RECT 28.620 144.095 28.790 144.445 ;
        RECT 28.960 144.265 29.340 144.665 ;
        RECT 27.775 143.925 29.360 144.095 ;
        RECT 29.530 143.990 29.805 144.335 ;
        RECT 30.035 144.205 30.280 144.665 ;
        RECT 29.190 143.755 29.360 143.925 ;
        RECT 26.805 143.425 27.460 143.755 ;
        RECT 25.555 142.285 26.090 142.905 ;
        RECT 26.295 142.115 26.635 143.190 ;
        RECT 26.805 142.830 27.045 143.425 ;
        RECT 27.240 142.965 27.560 143.255 ;
        RECT 27.730 143.135 28.470 143.755 ;
        RECT 28.640 143.425 29.020 143.755 ;
        RECT 29.190 143.425 29.465 143.755 ;
        RECT 29.190 143.255 29.360 143.425 ;
        RECT 29.635 143.255 29.805 143.990 ;
        RECT 29.975 143.425 30.290 144.035 ;
        RECT 30.460 143.675 30.710 144.485 ;
        RECT 30.880 144.140 31.140 144.665 ;
        RECT 31.310 144.015 31.570 144.470 ;
        RECT 31.740 144.185 32.000 144.665 ;
        RECT 32.170 144.015 32.430 144.470 ;
        RECT 32.600 144.185 32.860 144.665 ;
        RECT 33.030 144.015 33.290 144.470 ;
        RECT 33.460 144.185 33.720 144.665 ;
        RECT 33.890 144.015 34.150 144.470 ;
        RECT 34.320 144.185 34.620 144.665 ;
        RECT 35.315 144.035 35.695 144.485 ;
        RECT 31.310 143.845 34.620 144.015 ;
        RECT 30.460 143.425 33.480 143.675 ;
        RECT 28.700 143.085 29.360 143.255 ;
        RECT 28.700 142.965 28.870 143.085 ;
        RECT 27.240 142.795 28.870 142.965 ;
        RECT 26.815 142.455 28.870 142.625 ;
        RECT 26.820 142.335 28.870 142.455 ;
        RECT 29.040 142.115 29.320 142.915 ;
        RECT 29.530 142.285 29.805 143.255 ;
        RECT 29.985 142.115 30.280 143.225 ;
        RECT 30.460 142.290 30.710 143.425 ;
        RECT 33.650 143.255 34.620 143.845 ;
        RECT 30.880 142.115 31.140 143.225 ;
        RECT 31.310 143.015 34.620 143.255 ;
        RECT 35.055 143.085 35.285 143.775 ;
        RECT 35.465 143.585 35.695 144.035 ;
        RECT 35.875 143.885 36.105 144.665 ;
        RECT 36.285 143.955 36.715 144.485 ;
        RECT 36.285 143.705 36.530 143.955 ;
        RECT 36.895 143.755 37.105 144.375 ;
        RECT 37.275 143.935 37.605 144.665 ;
        RECT 37.795 143.940 38.085 144.665 ;
        RECT 38.265 144.175 38.595 144.665 ;
        RECT 38.765 144.070 39.385 144.495 ;
        RECT 31.310 142.290 31.570 143.015 ;
        RECT 31.740 142.115 32.000 142.845 ;
        RECT 32.170 142.290 32.430 143.015 ;
        RECT 32.600 142.115 32.860 142.845 ;
        RECT 33.030 142.290 33.290 143.015 ;
        RECT 33.460 142.115 33.720 142.845 ;
        RECT 33.890 142.290 34.150 143.015 ;
        RECT 35.465 142.905 35.805 143.585 ;
        RECT 34.320 142.115 34.615 142.845 ;
        RECT 35.045 142.705 35.805 142.905 ;
        RECT 35.995 143.405 36.530 143.705 ;
        RECT 36.710 143.405 37.105 143.755 ;
        RECT 37.300 143.405 37.590 143.755 ;
        RECT 38.255 143.425 38.595 144.005 ;
        RECT 38.765 143.735 39.125 144.070 ;
        RECT 39.845 143.975 40.175 144.665 ;
        RECT 41.015 143.990 41.275 144.495 ;
        RECT 41.455 144.285 41.785 144.665 ;
        RECT 41.965 144.115 42.135 144.495 ;
        RECT 38.765 143.455 40.185 143.735 ;
        RECT 35.045 142.315 35.305 142.705 ;
        RECT 35.475 142.115 35.805 142.525 ;
        RECT 35.995 142.295 36.325 143.405 ;
        RECT 36.495 143.025 37.535 143.225 ;
        RECT 36.495 142.295 36.685 143.025 ;
        RECT 36.855 142.115 37.185 142.845 ;
        RECT 37.365 142.295 37.535 143.025 ;
        RECT 37.795 142.115 38.085 143.280 ;
        RECT 38.265 142.115 38.595 143.255 ;
        RECT 38.765 142.285 39.125 143.455 ;
        RECT 39.325 142.115 39.655 143.285 ;
        RECT 39.855 142.285 40.185 143.455 ;
        RECT 40.385 142.115 40.715 143.285 ;
        RECT 41.015 143.190 41.185 143.990 ;
        RECT 41.470 143.945 42.135 144.115 ;
        RECT 41.470 143.690 41.640 143.945 ;
        RECT 43.325 143.855 43.595 144.665 ;
        RECT 43.765 143.855 44.095 144.495 ;
        RECT 44.265 143.855 44.505 144.665 ;
        RECT 44.695 143.895 46.365 144.665 ;
        RECT 41.355 143.360 41.640 143.690 ;
        RECT 41.875 143.395 42.205 143.765 ;
        RECT 43.315 143.425 43.665 143.675 ;
        RECT 41.470 143.215 41.640 143.360 ;
        RECT 43.835 143.255 44.005 143.855 ;
        RECT 44.175 143.425 44.525 143.675 ;
        RECT 44.695 143.375 45.445 143.895 ;
        RECT 47.005 143.855 47.275 144.665 ;
        RECT 47.445 143.855 47.775 144.495 ;
        RECT 47.945 143.855 48.185 144.665 ;
        RECT 48.380 144.265 48.715 144.665 ;
        RECT 48.885 144.095 49.090 144.495 ;
        RECT 49.300 144.185 49.575 144.665 ;
        RECT 49.785 144.165 50.045 144.495 ;
        RECT 48.405 143.925 49.090 144.095 ;
        RECT 41.015 142.285 41.285 143.190 ;
        RECT 41.470 143.045 42.135 143.215 ;
        RECT 41.455 142.115 41.785 142.875 ;
        RECT 41.965 142.285 42.135 143.045 ;
        RECT 43.325 142.115 43.655 143.255 ;
        RECT 43.835 143.085 44.515 143.255 ;
        RECT 45.615 143.205 46.365 143.725 ;
        RECT 46.995 143.425 47.345 143.675 ;
        RECT 47.515 143.255 47.685 143.855 ;
        RECT 47.855 143.425 48.205 143.675 ;
        RECT 44.185 142.300 44.515 143.085 ;
        RECT 44.695 142.115 46.365 143.205 ;
        RECT 47.005 142.115 47.335 143.255 ;
        RECT 47.515 143.085 48.195 143.255 ;
        RECT 47.865 142.300 48.195 143.085 ;
        RECT 48.405 142.895 48.745 143.925 ;
        RECT 48.915 143.255 49.165 143.755 ;
        RECT 49.345 143.425 49.705 144.005 ;
        RECT 49.875 143.255 50.045 144.165 ;
        RECT 50.265 144.010 50.595 144.445 ;
        RECT 50.765 144.055 50.935 144.665 ;
        RECT 48.915 143.085 50.045 143.255 ;
        RECT 50.215 143.925 50.595 144.010 ;
        RECT 51.105 143.925 51.435 144.450 ;
        RECT 51.695 144.135 51.905 144.665 ;
        RECT 52.180 144.215 52.965 144.385 ;
        RECT 53.135 144.215 53.540 144.385 ;
        RECT 50.215 143.885 50.440 143.925 ;
        RECT 50.215 143.305 50.385 143.885 ;
        RECT 51.105 143.755 51.305 143.925 ;
        RECT 52.180 143.755 52.350 144.215 ;
        RECT 50.555 143.425 51.305 143.755 ;
        RECT 51.475 143.425 52.350 143.755 ;
        RECT 50.215 143.255 50.430 143.305 ;
        RECT 50.215 143.175 50.605 143.255 ;
        RECT 48.405 142.720 49.070 142.895 ;
        RECT 48.380 142.115 48.715 142.540 ;
        RECT 48.885 142.315 49.070 142.720 ;
        RECT 49.275 142.115 49.605 142.895 ;
        RECT 49.775 142.315 50.045 143.085 ;
        RECT 50.275 142.330 50.605 143.175 ;
        RECT 51.115 143.220 51.305 143.425 ;
        RECT 50.775 142.115 50.945 143.125 ;
        RECT 51.115 142.845 52.010 143.220 ;
        RECT 51.115 142.285 51.455 142.845 ;
        RECT 51.685 142.115 52.000 142.615 ;
        RECT 52.180 142.585 52.350 143.425 ;
        RECT 52.520 143.715 52.985 144.045 ;
        RECT 53.370 143.985 53.540 144.215 ;
        RECT 53.720 144.165 54.090 144.665 ;
        RECT 54.410 144.215 55.085 144.385 ;
        RECT 55.280 144.215 55.615 144.385 ;
        RECT 52.520 142.755 52.840 143.715 ;
        RECT 53.370 143.685 54.200 143.985 ;
        RECT 53.010 142.785 53.200 143.505 ;
        RECT 53.370 142.615 53.540 143.685 ;
        RECT 54.000 143.655 54.200 143.685 ;
        RECT 53.710 143.435 53.880 143.505 ;
        RECT 54.410 143.435 54.580 144.215 ;
        RECT 55.445 144.075 55.615 144.215 ;
        RECT 55.785 144.205 56.035 144.665 ;
        RECT 53.710 143.265 54.580 143.435 ;
        RECT 54.750 143.795 55.275 144.015 ;
        RECT 55.445 143.945 55.670 144.075 ;
        RECT 53.710 143.175 54.220 143.265 ;
        RECT 52.180 142.415 53.065 142.585 ;
        RECT 53.290 142.285 53.540 142.615 ;
        RECT 53.710 142.115 53.880 142.915 ;
        RECT 54.050 142.560 54.220 143.175 ;
        RECT 54.750 143.095 54.920 143.795 ;
        RECT 54.390 142.730 54.920 143.095 ;
        RECT 55.090 143.030 55.330 143.625 ;
        RECT 55.500 142.840 55.670 143.945 ;
        RECT 55.840 143.085 56.120 144.035 ;
        RECT 55.365 142.710 55.670 142.840 ;
        RECT 54.050 142.390 55.155 142.560 ;
        RECT 55.365 142.285 55.615 142.710 ;
        RECT 55.785 142.115 56.050 142.575 ;
        RECT 56.290 142.285 56.475 144.405 ;
        RECT 56.645 144.285 56.975 144.665 ;
        RECT 57.145 144.115 57.315 144.405 ;
        RECT 56.650 143.945 57.315 144.115 ;
        RECT 56.650 142.955 56.880 143.945 ;
        RECT 57.050 143.125 57.400 143.775 ;
        RECT 56.650 142.785 57.315 142.955 ;
        RECT 56.645 142.115 56.975 142.615 ;
        RECT 57.145 142.285 57.315 142.785 ;
        RECT 58.495 142.285 58.775 144.385 ;
        RECT 59.005 144.205 59.175 144.665 ;
        RECT 59.445 144.275 60.695 144.455 ;
        RECT 59.830 144.035 60.195 144.105 ;
        RECT 58.945 143.855 60.195 144.035 ;
        RECT 60.365 144.055 60.695 144.275 ;
        RECT 60.865 144.225 61.035 144.665 ;
        RECT 61.205 144.055 61.545 144.470 ;
        RECT 60.365 143.885 61.545 144.055 ;
        RECT 61.715 143.895 63.385 144.665 ;
        RECT 63.555 143.940 63.845 144.665 ;
        RECT 58.945 143.255 59.220 143.855 ;
        RECT 59.390 143.425 59.745 143.675 ;
        RECT 59.940 143.645 60.405 143.675 ;
        RECT 59.935 143.475 60.405 143.645 ;
        RECT 59.940 143.425 60.405 143.475 ;
        RECT 60.575 143.425 60.905 143.675 ;
        RECT 61.080 143.475 61.545 143.675 ;
        RECT 60.725 143.305 60.905 143.425 ;
        RECT 61.715 143.375 62.465 143.895 ;
        RECT 58.945 143.045 60.555 143.255 ;
        RECT 60.725 143.135 61.055 143.305 ;
        RECT 60.145 142.945 60.555 143.045 ;
        RECT 58.965 142.115 59.750 142.875 ;
        RECT 60.145 142.285 60.530 142.945 ;
        RECT 60.855 142.345 61.055 143.135 ;
        RECT 61.225 142.115 61.545 143.295 ;
        RECT 62.635 143.205 63.385 143.725 ;
        RECT 64.015 143.720 64.355 144.495 ;
        RECT 64.525 144.205 64.695 144.665 ;
        RECT 64.935 144.230 65.295 144.495 ;
        RECT 64.935 144.225 65.290 144.230 ;
        RECT 64.935 144.215 65.285 144.225 ;
        RECT 64.935 144.210 65.280 144.215 ;
        RECT 64.935 144.200 65.275 144.210 ;
        RECT 65.925 144.205 66.095 144.665 ;
        RECT 64.935 144.195 65.270 144.200 ;
        RECT 64.935 144.185 65.260 144.195 ;
        RECT 64.935 144.175 65.250 144.185 ;
        RECT 64.935 144.035 65.235 144.175 ;
        RECT 64.525 143.845 65.235 144.035 ;
        RECT 65.425 144.035 65.755 144.115 ;
        RECT 66.265 144.035 66.605 144.495 ;
        RECT 65.425 143.845 66.605 144.035 ;
        RECT 66.775 143.895 68.445 144.665 ;
        RECT 68.705 144.115 68.875 144.405 ;
        RECT 69.045 144.285 69.375 144.665 ;
        RECT 68.705 143.945 69.370 144.115 ;
        RECT 61.715 142.115 63.385 143.205 ;
        RECT 63.555 142.115 63.845 143.280 ;
        RECT 64.015 142.285 64.295 143.720 ;
        RECT 64.525 143.275 64.810 143.845 ;
        RECT 64.995 143.445 65.465 143.675 ;
        RECT 65.635 143.655 65.965 143.675 ;
        RECT 65.635 143.475 66.085 143.655 ;
        RECT 66.275 143.475 66.605 143.675 ;
        RECT 64.525 143.060 65.675 143.275 ;
        RECT 64.465 142.115 65.175 142.890 ;
        RECT 65.345 142.285 65.675 143.060 ;
        RECT 65.870 142.360 66.085 143.475 ;
        RECT 66.375 143.135 66.605 143.475 ;
        RECT 66.775 143.375 67.525 143.895 ;
        RECT 67.695 143.205 68.445 143.725 ;
        RECT 66.265 142.115 66.595 142.835 ;
        RECT 66.775 142.115 68.445 143.205 ;
        RECT 68.620 143.125 68.970 143.775 ;
        RECT 69.140 142.955 69.370 143.945 ;
        RECT 68.705 142.785 69.370 142.955 ;
        RECT 68.705 142.285 68.875 142.785 ;
        RECT 69.045 142.115 69.375 142.615 ;
        RECT 69.545 142.285 69.730 144.405 ;
        RECT 69.985 144.205 70.235 144.665 ;
        RECT 70.405 144.215 70.740 144.385 ;
        RECT 70.935 144.215 71.610 144.385 ;
        RECT 70.405 144.075 70.575 144.215 ;
        RECT 69.900 143.085 70.180 144.035 ;
        RECT 70.350 143.945 70.575 144.075 ;
        RECT 70.350 142.840 70.520 143.945 ;
        RECT 70.745 143.795 71.270 144.015 ;
        RECT 70.690 143.030 70.930 143.625 ;
        RECT 71.100 143.095 71.270 143.795 ;
        RECT 71.440 143.435 71.610 144.215 ;
        RECT 71.930 144.165 72.300 144.665 ;
        RECT 72.480 144.215 72.885 144.385 ;
        RECT 73.055 144.215 73.840 144.385 ;
        RECT 72.480 143.985 72.650 144.215 ;
        RECT 71.820 143.685 72.650 143.985 ;
        RECT 73.035 143.715 73.500 144.045 ;
        RECT 71.820 143.655 72.020 143.685 ;
        RECT 72.140 143.435 72.310 143.505 ;
        RECT 71.440 143.265 72.310 143.435 ;
        RECT 71.800 143.175 72.310 143.265 ;
        RECT 70.350 142.710 70.655 142.840 ;
        RECT 71.100 142.730 71.630 143.095 ;
        RECT 69.970 142.115 70.235 142.575 ;
        RECT 70.405 142.285 70.655 142.710 ;
        RECT 71.800 142.560 71.970 143.175 ;
        RECT 70.865 142.390 71.970 142.560 ;
        RECT 72.140 142.115 72.310 142.915 ;
        RECT 72.480 142.615 72.650 143.685 ;
        RECT 72.820 142.785 73.010 143.505 ;
        RECT 73.180 142.755 73.500 143.715 ;
        RECT 73.670 143.755 73.840 144.215 ;
        RECT 74.115 144.135 74.325 144.665 ;
        RECT 74.585 143.925 74.915 144.450 ;
        RECT 75.085 144.055 75.255 144.665 ;
        RECT 75.425 144.010 75.755 144.445 ;
        RECT 75.975 144.120 81.320 144.665 ;
        RECT 81.495 144.120 86.840 144.665 ;
        RECT 75.425 143.925 75.805 144.010 ;
        RECT 74.715 143.755 74.915 143.925 ;
        RECT 75.580 143.885 75.805 143.925 ;
        RECT 73.670 143.425 74.545 143.755 ;
        RECT 74.715 143.425 75.465 143.755 ;
        RECT 72.480 142.285 72.730 142.615 ;
        RECT 73.670 142.585 73.840 143.425 ;
        RECT 74.715 143.220 74.905 143.425 ;
        RECT 75.635 143.305 75.805 143.885 ;
        RECT 75.590 143.255 75.805 143.305 ;
        RECT 77.560 143.290 77.900 144.120 ;
        RECT 74.010 142.845 74.905 143.220 ;
        RECT 75.415 143.175 75.805 143.255 ;
        RECT 72.955 142.415 73.840 142.585 ;
        RECT 74.020 142.115 74.335 142.615 ;
        RECT 74.565 142.285 74.905 142.845 ;
        RECT 75.075 142.115 75.245 143.125 ;
        RECT 75.415 142.330 75.745 143.175 ;
        RECT 79.380 142.550 79.730 143.800 ;
        RECT 83.080 143.290 83.420 144.120 ;
        RECT 87.015 143.895 88.685 144.665 ;
        RECT 89.315 143.915 90.525 144.665 ;
        RECT 84.900 142.550 85.250 143.800 ;
        RECT 87.015 143.375 87.765 143.895 ;
        RECT 87.935 143.205 88.685 143.725 ;
        RECT 75.975 142.115 81.320 142.550 ;
        RECT 81.495 142.115 86.840 142.550 ;
        RECT 87.015 142.115 88.685 143.205 ;
        RECT 89.315 143.205 89.835 143.745 ;
        RECT 90.005 143.375 90.525 143.915 ;
        RECT 100.140 144.320 100.810 146.580 ;
        RECT 101.480 146.010 105.520 146.180 ;
        RECT 101.140 144.950 101.310 145.950 ;
        RECT 105.690 144.950 105.860 145.950 ;
        RECT 101.480 144.720 105.520 144.890 ;
        RECT 106.200 144.320 106.370 146.580 ;
        RECT 100.140 144.150 106.370 144.320 ;
        RECT 89.315 142.115 90.525 143.205 ;
        RECT 11.950 141.945 90.610 142.115 ;
        RECT 12.035 140.855 13.245 141.945 ;
        RECT 13.415 140.855 16.925 141.945 ;
        RECT 17.645 141.275 17.815 141.775 ;
        RECT 17.985 141.445 18.315 141.945 ;
        RECT 17.645 141.105 18.310 141.275 ;
        RECT 12.035 140.145 12.555 140.685 ;
        RECT 12.725 140.315 13.245 140.855 ;
        RECT 13.415 140.165 15.065 140.685 ;
        RECT 15.235 140.335 16.925 140.855 ;
        RECT 17.560 140.285 17.910 140.935 ;
        RECT 12.035 139.395 13.245 140.145 ;
        RECT 13.415 139.395 16.925 140.165 ;
        RECT 18.080 140.115 18.310 141.105 ;
        RECT 17.645 139.945 18.310 140.115 ;
        RECT 17.645 139.655 17.815 139.945 ;
        RECT 17.985 139.395 18.315 139.775 ;
        RECT 18.485 139.655 18.670 141.775 ;
        RECT 18.910 141.485 19.175 141.945 ;
        RECT 19.345 141.350 19.595 141.775 ;
        RECT 19.805 141.500 20.910 141.670 ;
        RECT 19.290 141.220 19.595 141.350 ;
        RECT 18.840 140.025 19.120 140.975 ;
        RECT 19.290 140.115 19.460 141.220 ;
        RECT 19.630 140.435 19.870 141.030 ;
        RECT 20.040 140.965 20.570 141.330 ;
        RECT 20.040 140.265 20.210 140.965 ;
        RECT 20.740 140.885 20.910 141.500 ;
        RECT 21.080 141.145 21.250 141.945 ;
        RECT 21.420 141.445 21.670 141.775 ;
        RECT 21.895 141.475 22.780 141.645 ;
        RECT 20.740 140.795 21.250 140.885 ;
        RECT 19.290 139.985 19.515 140.115 ;
        RECT 19.685 140.045 20.210 140.265 ;
        RECT 20.380 140.625 21.250 140.795 ;
        RECT 18.925 139.395 19.175 139.855 ;
        RECT 19.345 139.845 19.515 139.985 ;
        RECT 20.380 139.845 20.550 140.625 ;
        RECT 21.080 140.555 21.250 140.625 ;
        RECT 20.760 140.375 20.960 140.405 ;
        RECT 21.420 140.375 21.590 141.445 ;
        RECT 21.760 140.555 21.950 141.275 ;
        RECT 20.760 140.075 21.590 140.375 ;
        RECT 22.120 140.345 22.440 141.305 ;
        RECT 19.345 139.675 19.680 139.845 ;
        RECT 19.875 139.675 20.550 139.845 ;
        RECT 20.870 139.395 21.240 139.895 ;
        RECT 21.420 139.845 21.590 140.075 ;
        RECT 21.975 140.015 22.440 140.345 ;
        RECT 22.610 140.635 22.780 141.475 ;
        RECT 22.960 141.445 23.275 141.945 ;
        RECT 23.505 141.215 23.845 141.775 ;
        RECT 22.950 140.840 23.845 141.215 ;
        RECT 24.015 140.935 24.185 141.945 ;
        RECT 23.655 140.635 23.845 140.840 ;
        RECT 24.355 140.885 24.685 141.730 ;
        RECT 24.355 140.805 24.745 140.885 ;
        RECT 24.530 140.755 24.745 140.805 ;
        RECT 24.915 140.780 25.205 141.945 ;
        RECT 25.835 140.975 26.105 141.745 ;
        RECT 26.275 141.165 26.605 141.945 ;
        RECT 26.810 141.340 26.995 141.745 ;
        RECT 27.165 141.520 27.500 141.945 ;
        RECT 26.810 141.165 27.475 141.340 ;
        RECT 25.835 140.805 26.965 140.975 ;
        RECT 22.610 140.305 23.485 140.635 ;
        RECT 23.655 140.305 24.405 140.635 ;
        RECT 22.610 139.845 22.780 140.305 ;
        RECT 23.655 140.135 23.855 140.305 ;
        RECT 24.575 140.175 24.745 140.755 ;
        RECT 24.520 140.135 24.745 140.175 ;
        RECT 21.420 139.675 21.825 139.845 ;
        RECT 21.995 139.675 22.780 139.845 ;
        RECT 23.055 139.395 23.265 139.925 ;
        RECT 23.525 139.610 23.855 140.135 ;
        RECT 24.365 140.050 24.745 140.135 ;
        RECT 24.025 139.395 24.195 140.005 ;
        RECT 24.365 139.615 24.695 140.050 ;
        RECT 24.915 139.395 25.205 140.120 ;
        RECT 25.835 139.895 26.005 140.805 ;
        RECT 26.175 140.055 26.535 140.635 ;
        RECT 26.715 140.305 26.965 140.805 ;
        RECT 27.135 140.135 27.475 141.165 ;
        RECT 27.735 140.885 28.065 141.730 ;
        RECT 28.235 140.935 28.405 141.945 ;
        RECT 28.575 141.215 28.915 141.775 ;
        RECT 29.145 141.445 29.460 141.945 ;
        RECT 29.640 141.475 30.525 141.645 ;
        RECT 26.790 139.965 27.475 140.135 ;
        RECT 27.675 140.805 28.065 140.885 ;
        RECT 28.575 140.840 29.470 141.215 ;
        RECT 27.675 140.755 27.890 140.805 ;
        RECT 27.675 140.175 27.845 140.755 ;
        RECT 28.575 140.635 28.765 140.840 ;
        RECT 29.640 140.635 29.810 141.475 ;
        RECT 30.750 141.445 31.000 141.775 ;
        RECT 28.015 140.305 28.765 140.635 ;
        RECT 28.935 140.305 29.810 140.635 ;
        RECT 27.675 140.135 27.900 140.175 ;
        RECT 28.565 140.135 28.765 140.305 ;
        RECT 27.675 140.050 28.055 140.135 ;
        RECT 25.835 139.565 26.095 139.895 ;
        RECT 26.305 139.395 26.580 139.875 ;
        RECT 26.790 139.565 26.995 139.965 ;
        RECT 27.165 139.395 27.500 139.795 ;
        RECT 27.725 139.615 28.055 140.050 ;
        RECT 28.225 139.395 28.395 140.005 ;
        RECT 28.565 139.610 28.895 140.135 ;
        RECT 29.155 139.395 29.365 139.925 ;
        RECT 29.640 139.845 29.810 140.305 ;
        RECT 29.980 140.345 30.300 141.305 ;
        RECT 30.470 140.555 30.660 141.275 ;
        RECT 30.830 140.375 31.000 141.445 ;
        RECT 31.170 141.145 31.340 141.945 ;
        RECT 31.510 141.500 32.615 141.670 ;
        RECT 31.510 140.885 31.680 141.500 ;
        RECT 32.825 141.350 33.075 141.775 ;
        RECT 33.245 141.485 33.510 141.945 ;
        RECT 31.850 140.965 32.380 141.330 ;
        RECT 32.825 141.220 33.130 141.350 ;
        RECT 31.170 140.795 31.680 140.885 ;
        RECT 31.170 140.625 32.040 140.795 ;
        RECT 31.170 140.555 31.340 140.625 ;
        RECT 31.460 140.375 31.660 140.405 ;
        RECT 29.980 140.015 30.445 140.345 ;
        RECT 30.830 140.075 31.660 140.375 ;
        RECT 30.830 139.845 31.000 140.075 ;
        RECT 29.640 139.675 30.425 139.845 ;
        RECT 30.595 139.675 31.000 139.845 ;
        RECT 31.180 139.395 31.550 139.895 ;
        RECT 31.870 139.845 32.040 140.625 ;
        RECT 32.210 140.265 32.380 140.965 ;
        RECT 32.550 140.435 32.790 141.030 ;
        RECT 32.210 140.045 32.735 140.265 ;
        RECT 32.960 140.115 33.130 141.220 ;
        RECT 32.905 139.985 33.130 140.115 ;
        RECT 33.300 140.025 33.580 140.975 ;
        RECT 32.905 139.845 33.075 139.985 ;
        RECT 31.870 139.675 32.545 139.845 ;
        RECT 32.740 139.675 33.075 139.845 ;
        RECT 33.245 139.395 33.495 139.855 ;
        RECT 33.750 139.655 33.935 141.775 ;
        RECT 34.105 141.445 34.435 141.945 ;
        RECT 34.605 141.275 34.775 141.775 ;
        RECT 34.110 141.105 34.775 141.275 ;
        RECT 34.110 140.115 34.340 141.105 ;
        RECT 34.510 140.285 34.860 140.935 ;
        RECT 35.035 140.805 35.420 141.775 ;
        RECT 35.590 141.485 35.915 141.945 ;
        RECT 36.435 141.315 36.715 141.775 ;
        RECT 35.590 141.095 36.715 141.315 ;
        RECT 35.035 140.135 35.315 140.805 ;
        RECT 35.590 140.635 36.040 141.095 ;
        RECT 36.905 140.925 37.305 141.775 ;
        RECT 37.705 141.485 37.975 141.945 ;
        RECT 38.145 141.315 38.430 141.775 ;
        RECT 35.485 140.305 36.040 140.635 ;
        RECT 36.210 140.365 37.305 140.925 ;
        RECT 35.590 140.195 36.040 140.305 ;
        RECT 34.110 139.945 34.775 140.115 ;
        RECT 34.105 139.395 34.435 139.775 ;
        RECT 34.605 139.655 34.775 139.945 ;
        RECT 35.035 139.565 35.420 140.135 ;
        RECT 35.590 140.025 36.715 140.195 ;
        RECT 35.590 139.395 35.915 139.855 ;
        RECT 36.435 139.565 36.715 140.025 ;
        RECT 36.905 139.565 37.305 140.365 ;
        RECT 37.475 141.095 38.430 141.315 ;
        RECT 37.475 140.195 37.685 141.095 ;
        RECT 37.855 140.365 38.545 140.925 ;
        RECT 38.715 140.855 40.385 141.945 ;
        RECT 40.645 141.275 40.815 141.775 ;
        RECT 40.985 141.445 41.315 141.945 ;
        RECT 40.645 141.105 41.310 141.275 ;
        RECT 37.475 140.025 38.430 140.195 ;
        RECT 37.705 139.395 37.975 139.855 ;
        RECT 38.145 139.565 38.430 140.025 ;
        RECT 38.715 140.165 39.465 140.685 ;
        RECT 39.635 140.335 40.385 140.855 ;
        RECT 40.560 140.285 40.910 140.935 ;
        RECT 38.715 139.395 40.385 140.165 ;
        RECT 41.080 140.115 41.310 141.105 ;
        RECT 40.645 139.945 41.310 140.115 ;
        RECT 40.645 139.655 40.815 139.945 ;
        RECT 40.985 139.395 41.315 139.775 ;
        RECT 41.485 139.655 41.670 141.775 ;
        RECT 41.910 141.485 42.175 141.945 ;
        RECT 42.345 141.350 42.595 141.775 ;
        RECT 42.805 141.500 43.910 141.670 ;
        RECT 42.290 141.220 42.595 141.350 ;
        RECT 41.840 140.025 42.120 140.975 ;
        RECT 42.290 140.115 42.460 141.220 ;
        RECT 42.630 140.435 42.870 141.030 ;
        RECT 43.040 140.965 43.570 141.330 ;
        RECT 43.040 140.265 43.210 140.965 ;
        RECT 43.740 140.885 43.910 141.500 ;
        RECT 44.080 141.145 44.250 141.945 ;
        RECT 44.420 141.445 44.670 141.775 ;
        RECT 44.895 141.475 45.780 141.645 ;
        RECT 43.740 140.795 44.250 140.885 ;
        RECT 42.290 139.985 42.515 140.115 ;
        RECT 42.685 140.045 43.210 140.265 ;
        RECT 43.380 140.625 44.250 140.795 ;
        RECT 41.925 139.395 42.175 139.855 ;
        RECT 42.345 139.845 42.515 139.985 ;
        RECT 43.380 139.845 43.550 140.625 ;
        RECT 44.080 140.555 44.250 140.625 ;
        RECT 43.760 140.375 43.960 140.405 ;
        RECT 44.420 140.375 44.590 141.445 ;
        RECT 44.760 140.555 44.950 141.275 ;
        RECT 43.760 140.075 44.590 140.375 ;
        RECT 45.120 140.345 45.440 141.305 ;
        RECT 42.345 139.675 42.680 139.845 ;
        RECT 42.875 139.675 43.550 139.845 ;
        RECT 43.870 139.395 44.240 139.895 ;
        RECT 44.420 139.845 44.590 140.075 ;
        RECT 44.975 140.015 45.440 140.345 ;
        RECT 45.610 140.635 45.780 141.475 ;
        RECT 45.960 141.445 46.275 141.945 ;
        RECT 46.505 141.215 46.845 141.775 ;
        RECT 45.950 140.840 46.845 141.215 ;
        RECT 47.015 140.935 47.185 141.945 ;
        RECT 46.655 140.635 46.845 140.840 ;
        RECT 47.355 140.885 47.685 141.730 ;
        RECT 48.375 141.390 48.980 141.945 ;
        RECT 49.155 141.435 49.635 141.775 ;
        RECT 49.805 141.400 50.060 141.945 ;
        RECT 48.375 141.290 48.990 141.390 ;
        RECT 48.805 141.265 48.990 141.290 ;
        RECT 47.355 140.805 47.745 140.885 ;
        RECT 47.530 140.755 47.745 140.805 ;
        RECT 45.610 140.305 46.485 140.635 ;
        RECT 46.655 140.305 47.405 140.635 ;
        RECT 45.610 139.845 45.780 140.305 ;
        RECT 46.655 140.135 46.855 140.305 ;
        RECT 47.575 140.175 47.745 140.755 ;
        RECT 48.375 140.670 48.635 141.120 ;
        RECT 48.805 141.020 49.135 141.265 ;
        RECT 49.305 140.945 50.060 141.195 ;
        RECT 50.230 141.075 50.505 141.775 ;
        RECT 49.290 140.910 50.060 140.945 ;
        RECT 49.275 140.900 50.060 140.910 ;
        RECT 49.270 140.885 50.165 140.900 ;
        RECT 49.250 140.870 50.165 140.885 ;
        RECT 49.230 140.860 50.165 140.870 ;
        RECT 49.205 140.850 50.165 140.860 ;
        RECT 49.135 140.820 50.165 140.850 ;
        RECT 49.115 140.790 50.165 140.820 ;
        RECT 49.095 140.760 50.165 140.790 ;
        RECT 49.065 140.735 50.165 140.760 ;
        RECT 49.030 140.700 50.165 140.735 ;
        RECT 49.000 140.695 50.165 140.700 ;
        RECT 49.000 140.690 49.390 140.695 ;
        RECT 49.000 140.680 49.365 140.690 ;
        RECT 49.000 140.675 49.350 140.680 ;
        RECT 49.000 140.670 49.335 140.675 ;
        RECT 48.375 140.665 49.335 140.670 ;
        RECT 48.375 140.655 49.325 140.665 ;
        RECT 48.375 140.650 49.315 140.655 ;
        RECT 48.375 140.640 49.305 140.650 ;
        RECT 48.375 140.630 49.300 140.640 ;
        RECT 48.375 140.625 49.295 140.630 ;
        RECT 48.375 140.610 49.285 140.625 ;
        RECT 48.375 140.595 49.280 140.610 ;
        RECT 48.375 140.570 49.270 140.595 ;
        RECT 48.375 140.500 49.265 140.570 ;
        RECT 47.520 140.135 47.745 140.175 ;
        RECT 44.420 139.675 44.825 139.845 ;
        RECT 44.995 139.675 45.780 139.845 ;
        RECT 46.055 139.395 46.265 139.925 ;
        RECT 46.525 139.610 46.855 140.135 ;
        RECT 47.365 140.050 47.745 140.135 ;
        RECT 47.025 139.395 47.195 140.005 ;
        RECT 47.365 139.615 47.695 140.050 ;
        RECT 48.375 139.945 48.925 140.330 ;
        RECT 49.095 139.775 49.265 140.500 ;
        RECT 48.375 139.605 49.265 139.775 ;
        RECT 49.435 140.100 49.765 140.525 ;
        RECT 49.935 140.300 50.165 140.695 ;
        RECT 49.435 140.075 49.685 140.100 ;
        RECT 49.435 139.615 49.655 140.075 ;
        RECT 50.335 140.045 50.505 141.075 ;
        RECT 50.675 140.780 50.965 141.945 ;
        RECT 51.220 141.325 51.395 141.775 ;
        RECT 51.565 141.505 51.895 141.945 ;
        RECT 52.200 141.355 52.370 141.775 ;
        RECT 52.605 141.535 53.275 141.945 ;
        RECT 53.490 141.355 53.660 141.775 ;
        RECT 53.860 141.535 54.190 141.945 ;
        RECT 51.220 141.155 51.850 141.325 ;
        RECT 51.135 140.305 51.500 140.985 ;
        RECT 51.680 140.635 51.850 141.155 ;
        RECT 52.200 141.185 54.215 141.355 ;
        RECT 51.680 140.305 52.030 140.635 ;
        RECT 51.680 140.135 51.850 140.305 ;
        RECT 49.825 139.395 50.075 139.935 ;
        RECT 50.245 139.565 50.505 140.045 ;
        RECT 50.675 139.395 50.965 140.120 ;
        RECT 51.220 139.965 51.850 140.135 ;
        RECT 51.220 139.565 51.395 139.965 ;
        RECT 52.200 139.895 52.370 141.185 ;
        RECT 51.565 139.395 51.895 139.775 ;
        RECT 52.140 139.565 52.370 139.895 ;
        RECT 52.570 139.730 52.850 141.005 ;
        RECT 53.075 139.905 53.345 141.005 ;
        RECT 53.535 139.975 53.875 141.005 ;
        RECT 54.045 140.635 54.215 141.185 ;
        RECT 54.385 140.805 54.645 141.775 ;
        RECT 54.825 140.995 55.100 141.765 ;
        RECT 55.270 141.335 55.600 141.765 ;
        RECT 55.770 141.505 55.965 141.945 ;
        RECT 56.145 141.335 56.475 141.765 ;
        RECT 55.270 141.165 56.475 141.335 ;
        RECT 56.905 141.215 57.200 141.945 ;
        RECT 54.825 140.805 55.410 140.995 ;
        RECT 55.580 140.835 56.475 141.165 ;
        RECT 57.370 141.045 57.630 141.770 ;
        RECT 57.800 141.215 58.060 141.945 ;
        RECT 58.230 141.045 58.490 141.770 ;
        RECT 58.660 141.215 58.920 141.945 ;
        RECT 59.090 141.045 59.350 141.770 ;
        RECT 59.520 141.215 59.780 141.945 ;
        RECT 59.950 141.045 60.210 141.770 ;
        RECT 54.045 140.305 54.305 140.635 ;
        RECT 54.475 140.115 54.645 140.805 ;
        RECT 53.035 139.735 53.345 139.905 ;
        RECT 53.075 139.730 53.345 139.735 ;
        RECT 53.805 139.395 54.135 139.775 ;
        RECT 54.305 139.650 54.645 140.115 ;
        RECT 54.825 139.985 55.065 140.635 ;
        RECT 55.235 140.135 55.410 140.805 ;
        RECT 56.900 140.805 60.210 141.045 ;
        RECT 60.380 140.835 60.640 141.945 ;
        RECT 55.580 140.305 55.995 140.635 ;
        RECT 56.175 140.305 56.470 140.635 ;
        RECT 55.235 139.955 55.565 140.135 ;
        RECT 54.305 139.605 54.640 139.650 ;
        RECT 54.840 139.395 55.170 139.785 ;
        RECT 55.340 139.575 55.565 139.955 ;
        RECT 55.765 139.685 55.995 140.305 ;
        RECT 56.900 140.215 57.870 140.805 ;
        RECT 60.810 140.635 61.060 141.770 ;
        RECT 61.240 140.835 61.535 141.945 ;
        RECT 61.715 140.855 62.925 141.945 ;
        RECT 58.040 140.385 61.060 140.635 ;
        RECT 56.175 139.395 56.475 140.125 ;
        RECT 56.900 140.045 60.210 140.215 ;
        RECT 56.900 139.395 57.200 139.875 ;
        RECT 57.370 139.590 57.630 140.045 ;
        RECT 57.800 139.395 58.060 139.875 ;
        RECT 58.230 139.590 58.490 140.045 ;
        RECT 58.660 139.395 58.920 139.875 ;
        RECT 59.090 139.590 59.350 140.045 ;
        RECT 59.520 139.395 59.780 139.875 ;
        RECT 59.950 139.590 60.210 140.045 ;
        RECT 60.380 139.395 60.640 139.920 ;
        RECT 60.810 139.575 61.060 140.385 ;
        RECT 61.230 140.025 61.545 140.635 ;
        RECT 61.715 140.145 62.235 140.685 ;
        RECT 62.405 140.315 62.925 140.855 ;
        RECT 63.095 141.515 63.435 141.775 ;
        RECT 61.240 139.395 61.485 139.855 ;
        RECT 61.715 139.395 62.925 140.145 ;
        RECT 63.095 140.115 63.355 141.515 ;
        RECT 63.605 141.145 63.935 141.945 ;
        RECT 64.400 140.975 64.650 141.775 ;
        RECT 64.835 141.225 65.165 141.945 ;
        RECT 65.385 140.975 65.635 141.775 ;
        RECT 65.805 141.565 66.140 141.945 ;
        RECT 66.315 141.510 71.660 141.945 ;
        RECT 63.545 140.805 65.735 140.975 ;
        RECT 63.545 140.635 63.860 140.805 ;
        RECT 63.530 140.385 63.860 140.635 ;
        RECT 63.095 139.605 63.435 140.115 ;
        RECT 63.605 139.395 63.875 140.195 ;
        RECT 64.055 139.665 64.335 140.635 ;
        RECT 64.515 139.665 64.815 140.635 ;
        RECT 64.995 139.670 65.345 140.635 ;
        RECT 65.565 139.895 65.735 140.805 ;
        RECT 65.905 140.075 66.145 141.385 ;
        RECT 67.900 139.940 68.240 140.770 ;
        RECT 69.720 140.260 70.070 141.510 ;
        RECT 71.835 140.855 75.345 141.945 ;
        RECT 71.835 140.165 73.485 140.685 ;
        RECT 73.655 140.335 75.345 140.855 ;
        RECT 76.435 140.780 76.725 141.945 ;
        RECT 76.895 141.510 82.240 141.945 ;
        RECT 82.415 141.510 87.760 141.945 ;
        RECT 65.565 139.565 66.060 139.895 ;
        RECT 66.315 139.395 71.660 139.940 ;
        RECT 71.835 139.395 75.345 140.165 ;
        RECT 76.435 139.395 76.725 140.120 ;
        RECT 78.480 139.940 78.820 140.770 ;
        RECT 80.300 140.260 80.650 141.510 ;
        RECT 84.000 139.940 84.340 140.770 ;
        RECT 85.820 140.260 86.170 141.510 ;
        RECT 87.935 140.855 89.145 141.945 ;
        RECT 87.935 140.145 88.455 140.685 ;
        RECT 88.625 140.315 89.145 140.855 ;
        RECT 89.315 140.855 90.525 141.945 ;
        RECT 100.140 140.890 100.810 144.150 ;
        RECT 101.480 143.580 105.520 143.750 ;
        RECT 101.140 141.520 101.310 143.520 ;
        RECT 105.690 141.520 105.860 143.520 ;
        RECT 101.480 141.290 105.520 141.460 ;
        RECT 106.200 140.890 106.370 144.150 ;
        RECT 89.315 140.315 89.835 140.855 ;
        RECT 100.140 140.720 106.370 140.890 ;
        RECT 90.005 140.145 90.525 140.685 ;
        RECT 76.895 139.395 82.240 139.940 ;
        RECT 82.415 139.395 87.760 139.940 ;
        RECT 87.935 139.395 89.145 140.145 ;
        RECT 89.315 139.395 90.525 140.145 ;
        RECT 11.950 139.225 90.610 139.395 ;
        RECT 12.035 138.475 13.245 139.225 ;
        RECT 12.035 137.935 12.555 138.475 ;
        RECT 13.420 138.385 13.680 139.225 ;
        RECT 13.855 138.480 14.110 139.055 ;
        RECT 14.280 138.845 14.610 139.225 ;
        RECT 14.825 138.675 14.995 139.055 ;
        RECT 14.280 138.505 14.995 138.675 ;
        RECT 12.725 137.765 13.245 138.305 ;
        RECT 12.035 136.675 13.245 137.765 ;
        RECT 13.420 136.675 13.680 137.825 ;
        RECT 13.855 137.750 14.025 138.480 ;
        RECT 14.280 138.315 14.450 138.505 ;
        RECT 15.255 138.455 18.765 139.225 ;
        RECT 19.855 138.575 20.115 139.055 ;
        RECT 20.285 138.765 20.615 139.225 ;
        RECT 20.805 138.585 21.005 139.005 ;
        RECT 14.195 137.985 14.450 138.315 ;
        RECT 14.280 137.775 14.450 137.985 ;
        RECT 14.730 137.955 15.085 138.325 ;
        RECT 15.255 137.935 16.905 138.455 ;
        RECT 13.855 136.845 14.110 137.750 ;
        RECT 14.280 137.605 14.995 137.775 ;
        RECT 17.075 137.765 18.765 138.285 ;
        RECT 14.280 136.675 14.610 137.435 ;
        RECT 14.825 136.845 14.995 137.605 ;
        RECT 15.255 136.675 18.765 137.765 ;
        RECT 19.855 137.545 20.025 138.575 ;
        RECT 20.195 137.885 20.425 138.315 ;
        RECT 20.595 138.065 21.005 138.585 ;
        RECT 21.175 138.740 21.965 139.005 ;
        RECT 21.175 137.885 21.430 138.740 ;
        RECT 22.145 138.405 22.475 138.825 ;
        RECT 22.645 138.405 22.905 139.225 ;
        RECT 23.075 138.475 24.285 139.225 ;
        RECT 24.620 138.715 24.860 139.225 ;
        RECT 25.040 138.715 25.320 139.045 ;
        RECT 25.550 138.715 25.765 139.225 ;
        RECT 22.145 138.315 22.395 138.405 ;
        RECT 21.600 138.065 22.395 138.315 ;
        RECT 20.195 137.715 21.985 137.885 ;
        RECT 19.855 136.845 20.130 137.545 ;
        RECT 20.300 137.420 21.015 137.715 ;
        RECT 21.235 137.355 21.565 137.545 ;
        RECT 20.340 136.675 20.555 137.220 ;
        RECT 20.725 136.845 21.200 137.185 ;
        RECT 21.370 137.180 21.565 137.355 ;
        RECT 21.735 137.350 21.985 137.715 ;
        RECT 21.370 136.675 21.985 137.180 ;
        RECT 22.225 136.845 22.395 138.065 ;
        RECT 22.565 137.355 22.905 138.235 ;
        RECT 23.075 137.935 23.595 138.475 ;
        RECT 23.765 137.765 24.285 138.305 ;
        RECT 24.515 137.985 24.870 138.545 ;
        RECT 25.040 137.815 25.210 138.715 ;
        RECT 25.380 137.985 25.645 138.545 ;
        RECT 25.935 138.485 26.550 139.055 ;
        RECT 26.755 138.845 27.645 139.015 ;
        RECT 25.895 137.815 26.065 138.315 ;
        RECT 22.645 136.675 22.905 137.185 ;
        RECT 23.075 136.675 24.285 137.765 ;
        RECT 24.640 137.645 26.065 137.815 ;
        RECT 24.640 137.470 25.030 137.645 ;
        RECT 25.515 136.675 25.845 137.475 ;
        RECT 26.235 137.465 26.550 138.485 ;
        RECT 26.755 138.290 27.305 138.675 ;
        RECT 27.475 138.120 27.645 138.845 ;
        RECT 26.755 138.050 27.645 138.120 ;
        RECT 27.815 138.520 28.035 139.005 ;
        RECT 28.205 138.685 28.455 139.225 ;
        RECT 28.625 138.575 28.885 139.055 ;
        RECT 27.815 138.095 28.145 138.520 ;
        RECT 26.755 138.025 27.650 138.050 ;
        RECT 26.755 138.010 27.660 138.025 ;
        RECT 26.755 137.995 27.665 138.010 ;
        RECT 26.755 137.990 27.675 137.995 ;
        RECT 26.755 137.980 27.680 137.990 ;
        RECT 26.755 137.970 27.685 137.980 ;
        RECT 26.755 137.965 27.695 137.970 ;
        RECT 26.755 137.955 27.705 137.965 ;
        RECT 26.755 137.950 27.715 137.955 ;
        RECT 26.755 137.500 27.015 137.950 ;
        RECT 27.380 137.945 27.715 137.950 ;
        RECT 27.380 137.940 27.730 137.945 ;
        RECT 27.380 137.930 27.745 137.940 ;
        RECT 27.380 137.925 27.770 137.930 ;
        RECT 28.315 137.925 28.545 138.320 ;
        RECT 27.380 137.920 28.545 137.925 ;
        RECT 27.410 137.885 28.545 137.920 ;
        RECT 27.445 137.860 28.545 137.885 ;
        RECT 27.475 137.830 28.545 137.860 ;
        RECT 27.495 137.800 28.545 137.830 ;
        RECT 27.515 137.770 28.545 137.800 ;
        RECT 27.585 137.760 28.545 137.770 ;
        RECT 27.610 137.750 28.545 137.760 ;
        RECT 27.630 137.735 28.545 137.750 ;
        RECT 27.650 137.720 28.545 137.735 ;
        RECT 27.655 137.710 28.440 137.720 ;
        RECT 27.670 137.675 28.440 137.710 ;
        RECT 26.015 136.845 26.550 137.465 ;
        RECT 27.185 137.355 27.515 137.600 ;
        RECT 27.685 137.425 28.440 137.675 ;
        RECT 28.715 137.545 28.885 138.575 ;
        RECT 29.145 138.675 29.315 138.965 ;
        RECT 29.485 138.845 29.815 139.225 ;
        RECT 29.145 138.505 29.810 138.675 ;
        RECT 29.060 137.685 29.410 138.335 ;
        RECT 27.185 137.330 27.370 137.355 ;
        RECT 26.755 137.230 27.370 137.330 ;
        RECT 26.755 136.675 27.360 137.230 ;
        RECT 27.535 136.845 28.015 137.185 ;
        RECT 28.185 136.675 28.440 137.220 ;
        RECT 28.610 136.845 28.885 137.545 ;
        RECT 29.580 137.515 29.810 138.505 ;
        RECT 29.145 137.345 29.810 137.515 ;
        RECT 29.145 136.845 29.315 137.345 ;
        RECT 29.485 136.675 29.815 137.175 ;
        RECT 29.985 136.845 30.170 138.965 ;
        RECT 30.425 138.765 30.675 139.225 ;
        RECT 30.845 138.775 31.180 138.945 ;
        RECT 31.375 138.775 32.050 138.945 ;
        RECT 30.845 138.635 31.015 138.775 ;
        RECT 30.340 137.645 30.620 138.595 ;
        RECT 30.790 138.505 31.015 138.635 ;
        RECT 30.790 137.400 30.960 138.505 ;
        RECT 31.185 138.355 31.710 138.575 ;
        RECT 31.130 137.590 31.370 138.185 ;
        RECT 31.540 137.655 31.710 138.355 ;
        RECT 31.880 137.995 32.050 138.775 ;
        RECT 32.370 138.725 32.740 139.225 ;
        RECT 32.920 138.775 33.325 138.945 ;
        RECT 33.495 138.775 34.280 138.945 ;
        RECT 32.920 138.545 33.090 138.775 ;
        RECT 32.260 138.245 33.090 138.545 ;
        RECT 33.475 138.275 33.940 138.605 ;
        RECT 32.260 138.215 32.460 138.245 ;
        RECT 32.580 137.995 32.750 138.065 ;
        RECT 31.880 137.825 32.750 137.995 ;
        RECT 32.240 137.735 32.750 137.825 ;
        RECT 30.790 137.270 31.095 137.400 ;
        RECT 31.540 137.290 32.070 137.655 ;
        RECT 30.410 136.675 30.675 137.135 ;
        RECT 30.845 136.845 31.095 137.270 ;
        RECT 32.240 137.120 32.410 137.735 ;
        RECT 31.305 136.950 32.410 137.120 ;
        RECT 32.580 136.675 32.750 137.475 ;
        RECT 32.920 137.175 33.090 138.245 ;
        RECT 33.260 137.345 33.450 138.065 ;
        RECT 33.620 137.315 33.940 138.275 ;
        RECT 34.110 138.315 34.280 138.775 ;
        RECT 34.555 138.695 34.765 139.225 ;
        RECT 35.025 138.485 35.355 139.010 ;
        RECT 35.525 138.615 35.695 139.225 ;
        RECT 35.865 138.570 36.195 139.005 ;
        RECT 35.865 138.485 36.245 138.570 ;
        RECT 35.155 138.315 35.355 138.485 ;
        RECT 36.020 138.445 36.245 138.485 ;
        RECT 34.110 137.985 34.985 138.315 ;
        RECT 35.155 137.985 35.905 138.315 ;
        RECT 32.920 136.845 33.170 137.175 ;
        RECT 34.110 137.145 34.280 137.985 ;
        RECT 35.155 137.780 35.345 137.985 ;
        RECT 36.075 137.865 36.245 138.445 ;
        RECT 36.415 138.475 37.625 139.225 ;
        RECT 37.795 138.500 38.085 139.225 ;
        RECT 39.235 138.765 39.480 139.225 ;
        RECT 36.415 137.935 36.935 138.475 ;
        RECT 36.030 137.815 36.245 137.865 ;
        RECT 34.450 137.405 35.345 137.780 ;
        RECT 35.855 137.735 36.245 137.815 ;
        RECT 37.105 137.765 37.625 138.305 ;
        RECT 39.175 137.985 39.490 138.595 ;
        RECT 39.660 138.235 39.910 139.045 ;
        RECT 40.080 138.700 40.340 139.225 ;
        RECT 40.510 138.575 40.770 139.030 ;
        RECT 40.940 138.745 41.200 139.225 ;
        RECT 41.370 138.575 41.630 139.030 ;
        RECT 41.800 138.745 42.060 139.225 ;
        RECT 42.230 138.575 42.490 139.030 ;
        RECT 42.660 138.745 42.920 139.225 ;
        RECT 43.090 138.575 43.350 139.030 ;
        RECT 43.520 138.745 43.820 139.225 ;
        RECT 44.240 138.970 44.575 139.015 ;
        RECT 40.510 138.405 43.820 138.575 ;
        RECT 39.660 137.985 42.680 138.235 ;
        RECT 33.395 136.975 34.280 137.145 ;
        RECT 34.460 136.675 34.775 137.175 ;
        RECT 35.005 136.845 35.345 137.405 ;
        RECT 35.515 136.675 35.685 137.685 ;
        RECT 35.855 136.890 36.185 137.735 ;
        RECT 36.415 136.675 37.625 137.765 ;
        RECT 37.795 136.675 38.085 137.840 ;
        RECT 39.185 136.675 39.480 137.785 ;
        RECT 39.660 136.850 39.910 137.985 ;
        RECT 42.850 137.815 43.820 138.405 ;
        RECT 40.080 136.675 40.340 137.785 ;
        RECT 40.510 137.575 43.820 137.815 ;
        RECT 44.235 138.505 44.575 138.970 ;
        RECT 44.745 138.845 45.075 139.225 ;
        RECT 45.535 138.885 45.805 138.890 ;
        RECT 45.535 138.715 45.845 138.885 ;
        RECT 44.235 137.815 44.405 138.505 ;
        RECT 44.575 137.985 44.835 138.315 ;
        RECT 40.510 136.850 40.770 137.575 ;
        RECT 40.940 136.675 41.200 137.405 ;
        RECT 41.370 136.850 41.630 137.575 ;
        RECT 41.800 136.675 42.060 137.405 ;
        RECT 42.230 136.850 42.490 137.575 ;
        RECT 42.660 136.675 42.920 137.405 ;
        RECT 43.090 136.850 43.350 137.575 ;
        RECT 43.520 136.675 43.815 137.405 ;
        RECT 44.235 136.845 44.495 137.815 ;
        RECT 44.665 137.435 44.835 137.985 ;
        RECT 45.005 137.615 45.345 138.645 ;
        RECT 45.535 137.615 45.805 138.715 ;
        RECT 46.030 137.615 46.310 138.890 ;
        RECT 46.510 138.725 46.740 139.055 ;
        RECT 46.985 138.845 47.315 139.225 ;
        RECT 46.510 137.435 46.680 138.725 ;
        RECT 47.485 138.655 47.660 139.055 ;
        RECT 47.030 138.485 47.660 138.655 ;
        RECT 47.915 138.505 48.255 139.015 ;
        RECT 47.030 138.315 47.200 138.485 ;
        RECT 46.850 137.985 47.200 138.315 ;
        RECT 44.665 137.265 46.680 137.435 ;
        RECT 47.030 137.465 47.200 137.985 ;
        RECT 47.380 137.635 47.745 138.315 ;
        RECT 47.030 137.295 47.660 137.465 ;
        RECT 44.690 136.675 45.020 137.085 ;
        RECT 45.220 136.845 45.390 137.265 ;
        RECT 45.605 136.675 46.275 137.085 ;
        RECT 46.510 136.845 46.680 137.265 ;
        RECT 46.985 136.675 47.315 137.115 ;
        RECT 47.485 136.845 47.660 137.295 ;
        RECT 47.915 137.105 48.175 138.505 ;
        RECT 48.425 138.425 48.695 139.225 ;
        RECT 48.350 137.985 48.680 138.235 ;
        RECT 48.875 137.985 49.155 138.955 ;
        RECT 49.335 137.985 49.635 138.955 ;
        RECT 49.815 137.985 50.165 138.950 ;
        RECT 50.385 138.725 50.880 139.055 ;
        RECT 48.365 137.815 48.680 137.985 ;
        RECT 50.385 137.815 50.555 138.725 ;
        RECT 48.365 137.645 50.555 137.815 ;
        RECT 47.915 136.845 48.255 137.105 ;
        RECT 48.425 136.675 48.755 137.475 ;
        RECT 49.220 136.845 49.470 137.645 ;
        RECT 49.655 136.675 49.985 137.395 ;
        RECT 50.205 136.845 50.455 137.645 ;
        RECT 50.725 137.235 50.965 138.545 ;
        RECT 51.145 138.415 51.415 139.225 ;
        RECT 51.585 138.415 51.915 139.055 ;
        RECT 52.085 138.415 52.325 139.225 ;
        RECT 52.515 138.455 56.025 139.225 ;
        RECT 56.700 138.765 56.965 139.225 ;
        RECT 57.335 138.585 57.505 139.055 ;
        RECT 57.755 138.765 57.925 139.225 ;
        RECT 58.175 138.585 58.345 139.055 ;
        RECT 58.595 138.765 58.765 139.225 ;
        RECT 59.015 138.585 59.185 139.055 ;
        RECT 59.355 138.760 59.605 139.225 ;
        RECT 51.135 137.985 51.485 138.235 ;
        RECT 51.655 137.815 51.825 138.415 ;
        RECT 51.995 137.985 52.345 138.235 ;
        RECT 52.515 137.935 54.165 138.455 ;
        RECT 57.335 138.405 59.705 138.585 ;
        RECT 50.625 136.675 50.960 137.055 ;
        RECT 51.145 136.675 51.475 137.815 ;
        RECT 51.655 137.645 52.335 137.815 ;
        RECT 54.335 137.765 56.025 138.285 ;
        RECT 56.675 137.985 59.185 138.235 ;
        RECT 59.355 137.815 59.705 138.405 ;
        RECT 59.875 138.455 63.385 139.225 ;
        RECT 63.555 138.500 63.845 139.225 ;
        RECT 64.015 138.455 65.685 139.225 ;
        RECT 59.875 137.935 61.525 138.455 ;
        RECT 52.005 136.860 52.335 137.645 ;
        RECT 52.515 136.675 56.025 137.765 ;
        RECT 56.700 136.675 56.995 137.815 ;
        RECT 57.255 137.645 59.705 137.815 ;
        RECT 61.695 137.765 63.385 138.285 ;
        RECT 64.015 137.935 64.765 138.455 ;
        RECT 65.865 138.415 66.135 139.225 ;
        RECT 66.305 138.415 66.635 139.055 ;
        RECT 66.805 138.415 67.045 139.225 ;
        RECT 67.235 138.475 68.445 139.225 ;
        RECT 68.700 138.655 68.875 139.055 ;
        RECT 69.045 138.845 69.375 139.225 ;
        RECT 69.620 138.725 69.850 139.055 ;
        RECT 68.700 138.485 69.330 138.655 ;
        RECT 57.255 136.845 57.585 137.645 ;
        RECT 57.755 136.675 57.925 137.475 ;
        RECT 58.095 136.845 58.425 137.645 ;
        RECT 58.935 137.625 59.705 137.645 ;
        RECT 58.595 136.675 58.765 137.475 ;
        RECT 58.935 136.845 59.265 137.625 ;
        RECT 59.435 136.675 59.605 137.135 ;
        RECT 59.875 136.675 63.385 137.765 ;
        RECT 63.555 136.675 63.845 137.840 ;
        RECT 64.935 137.765 65.685 138.285 ;
        RECT 65.855 137.985 66.205 138.235 ;
        RECT 66.375 137.815 66.545 138.415 ;
        RECT 66.715 137.985 67.065 138.235 ;
        RECT 67.235 137.935 67.755 138.475 ;
        RECT 69.160 138.315 69.330 138.485 ;
        RECT 64.015 136.675 65.685 137.765 ;
        RECT 65.865 136.675 66.195 137.815 ;
        RECT 66.375 137.645 67.055 137.815 ;
        RECT 67.925 137.765 68.445 138.305 ;
        RECT 66.725 136.860 67.055 137.645 ;
        RECT 67.235 136.675 68.445 137.765 ;
        RECT 68.615 137.635 68.980 138.315 ;
        RECT 69.160 137.985 69.510 138.315 ;
        RECT 69.160 137.465 69.330 137.985 ;
        RECT 68.700 137.295 69.330 137.465 ;
        RECT 69.680 137.435 69.850 138.725 ;
        RECT 70.050 137.615 70.330 138.890 ;
        RECT 70.555 138.885 70.825 138.890 ;
        RECT 70.515 138.715 70.825 138.885 ;
        RECT 71.285 138.845 71.615 139.225 ;
        RECT 71.785 138.970 72.120 139.015 ;
        RECT 70.555 137.615 70.825 138.715 ;
        RECT 71.015 137.615 71.355 138.645 ;
        RECT 71.785 138.505 72.125 138.970 ;
        RECT 72.345 138.570 72.675 139.005 ;
        RECT 72.845 138.615 73.015 139.225 ;
        RECT 71.525 137.985 71.785 138.315 ;
        RECT 71.525 137.435 71.695 137.985 ;
        RECT 71.955 137.815 72.125 138.505 ;
        RECT 68.700 136.845 68.875 137.295 ;
        RECT 69.680 137.265 71.695 137.435 ;
        RECT 69.045 136.675 69.375 137.115 ;
        RECT 69.680 136.845 69.850 137.265 ;
        RECT 70.085 136.675 70.755 137.085 ;
        RECT 70.970 136.845 71.140 137.265 ;
        RECT 71.340 136.675 71.670 137.085 ;
        RECT 71.865 136.845 72.125 137.815 ;
        RECT 72.295 138.485 72.675 138.570 ;
        RECT 73.185 138.485 73.515 139.010 ;
        RECT 73.775 138.695 73.985 139.225 ;
        RECT 74.260 138.775 75.045 138.945 ;
        RECT 75.215 138.775 75.620 138.945 ;
        RECT 72.295 138.445 72.520 138.485 ;
        RECT 72.295 137.865 72.465 138.445 ;
        RECT 73.185 138.315 73.385 138.485 ;
        RECT 74.260 138.315 74.430 138.775 ;
        RECT 72.635 137.985 73.385 138.315 ;
        RECT 73.555 137.985 74.430 138.315 ;
        RECT 72.295 137.815 72.510 137.865 ;
        RECT 72.295 137.735 72.685 137.815 ;
        RECT 72.355 136.890 72.685 137.735 ;
        RECT 73.195 137.780 73.385 137.985 ;
        RECT 72.855 136.675 73.025 137.685 ;
        RECT 73.195 137.405 74.090 137.780 ;
        RECT 73.195 136.845 73.535 137.405 ;
        RECT 73.765 136.675 74.080 137.175 ;
        RECT 74.260 137.145 74.430 137.985 ;
        RECT 74.600 138.275 75.065 138.605 ;
        RECT 75.450 138.545 75.620 138.775 ;
        RECT 75.800 138.725 76.170 139.225 ;
        RECT 76.490 138.775 77.165 138.945 ;
        RECT 77.360 138.775 77.695 138.945 ;
        RECT 74.600 137.315 74.920 138.275 ;
        RECT 75.450 138.245 76.280 138.545 ;
        RECT 75.090 137.345 75.280 138.065 ;
        RECT 75.450 137.175 75.620 138.245 ;
        RECT 76.080 138.215 76.280 138.245 ;
        RECT 75.790 137.995 75.960 138.065 ;
        RECT 76.490 137.995 76.660 138.775 ;
        RECT 77.525 138.635 77.695 138.775 ;
        RECT 77.865 138.765 78.115 139.225 ;
        RECT 75.790 137.825 76.660 137.995 ;
        RECT 76.830 138.355 77.355 138.575 ;
        RECT 77.525 138.505 77.750 138.635 ;
        RECT 75.790 137.735 76.300 137.825 ;
        RECT 74.260 136.975 75.145 137.145 ;
        RECT 75.370 136.845 75.620 137.175 ;
        RECT 75.790 136.675 75.960 137.475 ;
        RECT 76.130 137.120 76.300 137.735 ;
        RECT 76.830 137.655 77.000 138.355 ;
        RECT 76.470 137.290 77.000 137.655 ;
        RECT 77.170 137.590 77.410 138.185 ;
        RECT 77.580 137.400 77.750 138.505 ;
        RECT 77.920 137.645 78.200 138.595 ;
        RECT 77.445 137.270 77.750 137.400 ;
        RECT 76.130 136.950 77.235 137.120 ;
        RECT 77.445 136.845 77.695 137.270 ;
        RECT 77.865 136.675 78.130 137.135 ;
        RECT 78.370 136.845 78.555 138.965 ;
        RECT 78.725 138.845 79.055 139.225 ;
        RECT 79.225 138.675 79.395 138.965 ;
        RECT 79.655 138.680 85.000 139.225 ;
        RECT 78.730 138.505 79.395 138.675 ;
        RECT 78.730 137.515 78.960 138.505 ;
        RECT 79.130 137.685 79.480 138.335 ;
        RECT 81.240 137.850 81.580 138.680 ;
        RECT 85.175 138.455 88.685 139.225 ;
        RECT 89.315 138.475 90.525 139.225 ;
        RECT 78.730 137.345 79.395 137.515 ;
        RECT 78.725 136.675 79.055 137.175 ;
        RECT 79.225 136.845 79.395 137.345 ;
        RECT 83.060 137.110 83.410 138.360 ;
        RECT 85.175 137.935 86.825 138.455 ;
        RECT 86.995 137.765 88.685 138.285 ;
        RECT 79.655 136.675 85.000 137.110 ;
        RECT 85.175 136.675 88.685 137.765 ;
        RECT 89.315 137.765 89.835 138.305 ;
        RECT 90.005 137.935 90.525 138.475 ;
        RECT 89.315 136.675 90.525 137.765 ;
        RECT 100.140 137.460 100.810 140.720 ;
        RECT 101.480 140.150 105.520 140.320 ;
        RECT 101.140 138.090 101.310 140.090 ;
        RECT 105.690 138.090 105.860 140.090 ;
        RECT 101.480 137.860 105.520 138.030 ;
        RECT 106.200 137.460 106.370 140.720 ;
        RECT 100.140 137.450 106.370 137.460 ;
        RECT 107.960 146.720 117.790 146.760 ;
        RECT 120.510 146.740 126.250 146.750 ;
        RECT 107.960 146.590 118.590 146.720 ;
        RECT 107.960 144.330 108.130 146.590 ;
        RECT 108.855 146.020 116.895 146.190 ;
        RECT 108.470 144.960 108.640 145.960 ;
        RECT 117.110 144.960 117.280 145.960 ;
        RECT 108.855 144.730 116.895 144.900 ;
        RECT 117.620 144.330 118.590 146.590 ;
        RECT 107.960 144.160 118.590 144.330 ;
        RECT 107.960 140.900 108.130 144.160 ;
        RECT 108.855 143.590 116.895 143.760 ;
        RECT 108.470 141.530 108.640 143.530 ;
        RECT 117.110 141.530 117.280 143.530 ;
        RECT 108.855 141.300 116.895 141.470 ;
        RECT 117.620 140.900 118.590 144.160 ;
        RECT 107.960 140.730 118.590 140.900 ;
        RECT 107.960 137.470 108.130 140.730 ;
        RECT 108.855 140.160 116.895 140.330 ;
        RECT 108.470 138.100 108.640 140.100 ;
        RECT 117.110 138.100 117.280 140.100 ;
        RECT 108.855 137.870 116.895 138.040 ;
        RECT 117.620 137.470 118.590 140.730 ;
        RECT 100.140 137.350 106.380 137.450 ;
        RECT 100.130 136.790 106.380 137.350 ;
        RECT 100.130 136.770 105.300 136.790 ;
        RECT 100.130 136.700 104.120 136.770 ;
        RECT 11.950 136.505 90.610 136.675 ;
        RECT 12.035 135.415 13.245 136.505 ;
        RECT 13.415 136.070 18.760 136.505 ;
        RECT 18.935 136.070 24.280 136.505 ;
        RECT 12.035 134.705 12.555 135.245 ;
        RECT 12.725 134.875 13.245 135.415 ;
        RECT 12.035 133.955 13.245 134.705 ;
        RECT 15.000 134.500 15.340 135.330 ;
        RECT 16.820 134.820 17.170 136.070 ;
        RECT 20.520 134.500 20.860 135.330 ;
        RECT 22.340 134.820 22.690 136.070 ;
        RECT 24.915 135.340 25.205 136.505 ;
        RECT 25.375 135.415 28.885 136.505 ;
        RECT 25.375 134.725 27.025 135.245 ;
        RECT 27.195 134.895 28.885 135.415 ;
        RECT 29.985 135.365 30.315 136.505 ;
        RECT 13.415 133.955 18.760 134.500 ;
        RECT 18.935 133.955 24.280 134.500 ;
        RECT 24.915 133.955 25.205 134.680 ;
        RECT 25.375 133.955 28.885 134.725 ;
        RECT 29.975 134.615 30.315 135.195 ;
        RECT 30.485 135.165 30.845 136.335 ;
        RECT 31.045 135.335 31.375 136.505 ;
        RECT 31.575 135.165 31.905 136.335 ;
        RECT 32.105 135.335 32.435 136.505 ;
        RECT 32.745 135.555 33.020 136.325 ;
        RECT 33.190 135.895 33.520 136.325 ;
        RECT 33.690 136.065 33.885 136.505 ;
        RECT 34.065 135.895 34.395 136.325 ;
        RECT 33.190 135.725 34.395 135.895 ;
        RECT 32.745 135.365 33.330 135.555 ;
        RECT 33.500 135.395 34.395 135.725 ;
        RECT 34.575 135.415 36.245 136.505 ;
        RECT 36.965 135.835 37.135 136.335 ;
        RECT 37.305 136.005 37.635 136.505 ;
        RECT 36.965 135.665 37.630 135.835 ;
        RECT 30.485 134.885 31.905 135.165 ;
        RECT 30.485 134.550 30.845 134.885 ;
        RECT 29.985 133.955 30.315 134.445 ;
        RECT 30.485 134.125 31.105 134.550 ;
        RECT 31.565 133.955 31.895 134.645 ;
        RECT 32.745 134.545 32.985 135.195 ;
        RECT 33.155 134.695 33.330 135.365 ;
        RECT 33.500 134.865 33.915 135.195 ;
        RECT 34.095 134.865 34.390 135.195 ;
        RECT 33.155 134.515 33.485 134.695 ;
        RECT 32.760 133.955 33.090 134.345 ;
        RECT 33.260 134.135 33.485 134.515 ;
        RECT 33.685 134.245 33.915 134.865 ;
        RECT 34.575 134.725 35.325 135.245 ;
        RECT 35.495 134.895 36.245 135.415 ;
        RECT 36.880 134.845 37.230 135.495 ;
        RECT 34.095 133.955 34.395 134.685 ;
        RECT 34.575 133.955 36.245 134.725 ;
        RECT 37.400 134.675 37.630 135.665 ;
        RECT 36.965 134.505 37.630 134.675 ;
        RECT 36.965 134.215 37.135 134.505 ;
        RECT 37.305 133.955 37.635 134.335 ;
        RECT 37.805 134.215 37.990 136.335 ;
        RECT 38.230 136.045 38.495 136.505 ;
        RECT 38.665 135.910 38.915 136.335 ;
        RECT 39.125 136.060 40.230 136.230 ;
        RECT 38.610 135.780 38.915 135.910 ;
        RECT 38.160 134.585 38.440 135.535 ;
        RECT 38.610 134.675 38.780 135.780 ;
        RECT 38.950 134.995 39.190 135.590 ;
        RECT 39.360 135.525 39.890 135.890 ;
        RECT 39.360 134.825 39.530 135.525 ;
        RECT 40.060 135.445 40.230 136.060 ;
        RECT 40.400 135.705 40.570 136.505 ;
        RECT 40.740 136.005 40.990 136.335 ;
        RECT 41.215 136.035 42.100 136.205 ;
        RECT 40.060 135.355 40.570 135.445 ;
        RECT 38.610 134.545 38.835 134.675 ;
        RECT 39.005 134.605 39.530 134.825 ;
        RECT 39.700 135.185 40.570 135.355 ;
        RECT 38.245 133.955 38.495 134.415 ;
        RECT 38.665 134.405 38.835 134.545 ;
        RECT 39.700 134.405 39.870 135.185 ;
        RECT 40.400 135.115 40.570 135.185 ;
        RECT 40.080 134.935 40.280 134.965 ;
        RECT 40.740 134.935 40.910 136.005 ;
        RECT 41.080 135.115 41.270 135.835 ;
        RECT 40.080 134.635 40.910 134.935 ;
        RECT 41.440 134.905 41.760 135.865 ;
        RECT 38.665 134.235 39.000 134.405 ;
        RECT 39.195 134.235 39.870 134.405 ;
        RECT 40.190 133.955 40.560 134.455 ;
        RECT 40.740 134.405 40.910 134.635 ;
        RECT 41.295 134.575 41.760 134.905 ;
        RECT 41.930 135.195 42.100 136.035 ;
        RECT 42.280 136.005 42.595 136.505 ;
        RECT 42.825 135.775 43.165 136.335 ;
        RECT 42.270 135.400 43.165 135.775 ;
        RECT 43.335 135.495 43.505 136.505 ;
        RECT 42.975 135.195 43.165 135.400 ;
        RECT 43.675 135.445 44.005 136.290 ;
        RECT 44.235 136.070 49.580 136.505 ;
        RECT 43.675 135.365 44.065 135.445 ;
        RECT 43.850 135.315 44.065 135.365 ;
        RECT 41.930 134.865 42.805 135.195 ;
        RECT 42.975 134.865 43.725 135.195 ;
        RECT 41.930 134.405 42.100 134.865 ;
        RECT 42.975 134.695 43.175 134.865 ;
        RECT 43.895 134.735 44.065 135.315 ;
        RECT 43.840 134.695 44.065 134.735 ;
        RECT 40.740 134.235 41.145 134.405 ;
        RECT 41.315 134.235 42.100 134.405 ;
        RECT 42.375 133.955 42.585 134.485 ;
        RECT 42.845 134.170 43.175 134.695 ;
        RECT 43.685 134.610 44.065 134.695 ;
        RECT 43.345 133.955 43.515 134.565 ;
        RECT 43.685 134.175 44.015 134.610 ;
        RECT 45.820 134.500 46.160 135.330 ;
        RECT 47.640 134.820 47.990 136.070 ;
        RECT 50.675 135.340 50.965 136.505 ;
        RECT 51.140 136.080 51.475 136.505 ;
        RECT 51.645 135.900 51.830 136.305 ;
        RECT 51.165 135.725 51.830 135.900 ;
        RECT 52.035 135.725 52.365 136.505 ;
        RECT 51.165 134.695 51.505 135.725 ;
        RECT 52.535 135.535 52.805 136.305 ;
        RECT 51.675 135.365 52.805 135.535 ;
        RECT 52.975 135.415 56.485 136.505 ;
        RECT 56.740 135.885 56.915 136.335 ;
        RECT 57.085 136.065 57.415 136.505 ;
        RECT 57.720 135.915 57.890 136.335 ;
        RECT 58.125 136.095 58.795 136.505 ;
        RECT 59.010 135.915 59.180 136.335 ;
        RECT 59.380 136.095 59.710 136.505 ;
        RECT 56.740 135.715 57.370 135.885 ;
        RECT 51.675 134.865 51.925 135.365 ;
        RECT 44.235 133.955 49.580 134.500 ;
        RECT 50.675 133.955 50.965 134.680 ;
        RECT 51.165 134.525 51.850 134.695 ;
        RECT 52.105 134.615 52.465 135.195 ;
        RECT 51.140 133.955 51.475 134.355 ;
        RECT 51.645 134.125 51.850 134.525 ;
        RECT 52.635 134.455 52.805 135.365 ;
        RECT 52.060 133.955 52.335 134.435 ;
        RECT 52.545 134.125 52.805 134.455 ;
        RECT 52.975 134.725 54.625 135.245 ;
        RECT 54.795 134.895 56.485 135.415 ;
        RECT 56.655 134.865 57.020 135.545 ;
        RECT 57.200 135.195 57.370 135.715 ;
        RECT 57.720 135.745 59.735 135.915 ;
        RECT 57.200 134.865 57.550 135.195 ;
        RECT 52.975 133.955 56.485 134.725 ;
        RECT 57.200 134.695 57.370 134.865 ;
        RECT 56.740 134.525 57.370 134.695 ;
        RECT 56.740 134.125 56.915 134.525 ;
        RECT 57.720 134.455 57.890 135.745 ;
        RECT 57.085 133.955 57.415 134.335 ;
        RECT 57.660 134.125 57.890 134.455 ;
        RECT 58.090 134.290 58.370 135.565 ;
        RECT 58.595 135.485 58.865 135.565 ;
        RECT 58.555 135.315 58.865 135.485 ;
        RECT 58.595 134.290 58.865 135.315 ;
        RECT 59.055 134.535 59.395 135.565 ;
        RECT 59.565 135.195 59.735 135.745 ;
        RECT 59.905 135.365 60.165 136.335 ;
        RECT 60.345 135.365 60.675 136.505 ;
        RECT 61.205 135.535 61.535 136.320 ;
        RECT 60.855 135.365 61.535 135.535 ;
        RECT 62.185 135.365 62.515 136.505 ;
        RECT 63.045 135.535 63.375 136.320 ;
        RECT 62.695 135.365 63.375 135.535 ;
        RECT 64.475 135.635 64.750 136.335 ;
        RECT 64.920 135.960 65.175 136.505 ;
        RECT 65.345 135.995 65.825 136.335 ;
        RECT 66.000 135.950 66.605 136.505 ;
        RECT 65.990 135.850 66.605 135.950 ;
        RECT 65.990 135.825 66.175 135.850 ;
        RECT 59.565 134.865 59.825 135.195 ;
        RECT 59.995 134.675 60.165 135.365 ;
        RECT 60.335 134.945 60.685 135.195 ;
        RECT 60.855 134.765 61.025 135.365 ;
        RECT 61.195 134.945 61.545 135.195 ;
        RECT 62.175 134.945 62.525 135.195 ;
        RECT 62.695 134.765 62.865 135.365 ;
        RECT 63.035 134.945 63.385 135.195 ;
        RECT 59.325 133.955 59.655 134.335 ;
        RECT 59.825 134.210 60.165 134.675 ;
        RECT 59.825 134.165 60.160 134.210 ;
        RECT 60.345 133.955 60.615 134.765 ;
        RECT 60.785 134.125 61.115 134.765 ;
        RECT 61.285 133.955 61.525 134.765 ;
        RECT 62.185 133.955 62.455 134.765 ;
        RECT 62.625 134.125 62.955 134.765 ;
        RECT 63.125 133.955 63.365 134.765 ;
        RECT 64.475 134.605 64.645 135.635 ;
        RECT 64.920 135.505 65.675 135.755 ;
        RECT 65.845 135.580 66.175 135.825 ;
        RECT 64.920 135.470 65.690 135.505 ;
        RECT 64.920 135.460 65.705 135.470 ;
        RECT 64.815 135.445 65.710 135.460 ;
        RECT 64.815 135.430 65.730 135.445 ;
        RECT 64.815 135.420 65.750 135.430 ;
        RECT 64.815 135.410 65.775 135.420 ;
        RECT 64.815 135.380 65.845 135.410 ;
        RECT 64.815 135.350 65.865 135.380 ;
        RECT 64.815 135.320 65.885 135.350 ;
        RECT 64.815 135.295 65.915 135.320 ;
        RECT 64.815 135.260 65.950 135.295 ;
        RECT 64.815 135.255 65.980 135.260 ;
        RECT 64.815 134.860 65.045 135.255 ;
        RECT 65.590 135.250 65.980 135.255 ;
        RECT 65.615 135.240 65.980 135.250 ;
        RECT 65.630 135.235 65.980 135.240 ;
        RECT 65.645 135.230 65.980 135.235 ;
        RECT 66.345 135.230 66.605 135.680 ;
        RECT 66.785 135.555 67.060 136.325 ;
        RECT 67.230 135.895 67.560 136.325 ;
        RECT 67.730 136.065 67.925 136.505 ;
        RECT 68.105 135.895 68.435 136.325 ;
        RECT 67.230 135.725 68.435 135.895 ;
        RECT 66.785 135.365 67.370 135.555 ;
        RECT 67.540 135.395 68.435 135.725 ;
        RECT 69.535 135.655 69.915 136.335 ;
        RECT 70.505 135.655 70.675 136.505 ;
        RECT 70.845 135.825 71.175 136.335 ;
        RECT 71.345 135.995 71.515 136.505 ;
        RECT 71.685 135.825 72.085 136.335 ;
        RECT 70.845 135.655 72.085 135.825 ;
        RECT 65.645 135.225 66.605 135.230 ;
        RECT 65.655 135.215 66.605 135.225 ;
        RECT 65.665 135.210 66.605 135.215 ;
        RECT 65.675 135.200 66.605 135.210 ;
        RECT 65.680 135.190 66.605 135.200 ;
        RECT 65.685 135.185 66.605 135.190 ;
        RECT 65.695 135.170 66.605 135.185 ;
        RECT 65.700 135.155 66.605 135.170 ;
        RECT 65.710 135.130 66.605 135.155 ;
        RECT 65.215 134.660 65.545 135.085 ;
        RECT 64.475 134.125 64.735 134.605 ;
        RECT 64.905 133.955 65.155 134.495 ;
        RECT 65.325 134.175 65.545 134.660 ;
        RECT 65.715 135.060 66.605 135.130 ;
        RECT 65.715 134.335 65.885 135.060 ;
        RECT 66.055 134.505 66.605 134.890 ;
        RECT 66.785 134.545 67.025 135.195 ;
        RECT 67.195 134.695 67.370 135.365 ;
        RECT 67.540 134.865 67.955 135.195 ;
        RECT 68.135 134.865 68.430 135.195 ;
        RECT 67.195 134.515 67.525 134.695 ;
        RECT 65.715 134.165 66.605 134.335 ;
        RECT 66.800 133.955 67.130 134.345 ;
        RECT 67.300 134.135 67.525 134.515 ;
        RECT 67.725 134.245 67.955 134.865 ;
        RECT 69.535 134.695 69.705 135.655 ;
        RECT 69.875 135.315 71.180 135.485 ;
        RECT 72.265 135.405 72.585 136.335 ;
        RECT 72.755 135.415 76.265 136.505 ;
        RECT 69.875 134.865 70.120 135.315 ;
        RECT 70.290 134.945 70.840 135.145 ;
        RECT 71.010 135.115 71.180 135.315 ;
        RECT 71.955 135.235 72.585 135.405 ;
        RECT 71.010 134.945 71.385 135.115 ;
        RECT 71.555 134.695 71.785 135.195 ;
        RECT 68.135 133.955 68.435 134.685 ;
        RECT 69.535 134.525 71.785 134.695 ;
        RECT 69.585 133.955 69.915 134.345 ;
        RECT 70.085 134.205 70.255 134.525 ;
        RECT 71.955 134.355 72.125 135.235 ;
        RECT 70.425 133.955 70.755 134.345 ;
        RECT 71.170 134.185 72.125 134.355 ;
        RECT 72.295 133.955 72.585 134.790 ;
        RECT 72.755 134.725 74.405 135.245 ;
        RECT 74.575 134.895 76.265 135.415 ;
        RECT 76.435 135.340 76.725 136.505 ;
        RECT 76.895 136.070 82.240 136.505 ;
        RECT 82.415 136.070 87.760 136.505 ;
        RECT 72.755 133.955 76.265 134.725 ;
        RECT 76.435 133.955 76.725 134.680 ;
        RECT 78.480 134.500 78.820 135.330 ;
        RECT 80.300 134.820 80.650 136.070 ;
        RECT 84.000 134.500 84.340 135.330 ;
        RECT 85.820 134.820 86.170 136.070 ;
        RECT 87.935 135.415 89.145 136.505 ;
        RECT 87.935 134.705 88.455 135.245 ;
        RECT 88.625 134.875 89.145 135.415 ;
        RECT 89.315 135.415 90.525 136.505 ;
        RECT 100.130 135.430 102.050 136.700 ;
        RECT 103.560 136.690 104.120 136.700 ;
        RECT 103.790 135.600 104.120 136.690 ;
        RECT 104.490 136.220 105.530 136.390 ;
        RECT 104.490 135.780 105.530 135.950 ;
        RECT 105.700 135.920 105.870 136.250 ;
        RECT 89.315 134.875 89.835 135.415 ;
        RECT 103.950 135.380 104.120 135.600 ;
        RECT 106.210 135.380 106.380 136.790 ;
        RECT 90.005 134.705 90.525 135.245 ;
        RECT 103.950 135.210 106.380 135.380 ;
        RECT 107.960 137.300 118.590 137.470 ;
        RECT 120.020 146.580 126.250 146.740 ;
        RECT 120.020 144.320 120.690 146.580 ;
        RECT 121.360 146.010 125.400 146.180 ;
        RECT 121.020 144.950 121.190 145.950 ;
        RECT 125.570 144.950 125.740 145.950 ;
        RECT 121.360 144.720 125.400 144.890 ;
        RECT 126.080 144.320 126.250 146.580 ;
        RECT 120.020 144.150 126.250 144.320 ;
        RECT 120.020 140.890 120.690 144.150 ;
        RECT 121.360 143.580 125.400 143.750 ;
        RECT 121.020 141.520 121.190 143.520 ;
        RECT 125.570 141.520 125.740 143.520 ;
        RECT 121.360 141.290 125.400 141.460 ;
        RECT 126.080 140.890 126.250 144.150 ;
        RECT 120.020 140.720 126.250 140.890 ;
        RECT 120.020 137.460 120.690 140.720 ;
        RECT 121.360 140.150 125.400 140.320 ;
        RECT 121.020 138.090 121.190 140.090 ;
        RECT 125.570 138.090 125.740 140.090 ;
        RECT 121.360 137.860 125.400 138.030 ;
        RECT 126.080 137.460 126.250 140.720 ;
        RECT 120.020 137.450 126.250 137.460 ;
        RECT 127.840 146.720 137.670 146.760 ;
        RECT 140.540 146.740 146.280 146.750 ;
        RECT 127.840 146.590 138.470 146.720 ;
        RECT 127.840 144.330 128.010 146.590 ;
        RECT 128.735 146.020 136.775 146.190 ;
        RECT 128.350 144.960 128.520 145.960 ;
        RECT 136.990 144.960 137.160 145.960 ;
        RECT 128.735 144.730 136.775 144.900 ;
        RECT 137.500 144.330 138.470 146.590 ;
        RECT 127.840 144.160 138.470 144.330 ;
        RECT 127.840 140.900 128.010 144.160 ;
        RECT 128.735 143.590 136.775 143.760 ;
        RECT 128.350 141.530 128.520 143.530 ;
        RECT 136.990 141.530 137.160 143.530 ;
        RECT 128.735 141.300 136.775 141.470 ;
        RECT 137.500 140.900 138.470 144.160 ;
        RECT 127.840 140.730 138.470 140.900 ;
        RECT 127.840 137.470 128.010 140.730 ;
        RECT 128.735 140.160 136.775 140.330 ;
        RECT 128.350 138.100 128.520 140.100 ;
        RECT 136.990 138.100 137.160 140.100 ;
        RECT 128.735 137.870 136.775 138.040 ;
        RECT 137.500 137.470 138.470 140.730 ;
        RECT 120.020 137.350 126.260 137.450 ;
        RECT 107.960 135.040 108.130 137.300 ;
        RECT 108.855 136.730 116.895 136.900 ;
        RECT 108.470 135.670 108.640 136.670 ;
        RECT 117.110 135.670 117.280 136.670 ;
        RECT 108.855 135.440 116.895 135.610 ;
        RECT 117.620 135.040 118.590 137.300 ;
        RECT 120.010 136.790 126.260 137.350 ;
        RECT 120.010 136.770 125.180 136.790 ;
        RECT 120.010 136.700 124.000 136.770 ;
        RECT 120.010 135.430 121.930 136.700 ;
        RECT 123.440 136.690 124.000 136.700 ;
        RECT 123.670 135.600 124.000 136.690 ;
        RECT 124.370 136.220 125.410 136.390 ;
        RECT 124.370 135.780 125.410 135.950 ;
        RECT 125.580 135.920 125.750 136.250 ;
        RECT 123.830 135.380 124.000 135.600 ;
        RECT 126.090 135.380 126.260 136.790 ;
        RECT 123.830 135.210 126.260 135.380 ;
        RECT 127.840 137.300 138.470 137.470 ;
        RECT 140.050 146.580 146.280 146.740 ;
        RECT 140.050 144.320 140.720 146.580 ;
        RECT 141.390 146.010 145.430 146.180 ;
        RECT 141.050 144.950 141.220 145.950 ;
        RECT 145.600 144.950 145.770 145.950 ;
        RECT 141.390 144.720 145.430 144.890 ;
        RECT 146.110 144.320 146.280 146.580 ;
        RECT 140.050 144.150 146.280 144.320 ;
        RECT 140.050 140.890 140.720 144.150 ;
        RECT 141.390 143.580 145.430 143.750 ;
        RECT 141.050 141.520 141.220 143.520 ;
        RECT 145.600 141.520 145.770 143.520 ;
        RECT 141.390 141.290 145.430 141.460 ;
        RECT 146.110 140.890 146.280 144.150 ;
        RECT 140.050 140.720 146.280 140.890 ;
        RECT 140.050 137.460 140.720 140.720 ;
        RECT 141.390 140.150 145.430 140.320 ;
        RECT 141.050 138.090 141.220 140.090 ;
        RECT 145.600 138.090 145.770 140.090 ;
        RECT 141.390 137.860 145.430 138.030 ;
        RECT 146.110 137.460 146.280 140.720 ;
        RECT 140.050 137.450 146.280 137.460 ;
        RECT 147.870 146.720 157.700 146.760 ;
        RECT 147.870 146.590 158.500 146.720 ;
        RECT 147.870 144.330 148.040 146.590 ;
        RECT 148.765 146.020 156.805 146.190 ;
        RECT 148.380 144.960 148.550 145.960 ;
        RECT 157.020 144.960 157.190 145.960 ;
        RECT 148.765 144.730 156.805 144.900 ;
        RECT 157.530 144.330 158.500 146.590 ;
        RECT 147.870 144.160 158.500 144.330 ;
        RECT 147.870 140.900 148.040 144.160 ;
        RECT 148.765 143.590 156.805 143.760 ;
        RECT 148.380 141.530 148.550 143.530 ;
        RECT 157.020 141.530 157.190 143.530 ;
        RECT 148.765 141.300 156.805 141.470 ;
        RECT 157.530 140.900 158.500 144.160 ;
        RECT 147.870 140.730 158.500 140.900 ;
        RECT 147.870 137.470 148.040 140.730 ;
        RECT 148.765 140.160 156.805 140.330 ;
        RECT 148.380 138.100 148.550 140.100 ;
        RECT 157.020 138.100 157.190 140.100 ;
        RECT 148.765 137.870 156.805 138.040 ;
        RECT 157.530 137.470 158.500 140.730 ;
        RECT 140.050 137.350 146.290 137.450 ;
        RECT 107.960 135.010 118.590 135.040 ;
        RECT 127.840 135.040 128.010 137.300 ;
        RECT 128.735 136.730 136.775 136.900 ;
        RECT 128.350 135.670 128.520 136.670 ;
        RECT 136.990 135.670 137.160 136.670 ;
        RECT 128.735 135.440 136.775 135.610 ;
        RECT 137.500 135.040 138.470 137.300 ;
        RECT 140.040 136.790 146.290 137.350 ;
        RECT 140.040 136.770 145.210 136.790 ;
        RECT 140.040 136.700 144.030 136.770 ;
        RECT 140.040 135.430 141.960 136.700 ;
        RECT 143.470 136.690 144.030 136.700 ;
        RECT 143.700 135.600 144.030 136.690 ;
        RECT 144.400 136.220 145.440 136.390 ;
        RECT 144.400 135.780 145.440 135.950 ;
        RECT 145.610 135.920 145.780 136.250 ;
        RECT 143.860 135.380 144.030 135.600 ;
        RECT 146.120 135.380 146.290 136.790 ;
        RECT 143.860 135.210 146.290 135.380 ;
        RECT 147.870 137.300 158.500 137.470 ;
        RECT 127.840 135.010 138.470 135.040 ;
        RECT 147.870 135.040 148.040 137.300 ;
        RECT 148.765 136.730 156.805 136.900 ;
        RECT 148.380 135.670 148.550 136.670 ;
        RECT 157.020 135.670 157.190 136.670 ;
        RECT 148.765 135.440 156.805 135.610 ;
        RECT 157.530 135.040 158.500 137.300 ;
        RECT 147.870 135.010 158.500 135.040 ;
        RECT 107.930 134.900 118.590 135.010 ;
        RECT 127.810 134.900 138.470 135.010 ;
        RECT 147.840 134.900 158.500 135.010 ;
        RECT 106.180 134.850 118.590 134.900 ;
        RECT 126.060 134.850 138.470 134.900 ;
        RECT 146.090 134.850 158.500 134.900 ;
        RECT 76.895 133.955 82.240 134.500 ;
        RECT 82.415 133.955 87.760 134.500 ;
        RECT 87.935 133.955 89.145 134.705 ;
        RECT 89.315 133.955 90.525 134.705 ;
        RECT 101.840 134.680 118.590 134.850 ;
        RECT 11.950 133.785 90.610 133.955 ;
        RECT 12.035 133.035 13.245 133.785 ;
        RECT 13.415 133.240 18.760 133.785 ;
        RECT 18.935 133.240 24.280 133.785 ;
        RECT 12.035 132.495 12.555 133.035 ;
        RECT 12.725 132.325 13.245 132.865 ;
        RECT 15.000 132.410 15.340 133.240 ;
        RECT 12.035 131.235 13.245 132.325 ;
        RECT 16.820 131.670 17.170 132.920 ;
        RECT 20.520 132.410 20.860 133.240 ;
        RECT 24.455 133.035 25.665 133.785 ;
        RECT 25.835 133.135 26.095 133.615 ;
        RECT 26.265 133.325 26.595 133.785 ;
        RECT 26.785 133.145 26.985 133.565 ;
        RECT 22.340 131.670 22.690 132.920 ;
        RECT 24.455 132.495 24.975 133.035 ;
        RECT 25.145 132.325 25.665 132.865 ;
        RECT 13.415 131.235 18.760 131.670 ;
        RECT 18.935 131.235 24.280 131.670 ;
        RECT 24.455 131.235 25.665 132.325 ;
        RECT 25.835 132.105 26.005 133.135 ;
        RECT 26.175 132.445 26.405 132.875 ;
        RECT 26.575 132.625 26.985 133.145 ;
        RECT 27.155 133.300 27.945 133.565 ;
        RECT 27.155 132.445 27.410 133.300 ;
        RECT 28.125 132.965 28.455 133.385 ;
        RECT 28.625 132.965 28.885 133.785 ;
        RECT 29.630 133.155 29.915 133.615 ;
        RECT 30.085 133.325 30.355 133.785 ;
        RECT 29.630 132.985 30.585 133.155 ;
        RECT 28.125 132.875 28.375 132.965 ;
        RECT 27.580 132.625 28.375 132.875 ;
        RECT 26.175 132.275 27.965 132.445 ;
        RECT 25.835 131.405 26.110 132.105 ;
        RECT 26.280 131.980 26.995 132.275 ;
        RECT 27.215 131.915 27.545 132.105 ;
        RECT 26.320 131.235 26.535 131.780 ;
        RECT 26.705 131.405 27.180 131.745 ;
        RECT 27.350 131.740 27.545 131.915 ;
        RECT 27.715 131.910 27.965 132.275 ;
        RECT 27.350 131.235 27.965 131.740 ;
        RECT 28.205 131.405 28.375 132.625 ;
        RECT 28.545 131.915 28.885 132.795 ;
        RECT 29.515 132.255 30.205 132.815 ;
        RECT 30.375 132.085 30.585 132.985 ;
        RECT 29.630 131.865 30.585 132.085 ;
        RECT 30.755 132.815 31.155 133.615 ;
        RECT 31.345 133.155 31.625 133.615 ;
        RECT 32.145 133.325 32.470 133.785 ;
        RECT 31.345 132.985 32.470 133.155 ;
        RECT 32.640 133.045 33.025 133.615 ;
        RECT 32.020 132.875 32.470 132.985 ;
        RECT 30.755 132.255 31.850 132.815 ;
        RECT 32.020 132.545 32.575 132.875 ;
        RECT 28.625 131.235 28.885 131.745 ;
        RECT 29.630 131.405 29.915 131.865 ;
        RECT 30.085 131.235 30.355 131.695 ;
        RECT 30.755 131.405 31.155 132.255 ;
        RECT 32.020 132.085 32.470 132.545 ;
        RECT 32.745 132.375 33.025 133.045 ;
        RECT 34.230 133.155 34.515 133.615 ;
        RECT 34.685 133.325 34.955 133.785 ;
        RECT 34.230 132.985 35.185 133.155 ;
        RECT 31.345 131.865 32.470 132.085 ;
        RECT 31.345 131.405 31.625 131.865 ;
        RECT 32.145 131.235 32.470 131.695 ;
        RECT 32.640 131.405 33.025 132.375 ;
        RECT 34.115 132.255 34.805 132.815 ;
        RECT 34.975 132.085 35.185 132.985 ;
        RECT 34.230 131.865 35.185 132.085 ;
        RECT 35.355 132.815 35.755 133.615 ;
        RECT 35.945 133.155 36.225 133.615 ;
        RECT 36.745 133.325 37.070 133.785 ;
        RECT 35.945 132.985 37.070 133.155 ;
        RECT 37.240 133.045 37.625 133.615 ;
        RECT 37.795 133.060 38.085 133.785 ;
        RECT 38.280 133.395 38.610 133.785 ;
        RECT 38.780 133.225 39.005 133.605 ;
        RECT 36.620 132.875 37.070 132.985 ;
        RECT 35.355 132.255 36.450 132.815 ;
        RECT 36.620 132.545 37.175 132.875 ;
        RECT 34.230 131.405 34.515 131.865 ;
        RECT 34.685 131.235 34.955 131.695 ;
        RECT 35.355 131.405 35.755 132.255 ;
        RECT 36.620 132.085 37.070 132.545 ;
        RECT 37.345 132.375 37.625 133.045 ;
        RECT 38.265 132.545 38.505 133.195 ;
        RECT 38.675 133.045 39.005 133.225 ;
        RECT 35.945 131.865 37.070 132.085 ;
        RECT 35.945 131.405 36.225 131.865 ;
        RECT 36.745 131.235 37.070 131.695 ;
        RECT 37.240 131.405 37.625 132.375 ;
        RECT 37.795 131.235 38.085 132.400 ;
        RECT 38.675 132.375 38.850 133.045 ;
        RECT 39.205 132.875 39.435 133.495 ;
        RECT 39.615 133.055 39.915 133.785 ;
        RECT 40.095 133.035 41.305 133.785 ;
        RECT 41.475 133.045 41.860 133.615 ;
        RECT 42.030 133.325 42.355 133.785 ;
        RECT 42.875 133.155 43.155 133.615 ;
        RECT 39.020 132.545 39.435 132.875 ;
        RECT 39.615 132.545 39.910 132.875 ;
        RECT 40.095 132.495 40.615 133.035 ;
        RECT 38.265 132.185 38.850 132.375 ;
        RECT 38.265 131.415 38.540 132.185 ;
        RECT 39.020 132.015 39.915 132.345 ;
        RECT 40.785 132.325 41.305 132.865 ;
        RECT 38.710 131.845 39.915 132.015 ;
        RECT 38.710 131.415 39.040 131.845 ;
        RECT 39.210 131.235 39.405 131.675 ;
        RECT 39.585 131.415 39.915 131.845 ;
        RECT 40.095 131.235 41.305 132.325 ;
        RECT 41.475 132.375 41.755 133.045 ;
        RECT 42.030 132.985 43.155 133.155 ;
        RECT 42.030 132.875 42.480 132.985 ;
        RECT 41.925 132.545 42.480 132.875 ;
        RECT 43.345 132.815 43.745 133.615 ;
        RECT 44.145 133.325 44.415 133.785 ;
        RECT 44.585 133.155 44.870 133.615 ;
        RECT 41.475 131.405 41.860 132.375 ;
        RECT 42.030 132.085 42.480 132.545 ;
        RECT 42.650 132.255 43.745 132.815 ;
        RECT 42.030 131.865 43.155 132.085 ;
        RECT 42.030 131.235 42.355 131.695 ;
        RECT 42.875 131.405 43.155 131.865 ;
        RECT 43.345 131.405 43.745 132.255 ;
        RECT 43.915 132.985 44.870 133.155 ;
        RECT 45.155 132.985 45.850 133.615 ;
        RECT 46.055 132.985 46.365 133.785 ;
        RECT 47.505 133.395 47.835 133.785 ;
        RECT 48.005 133.215 48.175 133.535 ;
        RECT 48.345 133.395 48.675 133.785 ;
        RECT 49.090 133.385 50.045 133.555 ;
        RECT 47.455 133.045 49.705 133.215 ;
        RECT 43.915 132.085 44.125 132.985 ;
        RECT 44.295 132.255 44.985 132.815 ;
        RECT 45.175 132.545 45.510 132.795 ;
        RECT 45.680 132.385 45.850 132.985 ;
        RECT 46.020 132.545 46.355 132.815 ;
        RECT 43.915 131.865 44.870 132.085 ;
        RECT 44.145 131.235 44.415 131.695 ;
        RECT 44.585 131.405 44.870 131.865 ;
        RECT 45.155 131.235 45.415 132.375 ;
        RECT 45.585 131.405 45.915 132.385 ;
        RECT 46.085 131.235 46.365 132.375 ;
        RECT 47.455 132.085 47.625 133.045 ;
        RECT 47.795 132.425 48.040 132.875 ;
        RECT 48.210 132.595 48.760 132.795 ;
        RECT 48.930 132.625 49.305 132.795 ;
        RECT 48.930 132.425 49.100 132.625 ;
        RECT 49.475 132.545 49.705 133.045 ;
        RECT 47.795 132.255 49.100 132.425 ;
        RECT 49.875 132.505 50.045 133.385 ;
        RECT 50.215 132.950 50.505 133.785 ;
        RECT 50.760 133.215 50.935 133.615 ;
        RECT 51.105 133.405 51.435 133.785 ;
        RECT 51.680 133.285 51.910 133.615 ;
        RECT 50.760 133.045 51.390 133.215 ;
        RECT 51.220 132.875 51.390 133.045 ;
        RECT 49.875 132.335 50.505 132.505 ;
        RECT 47.455 131.405 47.835 132.085 ;
        RECT 48.425 131.235 48.595 132.085 ;
        RECT 48.765 131.915 50.005 132.085 ;
        RECT 48.765 131.405 49.095 131.915 ;
        RECT 49.265 131.235 49.435 131.745 ;
        RECT 49.605 131.405 50.005 131.915 ;
        RECT 50.185 131.405 50.505 132.335 ;
        RECT 50.675 132.195 51.040 132.875 ;
        RECT 51.220 132.545 51.570 132.875 ;
        RECT 51.220 132.025 51.390 132.545 ;
        RECT 50.760 131.855 51.390 132.025 ;
        RECT 51.740 131.995 51.910 133.285 ;
        RECT 52.110 132.175 52.390 133.450 ;
        RECT 52.615 133.445 52.885 133.450 ;
        RECT 52.575 133.275 52.885 133.445 ;
        RECT 53.345 133.405 53.675 133.785 ;
        RECT 53.845 133.530 54.180 133.575 ;
        RECT 52.615 132.175 52.885 133.275 ;
        RECT 53.075 132.175 53.415 133.205 ;
        RECT 53.845 133.065 54.185 133.530 ;
        RECT 53.585 132.545 53.845 132.875 ;
        RECT 53.585 131.995 53.755 132.545 ;
        RECT 54.015 132.375 54.185 133.065 ;
        RECT 54.355 133.015 56.025 133.785 ;
        RECT 56.285 133.235 56.455 133.525 ;
        RECT 56.625 133.405 56.955 133.785 ;
        RECT 56.285 133.065 56.950 133.235 ;
        RECT 54.355 132.495 55.105 133.015 ;
        RECT 50.760 131.405 50.935 131.855 ;
        RECT 51.740 131.825 53.755 131.995 ;
        RECT 51.105 131.235 51.435 131.675 ;
        RECT 51.740 131.405 51.910 131.825 ;
        RECT 52.145 131.235 52.815 131.645 ;
        RECT 53.030 131.405 53.200 131.825 ;
        RECT 53.400 131.235 53.730 131.645 ;
        RECT 53.925 131.405 54.185 132.375 ;
        RECT 55.275 132.325 56.025 132.845 ;
        RECT 54.355 131.235 56.025 132.325 ;
        RECT 56.200 132.245 56.550 132.895 ;
        RECT 56.720 132.075 56.950 133.065 ;
        RECT 56.285 131.905 56.950 132.075 ;
        RECT 56.285 131.405 56.455 131.905 ;
        RECT 56.625 131.235 56.955 131.735 ;
        RECT 57.125 131.405 57.310 133.525 ;
        RECT 57.565 133.325 57.815 133.785 ;
        RECT 57.985 133.335 58.320 133.505 ;
        RECT 58.515 133.335 59.190 133.505 ;
        RECT 57.985 133.195 58.155 133.335 ;
        RECT 57.480 132.205 57.760 133.155 ;
        RECT 57.930 133.065 58.155 133.195 ;
        RECT 57.930 131.960 58.100 133.065 ;
        RECT 58.325 132.915 58.850 133.135 ;
        RECT 58.270 132.150 58.510 132.745 ;
        RECT 58.680 132.215 58.850 132.915 ;
        RECT 59.020 132.555 59.190 133.335 ;
        RECT 59.510 133.285 59.880 133.785 ;
        RECT 60.060 133.335 60.465 133.505 ;
        RECT 60.635 133.335 61.420 133.505 ;
        RECT 60.060 133.105 60.230 133.335 ;
        RECT 59.400 132.805 60.230 133.105 ;
        RECT 60.615 132.835 61.080 133.165 ;
        RECT 59.400 132.775 59.600 132.805 ;
        RECT 59.720 132.555 59.890 132.625 ;
        RECT 59.020 132.385 59.890 132.555 ;
        RECT 59.380 132.295 59.890 132.385 ;
        RECT 57.930 131.830 58.235 131.960 ;
        RECT 58.680 131.850 59.210 132.215 ;
        RECT 57.550 131.235 57.815 131.695 ;
        RECT 57.985 131.405 58.235 131.830 ;
        RECT 59.380 131.680 59.550 132.295 ;
        RECT 58.445 131.510 59.550 131.680 ;
        RECT 59.720 131.235 59.890 132.035 ;
        RECT 60.060 131.735 60.230 132.805 ;
        RECT 60.400 131.905 60.590 132.625 ;
        RECT 60.760 131.875 61.080 132.835 ;
        RECT 61.250 132.875 61.420 133.335 ;
        RECT 61.695 133.255 61.905 133.785 ;
        RECT 62.165 133.045 62.495 133.570 ;
        RECT 62.665 133.175 62.835 133.785 ;
        RECT 63.005 133.130 63.335 133.565 ;
        RECT 63.005 133.045 63.385 133.130 ;
        RECT 63.555 133.060 63.845 133.785 ;
        RECT 65.025 133.235 65.195 133.525 ;
        RECT 65.365 133.405 65.695 133.785 ;
        RECT 65.025 133.065 65.690 133.235 ;
        RECT 62.295 132.875 62.495 133.045 ;
        RECT 63.160 133.005 63.385 133.045 ;
        RECT 61.250 132.545 62.125 132.875 ;
        RECT 62.295 132.545 63.045 132.875 ;
        RECT 60.060 131.405 60.310 131.735 ;
        RECT 61.250 131.705 61.420 132.545 ;
        RECT 62.295 132.340 62.485 132.545 ;
        RECT 63.215 132.425 63.385 133.005 ;
        RECT 63.170 132.375 63.385 132.425 ;
        RECT 61.590 131.965 62.485 132.340 ;
        RECT 62.995 132.295 63.385 132.375 ;
        RECT 60.535 131.535 61.420 131.705 ;
        RECT 61.600 131.235 61.915 131.735 ;
        RECT 62.145 131.405 62.485 131.965 ;
        RECT 62.655 131.235 62.825 132.245 ;
        RECT 62.995 131.450 63.325 132.295 ;
        RECT 63.555 131.235 63.845 132.400 ;
        RECT 64.940 132.245 65.290 132.895 ;
        RECT 65.460 132.075 65.690 133.065 ;
        RECT 65.025 131.905 65.690 132.075 ;
        RECT 65.025 131.405 65.195 131.905 ;
        RECT 65.365 131.235 65.695 131.735 ;
        RECT 65.865 131.405 66.050 133.525 ;
        RECT 66.305 133.325 66.555 133.785 ;
        RECT 66.725 133.335 67.060 133.505 ;
        RECT 67.255 133.335 67.930 133.505 ;
        RECT 66.725 133.195 66.895 133.335 ;
        RECT 66.220 132.205 66.500 133.155 ;
        RECT 66.670 133.065 66.895 133.195 ;
        RECT 66.670 131.960 66.840 133.065 ;
        RECT 67.065 132.915 67.590 133.135 ;
        RECT 67.010 132.150 67.250 132.745 ;
        RECT 67.420 132.215 67.590 132.915 ;
        RECT 67.760 132.555 67.930 133.335 ;
        RECT 68.250 133.285 68.620 133.785 ;
        RECT 68.800 133.335 69.205 133.505 ;
        RECT 69.375 133.335 70.160 133.505 ;
        RECT 68.800 133.105 68.970 133.335 ;
        RECT 68.140 132.805 68.970 133.105 ;
        RECT 69.355 132.835 69.820 133.165 ;
        RECT 68.140 132.775 68.340 132.805 ;
        RECT 68.460 132.555 68.630 132.625 ;
        RECT 67.760 132.385 68.630 132.555 ;
        RECT 68.120 132.295 68.630 132.385 ;
        RECT 66.670 131.830 66.975 131.960 ;
        RECT 67.420 131.850 67.950 132.215 ;
        RECT 66.290 131.235 66.555 131.695 ;
        RECT 66.725 131.405 66.975 131.830 ;
        RECT 68.120 131.680 68.290 132.295 ;
        RECT 67.185 131.510 68.290 131.680 ;
        RECT 68.460 131.235 68.630 132.035 ;
        RECT 68.800 131.735 68.970 132.805 ;
        RECT 69.140 131.905 69.330 132.625 ;
        RECT 69.500 131.875 69.820 132.835 ;
        RECT 69.990 132.875 70.160 133.335 ;
        RECT 70.435 133.255 70.645 133.785 ;
        RECT 70.905 133.045 71.235 133.570 ;
        RECT 71.405 133.175 71.575 133.785 ;
        RECT 71.745 133.130 72.075 133.565 ;
        RECT 72.295 133.240 77.640 133.785 ;
        RECT 77.815 133.240 83.160 133.785 ;
        RECT 83.335 133.240 88.680 133.785 ;
        RECT 71.745 133.045 72.125 133.130 ;
        RECT 71.035 132.875 71.235 133.045 ;
        RECT 71.900 133.005 72.125 133.045 ;
        RECT 69.990 132.545 70.865 132.875 ;
        RECT 71.035 132.545 71.785 132.875 ;
        RECT 68.800 131.405 69.050 131.735 ;
        RECT 69.990 131.705 70.160 132.545 ;
        RECT 71.035 132.340 71.225 132.545 ;
        RECT 71.955 132.425 72.125 133.005 ;
        RECT 71.910 132.375 72.125 132.425 ;
        RECT 73.880 132.410 74.220 133.240 ;
        RECT 70.330 131.965 71.225 132.340 ;
        RECT 71.735 132.295 72.125 132.375 ;
        RECT 69.275 131.535 70.160 131.705 ;
        RECT 70.340 131.235 70.655 131.735 ;
        RECT 70.885 131.405 71.225 131.965 ;
        RECT 71.395 131.235 71.565 132.245 ;
        RECT 71.735 131.450 72.065 132.295 ;
        RECT 75.700 131.670 76.050 132.920 ;
        RECT 79.400 132.410 79.740 133.240 ;
        RECT 81.220 131.670 81.570 132.920 ;
        RECT 84.920 132.410 85.260 133.240 ;
        RECT 89.315 133.035 90.525 133.785 ;
        RECT 101.840 133.270 102.010 134.680 ;
        RECT 102.380 134.110 105.420 134.280 ;
        RECT 102.380 133.670 105.420 133.840 ;
        RECT 105.635 133.810 105.805 134.140 ;
        RECT 106.140 133.920 118.590 134.680 ;
        RECT 121.720 134.680 138.470 134.850 ;
        RECT 106.140 133.910 118.480 133.920 ;
        RECT 106.140 133.900 112.020 133.910 ;
        RECT 106.140 133.880 106.710 133.900 ;
        RECT 107.930 133.890 112.020 133.900 ;
        RECT 106.150 133.270 106.320 133.880 ;
        RECT 101.840 133.100 106.320 133.270 ;
        RECT 121.720 133.270 121.890 134.680 ;
        RECT 122.260 134.110 125.300 134.280 ;
        RECT 122.260 133.670 125.300 133.840 ;
        RECT 125.515 133.810 125.685 134.140 ;
        RECT 126.020 133.920 138.470 134.680 ;
        RECT 141.750 134.680 158.500 134.850 ;
        RECT 126.020 133.910 138.360 133.920 ;
        RECT 126.020 133.900 131.900 133.910 ;
        RECT 126.020 133.880 126.590 133.900 ;
        RECT 127.810 133.890 131.900 133.900 ;
        RECT 126.030 133.270 126.200 133.880 ;
        RECT 121.720 133.100 126.200 133.270 ;
        RECT 141.750 133.270 141.920 134.680 ;
        RECT 142.290 134.110 145.330 134.280 ;
        RECT 142.290 133.670 145.330 133.840 ;
        RECT 145.545 133.810 145.715 134.140 ;
        RECT 146.050 133.920 158.500 134.680 ;
        RECT 146.050 133.910 158.390 133.920 ;
        RECT 146.050 133.900 151.930 133.910 ;
        RECT 146.050 133.880 146.620 133.900 ;
        RECT 147.840 133.890 151.930 133.900 ;
        RECT 146.060 133.270 146.230 133.880 ;
        RECT 141.750 133.100 146.230 133.270 ;
        RECT 86.740 131.670 87.090 132.920 ;
        RECT 89.315 132.325 89.835 132.865 ;
        RECT 90.005 132.495 90.525 133.035 ;
        RECT 72.295 131.235 77.640 131.670 ;
        RECT 77.815 131.235 83.160 131.670 ;
        RECT 83.335 131.235 88.680 131.670 ;
        RECT 89.315 131.235 90.525 132.325 ;
        RECT 120.510 131.800 126.250 131.810 ;
        RECT 100.630 131.740 106.370 131.750 ;
        RECT 100.140 131.580 106.370 131.740 ;
        RECT 11.950 131.065 90.610 131.235 ;
        RECT 12.035 129.975 13.245 131.065 ;
        RECT 13.415 130.630 18.760 131.065 ;
        RECT 18.935 130.630 24.280 131.065 ;
        RECT 12.035 129.265 12.555 129.805 ;
        RECT 12.725 129.435 13.245 129.975 ;
        RECT 12.035 128.515 13.245 129.265 ;
        RECT 15.000 129.060 15.340 129.890 ;
        RECT 16.820 129.380 17.170 130.630 ;
        RECT 20.520 129.060 20.860 129.890 ;
        RECT 22.340 129.380 22.690 130.630 ;
        RECT 24.915 129.900 25.205 131.065 ;
        RECT 25.435 130.005 25.765 130.850 ;
        RECT 25.935 130.055 26.105 131.065 ;
        RECT 26.275 130.335 26.615 130.895 ;
        RECT 26.845 130.565 27.160 131.065 ;
        RECT 27.340 130.595 28.225 130.765 ;
        RECT 25.375 129.925 25.765 130.005 ;
        RECT 26.275 129.960 27.170 130.335 ;
        RECT 25.375 129.875 25.590 129.925 ;
        RECT 25.375 129.295 25.545 129.875 ;
        RECT 26.275 129.755 26.465 129.960 ;
        RECT 27.340 129.755 27.510 130.595 ;
        RECT 28.450 130.565 28.700 130.895 ;
        RECT 25.715 129.425 26.465 129.755 ;
        RECT 26.635 129.425 27.510 129.755 ;
        RECT 25.375 129.255 25.600 129.295 ;
        RECT 26.265 129.255 26.465 129.425 ;
        RECT 13.415 128.515 18.760 129.060 ;
        RECT 18.935 128.515 24.280 129.060 ;
        RECT 24.915 128.515 25.205 129.240 ;
        RECT 25.375 129.170 25.755 129.255 ;
        RECT 25.425 128.735 25.755 129.170 ;
        RECT 25.925 128.515 26.095 129.125 ;
        RECT 26.265 128.730 26.595 129.255 ;
        RECT 26.855 128.515 27.065 129.045 ;
        RECT 27.340 128.965 27.510 129.425 ;
        RECT 27.680 129.465 28.000 130.425 ;
        RECT 28.170 129.675 28.360 130.395 ;
        RECT 28.530 129.495 28.700 130.565 ;
        RECT 28.870 130.265 29.040 131.065 ;
        RECT 29.210 130.620 30.315 130.790 ;
        RECT 29.210 130.005 29.380 130.620 ;
        RECT 30.525 130.470 30.775 130.895 ;
        RECT 30.945 130.605 31.210 131.065 ;
        RECT 29.550 130.085 30.080 130.450 ;
        RECT 30.525 130.340 30.830 130.470 ;
        RECT 28.870 129.915 29.380 130.005 ;
        RECT 28.870 129.745 29.740 129.915 ;
        RECT 28.870 129.675 29.040 129.745 ;
        RECT 29.160 129.495 29.360 129.525 ;
        RECT 27.680 129.135 28.145 129.465 ;
        RECT 28.530 129.195 29.360 129.495 ;
        RECT 28.530 128.965 28.700 129.195 ;
        RECT 27.340 128.795 28.125 128.965 ;
        RECT 28.295 128.795 28.700 128.965 ;
        RECT 28.880 128.515 29.250 129.015 ;
        RECT 29.570 128.965 29.740 129.745 ;
        RECT 29.910 129.385 30.080 130.085 ;
        RECT 30.250 129.555 30.490 130.150 ;
        RECT 29.910 129.165 30.435 129.385 ;
        RECT 30.660 129.235 30.830 130.340 ;
        RECT 30.605 129.105 30.830 129.235 ;
        RECT 31.000 129.145 31.280 130.095 ;
        RECT 30.605 128.965 30.775 129.105 ;
        RECT 29.570 128.795 30.245 128.965 ;
        RECT 30.440 128.795 30.775 128.965 ;
        RECT 30.945 128.515 31.195 128.975 ;
        RECT 31.450 128.775 31.635 130.895 ;
        RECT 31.805 130.565 32.135 131.065 ;
        RECT 32.305 130.395 32.475 130.895 ;
        RECT 31.810 130.225 32.475 130.395 ;
        RECT 32.770 130.275 33.305 130.895 ;
        RECT 31.810 129.235 32.040 130.225 ;
        RECT 32.210 129.405 32.560 130.055 ;
        RECT 32.770 129.255 33.085 130.275 ;
        RECT 33.475 130.265 33.805 131.065 ;
        RECT 35.125 130.395 35.295 130.895 ;
        RECT 35.465 130.565 35.795 131.065 ;
        RECT 34.290 130.095 34.680 130.270 ;
        RECT 35.125 130.225 35.790 130.395 ;
        RECT 33.255 129.925 34.680 130.095 ;
        RECT 33.255 129.425 33.425 129.925 ;
        RECT 31.810 129.065 32.475 129.235 ;
        RECT 31.805 128.515 32.135 128.895 ;
        RECT 32.305 128.775 32.475 129.065 ;
        RECT 32.770 128.685 33.385 129.255 ;
        RECT 33.675 129.195 33.940 129.755 ;
        RECT 34.110 129.025 34.280 129.925 ;
        RECT 34.450 129.195 34.805 129.755 ;
        RECT 35.040 129.405 35.390 130.055 ;
        RECT 35.560 129.235 35.790 130.225 ;
        RECT 35.125 129.065 35.790 129.235 ;
        RECT 33.555 128.515 33.770 129.025 ;
        RECT 34.000 128.695 34.280 129.025 ;
        RECT 34.460 128.515 34.700 129.025 ;
        RECT 35.125 128.775 35.295 129.065 ;
        RECT 35.465 128.515 35.795 128.895 ;
        RECT 35.965 128.775 36.150 130.895 ;
        RECT 36.390 130.605 36.655 131.065 ;
        RECT 36.825 130.470 37.075 130.895 ;
        RECT 37.285 130.620 38.390 130.790 ;
        RECT 36.770 130.340 37.075 130.470 ;
        RECT 36.320 129.145 36.600 130.095 ;
        RECT 36.770 129.235 36.940 130.340 ;
        RECT 37.110 129.555 37.350 130.150 ;
        RECT 37.520 130.085 38.050 130.450 ;
        RECT 37.520 129.385 37.690 130.085 ;
        RECT 38.220 130.005 38.390 130.620 ;
        RECT 38.560 130.265 38.730 131.065 ;
        RECT 38.900 130.565 39.150 130.895 ;
        RECT 39.375 130.595 40.260 130.765 ;
        RECT 38.220 129.915 38.730 130.005 ;
        RECT 36.770 129.105 36.995 129.235 ;
        RECT 37.165 129.165 37.690 129.385 ;
        RECT 37.860 129.745 38.730 129.915 ;
        RECT 36.405 128.515 36.655 128.975 ;
        RECT 36.825 128.965 36.995 129.105 ;
        RECT 37.860 128.965 38.030 129.745 ;
        RECT 38.560 129.675 38.730 129.745 ;
        RECT 38.240 129.495 38.440 129.525 ;
        RECT 38.900 129.495 39.070 130.565 ;
        RECT 39.240 129.675 39.430 130.395 ;
        RECT 38.240 129.195 39.070 129.495 ;
        RECT 39.600 129.465 39.920 130.425 ;
        RECT 36.825 128.795 37.160 128.965 ;
        RECT 37.355 128.795 38.030 128.965 ;
        RECT 38.350 128.515 38.720 129.015 ;
        RECT 38.900 128.965 39.070 129.195 ;
        RECT 39.455 129.135 39.920 129.465 ;
        RECT 40.090 129.755 40.260 130.595 ;
        RECT 40.440 130.565 40.755 131.065 ;
        RECT 40.985 130.335 41.325 130.895 ;
        RECT 40.430 129.960 41.325 130.335 ;
        RECT 41.495 130.055 41.665 131.065 ;
        RECT 41.135 129.755 41.325 129.960 ;
        RECT 41.835 130.005 42.165 130.850 ;
        RECT 42.475 130.435 42.655 130.895 ;
        RECT 42.825 130.605 43.075 131.065 ;
        RECT 43.245 130.685 43.575 130.855 ;
        RECT 43.745 130.800 44.000 130.895 ;
        RECT 43.245 130.435 43.415 130.685 ;
        RECT 43.745 130.630 44.885 130.800 ;
        RECT 45.145 130.665 45.475 131.065 ;
        RECT 43.745 130.495 44.000 130.630 ;
        RECT 42.475 130.265 43.415 130.435 ;
        RECT 43.590 130.325 44.000 130.495 ;
        RECT 44.715 130.405 44.885 130.630 ;
        RECT 41.835 129.925 42.225 130.005 ;
        RECT 42.010 129.875 42.225 129.925 ;
        RECT 40.090 129.425 40.965 129.755 ;
        RECT 41.135 129.425 41.885 129.755 ;
        RECT 40.090 128.965 40.260 129.425 ;
        RECT 41.135 129.255 41.335 129.425 ;
        RECT 42.055 129.295 42.225 129.875 ;
        RECT 42.000 129.255 42.225 129.295 ;
        RECT 38.900 128.795 39.305 128.965 ;
        RECT 39.475 128.795 40.260 128.965 ;
        RECT 40.535 128.515 40.745 129.045 ;
        RECT 41.005 128.730 41.335 129.255 ;
        RECT 41.845 129.170 42.225 129.255 ;
        RECT 42.450 129.195 42.710 130.085 ;
        RECT 42.910 129.785 43.390 130.085 ;
        RECT 42.910 129.195 43.170 129.785 ;
        RECT 43.590 129.300 43.760 130.325 ;
        RECT 44.280 130.145 44.450 130.335 ;
        RECT 44.715 130.235 45.475 130.405 ;
        RECT 41.505 128.515 41.675 129.125 ;
        RECT 41.845 128.735 42.175 129.170 ;
        RECT 43.410 129.130 43.760 129.300 ;
        RECT 43.930 129.975 44.450 130.145 ;
        RECT 43.930 129.255 44.100 129.975 ;
        RECT 44.290 129.425 44.580 129.805 ;
        RECT 44.750 129.425 45.080 130.045 ;
        RECT 45.305 129.755 45.475 130.235 ;
        RECT 45.645 129.955 45.905 130.895 ;
        RECT 45.305 129.425 45.560 129.755 ;
        RECT 42.435 128.515 42.835 129.025 ;
        RECT 43.410 128.685 43.580 129.130 ;
        RECT 43.930 129.085 44.810 129.255 ;
        RECT 45.730 129.240 45.905 129.955 ;
        RECT 43.750 128.515 44.470 128.915 ;
        RECT 44.640 128.685 44.810 129.085 ;
        RECT 45.045 128.515 45.475 128.960 ;
        RECT 45.645 128.685 45.905 129.240 ;
        RECT 46.075 129.925 46.460 130.895 ;
        RECT 46.630 130.605 46.955 131.065 ;
        RECT 47.475 130.435 47.755 130.895 ;
        RECT 46.630 130.215 47.755 130.435 ;
        RECT 46.075 129.255 46.355 129.925 ;
        RECT 46.630 129.755 47.080 130.215 ;
        RECT 47.945 130.045 48.345 130.895 ;
        RECT 48.745 130.605 49.015 131.065 ;
        RECT 49.185 130.435 49.470 130.895 ;
        RECT 46.525 129.425 47.080 129.755 ;
        RECT 47.250 129.485 48.345 130.045 ;
        RECT 46.630 129.315 47.080 129.425 ;
        RECT 46.075 128.685 46.460 129.255 ;
        RECT 46.630 129.145 47.755 129.315 ;
        RECT 46.630 128.515 46.955 128.975 ;
        RECT 47.475 128.685 47.755 129.145 ;
        RECT 47.945 128.685 48.345 129.485 ;
        RECT 48.515 130.215 49.470 130.435 ;
        RECT 48.515 129.315 48.725 130.215 ;
        RECT 48.895 129.485 49.585 130.045 ;
        RECT 50.675 129.900 50.965 131.065 ;
        RECT 51.135 129.925 51.395 131.065 ;
        RECT 51.565 129.915 51.895 130.895 ;
        RECT 52.065 129.925 52.345 131.065 ;
        RECT 52.605 130.395 52.775 130.895 ;
        RECT 52.945 130.565 53.275 131.065 ;
        RECT 52.605 130.225 53.270 130.395 ;
        RECT 51.155 129.505 51.490 129.755 ;
        RECT 51.660 129.315 51.830 129.915 ;
        RECT 52.000 129.485 52.335 129.755 ;
        RECT 52.520 129.405 52.870 130.055 ;
        RECT 48.515 129.145 49.470 129.315 ;
        RECT 48.745 128.515 49.015 128.975 ;
        RECT 49.185 128.685 49.470 129.145 ;
        RECT 50.675 128.515 50.965 129.240 ;
        RECT 51.135 128.685 51.830 129.315 ;
        RECT 52.035 128.515 52.345 129.315 ;
        RECT 53.040 129.235 53.270 130.225 ;
        RECT 52.605 129.065 53.270 129.235 ;
        RECT 52.605 128.775 52.775 129.065 ;
        RECT 52.945 128.515 53.275 128.895 ;
        RECT 53.445 128.775 53.630 130.895 ;
        RECT 53.870 130.605 54.135 131.065 ;
        RECT 54.305 130.470 54.555 130.895 ;
        RECT 54.765 130.620 55.870 130.790 ;
        RECT 54.250 130.340 54.555 130.470 ;
        RECT 53.800 129.145 54.080 130.095 ;
        RECT 54.250 129.235 54.420 130.340 ;
        RECT 54.590 129.555 54.830 130.150 ;
        RECT 55.000 130.085 55.530 130.450 ;
        RECT 55.000 129.385 55.170 130.085 ;
        RECT 55.700 130.005 55.870 130.620 ;
        RECT 56.040 130.265 56.210 131.065 ;
        RECT 56.380 130.565 56.630 130.895 ;
        RECT 56.855 130.595 57.740 130.765 ;
        RECT 55.700 129.915 56.210 130.005 ;
        RECT 54.250 129.105 54.475 129.235 ;
        RECT 54.645 129.165 55.170 129.385 ;
        RECT 55.340 129.745 56.210 129.915 ;
        RECT 53.885 128.515 54.135 128.975 ;
        RECT 54.305 128.965 54.475 129.105 ;
        RECT 55.340 128.965 55.510 129.745 ;
        RECT 56.040 129.675 56.210 129.745 ;
        RECT 55.720 129.495 55.920 129.525 ;
        RECT 56.380 129.495 56.550 130.565 ;
        RECT 56.720 129.675 56.910 130.395 ;
        RECT 55.720 129.195 56.550 129.495 ;
        RECT 57.080 129.465 57.400 130.425 ;
        RECT 54.305 128.795 54.640 128.965 ;
        RECT 54.835 128.795 55.510 128.965 ;
        RECT 55.830 128.515 56.200 129.015 ;
        RECT 56.380 128.965 56.550 129.195 ;
        RECT 56.935 129.135 57.400 129.465 ;
        RECT 57.570 129.755 57.740 130.595 ;
        RECT 57.920 130.565 58.235 131.065 ;
        RECT 58.465 130.335 58.805 130.895 ;
        RECT 57.910 129.960 58.805 130.335 ;
        RECT 58.975 130.055 59.145 131.065 ;
        RECT 58.615 129.755 58.805 129.960 ;
        RECT 59.315 130.005 59.645 130.850 ;
        RECT 59.315 129.925 59.705 130.005 ;
        RECT 59.875 129.975 63.385 131.065 ;
        RECT 64.100 130.445 64.275 130.895 ;
        RECT 64.445 130.625 64.775 131.065 ;
        RECT 65.080 130.475 65.250 130.895 ;
        RECT 65.485 130.655 66.155 131.065 ;
        RECT 66.370 130.475 66.540 130.895 ;
        RECT 66.740 130.655 67.070 131.065 ;
        RECT 64.100 130.275 64.730 130.445 ;
        RECT 59.490 129.875 59.705 129.925 ;
        RECT 57.570 129.425 58.445 129.755 ;
        RECT 58.615 129.425 59.365 129.755 ;
        RECT 57.570 128.965 57.740 129.425 ;
        RECT 58.615 129.255 58.815 129.425 ;
        RECT 59.535 129.295 59.705 129.875 ;
        RECT 59.480 129.255 59.705 129.295 ;
        RECT 56.380 128.795 56.785 128.965 ;
        RECT 56.955 128.795 57.740 128.965 ;
        RECT 58.015 128.515 58.225 129.045 ;
        RECT 58.485 128.730 58.815 129.255 ;
        RECT 59.325 129.170 59.705 129.255 ;
        RECT 59.875 129.285 61.525 129.805 ;
        RECT 61.695 129.455 63.385 129.975 ;
        RECT 64.015 129.425 64.380 130.105 ;
        RECT 64.560 129.755 64.730 130.275 ;
        RECT 65.080 130.305 67.095 130.475 ;
        RECT 64.560 129.425 64.910 129.755 ;
        RECT 58.985 128.515 59.155 129.125 ;
        RECT 59.325 128.735 59.655 129.170 ;
        RECT 59.875 128.515 63.385 129.285 ;
        RECT 64.560 129.255 64.730 129.425 ;
        RECT 64.100 129.085 64.730 129.255 ;
        RECT 64.100 128.685 64.275 129.085 ;
        RECT 65.080 129.015 65.250 130.305 ;
        RECT 64.445 128.515 64.775 128.895 ;
        RECT 65.020 128.685 65.250 129.015 ;
        RECT 65.450 128.850 65.730 130.125 ;
        RECT 65.955 129.025 66.225 130.125 ;
        RECT 66.415 129.095 66.755 130.125 ;
        RECT 66.925 129.755 67.095 130.305 ;
        RECT 67.265 129.925 67.525 130.895 ;
        RECT 67.695 130.630 73.040 131.065 ;
        RECT 66.925 129.425 67.185 129.755 ;
        RECT 67.355 129.235 67.525 129.925 ;
        RECT 65.915 128.855 66.225 129.025 ;
        RECT 65.955 128.850 66.225 128.855 ;
        RECT 66.685 128.515 67.015 128.895 ;
        RECT 67.185 128.770 67.525 129.235 ;
        RECT 69.280 129.060 69.620 129.890 ;
        RECT 71.100 129.380 71.450 130.630 ;
        RECT 73.215 129.975 75.805 131.065 ;
        RECT 73.215 129.285 74.425 129.805 ;
        RECT 74.595 129.455 75.805 129.975 ;
        RECT 76.435 129.900 76.725 131.065 ;
        RECT 76.895 130.630 82.240 131.065 ;
        RECT 82.415 130.630 87.760 131.065 ;
        RECT 67.185 128.725 67.520 128.770 ;
        RECT 67.695 128.515 73.040 129.060 ;
        RECT 73.215 128.515 75.805 129.285 ;
        RECT 76.435 128.515 76.725 129.240 ;
        RECT 78.480 129.060 78.820 129.890 ;
        RECT 80.300 129.380 80.650 130.630 ;
        RECT 84.000 129.060 84.340 129.890 ;
        RECT 85.820 129.380 86.170 130.630 ;
        RECT 87.935 129.975 89.145 131.065 ;
        RECT 87.935 129.265 88.455 129.805 ;
        RECT 88.625 129.435 89.145 129.975 ;
        RECT 89.315 129.975 90.525 131.065 ;
        RECT 89.315 129.435 89.835 129.975 ;
        RECT 90.005 129.265 90.525 129.805 ;
        RECT 76.895 128.515 82.240 129.060 ;
        RECT 82.415 128.515 87.760 129.060 ;
        RECT 87.935 128.515 89.145 129.265 ;
        RECT 89.315 128.515 90.525 129.265 ;
        RECT 100.140 129.320 100.810 131.580 ;
        RECT 101.480 131.010 105.520 131.180 ;
        RECT 101.140 129.950 101.310 130.950 ;
        RECT 105.690 129.950 105.860 130.950 ;
        RECT 101.480 129.720 105.520 129.890 ;
        RECT 106.200 129.320 106.370 131.580 ;
        RECT 100.140 129.150 106.370 129.320 ;
        RECT 11.950 128.345 90.610 128.515 ;
        RECT 12.035 127.595 13.245 128.345 ;
        RECT 13.415 127.800 18.760 128.345 ;
        RECT 18.935 127.800 24.280 128.345 ;
        RECT 12.035 127.055 12.555 127.595 ;
        RECT 12.725 126.885 13.245 127.425 ;
        RECT 15.000 126.970 15.340 127.800 ;
        RECT 12.035 125.795 13.245 126.885 ;
        RECT 16.820 126.230 17.170 127.480 ;
        RECT 20.520 126.970 20.860 127.800 ;
        RECT 24.455 127.575 27.045 128.345 ;
        RECT 27.265 127.690 27.595 128.125 ;
        RECT 27.765 127.735 27.935 128.345 ;
        RECT 27.215 127.605 27.595 127.690 ;
        RECT 28.105 127.605 28.435 128.130 ;
        RECT 28.695 127.815 28.905 128.345 ;
        RECT 29.180 127.895 29.965 128.065 ;
        RECT 30.135 127.895 30.540 128.065 ;
        RECT 22.340 126.230 22.690 127.480 ;
        RECT 24.455 127.055 25.665 127.575 ;
        RECT 27.215 127.565 27.440 127.605 ;
        RECT 25.835 126.885 27.045 127.405 ;
        RECT 13.415 125.795 18.760 126.230 ;
        RECT 18.935 125.795 24.280 126.230 ;
        RECT 24.455 125.795 27.045 126.885 ;
        RECT 27.215 126.985 27.385 127.565 ;
        RECT 28.105 127.435 28.305 127.605 ;
        RECT 29.180 127.435 29.350 127.895 ;
        RECT 27.555 127.105 28.305 127.435 ;
        RECT 28.475 127.105 29.350 127.435 ;
        RECT 27.215 126.935 27.430 126.985 ;
        RECT 27.215 126.855 27.605 126.935 ;
        RECT 27.275 126.010 27.605 126.855 ;
        RECT 28.115 126.900 28.305 127.105 ;
        RECT 27.775 125.795 27.945 126.805 ;
        RECT 28.115 126.525 29.010 126.900 ;
        RECT 28.115 125.965 28.455 126.525 ;
        RECT 28.685 125.795 29.000 126.295 ;
        RECT 29.180 126.265 29.350 127.105 ;
        RECT 29.520 127.395 29.985 127.725 ;
        RECT 30.370 127.665 30.540 127.895 ;
        RECT 30.720 127.845 31.090 128.345 ;
        RECT 31.410 127.895 32.085 128.065 ;
        RECT 32.280 127.895 32.615 128.065 ;
        RECT 29.520 126.435 29.840 127.395 ;
        RECT 30.370 127.365 31.200 127.665 ;
        RECT 30.010 126.465 30.200 127.185 ;
        RECT 30.370 126.295 30.540 127.365 ;
        RECT 31.000 127.335 31.200 127.365 ;
        RECT 30.710 127.115 30.880 127.185 ;
        RECT 31.410 127.115 31.580 127.895 ;
        RECT 32.445 127.755 32.615 127.895 ;
        RECT 32.785 127.885 33.035 128.345 ;
        RECT 30.710 126.945 31.580 127.115 ;
        RECT 31.750 127.475 32.275 127.695 ;
        RECT 32.445 127.625 32.670 127.755 ;
        RECT 30.710 126.855 31.220 126.945 ;
        RECT 29.180 126.095 30.065 126.265 ;
        RECT 30.290 125.965 30.540 126.295 ;
        RECT 30.710 125.795 30.880 126.595 ;
        RECT 31.050 126.240 31.220 126.855 ;
        RECT 31.750 126.775 31.920 127.475 ;
        RECT 31.390 126.410 31.920 126.775 ;
        RECT 32.090 126.710 32.330 127.305 ;
        RECT 32.500 126.520 32.670 127.625 ;
        RECT 32.840 126.765 33.120 127.715 ;
        RECT 32.365 126.390 32.670 126.520 ;
        RECT 31.050 126.070 32.155 126.240 ;
        RECT 32.365 125.965 32.615 126.390 ;
        RECT 32.785 125.795 33.050 126.255 ;
        RECT 33.290 125.965 33.475 128.085 ;
        RECT 33.645 127.965 33.975 128.345 ;
        RECT 34.145 127.795 34.315 128.085 ;
        RECT 33.650 127.625 34.315 127.795 ;
        RECT 33.650 126.635 33.880 127.625 ;
        RECT 34.575 127.605 34.895 128.085 ;
        RECT 35.065 127.775 35.295 128.175 ;
        RECT 35.465 127.955 35.815 128.345 ;
        RECT 35.065 127.695 35.575 127.775 ;
        RECT 35.985 127.695 36.315 128.175 ;
        RECT 35.065 127.605 36.315 127.695 ;
        RECT 34.050 126.805 34.400 127.455 ;
        RECT 34.575 126.675 34.745 127.605 ;
        RECT 35.405 127.525 36.315 127.605 ;
        RECT 36.485 127.525 36.655 128.345 ;
        RECT 37.160 127.605 37.625 128.150 ;
        RECT 37.795 127.620 38.085 128.345 ;
        RECT 39.290 127.715 39.575 128.175 ;
        RECT 39.745 127.885 40.015 128.345 ;
        RECT 34.915 127.015 35.085 127.435 ;
        RECT 35.315 127.185 35.915 127.355 ;
        RECT 34.915 126.845 35.575 127.015 ;
        RECT 33.650 126.465 34.315 126.635 ;
        RECT 34.575 126.475 35.235 126.675 ;
        RECT 35.405 126.645 35.575 126.845 ;
        RECT 35.745 126.985 35.915 127.185 ;
        RECT 36.085 127.155 36.780 127.355 ;
        RECT 37.040 126.985 37.285 127.435 ;
        RECT 35.745 126.815 37.285 126.985 ;
        RECT 37.455 126.645 37.625 127.605 ;
        RECT 39.290 127.545 40.245 127.715 ;
        RECT 35.405 126.475 37.625 126.645 ;
        RECT 33.645 125.795 33.975 126.295 ;
        RECT 34.145 125.965 34.315 126.465 ;
        RECT 35.065 126.305 35.235 126.475 ;
        RECT 34.595 125.795 34.895 126.305 ;
        RECT 35.065 126.135 35.445 126.305 ;
        RECT 36.025 125.795 36.655 126.305 ;
        RECT 36.825 125.965 37.155 126.475 ;
        RECT 37.325 125.795 37.625 126.305 ;
        RECT 37.795 125.795 38.085 126.960 ;
        RECT 39.175 126.815 39.865 127.375 ;
        RECT 40.035 126.645 40.245 127.545 ;
        RECT 39.290 126.425 40.245 126.645 ;
        RECT 40.415 127.375 40.815 128.175 ;
        RECT 41.005 127.715 41.285 128.175 ;
        RECT 41.805 127.885 42.130 128.345 ;
        RECT 41.005 127.545 42.130 127.715 ;
        RECT 42.300 127.605 42.685 128.175 ;
        RECT 42.895 127.835 43.295 128.345 ;
        RECT 43.870 127.730 44.040 128.175 ;
        RECT 44.210 127.945 44.930 128.345 ;
        RECT 45.100 127.775 45.270 128.175 ;
        RECT 45.505 127.900 45.935 128.345 ;
        RECT 41.680 127.435 42.130 127.545 ;
        RECT 40.415 126.815 41.510 127.375 ;
        RECT 41.680 127.105 42.235 127.435 ;
        RECT 39.290 125.965 39.575 126.425 ;
        RECT 39.745 125.795 40.015 126.255 ;
        RECT 40.415 125.965 40.815 126.815 ;
        RECT 41.680 126.645 42.130 127.105 ;
        RECT 42.405 126.935 42.685 127.605 ;
        RECT 41.005 126.425 42.130 126.645 ;
        RECT 41.005 125.965 41.285 126.425 ;
        RECT 41.805 125.795 42.130 126.255 ;
        RECT 42.300 125.965 42.685 126.935 ;
        RECT 42.910 126.775 43.170 127.665 ;
        RECT 43.370 127.075 43.630 127.665 ;
        RECT 43.870 127.560 44.220 127.730 ;
        RECT 43.370 126.775 43.850 127.075 ;
        RECT 42.935 126.425 43.875 126.595 ;
        RECT 42.935 125.965 43.115 126.425 ;
        RECT 43.285 125.795 43.535 126.255 ;
        RECT 43.705 126.175 43.875 126.425 ;
        RECT 44.050 126.535 44.220 127.560 ;
        RECT 44.390 127.605 45.270 127.775 ;
        RECT 46.105 127.620 46.365 128.175 ;
        RECT 46.625 127.795 46.795 128.085 ;
        RECT 46.965 127.965 47.295 128.345 ;
        RECT 46.625 127.625 47.290 127.795 ;
        RECT 44.390 126.885 44.560 127.605 ;
        RECT 44.750 127.055 45.040 127.435 ;
        RECT 44.390 126.715 44.910 126.885 ;
        RECT 45.210 126.815 45.540 127.435 ;
        RECT 45.765 127.105 46.020 127.435 ;
        RECT 44.050 126.365 44.460 126.535 ;
        RECT 44.740 126.525 44.910 126.715 ;
        RECT 45.765 126.625 45.935 127.105 ;
        RECT 46.190 126.905 46.365 127.620 ;
        RECT 44.205 126.230 44.460 126.365 ;
        RECT 45.175 126.455 45.935 126.625 ;
        RECT 45.175 126.230 45.345 126.455 ;
        RECT 43.705 126.005 44.035 126.175 ;
        RECT 44.205 126.060 45.345 126.230 ;
        RECT 44.205 125.965 44.460 126.060 ;
        RECT 45.605 125.795 45.935 126.195 ;
        RECT 46.105 125.965 46.365 126.905 ;
        RECT 46.540 126.805 46.890 127.455 ;
        RECT 47.060 126.635 47.290 127.625 ;
        RECT 46.625 126.465 47.290 126.635 ;
        RECT 46.625 125.965 46.795 126.465 ;
        RECT 46.965 125.795 47.295 126.295 ;
        RECT 47.465 125.965 47.650 128.085 ;
        RECT 47.905 127.885 48.155 128.345 ;
        RECT 48.325 127.895 48.660 128.065 ;
        RECT 48.855 127.895 49.530 128.065 ;
        RECT 48.325 127.755 48.495 127.895 ;
        RECT 47.820 126.765 48.100 127.715 ;
        RECT 48.270 127.625 48.495 127.755 ;
        RECT 48.270 126.520 48.440 127.625 ;
        RECT 48.665 127.475 49.190 127.695 ;
        RECT 48.610 126.710 48.850 127.305 ;
        RECT 49.020 126.775 49.190 127.475 ;
        RECT 49.360 127.115 49.530 127.895 ;
        RECT 49.850 127.845 50.220 128.345 ;
        RECT 50.400 127.895 50.805 128.065 ;
        RECT 50.975 127.895 51.760 128.065 ;
        RECT 50.400 127.665 50.570 127.895 ;
        RECT 49.740 127.365 50.570 127.665 ;
        RECT 50.955 127.395 51.420 127.725 ;
        RECT 49.740 127.335 49.940 127.365 ;
        RECT 50.060 127.115 50.230 127.185 ;
        RECT 49.360 126.945 50.230 127.115 ;
        RECT 49.720 126.855 50.230 126.945 ;
        RECT 48.270 126.390 48.575 126.520 ;
        RECT 49.020 126.410 49.550 126.775 ;
        RECT 47.890 125.795 48.155 126.255 ;
        RECT 48.325 125.965 48.575 126.390 ;
        RECT 49.720 126.240 49.890 126.855 ;
        RECT 48.785 126.070 49.890 126.240 ;
        RECT 50.060 125.795 50.230 126.595 ;
        RECT 50.400 126.295 50.570 127.365 ;
        RECT 50.740 126.465 50.930 127.185 ;
        RECT 51.100 126.435 51.420 127.395 ;
        RECT 51.590 127.435 51.760 127.895 ;
        RECT 52.035 127.815 52.245 128.345 ;
        RECT 52.505 127.605 52.835 128.130 ;
        RECT 53.005 127.735 53.175 128.345 ;
        RECT 53.345 127.690 53.675 128.125 ;
        RECT 53.895 127.800 59.240 128.345 ;
        RECT 53.345 127.605 53.725 127.690 ;
        RECT 52.635 127.435 52.835 127.605 ;
        RECT 53.500 127.565 53.725 127.605 ;
        RECT 51.590 127.105 52.465 127.435 ;
        RECT 52.635 127.105 53.385 127.435 ;
        RECT 50.400 125.965 50.650 126.295 ;
        RECT 51.590 126.265 51.760 127.105 ;
        RECT 52.635 126.900 52.825 127.105 ;
        RECT 53.555 126.985 53.725 127.565 ;
        RECT 53.510 126.935 53.725 126.985 ;
        RECT 55.480 126.970 55.820 127.800 ;
        RECT 59.415 127.575 62.925 128.345 ;
        RECT 63.555 127.620 63.845 128.345 ;
        RECT 64.015 127.800 69.360 128.345 ;
        RECT 69.535 127.800 74.880 128.345 ;
        RECT 75.055 127.800 80.400 128.345 ;
        RECT 80.575 127.800 85.920 128.345 ;
        RECT 51.930 126.525 52.825 126.900 ;
        RECT 53.335 126.855 53.725 126.935 ;
        RECT 50.875 126.095 51.760 126.265 ;
        RECT 51.940 125.795 52.255 126.295 ;
        RECT 52.485 125.965 52.825 126.525 ;
        RECT 52.995 125.795 53.165 126.805 ;
        RECT 53.335 126.010 53.665 126.855 ;
        RECT 57.300 126.230 57.650 127.480 ;
        RECT 59.415 127.055 61.065 127.575 ;
        RECT 61.235 126.885 62.925 127.405 ;
        RECT 65.600 126.970 65.940 127.800 ;
        RECT 53.895 125.795 59.240 126.230 ;
        RECT 59.415 125.795 62.925 126.885 ;
        RECT 63.555 125.795 63.845 126.960 ;
        RECT 67.420 126.230 67.770 127.480 ;
        RECT 71.120 126.970 71.460 127.800 ;
        RECT 72.940 126.230 73.290 127.480 ;
        RECT 76.640 126.970 76.980 127.800 ;
        RECT 78.460 126.230 78.810 127.480 ;
        RECT 82.160 126.970 82.500 127.800 ;
        RECT 86.095 127.575 88.685 128.345 ;
        RECT 89.315 127.595 90.525 128.345 ;
        RECT 83.980 126.230 84.330 127.480 ;
        RECT 86.095 127.055 87.305 127.575 ;
        RECT 87.475 126.885 88.685 127.405 ;
        RECT 64.015 125.795 69.360 126.230 ;
        RECT 69.535 125.795 74.880 126.230 ;
        RECT 75.055 125.795 80.400 126.230 ;
        RECT 80.575 125.795 85.920 126.230 ;
        RECT 86.095 125.795 88.685 126.885 ;
        RECT 89.315 126.885 89.835 127.425 ;
        RECT 90.005 127.055 90.525 127.595 ;
        RECT 89.315 125.795 90.525 126.885 ;
        RECT 100.140 125.890 100.810 129.150 ;
        RECT 101.480 128.580 105.520 128.750 ;
        RECT 101.140 126.520 101.310 128.520 ;
        RECT 105.690 126.520 105.860 128.520 ;
        RECT 101.480 126.290 105.520 126.460 ;
        RECT 106.200 125.890 106.370 129.150 ;
        RECT 11.950 125.625 90.610 125.795 ;
        RECT 100.140 125.720 106.370 125.890 ;
        RECT 12.035 124.535 13.245 125.625 ;
        RECT 13.415 125.190 18.760 125.625 ;
        RECT 18.935 125.190 24.280 125.625 ;
        RECT 12.035 123.825 12.555 124.365 ;
        RECT 12.725 123.995 13.245 124.535 ;
        RECT 12.035 123.075 13.245 123.825 ;
        RECT 15.000 123.620 15.340 124.450 ;
        RECT 16.820 123.940 17.170 125.190 ;
        RECT 20.520 123.620 20.860 124.450 ;
        RECT 22.340 123.940 22.690 125.190 ;
        RECT 24.915 124.460 25.205 125.625 ;
        RECT 25.375 124.535 26.585 125.625 ;
        RECT 26.870 124.995 27.155 125.455 ;
        RECT 27.325 125.165 27.595 125.625 ;
        RECT 26.870 124.775 27.825 124.995 ;
        RECT 25.375 123.825 25.895 124.365 ;
        RECT 26.065 123.995 26.585 124.535 ;
        RECT 26.755 124.045 27.445 124.605 ;
        RECT 27.615 123.875 27.825 124.775 ;
        RECT 13.415 123.075 18.760 123.620 ;
        RECT 18.935 123.075 24.280 123.620 ;
        RECT 24.915 123.075 25.205 123.800 ;
        RECT 25.375 123.075 26.585 123.825 ;
        RECT 26.870 123.705 27.825 123.875 ;
        RECT 27.995 124.605 28.395 125.455 ;
        RECT 28.585 124.995 28.865 125.455 ;
        RECT 29.385 125.165 29.710 125.625 ;
        RECT 28.585 124.775 29.710 124.995 ;
        RECT 27.995 124.045 29.090 124.605 ;
        RECT 29.260 124.315 29.710 124.775 ;
        RECT 29.880 124.485 30.265 125.455 ;
        RECT 30.435 124.535 33.025 125.625 ;
        RECT 26.870 123.245 27.155 123.705 ;
        RECT 27.325 123.075 27.595 123.535 ;
        RECT 27.995 123.245 28.395 124.045 ;
        RECT 29.260 123.985 29.815 124.315 ;
        RECT 29.260 123.875 29.710 123.985 ;
        RECT 28.585 123.705 29.710 123.875 ;
        RECT 29.985 123.815 30.265 124.485 ;
        RECT 28.585 123.245 28.865 123.705 ;
        RECT 29.385 123.075 29.710 123.535 ;
        RECT 29.880 123.245 30.265 123.815 ;
        RECT 30.435 123.845 31.645 124.365 ;
        RECT 31.815 124.015 33.025 124.535 ;
        RECT 33.655 124.060 34.005 125.455 ;
        RECT 34.175 124.825 34.580 125.625 ;
        RECT 34.750 125.285 36.285 125.455 ;
        RECT 34.750 124.655 34.920 125.285 ;
        RECT 34.175 124.485 34.920 124.655 ;
        RECT 30.435 123.075 33.025 123.845 ;
        RECT 33.655 123.245 33.925 124.060 ;
        RECT 34.175 123.985 34.345 124.485 ;
        RECT 35.090 124.315 35.360 125.060 ;
        RECT 34.515 123.985 34.850 124.315 ;
        RECT 35.020 123.985 35.360 124.315 ;
        RECT 35.550 124.315 35.785 125.060 ;
        RECT 35.955 124.655 36.285 125.285 ;
        RECT 36.470 124.825 36.705 125.625 ;
        RECT 36.875 124.655 37.165 125.455 ;
        RECT 35.955 124.485 37.165 124.655 ;
        RECT 37.335 125.035 38.035 125.455 ;
        RECT 38.235 125.265 38.565 125.625 ;
        RECT 38.735 125.035 39.065 125.435 ;
        RECT 37.335 124.805 39.065 125.035 ;
        RECT 35.550 123.985 35.840 124.315 ;
        RECT 36.010 123.985 36.410 124.315 ;
        RECT 36.580 123.815 36.750 124.485 ;
        RECT 36.920 123.985 37.165 124.315 ;
        RECT 37.335 123.835 37.540 124.805 ;
        RECT 37.710 124.065 38.040 124.605 ;
        RECT 38.215 124.315 38.540 124.605 ;
        RECT 38.735 124.585 39.065 124.805 ;
        RECT 39.235 124.315 39.405 125.285 ;
        RECT 39.585 124.565 39.915 125.625 ;
        RECT 40.185 124.955 40.355 125.455 ;
        RECT 40.525 125.125 40.855 125.625 ;
        RECT 40.185 124.785 40.850 124.955 ;
        RECT 38.215 123.985 38.710 124.315 ;
        RECT 39.030 123.985 39.405 124.315 ;
        RECT 39.615 123.985 39.925 124.315 ;
        RECT 40.100 123.965 40.450 124.615 ;
        RECT 34.095 123.075 34.765 123.815 ;
        RECT 34.935 123.645 36.330 123.815 ;
        RECT 34.935 123.300 35.230 123.645 ;
        RECT 35.410 123.075 35.785 123.475 ;
        RECT 36.000 123.300 36.330 123.645 ;
        RECT 36.580 123.245 37.165 123.815 ;
        RECT 37.335 123.245 38.045 123.835 ;
        RECT 38.555 123.605 39.915 123.815 ;
        RECT 40.620 123.795 40.850 124.785 ;
        RECT 38.555 123.245 38.885 123.605 ;
        RECT 39.085 123.075 39.415 123.435 ;
        RECT 39.585 123.245 39.915 123.605 ;
        RECT 40.185 123.625 40.850 123.795 ;
        RECT 40.185 123.335 40.355 123.625 ;
        RECT 40.525 123.075 40.855 123.455 ;
        RECT 41.025 123.335 41.210 125.455 ;
        RECT 41.450 125.165 41.715 125.625 ;
        RECT 41.885 125.030 42.135 125.455 ;
        RECT 42.345 125.180 43.450 125.350 ;
        RECT 41.830 124.900 42.135 125.030 ;
        RECT 41.380 123.705 41.660 124.655 ;
        RECT 41.830 123.795 42.000 124.900 ;
        RECT 42.170 124.115 42.410 124.710 ;
        RECT 42.580 124.645 43.110 125.010 ;
        RECT 42.580 123.945 42.750 124.645 ;
        RECT 43.280 124.565 43.450 125.180 ;
        RECT 43.620 124.825 43.790 125.625 ;
        RECT 43.960 125.125 44.210 125.455 ;
        RECT 44.435 125.155 45.320 125.325 ;
        RECT 43.280 124.475 43.790 124.565 ;
        RECT 41.830 123.665 42.055 123.795 ;
        RECT 42.225 123.725 42.750 123.945 ;
        RECT 42.920 124.305 43.790 124.475 ;
        RECT 41.465 123.075 41.715 123.535 ;
        RECT 41.885 123.525 42.055 123.665 ;
        RECT 42.920 123.525 43.090 124.305 ;
        RECT 43.620 124.235 43.790 124.305 ;
        RECT 43.300 124.055 43.500 124.085 ;
        RECT 43.960 124.055 44.130 125.125 ;
        RECT 44.300 124.235 44.490 124.955 ;
        RECT 43.300 123.755 44.130 124.055 ;
        RECT 44.660 124.025 44.980 124.985 ;
        RECT 41.885 123.355 42.220 123.525 ;
        RECT 42.415 123.355 43.090 123.525 ;
        RECT 43.410 123.075 43.780 123.575 ;
        RECT 43.960 123.525 44.130 123.755 ;
        RECT 44.515 123.695 44.980 124.025 ;
        RECT 45.150 124.315 45.320 125.155 ;
        RECT 45.500 125.125 45.815 125.625 ;
        RECT 46.045 124.895 46.385 125.455 ;
        RECT 45.490 124.520 46.385 124.895 ;
        RECT 46.555 124.615 46.725 125.625 ;
        RECT 46.195 124.315 46.385 124.520 ;
        RECT 46.895 124.565 47.225 125.410 ;
        RECT 47.455 125.115 48.645 125.405 ;
        RECT 47.475 124.775 48.645 124.945 ;
        RECT 48.815 124.825 49.095 125.625 ;
        RECT 46.895 124.485 47.285 124.565 ;
        RECT 47.475 124.485 47.800 124.775 ;
        RECT 48.475 124.655 48.645 124.775 ;
        RECT 47.070 124.435 47.285 124.485 ;
        RECT 45.150 123.985 46.025 124.315 ;
        RECT 46.195 123.985 46.945 124.315 ;
        RECT 45.150 123.525 45.320 123.985 ;
        RECT 46.195 123.815 46.395 123.985 ;
        RECT 47.115 123.855 47.285 124.435 ;
        RECT 47.970 124.315 48.165 124.605 ;
        RECT 48.475 124.485 49.135 124.655 ;
        RECT 49.305 124.485 49.580 125.455 ;
        RECT 48.965 124.315 49.135 124.485 ;
        RECT 47.455 123.985 47.800 124.315 ;
        RECT 47.970 123.985 48.795 124.315 ;
        RECT 48.965 123.985 49.240 124.315 ;
        RECT 47.060 123.815 47.285 123.855 ;
        RECT 48.965 123.815 49.135 123.985 ;
        RECT 43.960 123.355 44.365 123.525 ;
        RECT 44.535 123.355 45.320 123.525 ;
        RECT 45.595 123.075 45.805 123.605 ;
        RECT 46.065 123.290 46.395 123.815 ;
        RECT 46.905 123.730 47.285 123.815 ;
        RECT 46.565 123.075 46.735 123.685 ;
        RECT 46.905 123.295 47.235 123.730 ;
        RECT 47.470 123.645 49.135 123.815 ;
        RECT 49.410 123.750 49.580 124.485 ;
        RECT 50.675 124.460 50.965 125.625 ;
        RECT 51.135 124.655 51.445 125.455 ;
        RECT 51.615 124.825 51.925 125.625 ;
        RECT 52.095 124.995 52.355 125.455 ;
        RECT 52.525 125.165 52.780 125.625 ;
        RECT 52.955 124.995 53.215 125.455 ;
        RECT 52.095 124.825 53.215 124.995 ;
        RECT 52.575 124.775 52.745 124.825 ;
        RECT 51.135 124.485 52.165 124.655 ;
        RECT 47.470 123.295 47.725 123.645 ;
        RECT 47.895 123.075 48.225 123.475 ;
        RECT 48.395 123.295 48.565 123.645 ;
        RECT 48.735 123.075 49.115 123.475 ;
        RECT 49.305 123.405 49.580 123.750 ;
        RECT 50.675 123.075 50.965 123.800 ;
        RECT 51.135 123.575 51.305 124.485 ;
        RECT 51.475 123.745 51.825 124.315 ;
        RECT 51.995 124.235 52.165 124.485 ;
        RECT 52.955 124.575 53.215 124.825 ;
        RECT 53.385 124.755 53.670 125.625 ;
        RECT 52.955 124.405 53.710 124.575 ;
        RECT 53.895 124.535 55.565 125.625 ;
        RECT 51.995 124.065 53.135 124.235 ;
        RECT 53.305 123.895 53.710 124.405 ;
        RECT 52.060 123.725 53.710 123.895 ;
        RECT 53.895 123.845 54.645 124.365 ;
        RECT 54.815 124.015 55.565 124.535 ;
        RECT 55.735 124.485 56.120 125.455 ;
        RECT 56.290 125.165 56.615 125.625 ;
        RECT 57.135 124.995 57.415 125.455 ;
        RECT 56.290 124.775 57.415 124.995 ;
        RECT 51.135 123.245 51.435 123.575 ;
        RECT 51.605 123.075 51.880 123.555 ;
        RECT 52.060 123.335 52.355 123.725 ;
        RECT 52.525 123.075 52.780 123.555 ;
        RECT 52.955 123.335 53.215 123.725 ;
        RECT 53.385 123.075 53.665 123.555 ;
        RECT 53.895 123.075 55.565 123.845 ;
        RECT 55.735 123.815 56.015 124.485 ;
        RECT 56.290 124.315 56.740 124.775 ;
        RECT 57.605 124.605 58.005 125.455 ;
        RECT 58.405 125.165 58.675 125.625 ;
        RECT 58.845 124.995 59.130 125.455 ;
        RECT 56.185 123.985 56.740 124.315 ;
        RECT 56.910 124.045 58.005 124.605 ;
        RECT 56.290 123.875 56.740 123.985 ;
        RECT 55.735 123.245 56.120 123.815 ;
        RECT 56.290 123.705 57.415 123.875 ;
        RECT 56.290 123.075 56.615 123.535 ;
        RECT 57.135 123.245 57.415 123.705 ;
        RECT 57.605 123.245 58.005 124.045 ;
        RECT 58.175 124.775 59.130 124.995 ;
        RECT 58.175 123.875 58.385 124.775 ;
        RECT 58.555 124.045 59.245 124.605 ;
        RECT 59.415 124.535 61.085 125.625 ;
        RECT 58.175 123.705 59.130 123.875 ;
        RECT 58.405 123.075 58.675 123.535 ;
        RECT 58.845 123.245 59.130 123.705 ;
        RECT 59.415 123.845 60.165 124.365 ;
        RECT 60.335 124.015 61.085 124.535 ;
        RECT 61.255 124.485 61.640 125.455 ;
        RECT 61.810 125.165 62.135 125.625 ;
        RECT 62.655 124.995 62.935 125.455 ;
        RECT 61.810 124.775 62.935 124.995 ;
        RECT 59.415 123.075 61.085 123.845 ;
        RECT 61.255 123.815 61.535 124.485 ;
        RECT 61.810 124.315 62.260 124.775 ;
        RECT 63.125 124.605 63.525 125.455 ;
        RECT 63.925 125.165 64.195 125.625 ;
        RECT 64.365 124.995 64.650 125.455 ;
        RECT 61.705 123.985 62.260 124.315 ;
        RECT 62.430 124.045 63.525 124.605 ;
        RECT 61.810 123.875 62.260 123.985 ;
        RECT 61.255 123.245 61.640 123.815 ;
        RECT 61.810 123.705 62.935 123.875 ;
        RECT 61.810 123.075 62.135 123.535 ;
        RECT 62.655 123.245 62.935 123.705 ;
        RECT 63.125 123.245 63.525 124.045 ;
        RECT 63.695 124.775 64.650 124.995 ;
        RECT 63.695 123.875 63.905 124.775 ;
        RECT 64.075 124.045 64.765 124.605 ;
        RECT 64.935 124.485 65.275 125.455 ;
        RECT 65.445 124.485 65.615 125.625 ;
        RECT 65.885 124.825 66.135 125.625 ;
        RECT 66.780 124.655 67.110 125.455 ;
        RECT 67.410 124.825 67.740 125.625 ;
        RECT 67.910 124.655 68.240 125.455 ;
        RECT 68.615 125.190 73.960 125.625 ;
        RECT 65.805 124.485 68.240 124.655 ;
        RECT 64.935 124.435 65.165 124.485 ;
        RECT 64.935 123.875 65.110 124.435 ;
        RECT 65.805 124.235 65.975 124.485 ;
        RECT 65.280 124.065 65.975 124.235 ;
        RECT 66.150 124.065 66.570 124.265 ;
        RECT 66.740 124.065 67.070 124.265 ;
        RECT 67.240 124.065 67.570 124.265 ;
        RECT 63.695 123.705 64.650 123.875 ;
        RECT 63.925 123.075 64.195 123.535 ;
        RECT 64.365 123.245 64.650 123.705 ;
        RECT 64.935 123.245 65.275 123.875 ;
        RECT 65.445 123.075 65.695 123.875 ;
        RECT 65.885 123.725 67.110 123.895 ;
        RECT 65.885 123.245 66.215 123.725 ;
        RECT 66.385 123.075 66.610 123.535 ;
        RECT 66.780 123.245 67.110 123.725 ;
        RECT 67.740 123.855 67.910 124.485 ;
        RECT 68.095 124.065 68.445 124.315 ;
        RECT 67.740 123.245 68.240 123.855 ;
        RECT 70.200 123.620 70.540 124.450 ;
        RECT 72.020 123.940 72.370 125.190 ;
        RECT 74.135 124.535 75.805 125.625 ;
        RECT 74.135 123.845 74.885 124.365 ;
        RECT 75.055 124.015 75.805 124.535 ;
        RECT 76.435 124.460 76.725 125.625 ;
        RECT 76.895 125.190 82.240 125.625 ;
        RECT 82.415 125.190 87.760 125.625 ;
        RECT 68.615 123.075 73.960 123.620 ;
        RECT 74.135 123.075 75.805 123.845 ;
        RECT 76.435 123.075 76.725 123.800 ;
        RECT 78.480 123.620 78.820 124.450 ;
        RECT 80.300 123.940 80.650 125.190 ;
        RECT 84.000 123.620 84.340 124.450 ;
        RECT 85.820 123.940 86.170 125.190 ;
        RECT 87.935 124.535 89.145 125.625 ;
        RECT 87.935 123.825 88.455 124.365 ;
        RECT 88.625 123.995 89.145 124.535 ;
        RECT 89.315 124.535 90.525 125.625 ;
        RECT 89.315 123.995 89.835 124.535 ;
        RECT 90.005 123.825 90.525 124.365 ;
        RECT 76.895 123.075 82.240 123.620 ;
        RECT 82.415 123.075 87.760 123.620 ;
        RECT 87.935 123.075 89.145 123.825 ;
        RECT 89.315 123.075 90.525 123.825 ;
        RECT 11.950 122.905 90.610 123.075 ;
        RECT 12.035 122.155 13.245 122.905 ;
        RECT 13.415 122.360 18.760 122.905 ;
        RECT 12.035 121.615 12.555 122.155 ;
        RECT 12.725 121.445 13.245 121.985 ;
        RECT 15.000 121.530 15.340 122.360 ;
        RECT 18.935 122.135 21.525 122.905 ;
        RECT 21.785 122.355 21.955 122.645 ;
        RECT 22.125 122.525 22.455 122.905 ;
        RECT 21.785 122.185 22.450 122.355 ;
        RECT 12.035 120.355 13.245 121.445 ;
        RECT 16.820 120.790 17.170 122.040 ;
        RECT 18.935 121.615 20.145 122.135 ;
        RECT 20.315 121.445 21.525 121.965 ;
        RECT 13.415 120.355 18.760 120.790 ;
        RECT 18.935 120.355 21.525 121.445 ;
        RECT 21.700 121.365 22.050 122.015 ;
        RECT 22.220 121.195 22.450 122.185 ;
        RECT 21.785 121.025 22.450 121.195 ;
        RECT 21.785 120.525 21.955 121.025 ;
        RECT 22.125 120.355 22.455 120.855 ;
        RECT 22.625 120.525 22.810 122.645 ;
        RECT 23.065 122.445 23.315 122.905 ;
        RECT 23.485 122.455 23.820 122.625 ;
        RECT 24.015 122.455 24.690 122.625 ;
        RECT 23.485 122.315 23.655 122.455 ;
        RECT 22.980 121.325 23.260 122.275 ;
        RECT 23.430 122.185 23.655 122.315 ;
        RECT 23.430 121.080 23.600 122.185 ;
        RECT 23.825 122.035 24.350 122.255 ;
        RECT 23.770 121.270 24.010 121.865 ;
        RECT 24.180 121.335 24.350 122.035 ;
        RECT 24.520 121.675 24.690 122.455 ;
        RECT 25.010 122.405 25.380 122.905 ;
        RECT 25.560 122.455 25.965 122.625 ;
        RECT 26.135 122.455 26.920 122.625 ;
        RECT 25.560 122.225 25.730 122.455 ;
        RECT 24.900 121.925 25.730 122.225 ;
        RECT 26.115 121.955 26.580 122.285 ;
        RECT 24.900 121.895 25.100 121.925 ;
        RECT 25.220 121.675 25.390 121.745 ;
        RECT 24.520 121.505 25.390 121.675 ;
        RECT 24.880 121.415 25.390 121.505 ;
        RECT 23.430 120.950 23.735 121.080 ;
        RECT 24.180 120.970 24.710 121.335 ;
        RECT 23.050 120.355 23.315 120.815 ;
        RECT 23.485 120.525 23.735 120.950 ;
        RECT 24.880 120.800 25.050 121.415 ;
        RECT 23.945 120.630 25.050 120.800 ;
        RECT 25.220 120.355 25.390 121.155 ;
        RECT 25.560 120.855 25.730 121.925 ;
        RECT 25.900 121.025 26.090 121.745 ;
        RECT 26.260 120.995 26.580 121.955 ;
        RECT 26.750 121.995 26.920 122.455 ;
        RECT 27.195 122.375 27.405 122.905 ;
        RECT 27.665 122.165 27.995 122.690 ;
        RECT 28.165 122.295 28.335 122.905 ;
        RECT 28.505 122.250 28.835 122.685 ;
        RECT 29.055 122.360 34.400 122.905 ;
        RECT 28.505 122.165 28.885 122.250 ;
        RECT 27.795 121.995 27.995 122.165 ;
        RECT 28.660 122.125 28.885 122.165 ;
        RECT 26.750 121.665 27.625 121.995 ;
        RECT 27.795 121.665 28.545 121.995 ;
        RECT 25.560 120.525 25.810 120.855 ;
        RECT 26.750 120.825 26.920 121.665 ;
        RECT 27.795 121.460 27.985 121.665 ;
        RECT 28.715 121.545 28.885 122.125 ;
        RECT 28.670 121.495 28.885 121.545 ;
        RECT 30.640 121.530 30.980 122.360 ;
        RECT 34.575 122.135 37.165 122.905 ;
        RECT 37.795 122.180 38.085 122.905 ;
        RECT 38.255 122.360 43.600 122.905 ;
        RECT 27.090 121.085 27.985 121.460 ;
        RECT 28.495 121.415 28.885 121.495 ;
        RECT 26.035 120.655 26.920 120.825 ;
        RECT 27.100 120.355 27.415 120.855 ;
        RECT 27.645 120.525 27.985 121.085 ;
        RECT 28.155 120.355 28.325 121.365 ;
        RECT 28.495 120.570 28.825 121.415 ;
        RECT 32.460 120.790 32.810 122.040 ;
        RECT 34.575 121.615 35.785 122.135 ;
        RECT 35.955 121.445 37.165 121.965 ;
        RECT 39.840 121.530 40.180 122.360 ;
        RECT 43.810 122.165 44.425 122.735 ;
        RECT 44.595 122.395 44.810 122.905 ;
        RECT 45.040 122.395 45.320 122.725 ;
        RECT 45.500 122.395 45.740 122.905 ;
        RECT 29.055 120.355 34.400 120.790 ;
        RECT 34.575 120.355 37.165 121.445 ;
        RECT 37.795 120.355 38.085 121.520 ;
        RECT 41.660 120.790 42.010 122.040 ;
        RECT 43.810 121.145 44.125 122.165 ;
        RECT 44.295 121.495 44.465 121.995 ;
        RECT 44.715 121.665 44.980 122.225 ;
        RECT 45.150 121.495 45.320 122.395 ;
        RECT 45.490 121.665 45.845 122.225 ;
        RECT 46.135 122.085 46.345 122.905 ;
        RECT 46.515 122.105 46.845 122.735 ;
        RECT 46.515 121.505 46.765 122.105 ;
        RECT 47.015 122.085 47.245 122.905 ;
        RECT 47.465 122.095 47.735 122.905 ;
        RECT 47.905 122.095 48.235 122.735 ;
        RECT 48.405 122.095 48.645 122.905 ;
        RECT 48.835 122.135 52.345 122.905 ;
        RECT 52.515 122.155 53.725 122.905 ;
        RECT 53.985 122.355 54.155 122.645 ;
        RECT 54.325 122.525 54.655 122.905 ;
        RECT 53.985 122.185 54.650 122.355 ;
        RECT 46.935 121.665 47.265 121.915 ;
        RECT 47.455 121.665 47.805 121.915 ;
        RECT 44.295 121.325 45.720 121.495 ;
        RECT 38.255 120.355 43.600 120.790 ;
        RECT 43.810 120.525 44.345 121.145 ;
        RECT 44.515 120.355 44.845 121.155 ;
        RECT 45.330 121.150 45.720 121.325 ;
        RECT 46.135 120.355 46.345 121.495 ;
        RECT 46.515 120.525 46.845 121.505 ;
        RECT 47.975 121.495 48.145 122.095 ;
        RECT 48.315 121.665 48.665 121.915 ;
        RECT 48.835 121.615 50.485 122.135 ;
        RECT 47.015 120.355 47.245 121.495 ;
        RECT 47.465 120.355 47.795 121.495 ;
        RECT 47.975 121.325 48.655 121.495 ;
        RECT 50.655 121.445 52.345 121.965 ;
        RECT 52.515 121.615 53.035 122.155 ;
        RECT 53.205 121.445 53.725 121.985 ;
        RECT 48.325 120.540 48.655 121.325 ;
        RECT 48.835 120.355 52.345 121.445 ;
        RECT 52.515 120.355 53.725 121.445 ;
        RECT 53.900 121.365 54.250 122.015 ;
        RECT 54.420 121.195 54.650 122.185 ;
        RECT 53.985 121.025 54.650 121.195 ;
        RECT 53.985 120.525 54.155 121.025 ;
        RECT 54.325 120.355 54.655 120.855 ;
        RECT 54.825 120.525 55.010 122.645 ;
        RECT 55.265 122.445 55.515 122.905 ;
        RECT 55.685 122.455 56.020 122.625 ;
        RECT 56.215 122.455 56.890 122.625 ;
        RECT 55.685 122.315 55.855 122.455 ;
        RECT 55.180 121.325 55.460 122.275 ;
        RECT 55.630 122.185 55.855 122.315 ;
        RECT 55.630 121.080 55.800 122.185 ;
        RECT 56.025 122.035 56.550 122.255 ;
        RECT 55.970 121.270 56.210 121.865 ;
        RECT 56.380 121.335 56.550 122.035 ;
        RECT 56.720 121.675 56.890 122.455 ;
        RECT 57.210 122.405 57.580 122.905 ;
        RECT 57.760 122.455 58.165 122.625 ;
        RECT 58.335 122.455 59.120 122.625 ;
        RECT 57.760 122.225 57.930 122.455 ;
        RECT 57.100 121.925 57.930 122.225 ;
        RECT 58.315 121.955 58.780 122.285 ;
        RECT 57.100 121.895 57.300 121.925 ;
        RECT 57.420 121.675 57.590 121.745 ;
        RECT 56.720 121.505 57.590 121.675 ;
        RECT 57.080 121.415 57.590 121.505 ;
        RECT 55.630 120.950 55.935 121.080 ;
        RECT 56.380 120.970 56.910 121.335 ;
        RECT 55.250 120.355 55.515 120.815 ;
        RECT 55.685 120.525 55.935 120.950 ;
        RECT 57.080 120.800 57.250 121.415 ;
        RECT 56.145 120.630 57.250 120.800 ;
        RECT 57.420 120.355 57.590 121.155 ;
        RECT 57.760 120.855 57.930 121.925 ;
        RECT 58.100 121.025 58.290 121.745 ;
        RECT 58.460 120.995 58.780 121.955 ;
        RECT 58.950 121.995 59.120 122.455 ;
        RECT 59.395 122.375 59.605 122.905 ;
        RECT 59.865 122.165 60.195 122.690 ;
        RECT 60.365 122.295 60.535 122.905 ;
        RECT 60.705 122.250 61.035 122.685 ;
        RECT 60.705 122.165 61.085 122.250 ;
        RECT 59.995 121.995 60.195 122.165 ;
        RECT 60.860 122.125 61.085 122.165 ;
        RECT 58.950 121.665 59.825 121.995 ;
        RECT 59.995 121.665 60.745 121.995 ;
        RECT 57.760 120.525 58.010 120.855 ;
        RECT 58.950 120.825 59.120 121.665 ;
        RECT 59.995 121.460 60.185 121.665 ;
        RECT 60.915 121.545 61.085 122.125 ;
        RECT 61.275 122.095 61.515 122.905 ;
        RECT 61.685 122.095 62.015 122.735 ;
        RECT 62.185 122.095 62.455 122.905 ;
        RECT 63.555 122.180 63.845 122.905 ;
        RECT 64.015 122.135 65.685 122.905 ;
        RECT 65.905 122.250 66.235 122.685 ;
        RECT 66.405 122.295 66.575 122.905 ;
        RECT 65.855 122.165 66.235 122.250 ;
        RECT 66.745 122.165 67.075 122.690 ;
        RECT 67.335 122.375 67.545 122.905 ;
        RECT 67.820 122.455 68.605 122.625 ;
        RECT 68.775 122.455 69.180 122.625 ;
        RECT 61.255 121.665 61.605 121.915 ;
        RECT 60.870 121.495 61.085 121.545 ;
        RECT 61.775 121.495 61.945 122.095 ;
        RECT 62.115 121.665 62.465 121.915 ;
        RECT 64.015 121.615 64.765 122.135 ;
        RECT 65.855 122.125 66.080 122.165 ;
        RECT 59.290 121.085 60.185 121.460 ;
        RECT 60.695 121.415 61.085 121.495 ;
        RECT 58.235 120.655 59.120 120.825 ;
        RECT 59.300 120.355 59.615 120.855 ;
        RECT 59.845 120.525 60.185 121.085 ;
        RECT 60.355 120.355 60.525 121.365 ;
        RECT 60.695 120.570 61.025 121.415 ;
        RECT 61.265 121.325 61.945 121.495 ;
        RECT 61.265 120.540 61.595 121.325 ;
        RECT 62.125 120.355 62.455 121.495 ;
        RECT 63.555 120.355 63.845 121.520 ;
        RECT 64.935 121.445 65.685 121.965 ;
        RECT 64.015 120.355 65.685 121.445 ;
        RECT 65.855 121.545 66.025 122.125 ;
        RECT 66.745 121.995 66.945 122.165 ;
        RECT 67.820 121.995 67.990 122.455 ;
        RECT 66.195 121.665 66.945 121.995 ;
        RECT 67.115 121.665 67.990 121.995 ;
        RECT 65.855 121.495 66.070 121.545 ;
        RECT 65.855 121.415 66.245 121.495 ;
        RECT 65.915 120.570 66.245 121.415 ;
        RECT 66.755 121.460 66.945 121.665 ;
        RECT 66.415 120.355 66.585 121.365 ;
        RECT 66.755 121.085 67.650 121.460 ;
        RECT 66.755 120.525 67.095 121.085 ;
        RECT 67.325 120.355 67.640 120.855 ;
        RECT 67.820 120.825 67.990 121.665 ;
        RECT 68.160 121.955 68.625 122.285 ;
        RECT 69.010 122.225 69.180 122.455 ;
        RECT 69.360 122.405 69.730 122.905 ;
        RECT 70.050 122.455 70.725 122.625 ;
        RECT 70.920 122.455 71.255 122.625 ;
        RECT 68.160 120.995 68.480 121.955 ;
        RECT 69.010 121.925 69.840 122.225 ;
        RECT 68.650 121.025 68.840 121.745 ;
        RECT 69.010 120.855 69.180 121.925 ;
        RECT 69.640 121.895 69.840 121.925 ;
        RECT 69.350 121.675 69.520 121.745 ;
        RECT 70.050 121.675 70.220 122.455 ;
        RECT 71.085 122.315 71.255 122.455 ;
        RECT 71.425 122.445 71.675 122.905 ;
        RECT 69.350 121.505 70.220 121.675 ;
        RECT 70.390 122.035 70.915 122.255 ;
        RECT 71.085 122.185 71.310 122.315 ;
        RECT 69.350 121.415 69.860 121.505 ;
        RECT 67.820 120.655 68.705 120.825 ;
        RECT 68.930 120.525 69.180 120.855 ;
        RECT 69.350 120.355 69.520 121.155 ;
        RECT 69.690 120.800 69.860 121.415 ;
        RECT 70.390 121.335 70.560 122.035 ;
        RECT 70.030 120.970 70.560 121.335 ;
        RECT 70.730 121.270 70.970 121.865 ;
        RECT 71.140 121.080 71.310 122.185 ;
        RECT 71.480 121.325 71.760 122.275 ;
        RECT 71.005 120.950 71.310 121.080 ;
        RECT 69.690 120.630 70.795 120.800 ;
        RECT 71.005 120.525 71.255 120.950 ;
        RECT 71.425 120.355 71.690 120.815 ;
        RECT 71.930 120.525 72.115 122.645 ;
        RECT 72.285 122.525 72.615 122.905 ;
        RECT 72.785 122.355 72.955 122.645 ;
        RECT 73.215 122.360 78.560 122.905 ;
        RECT 78.735 122.360 84.080 122.905 ;
        RECT 72.290 122.185 72.955 122.355 ;
        RECT 72.290 121.195 72.520 122.185 ;
        RECT 72.690 121.365 73.040 122.015 ;
        RECT 74.800 121.530 75.140 122.360 ;
        RECT 72.290 121.025 72.955 121.195 ;
        RECT 72.285 120.355 72.615 120.855 ;
        RECT 72.785 120.525 72.955 121.025 ;
        RECT 76.620 120.790 76.970 122.040 ;
        RECT 80.320 121.530 80.660 122.360 ;
        RECT 84.255 122.135 87.765 122.905 ;
        RECT 87.935 122.155 89.145 122.905 ;
        RECT 89.315 122.155 90.525 122.905 ;
        RECT 100.140 122.460 100.810 125.720 ;
        RECT 101.480 125.150 105.520 125.320 ;
        RECT 101.140 123.090 101.310 125.090 ;
        RECT 105.690 123.090 105.860 125.090 ;
        RECT 101.480 122.860 105.520 123.030 ;
        RECT 106.200 122.460 106.370 125.720 ;
        RECT 100.140 122.450 106.370 122.460 ;
        RECT 107.960 131.720 117.790 131.760 ;
        RECT 107.960 131.590 118.590 131.720 ;
        RECT 107.960 129.330 108.130 131.590 ;
        RECT 108.855 131.020 116.895 131.190 ;
        RECT 108.470 129.960 108.640 130.960 ;
        RECT 117.110 129.960 117.280 130.960 ;
        RECT 108.855 129.730 116.895 129.900 ;
        RECT 117.620 129.330 118.590 131.590 ;
        RECT 107.960 129.160 118.590 129.330 ;
        RECT 107.960 125.900 108.130 129.160 ;
        RECT 108.855 128.590 116.895 128.760 ;
        RECT 108.470 126.530 108.640 128.530 ;
        RECT 117.110 126.530 117.280 128.530 ;
        RECT 108.855 126.300 116.895 126.470 ;
        RECT 117.620 125.900 118.590 129.160 ;
        RECT 107.960 125.730 118.590 125.900 ;
        RECT 107.960 122.470 108.130 125.730 ;
        RECT 108.855 125.160 116.895 125.330 ;
        RECT 108.470 123.100 108.640 125.100 ;
        RECT 117.110 123.100 117.280 125.100 ;
        RECT 108.855 122.870 116.895 123.040 ;
        RECT 117.620 122.470 118.590 125.730 ;
        RECT 100.140 122.350 106.380 122.450 ;
        RECT 82.140 120.790 82.490 122.040 ;
        RECT 84.255 121.615 85.905 122.135 ;
        RECT 86.075 121.445 87.765 121.965 ;
        RECT 87.935 121.615 88.455 122.155 ;
        RECT 88.625 121.445 89.145 121.985 ;
        RECT 73.215 120.355 78.560 120.790 ;
        RECT 78.735 120.355 84.080 120.790 ;
        RECT 84.255 120.355 87.765 121.445 ;
        RECT 87.935 120.355 89.145 121.445 ;
        RECT 89.315 121.445 89.835 121.985 ;
        RECT 90.005 121.615 90.525 122.155 ;
        RECT 100.130 121.790 106.380 122.350 ;
        RECT 100.130 121.770 105.300 121.790 ;
        RECT 100.130 121.700 104.120 121.770 ;
        RECT 89.315 120.355 90.525 121.445 ;
        RECT 100.130 120.430 102.050 121.700 ;
        RECT 103.560 121.690 104.120 121.700 ;
        RECT 103.790 120.600 104.120 121.690 ;
        RECT 104.490 121.220 105.530 121.390 ;
        RECT 104.490 120.780 105.530 120.950 ;
        RECT 105.700 120.920 105.870 121.250 ;
        RECT 103.950 120.380 104.120 120.600 ;
        RECT 106.210 120.380 106.380 121.790 ;
        RECT 11.950 120.185 90.610 120.355 ;
        RECT 103.950 120.210 106.380 120.380 ;
        RECT 107.960 122.300 118.590 122.470 ;
        RECT 120.020 131.640 126.250 131.800 ;
        RECT 120.020 129.380 120.690 131.640 ;
        RECT 121.360 131.070 125.400 131.240 ;
        RECT 121.020 130.010 121.190 131.010 ;
        RECT 125.570 130.010 125.740 131.010 ;
        RECT 121.360 129.780 125.400 129.950 ;
        RECT 126.080 129.380 126.250 131.640 ;
        RECT 120.020 129.210 126.250 129.380 ;
        RECT 120.020 125.950 120.690 129.210 ;
        RECT 121.360 128.640 125.400 128.810 ;
        RECT 121.020 126.580 121.190 128.580 ;
        RECT 125.570 126.580 125.740 128.580 ;
        RECT 121.360 126.350 125.400 126.520 ;
        RECT 126.080 125.950 126.250 129.210 ;
        RECT 120.020 125.780 126.250 125.950 ;
        RECT 120.020 122.520 120.690 125.780 ;
        RECT 121.360 125.210 125.400 125.380 ;
        RECT 121.020 123.150 121.190 125.150 ;
        RECT 125.570 123.150 125.740 125.150 ;
        RECT 121.360 122.920 125.400 123.090 ;
        RECT 126.080 122.520 126.250 125.780 ;
        RECT 120.020 122.510 126.250 122.520 ;
        RECT 127.840 131.780 137.670 131.820 ;
        RECT 140.540 131.800 146.280 131.810 ;
        RECT 127.840 131.650 138.470 131.780 ;
        RECT 127.840 129.390 128.010 131.650 ;
        RECT 128.735 131.080 136.775 131.250 ;
        RECT 128.350 130.020 128.520 131.020 ;
        RECT 136.990 130.020 137.160 131.020 ;
        RECT 128.735 129.790 136.775 129.960 ;
        RECT 137.500 129.390 138.470 131.650 ;
        RECT 127.840 129.220 138.470 129.390 ;
        RECT 127.840 125.960 128.010 129.220 ;
        RECT 128.735 128.650 136.775 128.820 ;
        RECT 128.350 126.590 128.520 128.590 ;
        RECT 136.990 126.590 137.160 128.590 ;
        RECT 128.735 126.360 136.775 126.530 ;
        RECT 137.500 125.960 138.470 129.220 ;
        RECT 127.840 125.790 138.470 125.960 ;
        RECT 127.840 122.530 128.010 125.790 ;
        RECT 128.735 125.220 136.775 125.390 ;
        RECT 128.350 123.160 128.520 125.160 ;
        RECT 136.990 123.160 137.160 125.160 ;
        RECT 128.735 122.930 136.775 123.100 ;
        RECT 137.500 122.530 138.470 125.790 ;
        RECT 120.020 122.410 126.260 122.510 ;
        RECT 12.035 119.095 13.245 120.185 ;
        RECT 13.415 119.095 14.625 120.185 ;
        RECT 14.855 119.125 15.185 119.970 ;
        RECT 15.355 119.175 15.525 120.185 ;
        RECT 15.695 119.455 16.035 120.015 ;
        RECT 16.265 119.685 16.580 120.185 ;
        RECT 16.760 119.715 17.645 119.885 ;
        RECT 12.035 118.385 12.555 118.925 ;
        RECT 12.725 118.555 13.245 119.095 ;
        RECT 13.415 118.385 13.935 118.925 ;
        RECT 14.105 118.555 14.625 119.095 ;
        RECT 14.795 119.045 15.185 119.125 ;
        RECT 15.695 119.080 16.590 119.455 ;
        RECT 14.795 118.995 15.010 119.045 ;
        RECT 14.795 118.415 14.965 118.995 ;
        RECT 15.695 118.875 15.885 119.080 ;
        RECT 16.760 118.875 16.930 119.715 ;
        RECT 17.870 119.685 18.120 120.015 ;
        RECT 15.135 118.545 15.885 118.875 ;
        RECT 16.055 118.545 16.930 118.875 ;
        RECT 12.035 117.635 13.245 118.385 ;
        RECT 13.415 117.635 14.625 118.385 ;
        RECT 14.795 118.375 15.020 118.415 ;
        RECT 15.685 118.375 15.885 118.545 ;
        RECT 14.795 118.290 15.175 118.375 ;
        RECT 14.845 117.855 15.175 118.290 ;
        RECT 15.345 117.635 15.515 118.245 ;
        RECT 15.685 117.850 16.015 118.375 ;
        RECT 16.275 117.635 16.485 118.165 ;
        RECT 16.760 118.085 16.930 118.545 ;
        RECT 17.100 118.585 17.420 119.545 ;
        RECT 17.590 118.795 17.780 119.515 ;
        RECT 17.950 118.615 18.120 119.685 ;
        RECT 18.290 119.385 18.460 120.185 ;
        RECT 18.630 119.740 19.735 119.910 ;
        RECT 18.630 119.125 18.800 119.740 ;
        RECT 19.945 119.590 20.195 120.015 ;
        RECT 20.365 119.725 20.630 120.185 ;
        RECT 18.970 119.205 19.500 119.570 ;
        RECT 19.945 119.460 20.250 119.590 ;
        RECT 18.290 119.035 18.800 119.125 ;
        RECT 18.290 118.865 19.160 119.035 ;
        RECT 18.290 118.795 18.460 118.865 ;
        RECT 18.580 118.615 18.780 118.645 ;
        RECT 17.100 118.255 17.565 118.585 ;
        RECT 17.950 118.315 18.780 118.615 ;
        RECT 17.950 118.085 18.120 118.315 ;
        RECT 16.760 117.915 17.545 118.085 ;
        RECT 17.715 117.915 18.120 118.085 ;
        RECT 18.300 117.635 18.670 118.135 ;
        RECT 18.990 118.085 19.160 118.865 ;
        RECT 19.330 118.505 19.500 119.205 ;
        RECT 19.670 118.675 19.910 119.270 ;
        RECT 19.330 118.285 19.855 118.505 ;
        RECT 20.080 118.355 20.250 119.460 ;
        RECT 20.025 118.225 20.250 118.355 ;
        RECT 20.420 118.265 20.700 119.215 ;
        RECT 20.025 118.085 20.195 118.225 ;
        RECT 18.990 117.915 19.665 118.085 ;
        RECT 19.860 117.915 20.195 118.085 ;
        RECT 20.365 117.635 20.615 118.095 ;
        RECT 20.870 117.895 21.055 120.015 ;
        RECT 21.225 119.685 21.555 120.185 ;
        RECT 21.725 119.515 21.895 120.015 ;
        RECT 21.230 119.345 21.895 119.515 ;
        RECT 21.230 118.355 21.460 119.345 ;
        RECT 21.630 118.525 21.980 119.175 ;
        RECT 22.155 118.580 22.435 120.015 ;
        RECT 22.605 119.410 23.315 120.185 ;
        RECT 23.485 119.240 23.815 120.015 ;
        RECT 22.665 119.025 23.815 119.240 ;
        RECT 21.230 118.185 21.895 118.355 ;
        RECT 21.225 117.635 21.555 118.015 ;
        RECT 21.725 117.895 21.895 118.185 ;
        RECT 22.155 117.805 22.495 118.580 ;
        RECT 22.665 118.455 22.950 119.025 ;
        RECT 23.135 118.625 23.605 118.855 ;
        RECT 24.010 118.825 24.225 119.940 ;
        RECT 24.405 119.465 24.735 120.185 ;
        RECT 24.515 118.825 24.745 119.165 ;
        RECT 24.915 119.020 25.205 120.185 ;
        RECT 25.465 119.515 25.635 120.015 ;
        RECT 25.805 119.685 26.135 120.185 ;
        RECT 25.465 119.345 26.130 119.515 ;
        RECT 23.775 118.645 24.225 118.825 ;
        RECT 23.775 118.625 24.105 118.645 ;
        RECT 24.415 118.625 24.745 118.825 ;
        RECT 25.380 118.525 25.730 119.175 ;
        RECT 22.665 118.265 23.375 118.455 ;
        RECT 23.075 118.125 23.375 118.265 ;
        RECT 23.565 118.265 24.745 118.455 ;
        RECT 23.565 118.185 23.895 118.265 ;
        RECT 23.075 118.115 23.390 118.125 ;
        RECT 23.075 118.105 23.400 118.115 ;
        RECT 23.075 118.100 23.410 118.105 ;
        RECT 22.665 117.635 22.835 118.095 ;
        RECT 23.075 118.090 23.415 118.100 ;
        RECT 23.075 118.085 23.420 118.090 ;
        RECT 23.075 118.075 23.425 118.085 ;
        RECT 23.075 118.070 23.430 118.075 ;
        RECT 23.075 117.805 23.435 118.070 ;
        RECT 24.065 117.635 24.235 118.095 ;
        RECT 24.405 117.805 24.745 118.265 ;
        RECT 24.915 117.635 25.205 118.360 ;
        RECT 25.900 118.355 26.130 119.345 ;
        RECT 25.465 118.185 26.130 118.355 ;
        RECT 25.465 117.895 25.635 118.185 ;
        RECT 25.805 117.635 26.135 118.015 ;
        RECT 26.305 117.895 26.490 120.015 ;
        RECT 26.730 119.725 26.995 120.185 ;
        RECT 27.165 119.590 27.415 120.015 ;
        RECT 27.625 119.740 28.730 119.910 ;
        RECT 27.110 119.460 27.415 119.590 ;
        RECT 26.660 118.265 26.940 119.215 ;
        RECT 27.110 118.355 27.280 119.460 ;
        RECT 27.450 118.675 27.690 119.270 ;
        RECT 27.860 119.205 28.390 119.570 ;
        RECT 27.860 118.505 28.030 119.205 ;
        RECT 28.560 119.125 28.730 119.740 ;
        RECT 28.900 119.385 29.070 120.185 ;
        RECT 29.240 119.685 29.490 120.015 ;
        RECT 29.715 119.715 30.600 119.885 ;
        RECT 28.560 119.035 29.070 119.125 ;
        RECT 27.110 118.225 27.335 118.355 ;
        RECT 27.505 118.285 28.030 118.505 ;
        RECT 28.200 118.865 29.070 119.035 ;
        RECT 26.745 117.635 26.995 118.095 ;
        RECT 27.165 118.085 27.335 118.225 ;
        RECT 28.200 118.085 28.370 118.865 ;
        RECT 28.900 118.795 29.070 118.865 ;
        RECT 28.580 118.615 28.780 118.645 ;
        RECT 29.240 118.615 29.410 119.685 ;
        RECT 29.580 118.795 29.770 119.515 ;
        RECT 28.580 118.315 29.410 118.615 ;
        RECT 29.940 118.585 30.260 119.545 ;
        RECT 27.165 117.915 27.500 118.085 ;
        RECT 27.695 117.915 28.370 118.085 ;
        RECT 28.690 117.635 29.060 118.135 ;
        RECT 29.240 118.085 29.410 118.315 ;
        RECT 29.795 118.255 30.260 118.585 ;
        RECT 30.430 118.875 30.600 119.715 ;
        RECT 30.780 119.685 31.095 120.185 ;
        RECT 31.325 119.455 31.665 120.015 ;
        RECT 30.770 119.080 31.665 119.455 ;
        RECT 31.835 119.175 32.005 120.185 ;
        RECT 31.475 118.875 31.665 119.080 ;
        RECT 32.175 119.125 32.505 119.970 ;
        RECT 32.175 119.045 32.565 119.125 ;
        RECT 32.350 118.995 32.565 119.045 ;
        RECT 30.430 118.545 31.305 118.875 ;
        RECT 31.475 118.545 32.225 118.875 ;
        RECT 30.430 118.085 30.600 118.545 ;
        RECT 31.475 118.375 31.675 118.545 ;
        RECT 32.395 118.415 32.565 118.995 ;
        RECT 32.340 118.375 32.565 118.415 ;
        RECT 29.240 117.915 29.645 118.085 ;
        RECT 29.815 117.915 30.600 118.085 ;
        RECT 30.875 117.635 31.085 118.165 ;
        RECT 31.345 117.850 31.675 118.375 ;
        RECT 32.185 118.290 32.565 118.375 ;
        RECT 32.735 119.045 33.120 120.015 ;
        RECT 33.290 119.725 33.615 120.185 ;
        RECT 34.135 119.555 34.415 120.015 ;
        RECT 33.290 119.335 34.415 119.555 ;
        RECT 32.735 118.375 33.015 119.045 ;
        RECT 33.290 118.875 33.740 119.335 ;
        RECT 34.605 119.165 35.005 120.015 ;
        RECT 35.405 119.725 35.675 120.185 ;
        RECT 35.845 119.555 36.130 120.015 ;
        RECT 33.185 118.545 33.740 118.875 ;
        RECT 33.910 118.605 35.005 119.165 ;
        RECT 33.290 118.435 33.740 118.545 ;
        RECT 31.845 117.635 32.015 118.245 ;
        RECT 32.185 117.855 32.515 118.290 ;
        RECT 32.735 117.805 33.120 118.375 ;
        RECT 33.290 118.265 34.415 118.435 ;
        RECT 33.290 117.635 33.615 118.095 ;
        RECT 34.135 117.805 34.415 118.265 ;
        RECT 34.605 117.805 35.005 118.605 ;
        RECT 35.175 119.335 36.130 119.555 ;
        RECT 35.175 118.435 35.385 119.335 ;
        RECT 35.555 118.605 36.245 119.165 ;
        RECT 36.875 119.045 37.260 120.015 ;
        RECT 37.430 119.725 37.755 120.185 ;
        RECT 38.275 119.555 38.555 120.015 ;
        RECT 37.430 119.335 38.555 119.555 ;
        RECT 35.175 118.265 36.130 118.435 ;
        RECT 35.405 117.635 35.675 118.095 ;
        RECT 35.845 117.805 36.130 118.265 ;
        RECT 36.875 118.375 37.155 119.045 ;
        RECT 37.430 118.875 37.880 119.335 ;
        RECT 38.745 119.165 39.145 120.015 ;
        RECT 39.545 119.725 39.815 120.185 ;
        RECT 39.985 119.555 40.270 120.015 ;
        RECT 40.555 119.750 45.900 120.185 ;
        RECT 37.325 118.545 37.880 118.875 ;
        RECT 38.050 118.605 39.145 119.165 ;
        RECT 37.430 118.435 37.880 118.545 ;
        RECT 36.875 117.805 37.260 118.375 ;
        RECT 37.430 118.265 38.555 118.435 ;
        RECT 37.430 117.635 37.755 118.095 ;
        RECT 38.275 117.805 38.555 118.265 ;
        RECT 38.745 117.805 39.145 118.605 ;
        RECT 39.315 119.335 40.270 119.555 ;
        RECT 39.315 118.435 39.525 119.335 ;
        RECT 39.695 118.605 40.385 119.165 ;
        RECT 39.315 118.265 40.270 118.435 ;
        RECT 39.545 117.635 39.815 118.095 ;
        RECT 39.985 117.805 40.270 118.265 ;
        RECT 42.140 118.180 42.480 119.010 ;
        RECT 43.960 118.500 44.310 119.750 ;
        RECT 46.075 119.095 49.585 120.185 ;
        RECT 46.075 118.405 47.725 118.925 ;
        RECT 47.895 118.575 49.585 119.095 ;
        RECT 50.675 119.020 50.965 120.185 ;
        RECT 51.225 119.515 51.395 120.015 ;
        RECT 51.565 119.685 51.895 120.185 ;
        RECT 51.225 119.345 51.890 119.515 ;
        RECT 51.140 118.525 51.490 119.175 ;
        RECT 40.555 117.635 45.900 118.180 ;
        RECT 46.075 117.635 49.585 118.405 ;
        RECT 50.675 117.635 50.965 118.360 ;
        RECT 51.660 118.355 51.890 119.345 ;
        RECT 51.225 118.185 51.890 118.355 ;
        RECT 51.225 117.895 51.395 118.185 ;
        RECT 51.565 117.635 51.895 118.015 ;
        RECT 52.065 117.895 52.250 120.015 ;
        RECT 52.490 119.725 52.755 120.185 ;
        RECT 52.925 119.590 53.175 120.015 ;
        RECT 53.385 119.740 54.490 119.910 ;
        RECT 52.870 119.460 53.175 119.590 ;
        RECT 52.420 118.265 52.700 119.215 ;
        RECT 52.870 118.355 53.040 119.460 ;
        RECT 53.210 118.675 53.450 119.270 ;
        RECT 53.620 119.205 54.150 119.570 ;
        RECT 53.620 118.505 53.790 119.205 ;
        RECT 54.320 119.125 54.490 119.740 ;
        RECT 54.660 119.385 54.830 120.185 ;
        RECT 55.000 119.685 55.250 120.015 ;
        RECT 55.475 119.715 56.360 119.885 ;
        RECT 54.320 119.035 54.830 119.125 ;
        RECT 52.870 118.225 53.095 118.355 ;
        RECT 53.265 118.285 53.790 118.505 ;
        RECT 53.960 118.865 54.830 119.035 ;
        RECT 52.505 117.635 52.755 118.095 ;
        RECT 52.925 118.085 53.095 118.225 ;
        RECT 53.960 118.085 54.130 118.865 ;
        RECT 54.660 118.795 54.830 118.865 ;
        RECT 54.340 118.615 54.540 118.645 ;
        RECT 55.000 118.615 55.170 119.685 ;
        RECT 55.340 118.795 55.530 119.515 ;
        RECT 54.340 118.315 55.170 118.615 ;
        RECT 55.700 118.585 56.020 119.545 ;
        RECT 52.925 117.915 53.260 118.085 ;
        RECT 53.455 117.915 54.130 118.085 ;
        RECT 54.450 117.635 54.820 118.135 ;
        RECT 55.000 118.085 55.170 118.315 ;
        RECT 55.555 118.255 56.020 118.585 ;
        RECT 56.190 118.875 56.360 119.715 ;
        RECT 56.540 119.685 56.855 120.185 ;
        RECT 57.085 119.455 57.425 120.015 ;
        RECT 56.530 119.080 57.425 119.455 ;
        RECT 57.595 119.175 57.765 120.185 ;
        RECT 57.235 118.875 57.425 119.080 ;
        RECT 57.935 119.125 58.265 119.970 ;
        RECT 59.045 119.515 59.215 120.015 ;
        RECT 59.385 119.685 59.715 120.185 ;
        RECT 59.045 119.345 59.710 119.515 ;
        RECT 57.935 119.045 58.325 119.125 ;
        RECT 58.110 118.995 58.325 119.045 ;
        RECT 56.190 118.545 57.065 118.875 ;
        RECT 57.235 118.545 57.985 118.875 ;
        RECT 56.190 118.085 56.360 118.545 ;
        RECT 57.235 118.375 57.435 118.545 ;
        RECT 58.155 118.415 58.325 118.995 ;
        RECT 58.960 118.525 59.310 119.175 ;
        RECT 58.100 118.375 58.325 118.415 ;
        RECT 55.000 117.915 55.405 118.085 ;
        RECT 55.575 117.915 56.360 118.085 ;
        RECT 56.635 117.635 56.845 118.165 ;
        RECT 57.105 117.850 57.435 118.375 ;
        RECT 57.945 118.290 58.325 118.375 ;
        RECT 59.480 118.355 59.710 119.345 ;
        RECT 57.605 117.635 57.775 118.245 ;
        RECT 57.945 117.855 58.275 118.290 ;
        RECT 59.045 118.185 59.710 118.355 ;
        RECT 59.045 117.895 59.215 118.185 ;
        RECT 59.385 117.635 59.715 118.015 ;
        RECT 59.885 117.895 60.070 120.015 ;
        RECT 60.310 119.725 60.575 120.185 ;
        RECT 60.745 119.590 60.995 120.015 ;
        RECT 61.205 119.740 62.310 119.910 ;
        RECT 60.690 119.460 60.995 119.590 ;
        RECT 60.240 118.265 60.520 119.215 ;
        RECT 60.690 118.355 60.860 119.460 ;
        RECT 61.030 118.675 61.270 119.270 ;
        RECT 61.440 119.205 61.970 119.570 ;
        RECT 61.440 118.505 61.610 119.205 ;
        RECT 62.140 119.125 62.310 119.740 ;
        RECT 62.480 119.385 62.650 120.185 ;
        RECT 62.820 119.685 63.070 120.015 ;
        RECT 63.295 119.715 64.180 119.885 ;
        RECT 62.140 119.035 62.650 119.125 ;
        RECT 60.690 118.225 60.915 118.355 ;
        RECT 61.085 118.285 61.610 118.505 ;
        RECT 61.780 118.865 62.650 119.035 ;
        RECT 60.325 117.635 60.575 118.095 ;
        RECT 60.745 118.085 60.915 118.225 ;
        RECT 61.780 118.085 61.950 118.865 ;
        RECT 62.480 118.795 62.650 118.865 ;
        RECT 62.160 118.615 62.360 118.645 ;
        RECT 62.820 118.615 62.990 119.685 ;
        RECT 63.160 118.795 63.350 119.515 ;
        RECT 62.160 118.315 62.990 118.615 ;
        RECT 63.520 118.585 63.840 119.545 ;
        RECT 60.745 117.915 61.080 118.085 ;
        RECT 61.275 117.915 61.950 118.085 ;
        RECT 62.270 117.635 62.640 118.135 ;
        RECT 62.820 118.085 62.990 118.315 ;
        RECT 63.375 118.255 63.840 118.585 ;
        RECT 64.010 118.875 64.180 119.715 ;
        RECT 64.360 119.685 64.675 120.185 ;
        RECT 64.905 119.455 65.245 120.015 ;
        RECT 64.350 119.080 65.245 119.455 ;
        RECT 65.415 119.175 65.585 120.185 ;
        RECT 65.055 118.875 65.245 119.080 ;
        RECT 65.755 119.125 66.085 119.970 ;
        RECT 65.755 119.045 66.145 119.125 ;
        RECT 65.930 118.995 66.145 119.045 ;
        RECT 64.010 118.545 64.885 118.875 ;
        RECT 65.055 118.545 65.805 118.875 ;
        RECT 64.010 118.085 64.180 118.545 ;
        RECT 65.055 118.375 65.255 118.545 ;
        RECT 65.975 118.415 66.145 118.995 ;
        RECT 65.920 118.375 66.145 118.415 ;
        RECT 62.820 117.915 63.225 118.085 ;
        RECT 63.395 117.915 64.180 118.085 ;
        RECT 64.455 117.635 64.665 118.165 ;
        RECT 64.925 117.850 65.255 118.375 ;
        RECT 65.765 118.290 66.145 118.375 ;
        RECT 66.315 119.045 66.700 120.015 ;
        RECT 66.870 119.725 67.195 120.185 ;
        RECT 67.715 119.555 67.995 120.015 ;
        RECT 66.870 119.335 67.995 119.555 ;
        RECT 66.315 118.375 66.595 119.045 ;
        RECT 66.870 118.875 67.320 119.335 ;
        RECT 68.185 119.165 68.585 120.015 ;
        RECT 68.985 119.725 69.255 120.185 ;
        RECT 69.425 119.555 69.710 120.015 ;
        RECT 66.765 118.545 67.320 118.875 ;
        RECT 67.490 118.605 68.585 119.165 ;
        RECT 66.870 118.435 67.320 118.545 ;
        RECT 65.425 117.635 65.595 118.245 ;
        RECT 65.765 117.855 66.095 118.290 ;
        RECT 66.315 117.805 66.700 118.375 ;
        RECT 66.870 118.265 67.995 118.435 ;
        RECT 66.870 117.635 67.195 118.095 ;
        RECT 67.715 117.805 67.995 118.265 ;
        RECT 68.185 117.805 68.585 118.605 ;
        RECT 68.755 119.335 69.710 119.555 ;
        RECT 70.000 119.795 70.335 120.015 ;
        RECT 71.340 119.805 71.695 120.185 ;
        RECT 68.755 118.435 68.965 119.335 ;
        RECT 70.000 119.175 70.255 119.795 ;
        RECT 70.505 119.635 70.735 119.675 ;
        RECT 71.865 119.635 72.115 120.015 ;
        RECT 70.505 119.435 72.115 119.635 ;
        RECT 70.505 119.345 70.690 119.435 ;
        RECT 71.280 119.425 72.115 119.435 ;
        RECT 72.365 119.405 72.615 120.185 ;
        RECT 72.785 119.335 73.045 120.015 ;
        RECT 70.845 119.235 71.175 119.265 ;
        RECT 70.845 119.175 72.645 119.235 ;
        RECT 69.135 118.605 69.825 119.165 ;
        RECT 70.000 119.065 72.705 119.175 ;
        RECT 70.000 119.005 71.175 119.065 ;
        RECT 72.505 119.030 72.705 119.065 ;
        RECT 69.995 118.625 70.485 118.825 ;
        RECT 70.675 118.625 71.150 118.835 ;
        RECT 68.755 118.265 69.710 118.435 ;
        RECT 68.985 117.635 69.255 118.095 ;
        RECT 69.425 117.805 69.710 118.265 ;
        RECT 70.000 117.635 70.455 118.400 ;
        RECT 70.930 118.225 71.150 118.625 ;
        RECT 71.395 118.625 71.725 118.835 ;
        RECT 71.395 118.225 71.605 118.625 ;
        RECT 71.895 118.590 72.305 118.895 ;
        RECT 72.535 118.455 72.705 119.030 ;
        RECT 72.435 118.335 72.705 118.455 ;
        RECT 71.860 118.290 72.705 118.335 ;
        RECT 71.860 118.165 72.615 118.290 ;
        RECT 71.860 118.015 72.030 118.165 ;
        RECT 72.875 118.135 73.045 119.335 ;
        RECT 73.215 119.095 75.805 120.185 ;
        RECT 70.730 117.805 72.030 118.015 ;
        RECT 72.285 117.635 72.615 117.995 ;
        RECT 72.785 117.805 73.045 118.135 ;
        RECT 73.215 118.405 74.425 118.925 ;
        RECT 74.595 118.575 75.805 119.095 ;
        RECT 76.435 119.020 76.725 120.185 ;
        RECT 76.895 119.750 82.240 120.185 ;
        RECT 82.415 119.750 87.760 120.185 ;
        RECT 73.215 117.635 75.805 118.405 ;
        RECT 76.435 117.635 76.725 118.360 ;
        RECT 78.480 118.180 78.820 119.010 ;
        RECT 80.300 118.500 80.650 119.750 ;
        RECT 84.000 118.180 84.340 119.010 ;
        RECT 85.820 118.500 86.170 119.750 ;
        RECT 87.935 119.095 89.145 120.185 ;
        RECT 87.935 118.385 88.455 118.925 ;
        RECT 88.625 118.555 89.145 119.095 ;
        RECT 89.315 119.095 90.525 120.185 ;
        RECT 107.960 120.040 108.130 122.300 ;
        RECT 108.855 121.730 116.895 121.900 ;
        RECT 108.470 120.670 108.640 121.670 ;
        RECT 117.110 120.670 117.280 121.670 ;
        RECT 108.855 120.440 116.895 120.610 ;
        RECT 117.620 120.040 118.590 122.300 ;
        RECT 120.010 121.850 126.260 122.410 ;
        RECT 120.010 121.830 125.180 121.850 ;
        RECT 120.010 121.760 124.000 121.830 ;
        RECT 120.010 120.490 121.930 121.760 ;
        RECT 123.440 121.750 124.000 121.760 ;
        RECT 123.670 120.660 124.000 121.750 ;
        RECT 124.370 121.280 125.410 121.450 ;
        RECT 124.370 120.840 125.410 121.010 ;
        RECT 125.580 120.980 125.750 121.310 ;
        RECT 123.830 120.440 124.000 120.660 ;
        RECT 126.090 120.440 126.260 121.850 ;
        RECT 123.830 120.270 126.260 120.440 ;
        RECT 127.840 122.360 138.470 122.530 ;
        RECT 140.050 131.640 146.280 131.800 ;
        RECT 140.050 129.380 140.720 131.640 ;
        RECT 141.390 131.070 145.430 131.240 ;
        RECT 141.050 130.010 141.220 131.010 ;
        RECT 145.600 130.010 145.770 131.010 ;
        RECT 141.390 129.780 145.430 129.950 ;
        RECT 146.110 129.380 146.280 131.640 ;
        RECT 140.050 129.210 146.280 129.380 ;
        RECT 140.050 125.950 140.720 129.210 ;
        RECT 141.390 128.640 145.430 128.810 ;
        RECT 141.050 126.580 141.220 128.580 ;
        RECT 145.600 126.580 145.770 128.580 ;
        RECT 141.390 126.350 145.430 126.520 ;
        RECT 146.110 125.950 146.280 129.210 ;
        RECT 140.050 125.780 146.280 125.950 ;
        RECT 140.050 122.520 140.720 125.780 ;
        RECT 141.390 125.210 145.430 125.380 ;
        RECT 141.050 123.150 141.220 125.150 ;
        RECT 145.600 123.150 145.770 125.150 ;
        RECT 141.390 122.920 145.430 123.090 ;
        RECT 146.110 122.520 146.280 125.780 ;
        RECT 140.050 122.510 146.280 122.520 ;
        RECT 147.870 131.780 157.700 131.820 ;
        RECT 147.870 131.650 158.500 131.780 ;
        RECT 147.870 129.390 148.040 131.650 ;
        RECT 148.765 131.080 156.805 131.250 ;
        RECT 148.380 130.020 148.550 131.020 ;
        RECT 157.020 130.020 157.190 131.020 ;
        RECT 148.765 129.790 156.805 129.960 ;
        RECT 157.530 129.390 158.500 131.650 ;
        RECT 147.870 129.220 158.500 129.390 ;
        RECT 147.870 125.960 148.040 129.220 ;
        RECT 148.765 128.650 156.805 128.820 ;
        RECT 148.380 126.590 148.550 128.590 ;
        RECT 157.020 126.590 157.190 128.590 ;
        RECT 148.765 126.360 156.805 126.530 ;
        RECT 157.530 125.960 158.500 129.220 ;
        RECT 147.870 125.790 158.500 125.960 ;
        RECT 147.870 122.530 148.040 125.790 ;
        RECT 148.765 125.220 156.805 125.390 ;
        RECT 148.380 123.160 148.550 125.160 ;
        RECT 157.020 123.160 157.190 125.160 ;
        RECT 148.765 122.930 156.805 123.100 ;
        RECT 157.530 122.530 158.500 125.790 ;
        RECT 140.050 122.410 146.290 122.510 ;
        RECT 127.840 120.100 128.010 122.360 ;
        RECT 128.735 121.790 136.775 121.960 ;
        RECT 128.350 120.730 128.520 121.730 ;
        RECT 136.990 120.730 137.160 121.730 ;
        RECT 128.735 120.500 136.775 120.670 ;
        RECT 137.500 120.100 138.470 122.360 ;
        RECT 140.040 121.850 146.290 122.410 ;
        RECT 140.040 121.830 145.210 121.850 ;
        RECT 140.040 121.760 144.030 121.830 ;
        RECT 140.040 120.490 141.960 121.760 ;
        RECT 143.470 121.750 144.030 121.760 ;
        RECT 143.700 120.660 144.030 121.750 ;
        RECT 144.400 121.280 145.440 121.450 ;
        RECT 144.400 120.840 145.440 121.010 ;
        RECT 145.610 120.980 145.780 121.310 ;
        RECT 143.860 120.440 144.030 120.660 ;
        RECT 146.120 120.440 146.290 121.850 ;
        RECT 143.860 120.270 146.290 120.440 ;
        RECT 147.870 122.360 158.500 122.530 ;
        RECT 127.840 120.070 138.470 120.100 ;
        RECT 147.870 120.100 148.040 122.360 ;
        RECT 148.765 121.790 156.805 121.960 ;
        RECT 148.380 120.730 148.550 121.730 ;
        RECT 157.020 120.730 157.190 121.730 ;
        RECT 148.765 120.500 156.805 120.670 ;
        RECT 157.530 120.100 158.500 122.360 ;
        RECT 147.870 120.070 158.500 120.100 ;
        RECT 107.960 120.010 118.590 120.040 ;
        RECT 107.930 119.900 118.590 120.010 ;
        RECT 127.810 119.960 138.470 120.070 ;
        RECT 147.840 119.960 158.500 120.070 ;
        RECT 126.060 119.910 138.470 119.960 ;
        RECT 146.090 119.910 158.500 119.960 ;
        RECT 106.180 119.850 118.590 119.900 ;
        RECT 101.840 119.680 118.590 119.850 ;
        RECT 89.315 118.555 89.835 119.095 ;
        RECT 90.005 118.385 90.525 118.925 ;
        RECT 76.895 117.635 82.240 118.180 ;
        RECT 82.415 117.635 87.760 118.180 ;
        RECT 87.935 117.635 89.145 118.385 ;
        RECT 89.315 117.635 90.525 118.385 ;
        RECT 101.840 118.270 102.010 119.680 ;
        RECT 102.380 119.110 105.420 119.280 ;
        RECT 102.380 118.670 105.420 118.840 ;
        RECT 105.635 118.810 105.805 119.140 ;
        RECT 106.140 118.920 118.590 119.680 ;
        RECT 121.720 119.740 138.470 119.910 ;
        RECT 106.140 118.910 118.480 118.920 ;
        RECT 106.140 118.900 112.020 118.910 ;
        RECT 106.140 118.880 106.710 118.900 ;
        RECT 107.930 118.890 112.020 118.900 ;
        RECT 106.150 118.270 106.320 118.880 ;
        RECT 101.840 118.100 106.320 118.270 ;
        RECT 121.720 118.330 121.890 119.740 ;
        RECT 122.260 119.170 125.300 119.340 ;
        RECT 122.260 118.730 125.300 118.900 ;
        RECT 125.515 118.870 125.685 119.200 ;
        RECT 126.020 118.980 138.470 119.740 ;
        RECT 141.750 119.740 158.500 119.910 ;
        RECT 126.020 118.970 138.360 118.980 ;
        RECT 126.020 118.960 131.900 118.970 ;
        RECT 126.020 118.940 126.590 118.960 ;
        RECT 127.810 118.950 131.900 118.960 ;
        RECT 126.030 118.330 126.200 118.940 ;
        RECT 121.720 118.160 126.200 118.330 ;
        RECT 141.750 118.330 141.920 119.740 ;
        RECT 142.290 119.170 145.330 119.340 ;
        RECT 142.290 118.730 145.330 118.900 ;
        RECT 145.545 118.870 145.715 119.200 ;
        RECT 146.050 118.980 158.500 119.740 ;
        RECT 146.050 118.970 158.390 118.980 ;
        RECT 146.050 118.960 151.930 118.970 ;
        RECT 146.050 118.940 146.620 118.960 ;
        RECT 147.840 118.950 151.930 118.960 ;
        RECT 146.060 118.330 146.230 118.940 ;
        RECT 141.750 118.160 146.230 118.330 ;
        RECT 11.950 117.465 90.610 117.635 ;
        RECT 12.035 116.715 13.245 117.465 ;
        RECT 13.415 116.965 13.675 117.295 ;
        RECT 13.885 116.985 14.160 117.465 ;
        RECT 12.035 116.175 12.555 116.715 ;
        RECT 12.725 116.005 13.245 116.545 ;
        RECT 12.035 114.915 13.245 116.005 ;
        RECT 13.415 116.055 13.585 116.965 ;
        RECT 14.370 116.895 14.575 117.295 ;
        RECT 14.745 117.065 15.080 117.465 ;
        RECT 15.255 116.920 20.600 117.465 ;
        RECT 13.755 116.225 14.115 116.805 ;
        RECT 14.370 116.725 15.055 116.895 ;
        RECT 14.295 116.055 14.545 116.555 ;
        RECT 13.415 115.885 14.545 116.055 ;
        RECT 13.415 115.115 13.685 115.885 ;
        RECT 14.715 115.695 15.055 116.725 ;
        RECT 16.840 116.090 17.180 116.920 ;
        RECT 20.775 116.695 22.445 117.465 ;
        RECT 22.640 117.075 22.970 117.465 ;
        RECT 23.140 116.905 23.365 117.285 ;
        RECT 13.855 114.915 14.185 115.695 ;
        RECT 14.390 115.520 15.055 115.695 ;
        RECT 14.390 115.115 14.575 115.520 ;
        RECT 18.660 115.350 19.010 116.600 ;
        RECT 20.775 116.175 21.525 116.695 ;
        RECT 21.695 116.005 22.445 116.525 ;
        RECT 22.625 116.225 22.865 116.875 ;
        RECT 23.035 116.725 23.365 116.905 ;
        RECT 23.035 116.055 23.210 116.725 ;
        RECT 23.565 116.555 23.795 117.175 ;
        RECT 23.975 116.735 24.275 117.465 ;
        RECT 24.455 116.815 24.715 117.295 ;
        RECT 24.885 116.925 25.135 117.465 ;
        RECT 23.380 116.225 23.795 116.555 ;
        RECT 23.975 116.225 24.270 116.555 ;
        RECT 14.745 114.915 15.080 115.340 ;
        RECT 15.255 114.915 20.600 115.350 ;
        RECT 20.775 114.915 22.445 116.005 ;
        RECT 22.625 115.865 23.210 116.055 ;
        RECT 22.625 115.095 22.900 115.865 ;
        RECT 23.380 115.695 24.275 116.025 ;
        RECT 23.070 115.525 24.275 115.695 ;
        RECT 23.070 115.095 23.400 115.525 ;
        RECT 23.570 114.915 23.765 115.355 ;
        RECT 23.945 115.095 24.275 115.525 ;
        RECT 24.455 115.785 24.625 116.815 ;
        RECT 25.305 116.760 25.525 117.245 ;
        RECT 24.795 116.165 25.025 116.560 ;
        RECT 25.195 116.335 25.525 116.760 ;
        RECT 25.695 117.085 26.585 117.255 ;
        RECT 25.695 116.360 25.865 117.085 ;
        RECT 26.035 116.530 26.585 116.915 ;
        RECT 26.755 116.725 27.140 117.295 ;
        RECT 27.310 117.005 27.635 117.465 ;
        RECT 28.155 116.835 28.435 117.295 ;
        RECT 25.695 116.290 26.585 116.360 ;
        RECT 25.690 116.265 26.585 116.290 ;
        RECT 25.680 116.250 26.585 116.265 ;
        RECT 25.675 116.235 26.585 116.250 ;
        RECT 25.665 116.230 26.585 116.235 ;
        RECT 25.660 116.220 26.585 116.230 ;
        RECT 25.655 116.210 26.585 116.220 ;
        RECT 25.645 116.205 26.585 116.210 ;
        RECT 25.635 116.195 26.585 116.205 ;
        RECT 25.625 116.190 26.585 116.195 ;
        RECT 25.625 116.185 25.960 116.190 ;
        RECT 25.610 116.180 25.960 116.185 ;
        RECT 25.595 116.170 25.960 116.180 ;
        RECT 25.570 116.165 25.960 116.170 ;
        RECT 24.795 116.160 25.960 116.165 ;
        RECT 24.795 116.125 25.930 116.160 ;
        RECT 24.795 116.100 25.895 116.125 ;
        RECT 24.795 116.070 25.865 116.100 ;
        RECT 24.795 116.040 25.845 116.070 ;
        RECT 24.795 116.010 25.825 116.040 ;
        RECT 24.795 116.000 25.755 116.010 ;
        RECT 24.795 115.990 25.730 116.000 ;
        RECT 24.795 115.975 25.710 115.990 ;
        RECT 24.795 115.960 25.690 115.975 ;
        RECT 24.900 115.950 25.685 115.960 ;
        RECT 24.900 115.915 25.670 115.950 ;
        RECT 24.455 115.085 24.730 115.785 ;
        RECT 24.900 115.665 25.655 115.915 ;
        RECT 25.825 115.595 26.155 115.840 ;
        RECT 26.325 115.740 26.585 116.190 ;
        RECT 26.755 116.055 27.035 116.725 ;
        RECT 27.310 116.665 28.435 116.835 ;
        RECT 27.310 116.555 27.760 116.665 ;
        RECT 27.205 116.225 27.760 116.555 ;
        RECT 28.625 116.495 29.025 117.295 ;
        RECT 29.425 117.005 29.695 117.465 ;
        RECT 29.865 116.835 30.150 117.295 ;
        RECT 25.970 115.570 26.155 115.595 ;
        RECT 25.970 115.470 26.585 115.570 ;
        RECT 24.900 114.915 25.155 115.460 ;
        RECT 25.325 115.085 25.805 115.425 ;
        RECT 25.980 114.915 26.585 115.470 ;
        RECT 26.755 115.085 27.140 116.055 ;
        RECT 27.310 115.765 27.760 116.225 ;
        RECT 27.930 115.935 29.025 116.495 ;
        RECT 27.310 115.545 28.435 115.765 ;
        RECT 27.310 114.915 27.635 115.375 ;
        RECT 28.155 115.085 28.435 115.545 ;
        RECT 28.625 115.085 29.025 115.935 ;
        RECT 29.195 116.665 30.150 116.835 ;
        RECT 29.195 115.765 29.405 116.665 ;
        RECT 30.455 116.655 30.695 117.465 ;
        RECT 30.865 116.655 31.195 117.295 ;
        RECT 31.365 116.655 31.635 117.465 ;
        RECT 31.815 116.695 34.405 117.465 ;
        RECT 34.585 116.740 34.915 117.250 ;
        RECT 35.085 117.065 35.415 117.465 ;
        RECT 36.465 116.895 36.795 117.235 ;
        RECT 36.965 117.065 37.295 117.465 ;
        RECT 29.575 115.935 30.265 116.495 ;
        RECT 30.435 116.225 30.785 116.475 ;
        RECT 30.955 116.055 31.125 116.655 ;
        RECT 31.295 116.225 31.645 116.475 ;
        RECT 31.815 116.175 33.025 116.695 ;
        RECT 30.445 115.885 31.125 116.055 ;
        RECT 29.195 115.545 30.150 115.765 ;
        RECT 29.425 114.915 29.695 115.375 ;
        RECT 29.865 115.085 30.150 115.545 ;
        RECT 30.445 115.100 30.775 115.885 ;
        RECT 31.305 114.915 31.635 116.055 ;
        RECT 33.195 116.005 34.405 116.525 ;
        RECT 31.815 114.915 34.405 116.005 ;
        RECT 34.585 115.975 34.775 116.740 ;
        RECT 35.085 116.725 37.450 116.895 ;
        RECT 37.795 116.740 38.085 117.465 ;
        RECT 35.085 116.555 35.255 116.725 ;
        RECT 34.945 116.225 35.255 116.555 ;
        RECT 35.425 116.225 35.730 116.555 ;
        RECT 34.585 115.125 34.915 115.975 ;
        RECT 35.085 114.915 35.335 116.055 ;
        RECT 35.515 115.895 35.730 116.225 ;
        RECT 35.905 115.895 36.190 116.555 ;
        RECT 36.385 115.895 36.650 116.555 ;
        RECT 36.865 115.895 37.110 116.555 ;
        RECT 37.280 115.725 37.450 116.725 ;
        RECT 38.715 116.665 39.410 117.295 ;
        RECT 39.615 116.665 39.925 117.465 ;
        RECT 40.210 116.835 40.495 117.295 ;
        RECT 40.665 117.005 40.935 117.465 ;
        RECT 40.210 116.665 41.165 116.835 ;
        RECT 38.735 116.225 39.070 116.475 ;
        RECT 35.525 115.555 36.815 115.725 ;
        RECT 35.525 115.135 35.775 115.555 ;
        RECT 36.005 114.915 36.335 115.385 ;
        RECT 36.565 115.135 36.815 115.555 ;
        RECT 36.995 115.555 37.450 115.725 ;
        RECT 36.995 115.125 37.325 115.555 ;
        RECT 37.795 114.915 38.085 116.080 ;
        RECT 39.240 116.065 39.410 116.665 ;
        RECT 39.580 116.225 39.915 116.495 ;
        RECT 38.715 114.915 38.975 116.055 ;
        RECT 39.145 115.085 39.475 116.065 ;
        RECT 39.645 114.915 39.925 116.055 ;
        RECT 40.095 115.935 40.785 116.495 ;
        RECT 40.955 115.765 41.165 116.665 ;
        RECT 40.210 115.545 41.165 115.765 ;
        RECT 41.335 116.495 41.735 117.295 ;
        RECT 41.925 116.835 42.205 117.295 ;
        RECT 42.725 117.005 43.050 117.465 ;
        RECT 41.925 116.665 43.050 116.835 ;
        RECT 43.220 116.725 43.605 117.295 ;
        RECT 42.600 116.555 43.050 116.665 ;
        RECT 41.335 115.935 42.430 116.495 ;
        RECT 42.600 116.225 43.155 116.555 ;
        RECT 40.210 115.085 40.495 115.545 ;
        RECT 40.665 114.915 40.935 115.375 ;
        RECT 41.335 115.085 41.735 115.935 ;
        RECT 42.600 115.765 43.050 116.225 ;
        RECT 43.325 116.055 43.605 116.725 ;
        RECT 43.775 116.665 44.085 117.465 ;
        RECT 44.290 116.665 44.985 117.295 ;
        RECT 45.155 116.725 45.540 117.295 ;
        RECT 45.710 117.005 46.035 117.465 ;
        RECT 46.555 116.835 46.835 117.295 ;
        RECT 43.785 116.225 44.120 116.495 ;
        RECT 44.290 116.065 44.460 116.665 ;
        RECT 44.630 116.225 44.965 116.475 ;
        RECT 41.925 115.545 43.050 115.765 ;
        RECT 41.925 115.085 42.205 115.545 ;
        RECT 42.725 114.915 43.050 115.375 ;
        RECT 43.220 115.085 43.605 116.055 ;
        RECT 43.775 114.915 44.055 116.055 ;
        RECT 44.225 115.085 44.555 116.065 ;
        RECT 45.155 116.055 45.435 116.725 ;
        RECT 45.710 116.665 46.835 116.835 ;
        RECT 45.710 116.555 46.160 116.665 ;
        RECT 45.605 116.225 46.160 116.555 ;
        RECT 47.025 116.495 47.425 117.295 ;
        RECT 47.825 117.005 48.095 117.465 ;
        RECT 48.265 116.835 48.550 117.295 ;
        RECT 44.725 114.915 44.985 116.055 ;
        RECT 45.155 115.085 45.540 116.055 ;
        RECT 45.710 115.765 46.160 116.225 ;
        RECT 46.330 115.935 47.425 116.495 ;
        RECT 45.710 115.545 46.835 115.765 ;
        RECT 45.710 114.915 46.035 115.375 ;
        RECT 46.555 115.085 46.835 115.545 ;
        RECT 47.025 115.085 47.425 115.935 ;
        RECT 47.595 116.665 48.550 116.835 ;
        RECT 48.925 116.915 49.095 117.205 ;
        RECT 49.265 117.085 49.595 117.465 ;
        RECT 48.925 116.745 49.590 116.915 ;
        RECT 47.595 115.765 47.805 116.665 ;
        RECT 47.975 115.935 48.665 116.495 ;
        RECT 48.840 115.925 49.190 116.575 ;
        RECT 47.595 115.545 48.550 115.765 ;
        RECT 49.360 115.755 49.590 116.745 ;
        RECT 47.825 114.915 48.095 115.375 ;
        RECT 48.265 115.085 48.550 115.545 ;
        RECT 48.925 115.585 49.590 115.755 ;
        RECT 48.925 115.085 49.095 115.585 ;
        RECT 49.265 114.915 49.595 115.415 ;
        RECT 49.765 115.085 49.950 117.205 ;
        RECT 50.205 117.005 50.455 117.465 ;
        RECT 50.625 117.015 50.960 117.185 ;
        RECT 51.155 117.015 51.830 117.185 ;
        RECT 50.625 116.875 50.795 117.015 ;
        RECT 50.120 115.885 50.400 116.835 ;
        RECT 50.570 116.745 50.795 116.875 ;
        RECT 50.570 115.640 50.740 116.745 ;
        RECT 50.965 116.595 51.490 116.815 ;
        RECT 50.910 115.830 51.150 116.425 ;
        RECT 51.320 115.895 51.490 116.595 ;
        RECT 51.660 116.235 51.830 117.015 ;
        RECT 52.150 116.965 52.520 117.465 ;
        RECT 52.700 117.015 53.105 117.185 ;
        RECT 53.275 117.015 54.060 117.185 ;
        RECT 52.700 116.785 52.870 117.015 ;
        RECT 52.040 116.485 52.870 116.785 ;
        RECT 53.255 116.515 53.720 116.845 ;
        RECT 52.040 116.455 52.240 116.485 ;
        RECT 52.360 116.235 52.530 116.305 ;
        RECT 51.660 116.065 52.530 116.235 ;
        RECT 52.020 115.975 52.530 116.065 ;
        RECT 50.570 115.510 50.875 115.640 ;
        RECT 51.320 115.530 51.850 115.895 ;
        RECT 50.190 114.915 50.455 115.375 ;
        RECT 50.625 115.085 50.875 115.510 ;
        RECT 52.020 115.360 52.190 115.975 ;
        RECT 51.085 115.190 52.190 115.360 ;
        RECT 52.360 114.915 52.530 115.715 ;
        RECT 52.700 115.415 52.870 116.485 ;
        RECT 53.040 115.585 53.230 116.305 ;
        RECT 53.400 115.555 53.720 116.515 ;
        RECT 53.890 116.555 54.060 117.015 ;
        RECT 54.335 116.935 54.545 117.465 ;
        RECT 54.805 116.725 55.135 117.250 ;
        RECT 55.305 116.855 55.475 117.465 ;
        RECT 55.645 116.810 55.975 117.245 ;
        RECT 56.195 116.920 61.540 117.465 ;
        RECT 55.645 116.725 56.025 116.810 ;
        RECT 54.935 116.555 55.135 116.725 ;
        RECT 55.800 116.685 56.025 116.725 ;
        RECT 53.890 116.225 54.765 116.555 ;
        RECT 54.935 116.225 55.685 116.555 ;
        RECT 52.700 115.085 52.950 115.415 ;
        RECT 53.890 115.385 54.060 116.225 ;
        RECT 54.935 116.020 55.125 116.225 ;
        RECT 55.855 116.105 56.025 116.685 ;
        RECT 55.810 116.055 56.025 116.105 ;
        RECT 57.780 116.090 58.120 116.920 ;
        RECT 61.715 116.695 63.385 117.465 ;
        RECT 63.555 116.740 63.845 117.465 ;
        RECT 54.230 115.645 55.125 116.020 ;
        RECT 55.635 115.975 56.025 116.055 ;
        RECT 53.175 115.215 54.060 115.385 ;
        RECT 54.240 114.915 54.555 115.415 ;
        RECT 54.785 115.085 55.125 115.645 ;
        RECT 55.295 114.915 55.465 115.925 ;
        RECT 55.635 115.130 55.965 115.975 ;
        RECT 59.600 115.350 59.950 116.600 ;
        RECT 61.715 116.175 62.465 116.695 ;
        RECT 64.475 116.665 65.170 117.295 ;
        RECT 65.375 116.665 65.685 117.465 ;
        RECT 65.855 116.715 67.065 117.465 ;
        RECT 62.635 116.005 63.385 116.525 ;
        RECT 64.495 116.225 64.830 116.475 ;
        RECT 56.195 114.915 61.540 115.350 ;
        RECT 61.715 114.915 63.385 116.005 ;
        RECT 63.555 114.915 63.845 116.080 ;
        RECT 65.000 116.065 65.170 116.665 ;
        RECT 65.340 116.225 65.675 116.495 ;
        RECT 65.855 116.175 66.375 116.715 ;
        RECT 67.255 116.655 67.495 117.465 ;
        RECT 67.665 116.655 67.995 117.295 ;
        RECT 68.165 116.655 68.435 117.465 ;
        RECT 68.615 116.695 70.285 117.465 ;
        RECT 70.920 116.960 71.255 117.465 ;
        RECT 71.425 116.895 71.665 117.270 ;
        RECT 71.945 117.135 72.115 117.280 ;
        RECT 71.945 116.940 72.320 117.135 ;
        RECT 72.680 116.970 73.075 117.465 ;
        RECT 64.475 114.915 64.735 116.055 ;
        RECT 64.905 115.085 65.235 116.065 ;
        RECT 65.405 114.915 65.685 116.055 ;
        RECT 66.545 116.005 67.065 116.545 ;
        RECT 67.235 116.225 67.585 116.475 ;
        RECT 67.755 116.055 67.925 116.655 ;
        RECT 68.095 116.225 68.445 116.475 ;
        RECT 68.615 116.175 69.365 116.695 ;
        RECT 65.855 114.915 67.065 116.005 ;
        RECT 67.245 115.885 67.925 116.055 ;
        RECT 67.245 115.100 67.575 115.885 ;
        RECT 68.105 114.915 68.435 116.055 ;
        RECT 69.535 116.005 70.285 116.525 ;
        RECT 68.615 114.915 70.285 116.005 ;
        RECT 70.975 115.935 71.275 116.785 ;
        RECT 71.445 116.745 71.665 116.895 ;
        RECT 71.445 116.415 71.980 116.745 ;
        RECT 72.150 116.605 72.320 116.940 ;
        RECT 73.245 116.775 73.485 117.295 ;
        RECT 73.675 116.920 79.020 117.465 ;
        RECT 79.195 116.920 84.540 117.465 ;
        RECT 71.445 115.765 71.680 116.415 ;
        RECT 72.150 116.245 73.135 116.605 ;
        RECT 71.005 115.535 71.680 115.765 ;
        RECT 71.850 116.225 73.135 116.245 ;
        RECT 71.850 116.075 72.710 116.225 ;
        RECT 71.005 115.105 71.175 115.535 ;
        RECT 71.345 114.915 71.675 115.365 ;
        RECT 71.850 115.130 72.135 116.075 ;
        RECT 73.310 115.970 73.485 116.775 ;
        RECT 75.260 116.090 75.600 116.920 ;
        RECT 72.310 115.595 73.005 115.905 ;
        RECT 72.315 114.915 73.000 115.385 ;
        RECT 73.180 115.185 73.485 115.970 ;
        RECT 77.080 115.350 77.430 116.600 ;
        RECT 80.780 116.090 81.120 116.920 ;
        RECT 84.715 116.695 87.305 117.465 ;
        RECT 87.565 116.915 87.735 117.295 ;
        RECT 87.950 117.085 88.280 117.465 ;
        RECT 87.565 116.745 88.280 116.915 ;
        RECT 82.600 115.350 82.950 116.600 ;
        RECT 84.715 116.175 85.925 116.695 ;
        RECT 86.095 116.005 87.305 116.525 ;
        RECT 87.475 116.195 87.830 116.565 ;
        RECT 88.110 116.555 88.280 116.745 ;
        RECT 88.450 116.720 88.705 117.295 ;
        RECT 88.110 116.225 88.365 116.555 ;
        RECT 88.110 116.015 88.280 116.225 ;
        RECT 73.675 114.915 79.020 115.350 ;
        RECT 79.195 114.915 84.540 115.350 ;
        RECT 84.715 114.915 87.305 116.005 ;
        RECT 87.565 115.845 88.280 116.015 ;
        RECT 88.535 115.990 88.705 116.720 ;
        RECT 88.880 116.625 89.140 117.465 ;
        RECT 89.315 116.715 90.525 117.465 ;
        RECT 100.580 116.800 106.320 116.810 ;
        RECT 87.565 115.085 87.735 115.845 ;
        RECT 87.950 114.915 88.280 115.675 ;
        RECT 88.450 115.085 88.705 115.990 ;
        RECT 88.880 114.915 89.140 116.065 ;
        RECT 89.315 116.005 89.835 116.545 ;
        RECT 90.005 116.175 90.525 116.715 ;
        RECT 100.090 116.640 106.320 116.800 ;
        RECT 89.315 114.915 90.525 116.005 ;
        RECT 11.950 114.745 90.610 114.915 ;
        RECT 12.035 113.655 13.245 114.745 ;
        RECT 13.415 114.150 13.850 114.575 ;
        RECT 14.020 114.320 14.405 114.745 ;
        RECT 13.415 113.980 14.405 114.150 ;
        RECT 12.035 112.945 12.555 113.485 ;
        RECT 12.725 113.115 13.245 113.655 ;
        RECT 13.415 113.105 13.900 113.810 ;
        RECT 14.070 113.435 14.405 113.980 ;
        RECT 14.575 113.785 15.000 114.575 ;
        RECT 15.170 114.150 15.445 114.575 ;
        RECT 15.615 114.320 16.000 114.745 ;
        RECT 15.170 113.955 16.000 114.150 ;
        RECT 14.575 113.605 15.480 113.785 ;
        RECT 14.070 113.105 14.480 113.435 ;
        RECT 14.650 113.105 15.480 113.605 ;
        RECT 15.650 113.435 16.000 113.955 ;
        RECT 16.170 113.785 16.415 114.575 ;
        RECT 16.605 114.150 16.860 114.575 ;
        RECT 17.030 114.320 17.415 114.745 ;
        RECT 16.605 113.955 17.415 114.150 ;
        RECT 16.170 113.605 16.895 113.785 ;
        RECT 15.650 113.105 16.075 113.435 ;
        RECT 16.245 113.105 16.895 113.605 ;
        RECT 17.065 113.435 17.415 113.955 ;
        RECT 17.585 113.605 17.845 114.575 ;
        RECT 17.065 113.105 17.490 113.435 ;
        RECT 12.035 112.195 13.245 112.945 ;
        RECT 14.070 112.935 14.405 113.105 ;
        RECT 14.650 112.935 15.000 113.105 ;
        RECT 15.650 112.935 16.000 113.105 ;
        RECT 16.245 112.935 16.415 113.105 ;
        RECT 17.065 112.935 17.415 113.105 ;
        RECT 17.660 112.935 17.845 113.605 ;
        RECT 13.415 112.765 14.405 112.935 ;
        RECT 13.415 112.365 13.850 112.765 ;
        RECT 14.020 112.195 14.405 112.595 ;
        RECT 14.575 112.365 15.000 112.935 ;
        RECT 15.190 112.765 16.000 112.935 ;
        RECT 15.190 112.365 15.445 112.765 ;
        RECT 15.615 112.195 16.000 112.595 ;
        RECT 16.170 112.365 16.415 112.935 ;
        RECT 16.605 112.765 17.415 112.935 ;
        RECT 16.605 112.365 16.860 112.765 ;
        RECT 17.030 112.195 17.415 112.595 ;
        RECT 17.585 112.365 17.845 112.935 ;
        RECT 18.015 113.605 18.400 114.575 ;
        RECT 18.570 114.285 18.895 114.745 ;
        RECT 19.415 114.115 19.695 114.575 ;
        RECT 18.570 113.895 19.695 114.115 ;
        RECT 18.015 112.935 18.295 113.605 ;
        RECT 18.570 113.435 19.020 113.895 ;
        RECT 19.885 113.725 20.285 114.575 ;
        RECT 20.685 114.285 20.955 114.745 ;
        RECT 21.125 114.115 21.410 114.575 ;
        RECT 18.465 113.105 19.020 113.435 ;
        RECT 19.190 113.165 20.285 113.725 ;
        RECT 18.570 112.995 19.020 113.105 ;
        RECT 18.015 112.365 18.400 112.935 ;
        RECT 18.570 112.825 19.695 112.995 ;
        RECT 18.570 112.195 18.895 112.655 ;
        RECT 19.415 112.365 19.695 112.825 ;
        RECT 19.885 112.365 20.285 113.165 ;
        RECT 20.455 113.895 21.410 114.115 ;
        RECT 20.455 112.995 20.665 113.895 ;
        RECT 20.835 113.165 21.525 113.725 ;
        RECT 21.695 113.655 24.285 114.745 ;
        RECT 20.455 112.825 21.410 112.995 ;
        RECT 20.685 112.195 20.955 112.655 ;
        RECT 21.125 112.365 21.410 112.825 ;
        RECT 21.695 112.965 22.905 113.485 ;
        RECT 23.075 113.135 24.285 113.655 ;
        RECT 24.915 113.580 25.205 114.745 ;
        RECT 25.375 114.310 30.720 114.745 ;
        RECT 21.695 112.195 24.285 112.965 ;
        RECT 24.915 112.195 25.205 112.920 ;
        RECT 26.960 112.740 27.300 113.570 ;
        RECT 28.780 113.060 29.130 114.310 ;
        RECT 30.895 113.655 32.565 114.745 ;
        RECT 33.285 114.075 33.455 114.575 ;
        RECT 33.625 114.245 33.955 114.745 ;
        RECT 33.285 113.905 33.950 114.075 ;
        RECT 30.895 112.965 31.645 113.485 ;
        RECT 31.815 113.135 32.565 113.655 ;
        RECT 33.200 113.085 33.550 113.735 ;
        RECT 25.375 112.195 30.720 112.740 ;
        RECT 30.895 112.195 32.565 112.965 ;
        RECT 33.720 112.915 33.950 113.905 ;
        RECT 33.285 112.745 33.950 112.915 ;
        RECT 33.285 112.455 33.455 112.745 ;
        RECT 33.625 112.195 33.955 112.575 ;
        RECT 34.125 112.455 34.310 114.575 ;
        RECT 34.550 114.285 34.815 114.745 ;
        RECT 34.985 114.150 35.235 114.575 ;
        RECT 35.445 114.300 36.550 114.470 ;
        RECT 34.930 114.020 35.235 114.150 ;
        RECT 34.480 112.825 34.760 113.775 ;
        RECT 34.930 112.915 35.100 114.020 ;
        RECT 35.270 113.235 35.510 113.830 ;
        RECT 35.680 113.765 36.210 114.130 ;
        RECT 35.680 113.065 35.850 113.765 ;
        RECT 36.380 113.685 36.550 114.300 ;
        RECT 36.720 113.945 36.890 114.745 ;
        RECT 37.060 114.245 37.310 114.575 ;
        RECT 37.535 114.275 38.420 114.445 ;
        RECT 36.380 113.595 36.890 113.685 ;
        RECT 34.930 112.785 35.155 112.915 ;
        RECT 35.325 112.845 35.850 113.065 ;
        RECT 36.020 113.425 36.890 113.595 ;
        RECT 34.565 112.195 34.815 112.655 ;
        RECT 34.985 112.645 35.155 112.785 ;
        RECT 36.020 112.645 36.190 113.425 ;
        RECT 36.720 113.355 36.890 113.425 ;
        RECT 36.400 113.175 36.600 113.205 ;
        RECT 37.060 113.175 37.230 114.245 ;
        RECT 37.400 113.355 37.590 114.075 ;
        RECT 36.400 112.875 37.230 113.175 ;
        RECT 37.760 113.145 38.080 114.105 ;
        RECT 34.985 112.475 35.320 112.645 ;
        RECT 35.515 112.475 36.190 112.645 ;
        RECT 36.510 112.195 36.880 112.695 ;
        RECT 37.060 112.645 37.230 112.875 ;
        RECT 37.615 112.815 38.080 113.145 ;
        RECT 38.250 113.435 38.420 114.275 ;
        RECT 38.600 114.245 38.915 114.745 ;
        RECT 39.145 114.015 39.485 114.575 ;
        RECT 38.590 113.640 39.485 114.015 ;
        RECT 39.655 113.735 39.825 114.745 ;
        RECT 39.295 113.435 39.485 113.640 ;
        RECT 39.995 113.685 40.325 114.530 ;
        RECT 39.995 113.605 40.385 113.685 ;
        RECT 40.170 113.555 40.385 113.605 ;
        RECT 38.250 113.105 39.125 113.435 ;
        RECT 39.295 113.105 40.045 113.435 ;
        RECT 38.250 112.645 38.420 113.105 ;
        RECT 39.295 112.935 39.495 113.105 ;
        RECT 40.215 112.975 40.385 113.555 ;
        RECT 40.160 112.935 40.385 112.975 ;
        RECT 37.060 112.475 37.465 112.645 ;
        RECT 37.635 112.475 38.420 112.645 ;
        RECT 38.695 112.195 38.905 112.725 ;
        RECT 39.165 112.410 39.495 112.935 ;
        RECT 40.005 112.850 40.385 112.935 ;
        RECT 39.665 112.195 39.835 112.805 ;
        RECT 40.005 112.415 40.335 112.850 ;
        RECT 40.565 112.375 40.825 114.565 ;
        RECT 40.995 114.015 41.335 114.745 ;
        RECT 41.515 113.835 41.785 114.565 ;
        RECT 41.015 113.615 41.785 113.835 ;
        RECT 41.965 113.855 42.195 114.565 ;
        RECT 42.365 114.035 42.695 114.745 ;
        RECT 42.865 113.855 43.125 114.565 ;
        RECT 43.405 114.075 43.575 114.575 ;
        RECT 43.745 114.245 44.075 114.745 ;
        RECT 43.405 113.905 44.070 114.075 ;
        RECT 41.965 113.615 43.125 113.855 ;
        RECT 41.015 112.945 41.305 113.615 ;
        RECT 41.485 113.125 41.950 113.435 ;
        RECT 42.130 113.125 42.655 113.435 ;
        RECT 41.015 112.745 42.245 112.945 ;
        RECT 41.085 112.195 41.755 112.565 ;
        RECT 41.935 112.375 42.245 112.745 ;
        RECT 42.425 112.485 42.655 113.125 ;
        RECT 42.835 113.105 43.135 113.435 ;
        RECT 43.320 113.085 43.670 113.735 ;
        RECT 42.835 112.195 43.125 112.925 ;
        RECT 43.840 112.915 44.070 113.905 ;
        RECT 43.405 112.745 44.070 112.915 ;
        RECT 43.405 112.455 43.575 112.745 ;
        RECT 43.745 112.195 44.075 112.575 ;
        RECT 44.245 112.455 44.430 114.575 ;
        RECT 44.670 114.285 44.935 114.745 ;
        RECT 45.105 114.150 45.355 114.575 ;
        RECT 45.565 114.300 46.670 114.470 ;
        RECT 45.050 114.020 45.355 114.150 ;
        RECT 44.600 112.825 44.880 113.775 ;
        RECT 45.050 112.915 45.220 114.020 ;
        RECT 45.390 113.235 45.630 113.830 ;
        RECT 45.800 113.765 46.330 114.130 ;
        RECT 45.800 113.065 45.970 113.765 ;
        RECT 46.500 113.685 46.670 114.300 ;
        RECT 46.840 113.945 47.010 114.745 ;
        RECT 47.180 114.245 47.430 114.575 ;
        RECT 47.655 114.275 48.540 114.445 ;
        RECT 46.500 113.595 47.010 113.685 ;
        RECT 45.050 112.785 45.275 112.915 ;
        RECT 45.445 112.845 45.970 113.065 ;
        RECT 46.140 113.425 47.010 113.595 ;
        RECT 44.685 112.195 44.935 112.655 ;
        RECT 45.105 112.645 45.275 112.785 ;
        RECT 46.140 112.645 46.310 113.425 ;
        RECT 46.840 113.355 47.010 113.425 ;
        RECT 46.520 113.175 46.720 113.205 ;
        RECT 47.180 113.175 47.350 114.245 ;
        RECT 47.520 113.355 47.710 114.075 ;
        RECT 46.520 112.875 47.350 113.175 ;
        RECT 47.880 113.145 48.200 114.105 ;
        RECT 45.105 112.475 45.440 112.645 ;
        RECT 45.635 112.475 46.310 112.645 ;
        RECT 46.630 112.195 47.000 112.695 ;
        RECT 47.180 112.645 47.350 112.875 ;
        RECT 47.735 112.815 48.200 113.145 ;
        RECT 48.370 113.435 48.540 114.275 ;
        RECT 48.720 114.245 49.035 114.745 ;
        RECT 49.265 114.015 49.605 114.575 ;
        RECT 48.710 113.640 49.605 114.015 ;
        RECT 49.775 113.735 49.945 114.745 ;
        RECT 49.415 113.435 49.605 113.640 ;
        RECT 50.115 113.685 50.445 114.530 ;
        RECT 50.115 113.605 50.505 113.685 ;
        RECT 50.290 113.555 50.505 113.605 ;
        RECT 50.675 113.580 50.965 114.745 ;
        RECT 51.135 113.655 53.725 114.745 ;
        RECT 53.895 114.235 54.155 114.745 ;
        RECT 48.370 113.105 49.245 113.435 ;
        RECT 49.415 113.105 50.165 113.435 ;
        RECT 48.370 112.645 48.540 113.105 ;
        RECT 49.415 112.935 49.615 113.105 ;
        RECT 50.335 112.975 50.505 113.555 ;
        RECT 50.280 112.935 50.505 112.975 ;
        RECT 47.180 112.475 47.585 112.645 ;
        RECT 47.755 112.475 48.540 112.645 ;
        RECT 48.815 112.195 49.025 112.725 ;
        RECT 49.285 112.410 49.615 112.935 ;
        RECT 50.125 112.850 50.505 112.935 ;
        RECT 51.135 112.965 52.345 113.485 ;
        RECT 52.515 113.135 53.725 113.655 ;
        RECT 53.895 113.185 54.235 114.065 ;
        RECT 54.405 113.355 54.575 114.575 ;
        RECT 54.815 114.240 55.430 114.745 ;
        RECT 54.815 113.705 55.065 114.070 ;
        RECT 55.235 114.065 55.430 114.240 ;
        RECT 55.600 114.235 56.075 114.575 ;
        RECT 56.245 114.200 56.460 114.745 ;
        RECT 55.235 113.875 55.565 114.065 ;
        RECT 55.785 113.705 56.500 114.000 ;
        RECT 56.670 113.875 56.945 114.575 ;
        RECT 57.205 114.075 57.375 114.575 ;
        RECT 57.545 114.245 57.875 114.745 ;
        RECT 57.205 113.905 57.870 114.075 ;
        RECT 54.815 113.535 56.605 113.705 ;
        RECT 54.405 113.105 55.200 113.355 ;
        RECT 54.405 113.015 54.655 113.105 ;
        RECT 49.785 112.195 49.955 112.805 ;
        RECT 50.125 112.415 50.455 112.850 ;
        RECT 50.675 112.195 50.965 112.920 ;
        RECT 51.135 112.195 53.725 112.965 ;
        RECT 53.895 112.195 54.155 113.015 ;
        RECT 54.325 112.595 54.655 113.015 ;
        RECT 55.370 112.680 55.625 113.535 ;
        RECT 54.835 112.415 55.625 112.680 ;
        RECT 55.795 112.835 56.205 113.355 ;
        RECT 56.375 113.105 56.605 113.535 ;
        RECT 56.775 112.845 56.945 113.875 ;
        RECT 57.120 113.085 57.470 113.735 ;
        RECT 57.640 112.915 57.870 113.905 ;
        RECT 55.795 112.415 55.995 112.835 ;
        RECT 56.185 112.195 56.515 112.655 ;
        RECT 56.685 112.365 56.945 112.845 ;
        RECT 57.205 112.745 57.870 112.915 ;
        RECT 57.205 112.455 57.375 112.745 ;
        RECT 57.545 112.195 57.875 112.575 ;
        RECT 58.045 112.455 58.230 114.575 ;
        RECT 58.470 114.285 58.735 114.745 ;
        RECT 58.905 114.150 59.155 114.575 ;
        RECT 59.365 114.300 60.470 114.470 ;
        RECT 58.850 114.020 59.155 114.150 ;
        RECT 58.400 112.825 58.680 113.775 ;
        RECT 58.850 112.915 59.020 114.020 ;
        RECT 59.190 113.235 59.430 113.830 ;
        RECT 59.600 113.765 60.130 114.130 ;
        RECT 59.600 113.065 59.770 113.765 ;
        RECT 60.300 113.685 60.470 114.300 ;
        RECT 60.640 113.945 60.810 114.745 ;
        RECT 60.980 114.245 61.230 114.575 ;
        RECT 61.455 114.275 62.340 114.445 ;
        RECT 60.300 113.595 60.810 113.685 ;
        RECT 58.850 112.785 59.075 112.915 ;
        RECT 59.245 112.845 59.770 113.065 ;
        RECT 59.940 113.425 60.810 113.595 ;
        RECT 58.485 112.195 58.735 112.655 ;
        RECT 58.905 112.645 59.075 112.785 ;
        RECT 59.940 112.645 60.110 113.425 ;
        RECT 60.640 113.355 60.810 113.425 ;
        RECT 60.320 113.175 60.520 113.205 ;
        RECT 60.980 113.175 61.150 114.245 ;
        RECT 61.320 113.355 61.510 114.075 ;
        RECT 60.320 112.875 61.150 113.175 ;
        RECT 61.680 113.145 62.000 114.105 ;
        RECT 58.905 112.475 59.240 112.645 ;
        RECT 59.435 112.475 60.110 112.645 ;
        RECT 60.430 112.195 60.800 112.695 ;
        RECT 60.980 112.645 61.150 112.875 ;
        RECT 61.535 112.815 62.000 113.145 ;
        RECT 62.170 113.435 62.340 114.275 ;
        RECT 62.520 114.245 62.835 114.745 ;
        RECT 63.065 114.015 63.405 114.575 ;
        RECT 62.510 113.640 63.405 114.015 ;
        RECT 63.575 113.735 63.745 114.745 ;
        RECT 63.215 113.435 63.405 113.640 ;
        RECT 63.915 113.685 64.245 114.530 ;
        RECT 64.485 113.775 64.815 114.560 ;
        RECT 63.915 113.605 64.305 113.685 ;
        RECT 64.485 113.605 65.165 113.775 ;
        RECT 65.345 113.605 65.675 114.745 ;
        RECT 65.855 113.655 67.065 114.745 ;
        RECT 64.090 113.555 64.305 113.605 ;
        RECT 62.170 113.105 63.045 113.435 ;
        RECT 63.215 113.105 63.965 113.435 ;
        RECT 62.170 112.645 62.340 113.105 ;
        RECT 63.215 112.935 63.415 113.105 ;
        RECT 64.135 112.975 64.305 113.555 ;
        RECT 64.475 113.185 64.825 113.435 ;
        RECT 64.995 113.005 65.165 113.605 ;
        RECT 65.335 113.185 65.685 113.435 ;
        RECT 64.080 112.935 64.305 112.975 ;
        RECT 60.980 112.475 61.385 112.645 ;
        RECT 61.555 112.475 62.340 112.645 ;
        RECT 62.615 112.195 62.825 112.725 ;
        RECT 63.085 112.410 63.415 112.935 ;
        RECT 63.925 112.850 64.305 112.935 ;
        RECT 63.585 112.195 63.755 112.805 ;
        RECT 63.925 112.415 64.255 112.850 ;
        RECT 64.495 112.195 64.735 113.005 ;
        RECT 64.905 112.365 65.235 113.005 ;
        RECT 65.405 112.195 65.675 113.005 ;
        RECT 65.855 112.945 66.375 113.485 ;
        RECT 66.545 113.115 67.065 113.655 ;
        RECT 67.295 113.605 67.505 114.745 ;
        RECT 67.675 113.595 68.005 114.575 ;
        RECT 68.175 113.605 68.405 114.745 ;
        RECT 68.675 113.685 69.005 114.530 ;
        RECT 69.175 113.735 69.345 114.745 ;
        RECT 69.515 114.015 69.855 114.575 ;
        RECT 70.085 114.245 70.400 114.745 ;
        RECT 70.580 114.275 71.465 114.445 ;
        RECT 68.615 113.605 69.005 113.685 ;
        RECT 69.515 113.640 70.410 114.015 ;
        RECT 65.855 112.195 67.065 112.945 ;
        RECT 67.295 112.195 67.505 113.015 ;
        RECT 67.675 112.995 67.925 113.595 ;
        RECT 68.615 113.555 68.830 113.605 ;
        RECT 68.095 113.185 68.425 113.435 ;
        RECT 67.675 112.365 68.005 112.995 ;
        RECT 68.175 112.195 68.405 113.015 ;
        RECT 68.615 112.975 68.785 113.555 ;
        RECT 69.515 113.435 69.705 113.640 ;
        RECT 70.580 113.435 70.750 114.275 ;
        RECT 71.690 114.245 71.940 114.575 ;
        RECT 68.955 113.105 69.705 113.435 ;
        RECT 69.875 113.105 70.750 113.435 ;
        RECT 68.615 112.935 68.840 112.975 ;
        RECT 69.505 112.935 69.705 113.105 ;
        RECT 68.615 112.850 68.995 112.935 ;
        RECT 68.665 112.415 68.995 112.850 ;
        RECT 69.165 112.195 69.335 112.805 ;
        RECT 69.505 112.410 69.835 112.935 ;
        RECT 70.095 112.195 70.305 112.725 ;
        RECT 70.580 112.645 70.750 113.105 ;
        RECT 70.920 113.145 71.240 114.105 ;
        RECT 71.410 113.355 71.600 114.075 ;
        RECT 71.770 113.175 71.940 114.245 ;
        RECT 72.110 113.945 72.280 114.745 ;
        RECT 72.450 114.300 73.555 114.470 ;
        RECT 72.450 113.685 72.620 114.300 ;
        RECT 73.765 114.150 74.015 114.575 ;
        RECT 74.185 114.285 74.450 114.745 ;
        RECT 72.790 113.765 73.320 114.130 ;
        RECT 73.765 114.020 74.070 114.150 ;
        RECT 72.110 113.595 72.620 113.685 ;
        RECT 72.110 113.425 72.980 113.595 ;
        RECT 72.110 113.355 72.280 113.425 ;
        RECT 72.400 113.175 72.600 113.205 ;
        RECT 70.920 112.815 71.385 113.145 ;
        RECT 71.770 112.875 72.600 113.175 ;
        RECT 71.770 112.645 71.940 112.875 ;
        RECT 70.580 112.475 71.365 112.645 ;
        RECT 71.535 112.475 71.940 112.645 ;
        RECT 72.120 112.195 72.490 112.695 ;
        RECT 72.810 112.645 72.980 113.425 ;
        RECT 73.150 113.065 73.320 113.765 ;
        RECT 73.490 113.235 73.730 113.830 ;
        RECT 73.150 112.845 73.675 113.065 ;
        RECT 73.900 112.915 74.070 114.020 ;
        RECT 73.845 112.785 74.070 112.915 ;
        RECT 74.240 112.825 74.520 113.775 ;
        RECT 73.845 112.645 74.015 112.785 ;
        RECT 72.810 112.475 73.485 112.645 ;
        RECT 73.680 112.475 74.015 112.645 ;
        RECT 74.185 112.195 74.435 112.655 ;
        RECT 74.690 112.455 74.875 114.575 ;
        RECT 75.045 114.245 75.375 114.745 ;
        RECT 75.545 114.075 75.715 114.575 ;
        RECT 75.050 113.905 75.715 114.075 ;
        RECT 75.050 112.915 75.280 113.905 ;
        RECT 75.450 113.085 75.800 113.735 ;
        RECT 76.435 113.580 76.725 114.745 ;
        RECT 76.895 114.310 82.240 114.745 ;
        RECT 75.050 112.745 75.715 112.915 ;
        RECT 75.045 112.195 75.375 112.575 ;
        RECT 75.545 112.455 75.715 112.745 ;
        RECT 76.435 112.195 76.725 112.920 ;
        RECT 78.480 112.740 78.820 113.570 ;
        RECT 80.300 113.060 80.650 114.310 ;
        RECT 82.415 113.655 85.925 114.745 ;
        RECT 82.415 112.965 84.065 113.485 ;
        RECT 84.235 113.135 85.925 113.655 ;
        RECT 86.185 113.815 86.355 114.575 ;
        RECT 86.535 113.985 86.865 114.745 ;
        RECT 86.185 113.645 86.850 113.815 ;
        RECT 87.035 113.670 87.305 114.575 ;
        RECT 86.680 113.500 86.850 113.645 ;
        RECT 86.115 113.095 86.445 113.465 ;
        RECT 86.680 113.170 86.965 113.500 ;
        RECT 76.895 112.195 82.240 112.740 ;
        RECT 82.415 112.195 85.925 112.965 ;
        RECT 86.680 112.915 86.850 113.170 ;
        RECT 86.185 112.745 86.850 112.915 ;
        RECT 87.135 112.870 87.305 113.670 ;
        RECT 87.565 113.815 87.735 114.575 ;
        RECT 87.950 113.985 88.280 114.745 ;
        RECT 87.565 113.645 88.280 113.815 ;
        RECT 88.450 113.670 88.705 114.575 ;
        RECT 87.475 113.095 87.830 113.465 ;
        RECT 88.110 113.435 88.280 113.645 ;
        RECT 88.110 113.105 88.365 113.435 ;
        RECT 88.110 112.915 88.280 113.105 ;
        RECT 88.535 112.940 88.705 113.670 ;
        RECT 88.880 113.595 89.140 114.745 ;
        RECT 89.315 113.655 90.525 114.745 ;
        RECT 100.090 114.380 100.760 116.640 ;
        RECT 101.430 116.070 105.470 116.240 ;
        RECT 101.090 115.010 101.260 116.010 ;
        RECT 105.640 115.010 105.810 116.010 ;
        RECT 101.430 114.780 105.470 114.950 ;
        RECT 106.150 114.380 106.320 116.640 ;
        RECT 100.090 114.210 106.320 114.380 ;
        RECT 89.315 113.115 89.835 113.655 ;
        RECT 86.185 112.365 86.355 112.745 ;
        RECT 86.535 112.195 86.865 112.575 ;
        RECT 87.045 112.365 87.305 112.870 ;
        RECT 87.565 112.745 88.280 112.915 ;
        RECT 87.565 112.365 87.735 112.745 ;
        RECT 87.950 112.195 88.280 112.575 ;
        RECT 88.450 112.365 88.705 112.940 ;
        RECT 88.880 112.195 89.140 113.035 ;
        RECT 90.005 112.945 90.525 113.485 ;
        RECT 89.315 112.195 90.525 112.945 ;
        RECT 11.950 112.025 90.610 112.195 ;
        RECT 12.035 111.275 13.245 112.025 ;
        RECT 13.415 111.275 14.625 112.025 ;
        RECT 14.800 111.495 15.090 111.845 ;
        RECT 15.285 111.665 15.615 112.025 ;
        RECT 15.785 111.495 16.015 111.800 ;
        RECT 14.800 111.325 16.015 111.495 ;
        RECT 12.035 110.735 12.555 111.275 ;
        RECT 12.725 110.565 13.245 111.105 ;
        RECT 13.415 110.735 13.935 111.275 ;
        RECT 16.205 111.155 16.375 111.720 ;
        RECT 16.750 111.395 17.035 111.855 ;
        RECT 17.205 111.565 17.475 112.025 ;
        RECT 16.750 111.225 17.705 111.395 ;
        RECT 14.105 110.565 14.625 111.105 ;
        RECT 14.860 111.005 15.120 111.115 ;
        RECT 14.855 110.835 15.120 111.005 ;
        RECT 14.860 110.785 15.120 110.835 ;
        RECT 15.300 110.785 15.685 111.115 ;
        RECT 15.855 110.985 16.375 111.155 ;
        RECT 12.035 109.475 13.245 110.565 ;
        RECT 13.415 109.475 14.625 110.565 ;
        RECT 14.800 109.475 15.120 110.615 ;
        RECT 15.300 109.735 15.495 110.785 ;
        RECT 15.855 110.605 16.025 110.985 ;
        RECT 15.675 110.325 16.025 110.605 ;
        RECT 16.215 110.455 16.460 110.815 ;
        RECT 16.635 110.495 17.325 111.055 ;
        RECT 17.495 110.325 17.705 111.225 ;
        RECT 15.675 109.645 16.005 110.325 ;
        RECT 16.205 109.475 16.460 110.275 ;
        RECT 16.750 110.105 17.705 110.325 ;
        RECT 17.875 111.055 18.275 111.855 ;
        RECT 18.465 111.395 18.745 111.855 ;
        RECT 19.265 111.565 19.590 112.025 ;
        RECT 18.465 111.225 19.590 111.395 ;
        RECT 19.760 111.285 20.145 111.855 ;
        RECT 20.405 111.475 20.575 111.765 ;
        RECT 20.745 111.645 21.075 112.025 ;
        RECT 20.405 111.305 21.070 111.475 ;
        RECT 19.140 111.115 19.590 111.225 ;
        RECT 17.875 110.495 18.970 111.055 ;
        RECT 19.140 110.785 19.695 111.115 ;
        RECT 16.750 109.645 17.035 110.105 ;
        RECT 17.205 109.475 17.475 109.935 ;
        RECT 17.875 109.645 18.275 110.495 ;
        RECT 19.140 110.325 19.590 110.785 ;
        RECT 19.865 110.615 20.145 111.285 ;
        RECT 18.465 110.105 19.590 110.325 ;
        RECT 18.465 109.645 18.745 110.105 ;
        RECT 19.265 109.475 19.590 109.935 ;
        RECT 19.760 109.645 20.145 110.615 ;
        RECT 20.320 110.485 20.670 111.135 ;
        RECT 20.840 110.315 21.070 111.305 ;
        RECT 20.405 110.145 21.070 110.315 ;
        RECT 20.405 109.645 20.575 110.145 ;
        RECT 20.745 109.475 21.075 109.975 ;
        RECT 21.245 109.645 21.430 111.765 ;
        RECT 21.685 111.565 21.935 112.025 ;
        RECT 22.105 111.575 22.440 111.745 ;
        RECT 22.635 111.575 23.310 111.745 ;
        RECT 22.105 111.435 22.275 111.575 ;
        RECT 21.600 110.445 21.880 111.395 ;
        RECT 22.050 111.305 22.275 111.435 ;
        RECT 22.050 110.200 22.220 111.305 ;
        RECT 22.445 111.155 22.970 111.375 ;
        RECT 22.390 110.390 22.630 110.985 ;
        RECT 22.800 110.455 22.970 111.155 ;
        RECT 23.140 110.795 23.310 111.575 ;
        RECT 23.630 111.525 24.000 112.025 ;
        RECT 24.180 111.575 24.585 111.745 ;
        RECT 24.755 111.575 25.540 111.745 ;
        RECT 24.180 111.345 24.350 111.575 ;
        RECT 23.520 111.045 24.350 111.345 ;
        RECT 24.735 111.075 25.200 111.405 ;
        RECT 23.520 111.015 23.720 111.045 ;
        RECT 23.840 110.795 24.010 110.865 ;
        RECT 23.140 110.625 24.010 110.795 ;
        RECT 23.500 110.535 24.010 110.625 ;
        RECT 22.050 110.070 22.355 110.200 ;
        RECT 22.800 110.090 23.330 110.455 ;
        RECT 21.670 109.475 21.935 109.935 ;
        RECT 22.105 109.645 22.355 110.070 ;
        RECT 23.500 109.920 23.670 110.535 ;
        RECT 22.565 109.750 23.670 109.920 ;
        RECT 23.840 109.475 24.010 110.275 ;
        RECT 24.180 109.975 24.350 111.045 ;
        RECT 24.520 110.145 24.710 110.865 ;
        RECT 24.880 110.115 25.200 111.075 ;
        RECT 25.370 111.115 25.540 111.575 ;
        RECT 25.815 111.495 26.025 112.025 ;
        RECT 26.285 111.285 26.615 111.810 ;
        RECT 26.785 111.415 26.955 112.025 ;
        RECT 27.125 111.370 27.455 111.805 ;
        RECT 27.125 111.285 27.505 111.370 ;
        RECT 26.415 111.115 26.615 111.285 ;
        RECT 27.280 111.245 27.505 111.285 ;
        RECT 25.370 110.785 26.245 111.115 ;
        RECT 26.415 110.785 27.165 111.115 ;
        RECT 24.180 109.645 24.430 109.975 ;
        RECT 25.370 109.945 25.540 110.785 ;
        RECT 26.415 110.580 26.605 110.785 ;
        RECT 27.335 110.665 27.505 111.245 ;
        RECT 27.695 111.215 27.935 112.025 ;
        RECT 28.105 111.215 28.435 111.855 ;
        RECT 28.605 111.215 28.875 112.025 ;
        RECT 30.065 111.475 30.235 111.765 ;
        RECT 30.405 111.645 30.735 112.025 ;
        RECT 30.065 111.305 30.730 111.475 ;
        RECT 27.675 110.785 28.025 111.035 ;
        RECT 27.290 110.615 27.505 110.665 ;
        RECT 28.195 110.615 28.365 111.215 ;
        RECT 28.535 110.785 28.885 111.035 ;
        RECT 25.710 110.205 26.605 110.580 ;
        RECT 27.115 110.535 27.505 110.615 ;
        RECT 24.655 109.775 25.540 109.945 ;
        RECT 25.720 109.475 26.035 109.975 ;
        RECT 26.265 109.645 26.605 110.205 ;
        RECT 26.775 109.475 26.945 110.485 ;
        RECT 27.115 109.690 27.445 110.535 ;
        RECT 27.685 110.445 28.365 110.615 ;
        RECT 27.685 109.660 28.015 110.445 ;
        RECT 28.545 109.475 28.875 110.615 ;
        RECT 29.980 110.485 30.330 111.135 ;
        RECT 30.500 110.315 30.730 111.305 ;
        RECT 30.065 110.145 30.730 110.315 ;
        RECT 30.065 109.645 30.235 110.145 ;
        RECT 30.405 109.475 30.735 109.975 ;
        RECT 30.905 109.645 31.090 111.765 ;
        RECT 31.345 111.565 31.595 112.025 ;
        RECT 31.765 111.575 32.100 111.745 ;
        RECT 32.295 111.575 32.970 111.745 ;
        RECT 31.765 111.435 31.935 111.575 ;
        RECT 31.260 110.445 31.540 111.395 ;
        RECT 31.710 111.305 31.935 111.435 ;
        RECT 31.710 110.200 31.880 111.305 ;
        RECT 32.105 111.155 32.630 111.375 ;
        RECT 32.050 110.390 32.290 110.985 ;
        RECT 32.460 110.455 32.630 111.155 ;
        RECT 32.800 110.795 32.970 111.575 ;
        RECT 33.290 111.525 33.660 112.025 ;
        RECT 33.840 111.575 34.245 111.745 ;
        RECT 34.415 111.575 35.200 111.745 ;
        RECT 33.840 111.345 34.010 111.575 ;
        RECT 33.180 111.045 34.010 111.345 ;
        RECT 34.395 111.075 34.860 111.405 ;
        RECT 33.180 111.015 33.380 111.045 ;
        RECT 33.500 110.795 33.670 110.865 ;
        RECT 32.800 110.625 33.670 110.795 ;
        RECT 33.160 110.535 33.670 110.625 ;
        RECT 31.710 110.070 32.015 110.200 ;
        RECT 32.460 110.090 32.990 110.455 ;
        RECT 31.330 109.475 31.595 109.935 ;
        RECT 31.765 109.645 32.015 110.070 ;
        RECT 33.160 109.920 33.330 110.535 ;
        RECT 32.225 109.750 33.330 109.920 ;
        RECT 33.500 109.475 33.670 110.275 ;
        RECT 33.840 109.975 34.010 111.045 ;
        RECT 34.180 110.145 34.370 110.865 ;
        RECT 34.540 110.115 34.860 111.075 ;
        RECT 35.030 111.115 35.200 111.575 ;
        RECT 35.475 111.495 35.685 112.025 ;
        RECT 35.945 111.285 36.275 111.810 ;
        RECT 36.445 111.415 36.615 112.025 ;
        RECT 36.785 111.370 37.115 111.805 ;
        RECT 36.785 111.285 37.165 111.370 ;
        RECT 37.795 111.300 38.085 112.025 ;
        RECT 38.270 111.455 38.525 111.805 ;
        RECT 38.695 111.625 39.025 112.025 ;
        RECT 39.195 111.455 39.365 111.805 ;
        RECT 39.535 111.625 39.915 112.025 ;
        RECT 38.270 111.285 39.935 111.455 ;
        RECT 40.105 111.350 40.380 111.695 ;
        RECT 41.180 111.515 41.420 112.025 ;
        RECT 41.600 111.515 41.880 111.845 ;
        RECT 42.110 111.515 42.325 112.025 ;
        RECT 36.075 111.115 36.275 111.285 ;
        RECT 36.940 111.245 37.165 111.285 ;
        RECT 35.030 110.785 35.905 111.115 ;
        RECT 36.075 110.785 36.825 111.115 ;
        RECT 33.840 109.645 34.090 109.975 ;
        RECT 35.030 109.945 35.200 110.785 ;
        RECT 36.075 110.580 36.265 110.785 ;
        RECT 36.995 110.665 37.165 111.245 ;
        RECT 39.765 111.115 39.935 111.285 ;
        RECT 38.255 110.785 38.600 111.115 ;
        RECT 38.770 110.785 39.595 111.115 ;
        RECT 39.765 110.785 40.040 111.115 ;
        RECT 36.950 110.615 37.165 110.665 ;
        RECT 35.370 110.205 36.265 110.580 ;
        RECT 36.775 110.535 37.165 110.615 ;
        RECT 34.315 109.775 35.200 109.945 ;
        RECT 35.380 109.475 35.695 109.975 ;
        RECT 35.925 109.645 36.265 110.205 ;
        RECT 36.435 109.475 36.605 110.485 ;
        RECT 36.775 109.690 37.105 110.535 ;
        RECT 37.795 109.475 38.085 110.640 ;
        RECT 38.275 110.325 38.600 110.615 ;
        RECT 38.770 110.495 38.965 110.785 ;
        RECT 39.765 110.615 39.935 110.785 ;
        RECT 40.210 110.615 40.380 111.350 ;
        RECT 41.075 110.785 41.430 111.345 ;
        RECT 41.600 110.615 41.770 111.515 ;
        RECT 41.940 110.785 42.205 111.345 ;
        RECT 42.495 111.285 43.110 111.855 ;
        RECT 43.320 111.495 43.610 111.845 ;
        RECT 43.805 111.665 44.135 112.025 ;
        RECT 44.305 111.495 44.535 111.800 ;
        RECT 43.320 111.325 44.535 111.495 ;
        RECT 44.725 111.685 44.895 111.720 ;
        RECT 44.725 111.515 44.925 111.685 ;
        RECT 42.455 110.615 42.625 111.115 ;
        RECT 39.275 110.445 39.935 110.615 ;
        RECT 39.275 110.325 39.445 110.445 ;
        RECT 38.275 110.155 39.445 110.325 ;
        RECT 38.255 109.695 39.445 109.985 ;
        RECT 39.615 109.475 39.895 110.275 ;
        RECT 40.105 109.645 40.380 110.615 ;
        RECT 41.200 110.445 42.625 110.615 ;
        RECT 41.200 110.270 41.590 110.445 ;
        RECT 42.075 109.475 42.405 110.275 ;
        RECT 42.795 110.265 43.110 111.285 ;
        RECT 44.725 111.155 44.895 111.515 ;
        RECT 45.195 111.205 45.425 112.025 ;
        RECT 45.595 111.225 45.925 111.855 ;
        RECT 43.380 111.005 43.640 111.115 ;
        RECT 43.375 110.835 43.640 111.005 ;
        RECT 43.380 110.785 43.640 110.835 ;
        RECT 43.820 110.785 44.205 111.115 ;
        RECT 44.375 110.985 44.895 111.155 ;
        RECT 42.575 109.645 43.110 110.265 ;
        RECT 43.320 109.475 43.640 110.615 ;
        RECT 43.820 109.735 44.015 110.785 ;
        RECT 44.375 110.605 44.545 110.985 ;
        RECT 44.195 110.325 44.545 110.605 ;
        RECT 44.735 110.455 44.980 110.815 ;
        RECT 45.175 110.785 45.505 111.035 ;
        RECT 45.675 110.625 45.925 111.225 ;
        RECT 46.095 111.205 46.305 112.025 ;
        RECT 46.535 111.480 51.880 112.025 ;
        RECT 48.120 110.650 48.460 111.480 ;
        RECT 52.055 111.255 53.725 112.025 ;
        RECT 54.360 111.455 54.680 111.855 ;
        RECT 44.195 109.645 44.525 110.325 ;
        RECT 44.725 109.475 44.980 110.275 ;
        RECT 45.195 109.475 45.425 110.615 ;
        RECT 45.595 109.645 45.925 110.625 ;
        RECT 46.095 109.475 46.305 110.615 ;
        RECT 49.940 109.910 50.290 111.160 ;
        RECT 52.055 110.735 52.805 111.255 ;
        RECT 52.975 110.565 53.725 111.085 ;
        RECT 46.535 109.475 51.880 109.910 ;
        RECT 52.055 109.475 53.725 110.565 ;
        RECT 54.360 110.665 54.530 111.455 ;
        RECT 54.850 111.205 55.160 112.025 ;
        RECT 55.330 111.395 55.660 111.855 ;
        RECT 55.830 111.565 56.080 112.025 ;
        RECT 56.270 111.645 58.320 111.855 ;
        RECT 56.270 111.395 57.020 111.475 ;
        RECT 55.330 111.205 57.020 111.395 ;
        RECT 57.190 111.205 57.360 111.645 ;
        RECT 57.530 111.205 58.320 111.475 ;
        RECT 54.700 110.835 55.050 111.035 ;
        RECT 55.330 110.835 56.010 111.035 ;
        RECT 56.220 110.835 57.410 111.035 ;
        RECT 57.590 110.665 57.920 111.035 ;
        RECT 54.360 110.495 57.920 110.665 ;
        RECT 54.360 110.045 54.530 110.495 ;
        RECT 58.120 110.325 58.320 111.205 ;
        RECT 58.495 111.255 60.165 112.025 ;
        RECT 60.795 111.395 61.135 111.855 ;
        RECT 61.305 111.565 61.475 112.025 ;
        RECT 62.105 111.590 62.465 111.855 ;
        RECT 62.110 111.585 62.465 111.590 ;
        RECT 62.115 111.575 62.465 111.585 ;
        RECT 62.120 111.570 62.465 111.575 ;
        RECT 62.125 111.560 62.465 111.570 ;
        RECT 62.705 111.565 62.875 112.025 ;
        RECT 62.130 111.555 62.465 111.560 ;
        RECT 62.140 111.545 62.465 111.555 ;
        RECT 62.150 111.535 62.465 111.545 ;
        RECT 61.645 111.395 61.975 111.475 ;
        RECT 58.495 110.735 59.245 111.255 ;
        RECT 60.795 111.205 61.975 111.395 ;
        RECT 62.165 111.395 62.465 111.535 ;
        RECT 62.165 111.205 62.875 111.395 ;
        RECT 59.415 110.565 60.165 111.085 ;
        RECT 54.360 109.645 54.680 110.045 ;
        RECT 54.850 109.475 55.160 110.275 ;
        RECT 55.330 110.155 58.320 110.325 ;
        RECT 55.330 110.105 56.500 110.155 ;
        RECT 55.330 109.645 55.660 110.105 ;
        RECT 55.830 109.475 56.000 109.935 ;
        RECT 56.170 109.645 56.500 110.105 ;
        RECT 57.530 110.105 58.320 110.155 ;
        RECT 56.670 109.475 56.920 109.935 ;
        RECT 57.110 109.475 57.360 109.935 ;
        RECT 57.530 109.645 57.780 110.105 ;
        RECT 58.030 109.475 58.320 109.935 ;
        RECT 58.495 109.475 60.165 110.565 ;
        RECT 60.795 110.835 61.125 111.035 ;
        RECT 61.435 111.015 61.765 111.035 ;
        RECT 61.315 110.835 61.765 111.015 ;
        RECT 60.795 110.495 61.025 110.835 ;
        RECT 60.805 109.475 61.135 110.195 ;
        RECT 61.315 109.720 61.530 110.835 ;
        RECT 61.935 110.805 62.405 111.035 ;
        RECT 62.590 110.635 62.875 111.205 ;
        RECT 63.045 111.080 63.385 111.855 ;
        RECT 63.555 111.300 63.845 112.025 ;
        RECT 64.100 111.455 64.275 111.855 ;
        RECT 64.445 111.645 64.775 112.025 ;
        RECT 65.020 111.525 65.250 111.855 ;
        RECT 64.100 111.285 64.730 111.455 ;
        RECT 64.560 111.115 64.730 111.285 ;
        RECT 61.725 110.420 62.875 110.635 ;
        RECT 61.725 109.645 62.055 110.420 ;
        RECT 62.225 109.475 62.935 110.250 ;
        RECT 63.105 109.645 63.385 111.080 ;
        RECT 63.555 109.475 63.845 110.640 ;
        RECT 64.015 110.435 64.380 111.115 ;
        RECT 64.560 110.785 64.910 111.115 ;
        RECT 64.560 110.265 64.730 110.785 ;
        RECT 64.100 110.095 64.730 110.265 ;
        RECT 65.080 110.235 65.250 111.525 ;
        RECT 65.450 110.415 65.730 111.690 ;
        RECT 65.955 111.685 66.225 111.690 ;
        RECT 65.915 111.515 66.225 111.685 ;
        RECT 66.685 111.645 67.015 112.025 ;
        RECT 67.185 111.770 67.520 111.815 ;
        RECT 65.955 110.415 66.225 111.515 ;
        RECT 66.415 110.415 66.755 111.445 ;
        RECT 67.185 111.305 67.525 111.770 ;
        RECT 66.925 110.785 67.185 111.115 ;
        RECT 66.925 110.235 67.095 110.785 ;
        RECT 67.355 110.615 67.525 111.305 ;
        RECT 64.100 109.645 64.275 110.095 ;
        RECT 65.080 110.065 67.095 110.235 ;
        RECT 64.445 109.475 64.775 109.915 ;
        RECT 65.080 109.645 65.250 110.065 ;
        RECT 65.485 109.475 66.155 109.885 ;
        RECT 66.370 109.645 66.540 110.065 ;
        RECT 66.740 109.475 67.070 109.885 ;
        RECT 67.265 109.645 67.525 110.615 ;
        RECT 68.615 111.285 69.000 111.855 ;
        RECT 69.170 111.565 69.495 112.025 ;
        RECT 70.015 111.395 70.295 111.855 ;
        RECT 68.615 110.615 68.895 111.285 ;
        RECT 69.170 111.225 70.295 111.395 ;
        RECT 69.170 111.115 69.620 111.225 ;
        RECT 69.065 110.785 69.620 111.115 ;
        RECT 70.485 111.055 70.885 111.855 ;
        RECT 71.285 111.565 71.555 112.025 ;
        RECT 71.725 111.395 72.010 111.855 ;
        RECT 72.295 111.635 73.555 111.815 ;
        RECT 68.615 109.645 69.000 110.615 ;
        RECT 69.170 110.325 69.620 110.785 ;
        RECT 69.790 110.495 70.885 111.055 ;
        RECT 69.170 110.105 70.295 110.325 ;
        RECT 69.170 109.475 69.495 109.935 ;
        RECT 70.015 109.645 70.295 110.105 ;
        RECT 70.485 109.645 70.885 110.495 ;
        RECT 71.055 111.225 72.010 111.395 ;
        RECT 71.055 110.325 71.265 111.225 ;
        RECT 71.435 110.495 72.125 111.055 ;
        RECT 71.055 110.105 72.010 110.325 ;
        RECT 72.295 110.120 72.535 111.445 ;
        RECT 72.705 111.285 73.055 111.465 ;
        RECT 73.225 111.415 73.555 111.635 ;
        RECT 73.745 111.585 73.915 112.025 ;
        RECT 74.085 111.415 74.425 111.830 ;
        RECT 73.225 111.285 74.425 111.415 ;
        RECT 72.705 110.275 72.875 111.285 ;
        RECT 73.395 111.245 74.425 111.285 ;
        RECT 74.595 111.255 78.105 112.025 ;
        RECT 78.365 111.475 78.535 111.765 ;
        RECT 78.705 111.645 79.035 112.025 ;
        RECT 78.365 111.305 79.030 111.475 ;
        RECT 73.045 110.695 73.215 111.115 ;
        RECT 73.430 110.865 73.795 111.035 ;
        RECT 73.045 110.445 73.445 110.695 ;
        RECT 73.615 110.665 73.795 110.865 ;
        RECT 73.965 110.835 74.425 111.035 ;
        RECT 74.595 110.735 76.245 111.255 ;
        RECT 73.615 110.495 73.935 110.665 ;
        RECT 71.285 109.475 71.555 109.935 ;
        RECT 71.725 109.645 72.010 110.105 ;
        RECT 72.705 110.065 73.545 110.275 ;
        RECT 72.345 109.475 72.555 109.935 ;
        RECT 73.045 109.645 73.545 110.065 ;
        RECT 73.735 109.705 73.935 110.495 ;
        RECT 74.105 109.475 74.425 110.655 ;
        RECT 76.415 110.565 78.105 111.085 ;
        RECT 74.595 109.475 78.105 110.565 ;
        RECT 78.280 110.485 78.630 111.135 ;
        RECT 78.800 110.315 79.030 111.305 ;
        RECT 78.365 110.145 79.030 110.315 ;
        RECT 78.365 109.645 78.535 110.145 ;
        RECT 78.705 109.475 79.035 109.975 ;
        RECT 79.205 109.645 79.390 111.765 ;
        RECT 79.645 111.565 79.895 112.025 ;
        RECT 80.065 111.575 80.400 111.745 ;
        RECT 80.595 111.575 81.270 111.745 ;
        RECT 80.065 111.435 80.235 111.575 ;
        RECT 79.560 110.445 79.840 111.395 ;
        RECT 80.010 111.305 80.235 111.435 ;
        RECT 80.010 110.200 80.180 111.305 ;
        RECT 80.405 111.155 80.930 111.375 ;
        RECT 80.350 110.390 80.590 110.985 ;
        RECT 80.760 110.455 80.930 111.155 ;
        RECT 81.100 110.795 81.270 111.575 ;
        RECT 81.590 111.525 81.960 112.025 ;
        RECT 82.140 111.575 82.545 111.745 ;
        RECT 82.715 111.575 83.500 111.745 ;
        RECT 82.140 111.345 82.310 111.575 ;
        RECT 81.480 111.045 82.310 111.345 ;
        RECT 82.695 111.075 83.160 111.405 ;
        RECT 81.480 111.015 81.680 111.045 ;
        RECT 81.800 110.795 81.970 110.865 ;
        RECT 81.100 110.625 81.970 110.795 ;
        RECT 81.460 110.535 81.970 110.625 ;
        RECT 80.010 110.070 80.315 110.200 ;
        RECT 80.760 110.090 81.290 110.455 ;
        RECT 79.630 109.475 79.895 109.935 ;
        RECT 80.065 109.645 80.315 110.070 ;
        RECT 81.460 109.920 81.630 110.535 ;
        RECT 80.525 109.750 81.630 109.920 ;
        RECT 81.800 109.475 81.970 110.275 ;
        RECT 82.140 109.975 82.310 111.045 ;
        RECT 82.480 110.145 82.670 110.865 ;
        RECT 82.840 110.115 83.160 111.075 ;
        RECT 83.330 111.115 83.500 111.575 ;
        RECT 83.775 111.495 83.985 112.025 ;
        RECT 84.245 111.285 84.575 111.810 ;
        RECT 84.745 111.415 84.915 112.025 ;
        RECT 85.085 111.370 85.415 111.805 ;
        RECT 85.085 111.285 85.465 111.370 ;
        RECT 84.375 111.115 84.575 111.285 ;
        RECT 85.240 111.245 85.465 111.285 ;
        RECT 83.330 110.785 84.205 111.115 ;
        RECT 84.375 110.785 85.125 111.115 ;
        RECT 82.140 109.645 82.390 109.975 ;
        RECT 83.330 109.945 83.500 110.785 ;
        RECT 84.375 110.580 84.565 110.785 ;
        RECT 85.295 110.665 85.465 111.245 ;
        RECT 85.250 110.615 85.465 110.665 ;
        RECT 83.670 110.205 84.565 110.580 ;
        RECT 85.075 110.535 85.465 110.615 ;
        RECT 85.635 111.285 86.020 111.855 ;
        RECT 86.190 111.565 86.515 112.025 ;
        RECT 87.035 111.395 87.315 111.855 ;
        RECT 85.635 110.615 85.915 111.285 ;
        RECT 86.190 111.225 87.315 111.395 ;
        RECT 86.190 111.115 86.640 111.225 ;
        RECT 86.085 110.785 86.640 111.115 ;
        RECT 87.505 111.055 87.905 111.855 ;
        RECT 88.305 111.565 88.575 112.025 ;
        RECT 88.745 111.395 89.030 111.855 ;
        RECT 82.615 109.775 83.500 109.945 ;
        RECT 83.680 109.475 83.995 109.975 ;
        RECT 84.225 109.645 84.565 110.205 ;
        RECT 84.735 109.475 84.905 110.485 ;
        RECT 85.075 109.690 85.405 110.535 ;
        RECT 85.635 109.645 86.020 110.615 ;
        RECT 86.190 110.325 86.640 110.785 ;
        RECT 86.810 110.495 87.905 111.055 ;
        RECT 86.190 110.105 87.315 110.325 ;
        RECT 86.190 109.475 86.515 109.935 ;
        RECT 87.035 109.645 87.315 110.105 ;
        RECT 87.505 109.645 87.905 110.495 ;
        RECT 88.075 111.225 89.030 111.395 ;
        RECT 89.315 111.275 90.525 112.025 ;
        RECT 88.075 110.325 88.285 111.225 ;
        RECT 88.455 110.495 89.145 111.055 ;
        RECT 89.315 110.565 89.835 111.105 ;
        RECT 90.005 110.735 90.525 111.275 ;
        RECT 100.090 110.950 100.760 114.210 ;
        RECT 101.430 113.640 105.470 113.810 ;
        RECT 101.090 111.580 101.260 113.580 ;
        RECT 105.640 111.580 105.810 113.580 ;
        RECT 101.430 111.350 105.470 111.520 ;
        RECT 106.150 110.950 106.320 114.210 ;
        RECT 100.090 110.780 106.320 110.950 ;
        RECT 88.075 110.105 89.030 110.325 ;
        RECT 88.305 109.475 88.575 109.935 ;
        RECT 88.745 109.645 89.030 110.105 ;
        RECT 89.315 109.475 90.525 110.565 ;
        RECT 11.950 109.305 90.610 109.475 ;
        RECT 12.035 108.215 13.245 109.305 ;
        RECT 13.505 108.635 13.675 109.135 ;
        RECT 13.845 108.805 14.175 109.305 ;
        RECT 13.505 108.465 14.170 108.635 ;
        RECT 12.035 107.505 12.555 108.045 ;
        RECT 12.725 107.675 13.245 108.215 ;
        RECT 13.420 107.645 13.770 108.295 ;
        RECT 12.035 106.755 13.245 107.505 ;
        RECT 13.940 107.475 14.170 108.465 ;
        RECT 13.505 107.305 14.170 107.475 ;
        RECT 13.505 107.015 13.675 107.305 ;
        RECT 13.845 106.755 14.175 107.135 ;
        RECT 14.345 107.015 14.530 109.135 ;
        RECT 14.770 108.845 15.035 109.305 ;
        RECT 15.205 108.710 15.455 109.135 ;
        RECT 15.665 108.860 16.770 109.030 ;
        RECT 15.150 108.580 15.455 108.710 ;
        RECT 14.700 107.385 14.980 108.335 ;
        RECT 15.150 107.475 15.320 108.580 ;
        RECT 15.490 107.795 15.730 108.390 ;
        RECT 15.900 108.325 16.430 108.690 ;
        RECT 15.900 107.625 16.070 108.325 ;
        RECT 16.600 108.245 16.770 108.860 ;
        RECT 16.940 108.505 17.110 109.305 ;
        RECT 17.280 108.805 17.530 109.135 ;
        RECT 17.755 108.835 18.640 109.005 ;
        RECT 16.600 108.155 17.110 108.245 ;
        RECT 15.150 107.345 15.375 107.475 ;
        RECT 15.545 107.405 16.070 107.625 ;
        RECT 16.240 107.985 17.110 108.155 ;
        RECT 14.785 106.755 15.035 107.215 ;
        RECT 15.205 107.205 15.375 107.345 ;
        RECT 16.240 107.205 16.410 107.985 ;
        RECT 16.940 107.915 17.110 107.985 ;
        RECT 16.620 107.735 16.820 107.765 ;
        RECT 17.280 107.735 17.450 108.805 ;
        RECT 17.620 107.915 17.810 108.635 ;
        RECT 16.620 107.435 17.450 107.735 ;
        RECT 17.980 107.705 18.300 108.665 ;
        RECT 15.205 107.035 15.540 107.205 ;
        RECT 15.735 107.035 16.410 107.205 ;
        RECT 16.730 106.755 17.100 107.255 ;
        RECT 17.280 107.205 17.450 107.435 ;
        RECT 17.835 107.375 18.300 107.705 ;
        RECT 18.470 107.995 18.640 108.835 ;
        RECT 18.820 108.805 19.135 109.305 ;
        RECT 19.365 108.575 19.705 109.135 ;
        RECT 18.810 108.200 19.705 108.575 ;
        RECT 19.875 108.295 20.045 109.305 ;
        RECT 19.515 107.995 19.705 108.200 ;
        RECT 20.215 108.245 20.545 109.090 ;
        RECT 20.215 108.165 20.605 108.245 ;
        RECT 20.780 108.165 21.100 109.305 ;
        RECT 20.390 108.115 20.605 108.165 ;
        RECT 18.470 107.665 19.345 107.995 ;
        RECT 19.515 107.665 20.265 107.995 ;
        RECT 18.470 107.205 18.640 107.665 ;
        RECT 19.515 107.495 19.715 107.665 ;
        RECT 20.435 107.535 20.605 108.115 ;
        RECT 21.280 107.995 21.475 109.045 ;
        RECT 21.655 108.455 21.985 109.135 ;
        RECT 22.185 108.505 22.440 109.305 ;
        RECT 22.650 108.515 23.185 109.135 ;
        RECT 21.655 108.175 22.005 108.455 ;
        RECT 20.840 107.945 21.100 107.995 ;
        RECT 20.835 107.775 21.100 107.945 ;
        RECT 20.840 107.665 21.100 107.775 ;
        RECT 21.280 107.665 21.665 107.995 ;
        RECT 21.835 107.795 22.005 108.175 ;
        RECT 22.195 107.965 22.440 108.325 ;
        RECT 21.835 107.625 22.355 107.795 ;
        RECT 20.380 107.495 20.605 107.535 ;
        RECT 17.280 107.035 17.685 107.205 ;
        RECT 17.855 107.035 18.640 107.205 ;
        RECT 18.915 106.755 19.125 107.285 ;
        RECT 19.385 106.970 19.715 107.495 ;
        RECT 20.225 107.410 20.605 107.495 ;
        RECT 19.885 106.755 20.055 107.365 ;
        RECT 20.225 106.975 20.555 107.410 ;
        RECT 20.780 107.285 21.995 107.455 ;
        RECT 20.780 106.935 21.070 107.285 ;
        RECT 21.265 106.755 21.595 107.115 ;
        RECT 21.765 106.980 21.995 107.285 ;
        RECT 22.185 107.060 22.355 107.625 ;
        RECT 22.650 107.495 22.965 108.515 ;
        RECT 23.355 108.505 23.685 109.305 ;
        RECT 24.170 108.335 24.560 108.510 ;
        RECT 23.135 108.165 24.560 108.335 ;
        RECT 23.135 107.665 23.305 108.165 ;
        RECT 22.650 106.925 23.265 107.495 ;
        RECT 23.555 107.435 23.820 107.995 ;
        RECT 23.990 107.265 24.160 108.165 ;
        RECT 24.915 108.140 25.205 109.305 ;
        RECT 26.295 108.795 27.495 109.035 ;
        RECT 27.675 108.880 28.005 109.305 ;
        RECT 28.520 108.880 28.880 109.305 ;
        RECT 29.085 108.710 29.345 108.890 ;
        RECT 27.710 108.625 29.345 108.710 ;
        RECT 26.295 108.165 26.600 108.595 ;
        RECT 26.770 108.540 29.345 108.625 ;
        RECT 26.770 108.455 27.880 108.540 ;
        RECT 28.665 108.480 29.345 108.540 ;
        RECT 24.330 107.435 24.685 107.995 ;
        RECT 26.295 107.495 26.465 108.165 ;
        RECT 26.770 107.995 26.940 108.455 ;
        RECT 26.640 107.665 26.940 107.995 ;
        RECT 27.200 107.745 27.735 108.285 ;
        RECT 28.100 108.165 28.495 108.370 ;
        RECT 27.985 107.605 28.155 107.995 ;
        RECT 27.835 107.575 28.155 107.605 ;
        RECT 27.270 107.495 28.155 107.575 ;
        RECT 23.435 106.755 23.650 107.265 ;
        RECT 23.880 106.935 24.160 107.265 ;
        RECT 24.340 106.755 24.580 107.265 ;
        RECT 24.915 106.755 25.205 107.480 ;
        RECT 26.295 107.435 28.155 107.495 ;
        RECT 26.295 107.405 28.005 107.435 ;
        RECT 26.295 107.325 27.440 107.405 ;
        RECT 26.295 107.275 26.600 107.325 ;
        RECT 26.345 106.975 26.600 107.275 ;
        RECT 26.770 106.755 27.100 107.155 ;
        RECT 27.270 106.975 27.440 107.325 ;
        RECT 28.325 107.265 28.495 108.165 ;
        RECT 28.665 107.575 28.835 108.480 ;
        RECT 29.005 107.745 29.345 108.310 ;
        RECT 29.520 108.165 29.795 109.135 ;
        RECT 30.005 108.505 30.285 109.305 ;
        RECT 30.455 108.795 31.645 109.085 ;
        RECT 30.455 108.455 31.625 108.625 ;
        RECT 30.455 108.335 30.625 108.455 ;
        RECT 29.965 108.165 30.625 108.335 ;
        RECT 28.665 107.405 29.345 107.575 ;
        RECT 27.740 106.755 27.910 107.235 ;
        RECT 28.145 106.935 28.495 107.265 ;
        RECT 28.665 106.755 28.835 107.235 ;
        RECT 29.085 106.960 29.345 107.405 ;
        RECT 29.520 107.430 29.690 108.165 ;
        RECT 29.965 107.995 30.135 108.165 ;
        RECT 30.935 107.995 31.130 108.285 ;
        RECT 31.300 108.165 31.625 108.455 ;
        RECT 31.815 108.215 33.485 109.305 ;
        RECT 29.860 107.665 30.135 107.995 ;
        RECT 30.305 107.665 31.130 107.995 ;
        RECT 31.300 107.665 31.645 107.995 ;
        RECT 29.965 107.495 30.135 107.665 ;
        RECT 31.815 107.525 32.565 108.045 ;
        RECT 32.735 107.695 33.485 108.215 ;
        RECT 34.115 108.165 34.395 109.305 ;
        RECT 34.565 108.155 34.895 109.135 ;
        RECT 35.065 108.165 35.325 109.305 ;
        RECT 35.495 108.165 35.770 109.135 ;
        RECT 35.980 108.505 36.260 109.305 ;
        RECT 36.430 108.795 38.045 109.125 ;
        RECT 36.430 108.455 37.605 108.625 ;
        RECT 36.430 108.335 36.600 108.455 ;
        RECT 35.940 108.165 36.600 108.335 ;
        RECT 34.125 107.725 34.460 107.995 ;
        RECT 34.630 107.555 34.800 108.155 ;
        RECT 34.970 107.745 35.305 107.995 ;
        RECT 29.520 107.085 29.795 107.430 ;
        RECT 29.965 107.325 31.630 107.495 ;
        RECT 29.985 106.755 30.365 107.155 ;
        RECT 30.535 106.975 30.705 107.325 ;
        RECT 30.875 106.755 31.205 107.155 ;
        RECT 31.375 106.975 31.630 107.325 ;
        RECT 31.815 106.755 33.485 107.525 ;
        RECT 34.115 106.755 34.425 107.555 ;
        RECT 34.630 106.925 35.325 107.555 ;
        RECT 35.495 107.430 35.665 108.165 ;
        RECT 35.940 107.995 36.110 108.165 ;
        RECT 36.860 107.995 37.105 108.285 ;
        RECT 37.275 108.165 37.605 108.455 ;
        RECT 37.865 107.995 38.035 108.555 ;
        RECT 38.285 108.165 38.545 109.305 ;
        RECT 38.715 108.165 39.100 109.135 ;
        RECT 39.270 108.845 39.595 109.305 ;
        RECT 40.115 108.675 40.395 109.135 ;
        RECT 39.270 108.455 40.395 108.675 ;
        RECT 35.835 107.665 36.110 107.995 ;
        RECT 36.280 107.665 37.105 107.995 ;
        RECT 37.320 107.665 38.035 107.995 ;
        RECT 38.205 107.745 38.540 107.995 ;
        RECT 35.940 107.495 36.110 107.665 ;
        RECT 37.785 107.575 38.035 107.665 ;
        RECT 35.495 107.085 35.770 107.430 ;
        RECT 35.940 107.325 37.605 107.495 ;
        RECT 35.960 106.755 36.335 107.155 ;
        RECT 36.505 106.975 36.675 107.325 ;
        RECT 36.845 106.755 37.175 107.155 ;
        RECT 37.345 106.925 37.605 107.325 ;
        RECT 37.785 107.155 38.115 107.575 ;
        RECT 38.285 106.755 38.545 107.575 ;
        RECT 38.715 107.495 38.995 108.165 ;
        RECT 39.270 107.995 39.720 108.455 ;
        RECT 40.585 108.285 40.985 109.135 ;
        RECT 41.385 108.845 41.655 109.305 ;
        RECT 41.825 108.675 42.110 109.135 ;
        RECT 39.165 107.665 39.720 107.995 ;
        RECT 39.890 107.725 40.985 108.285 ;
        RECT 39.270 107.555 39.720 107.665 ;
        RECT 38.715 106.925 39.100 107.495 ;
        RECT 39.270 107.385 40.395 107.555 ;
        RECT 39.270 106.755 39.595 107.215 ;
        RECT 40.115 106.925 40.395 107.385 ;
        RECT 40.585 106.925 40.985 107.725 ;
        RECT 41.155 108.455 42.110 108.675 ;
        RECT 42.595 108.635 42.875 109.305 ;
        RECT 41.155 107.555 41.365 108.455 ;
        RECT 43.045 108.415 43.345 108.965 ;
        RECT 43.545 108.585 43.875 109.305 ;
        RECT 44.065 108.585 44.525 109.135 ;
        RECT 41.535 107.725 42.225 108.285 ;
        RECT 42.410 107.995 42.675 108.355 ;
        RECT 43.045 108.245 43.985 108.415 ;
        RECT 43.815 107.995 43.985 108.245 ;
        RECT 42.410 107.745 43.085 107.995 ;
        RECT 43.305 107.745 43.645 107.995 ;
        RECT 43.815 107.665 44.105 107.995 ;
        RECT 43.815 107.575 43.985 107.665 ;
        RECT 41.155 107.385 42.110 107.555 ;
        RECT 41.385 106.755 41.655 107.215 ;
        RECT 41.825 106.925 42.110 107.385 ;
        RECT 42.595 107.385 43.985 107.575 ;
        RECT 42.595 107.025 42.925 107.385 ;
        RECT 44.275 107.215 44.525 108.585 ;
        RECT 44.695 108.215 48.205 109.305 ;
        RECT 48.375 108.750 48.980 109.305 ;
        RECT 49.155 108.795 49.635 109.135 ;
        RECT 49.805 108.760 50.060 109.305 ;
        RECT 48.375 108.650 48.990 108.750 ;
        RECT 48.805 108.625 48.990 108.650 ;
        RECT 43.545 106.755 43.795 107.215 ;
        RECT 43.965 106.925 44.525 107.215 ;
        RECT 44.695 107.525 46.345 108.045 ;
        RECT 46.515 107.695 48.205 108.215 ;
        RECT 48.375 108.030 48.635 108.480 ;
        RECT 48.805 108.380 49.135 108.625 ;
        RECT 49.305 108.305 50.060 108.555 ;
        RECT 50.230 108.435 50.505 109.135 ;
        RECT 49.290 108.270 50.060 108.305 ;
        RECT 49.275 108.260 50.060 108.270 ;
        RECT 49.270 108.245 50.165 108.260 ;
        RECT 49.250 108.230 50.165 108.245 ;
        RECT 49.230 108.220 50.165 108.230 ;
        RECT 49.205 108.210 50.165 108.220 ;
        RECT 49.135 108.180 50.165 108.210 ;
        RECT 49.115 108.150 50.165 108.180 ;
        RECT 49.095 108.120 50.165 108.150 ;
        RECT 49.065 108.095 50.165 108.120 ;
        RECT 49.030 108.060 50.165 108.095 ;
        RECT 49.000 108.055 50.165 108.060 ;
        RECT 49.000 108.050 49.390 108.055 ;
        RECT 49.000 108.040 49.365 108.050 ;
        RECT 49.000 108.035 49.350 108.040 ;
        RECT 49.000 108.030 49.335 108.035 ;
        RECT 48.375 108.025 49.335 108.030 ;
        RECT 48.375 108.015 49.325 108.025 ;
        RECT 48.375 108.010 49.315 108.015 ;
        RECT 48.375 108.000 49.305 108.010 ;
        RECT 48.375 107.990 49.300 108.000 ;
        RECT 48.375 107.985 49.295 107.990 ;
        RECT 48.375 107.970 49.285 107.985 ;
        RECT 48.375 107.955 49.280 107.970 ;
        RECT 48.375 107.930 49.270 107.955 ;
        RECT 48.375 107.860 49.265 107.930 ;
        RECT 44.695 106.755 48.205 107.525 ;
        RECT 48.375 107.305 48.925 107.690 ;
        RECT 49.095 107.135 49.265 107.860 ;
        RECT 48.375 106.965 49.265 107.135 ;
        RECT 49.435 107.460 49.765 107.885 ;
        RECT 49.935 107.660 50.165 108.055 ;
        RECT 49.435 106.975 49.655 107.460 ;
        RECT 50.335 107.405 50.505 108.435 ;
        RECT 50.675 108.140 50.965 109.305 ;
        RECT 51.145 108.495 51.440 109.305 ;
        RECT 51.620 107.995 51.865 109.135 ;
        RECT 52.040 108.495 52.300 109.305 ;
        RECT 52.900 109.300 59.175 109.305 ;
        RECT 52.480 107.995 52.730 109.130 ;
        RECT 52.900 108.505 53.160 109.300 ;
        RECT 53.330 108.405 53.590 109.130 ;
        RECT 53.760 108.575 54.020 109.300 ;
        RECT 54.190 108.405 54.450 109.130 ;
        RECT 54.620 108.575 54.880 109.300 ;
        RECT 55.050 108.405 55.310 109.130 ;
        RECT 55.480 108.575 55.740 109.300 ;
        RECT 55.910 108.405 56.170 109.130 ;
        RECT 56.340 108.575 56.585 109.300 ;
        RECT 56.755 108.405 57.015 109.130 ;
        RECT 57.200 108.575 57.445 109.300 ;
        RECT 57.615 108.405 57.875 109.130 ;
        RECT 58.060 108.575 58.305 109.300 ;
        RECT 58.475 108.405 58.735 109.130 ;
        RECT 58.920 108.575 59.175 109.300 ;
        RECT 53.330 108.390 58.735 108.405 ;
        RECT 59.345 108.390 59.635 109.130 ;
        RECT 59.805 108.560 60.075 109.305 ;
        RECT 53.330 108.165 60.075 108.390 ;
        RECT 60.335 108.215 63.845 109.305 ;
        RECT 49.825 106.755 50.075 107.295 ;
        RECT 50.245 106.925 50.505 107.405 ;
        RECT 50.675 106.755 50.965 107.480 ;
        RECT 51.135 107.435 51.450 107.995 ;
        RECT 51.620 107.745 58.740 107.995 ;
        RECT 51.135 106.755 51.440 107.265 ;
        RECT 51.620 106.935 51.870 107.745 ;
        RECT 52.040 106.755 52.300 107.280 ;
        RECT 52.480 106.935 52.730 107.745 ;
        RECT 58.910 107.575 60.075 108.165 ;
        RECT 53.330 107.405 60.075 107.575 ;
        RECT 60.335 107.525 61.985 108.045 ;
        RECT 62.155 107.695 63.845 108.215 ;
        RECT 64.975 108.165 65.205 109.305 ;
        RECT 65.375 108.155 65.705 109.135 ;
        RECT 65.875 108.165 66.085 109.305 ;
        RECT 66.315 108.215 67.525 109.305 ;
        RECT 64.955 107.745 65.285 107.995 ;
        RECT 52.900 106.755 53.160 107.315 ;
        RECT 53.330 106.950 53.590 107.405 ;
        RECT 53.760 106.755 54.020 107.235 ;
        RECT 54.190 106.950 54.450 107.405 ;
        RECT 54.620 106.755 54.880 107.235 ;
        RECT 55.050 106.950 55.310 107.405 ;
        RECT 55.480 106.755 55.725 107.235 ;
        RECT 55.895 106.950 56.170 107.405 ;
        RECT 56.340 106.755 56.585 107.235 ;
        RECT 56.755 106.950 57.015 107.405 ;
        RECT 57.195 106.755 57.445 107.235 ;
        RECT 57.615 106.950 57.875 107.405 ;
        RECT 58.055 106.755 58.305 107.235 ;
        RECT 58.475 106.950 58.735 107.405 ;
        RECT 58.915 106.755 59.175 107.235 ;
        RECT 59.345 106.950 59.605 107.405 ;
        RECT 59.775 106.755 60.075 107.235 ;
        RECT 60.335 106.755 63.845 107.525 ;
        RECT 64.975 106.755 65.205 107.575 ;
        RECT 65.455 107.555 65.705 108.155 ;
        RECT 65.375 106.925 65.705 107.555 ;
        RECT 65.875 106.755 66.085 107.575 ;
        RECT 66.315 107.505 66.835 108.045 ;
        RECT 67.005 107.675 67.525 108.215 ;
        RECT 67.695 108.435 67.970 109.135 ;
        RECT 68.180 108.760 68.395 109.305 ;
        RECT 68.565 108.795 69.040 109.135 ;
        RECT 69.210 108.800 69.825 109.305 ;
        RECT 69.210 108.625 69.405 108.800 ;
        RECT 66.315 106.755 67.525 107.505 ;
        RECT 67.695 107.405 67.865 108.435 ;
        RECT 68.140 108.265 68.855 108.560 ;
        RECT 69.075 108.435 69.405 108.625 ;
        RECT 69.575 108.265 69.825 108.630 ;
        RECT 68.035 108.095 69.825 108.265 ;
        RECT 68.035 107.665 68.265 108.095 ;
        RECT 67.695 106.925 67.955 107.405 ;
        RECT 68.435 107.395 68.845 107.915 ;
        RECT 68.125 106.755 68.455 107.215 ;
        RECT 68.645 106.975 68.845 107.395 ;
        RECT 69.015 107.240 69.270 108.095 ;
        RECT 70.065 107.915 70.235 109.135 ;
        RECT 70.485 108.795 70.745 109.305 ;
        RECT 70.915 108.795 72.105 109.085 ;
        RECT 69.440 107.665 70.235 107.915 ;
        RECT 70.405 107.745 70.745 108.625 ;
        RECT 70.935 108.455 72.105 108.625 ;
        RECT 72.275 108.505 72.555 109.305 ;
        RECT 70.935 108.165 71.260 108.455 ;
        RECT 71.935 108.335 72.105 108.455 ;
        RECT 71.430 107.995 71.625 108.285 ;
        RECT 71.935 108.165 72.595 108.335 ;
        RECT 72.765 108.165 73.040 109.135 ;
        RECT 73.215 108.165 73.475 109.305 ;
        RECT 73.645 108.335 73.975 109.135 ;
        RECT 74.145 108.505 74.315 109.305 ;
        RECT 74.485 108.335 74.815 109.135 ;
        RECT 74.985 108.505 75.240 109.305 ;
        RECT 73.645 108.165 75.345 108.335 ;
        RECT 72.425 107.995 72.595 108.165 ;
        RECT 70.915 107.665 71.260 107.995 ;
        RECT 71.430 107.665 72.255 107.995 ;
        RECT 72.425 107.665 72.700 107.995 ;
        RECT 69.985 107.575 70.235 107.665 ;
        RECT 69.015 106.975 69.805 107.240 ;
        RECT 69.985 107.155 70.315 107.575 ;
        RECT 70.485 106.755 70.745 107.575 ;
        RECT 72.425 107.495 72.595 107.665 ;
        RECT 70.930 107.325 72.595 107.495 ;
        RECT 72.870 107.430 73.040 108.165 ;
        RECT 73.215 107.745 73.975 107.995 ;
        RECT 74.145 107.745 74.895 107.995 ;
        RECT 75.065 107.575 75.345 108.165 ;
        RECT 76.435 108.140 76.725 109.305 ;
        RECT 77.390 108.505 77.640 109.305 ;
        RECT 77.810 108.675 78.140 109.135 ;
        RECT 78.310 108.845 78.525 109.305 ;
        RECT 77.810 108.505 78.980 108.675 ;
        RECT 76.900 108.335 77.180 108.495 ;
        RECT 76.900 108.165 78.235 108.335 ;
        RECT 78.065 107.995 78.235 108.165 ;
        RECT 76.900 107.745 77.250 107.985 ;
        RECT 77.420 107.745 77.895 107.985 ;
        RECT 78.065 107.745 78.440 107.995 ;
        RECT 78.065 107.575 78.235 107.745 ;
        RECT 70.930 106.975 71.185 107.325 ;
        RECT 71.355 106.755 71.685 107.155 ;
        RECT 71.855 106.975 72.025 107.325 ;
        RECT 72.195 106.755 72.575 107.155 ;
        RECT 72.765 107.085 73.040 107.430 ;
        RECT 73.215 107.385 74.315 107.555 ;
        RECT 73.215 106.925 73.555 107.385 ;
        RECT 73.725 106.755 73.895 107.215 ;
        RECT 74.065 107.135 74.315 107.385 ;
        RECT 74.485 107.325 75.345 107.575 ;
        RECT 74.905 107.135 75.235 107.155 ;
        RECT 74.065 106.925 75.235 107.135 ;
        RECT 76.435 106.755 76.725 107.480 ;
        RECT 76.900 107.405 78.235 107.575 ;
        RECT 76.900 107.195 77.170 107.405 ;
        RECT 78.610 107.215 78.980 108.505 ;
        RECT 79.195 108.215 80.405 109.305 ;
        RECT 77.390 106.755 77.720 107.215 ;
        RECT 78.230 106.925 78.980 107.215 ;
        RECT 79.195 107.505 79.715 108.045 ;
        RECT 79.885 107.675 80.405 108.215 ;
        RECT 80.580 108.165 80.915 109.135 ;
        RECT 81.085 108.165 81.255 109.305 ;
        RECT 81.425 108.965 83.455 109.135 ;
        RECT 79.195 106.755 80.405 107.505 ;
        RECT 80.580 107.495 80.750 108.165 ;
        RECT 81.425 107.995 81.595 108.965 ;
        RECT 80.920 107.665 81.175 107.995 ;
        RECT 81.400 107.665 81.595 107.995 ;
        RECT 81.765 108.625 82.890 108.795 ;
        RECT 81.005 107.495 81.175 107.665 ;
        RECT 81.765 107.495 81.935 108.625 ;
        RECT 80.580 106.925 80.835 107.495 ;
        RECT 81.005 107.325 81.935 107.495 ;
        RECT 82.105 108.285 83.115 108.455 ;
        RECT 82.105 107.485 82.275 108.285 ;
        RECT 82.480 107.945 82.755 108.085 ;
        RECT 82.475 107.775 82.755 107.945 ;
        RECT 81.760 107.290 81.935 107.325 ;
        RECT 81.005 106.755 81.335 107.155 ;
        RECT 81.760 106.925 82.290 107.290 ;
        RECT 82.480 106.925 82.755 107.775 ;
        RECT 82.925 106.925 83.115 108.285 ;
        RECT 83.285 108.300 83.455 108.965 ;
        RECT 83.625 108.545 83.795 109.305 ;
        RECT 84.030 108.545 84.545 108.955 ;
        RECT 83.285 108.110 84.035 108.300 ;
        RECT 84.205 107.735 84.545 108.545 ;
        RECT 84.715 108.215 85.925 109.305 ;
        RECT 83.315 107.565 84.545 107.735 ;
        RECT 83.295 106.755 83.805 107.290 ;
        RECT 84.025 106.960 84.270 107.565 ;
        RECT 84.715 107.505 85.235 108.045 ;
        RECT 85.405 107.675 85.925 108.215 ;
        RECT 86.185 108.375 86.355 109.135 ;
        RECT 86.535 108.545 86.865 109.305 ;
        RECT 86.185 108.205 86.850 108.375 ;
        RECT 87.035 108.230 87.305 109.135 ;
        RECT 86.680 108.060 86.850 108.205 ;
        RECT 86.115 107.655 86.445 108.025 ;
        RECT 86.680 107.730 86.965 108.060 ;
        RECT 84.715 106.755 85.925 107.505 ;
        RECT 86.680 107.475 86.850 107.730 ;
        RECT 86.185 107.305 86.850 107.475 ;
        RECT 87.135 107.430 87.305 108.230 ;
        RECT 87.475 108.215 89.145 109.305 ;
        RECT 86.185 106.925 86.355 107.305 ;
        RECT 86.535 106.755 86.865 107.135 ;
        RECT 87.045 106.925 87.305 107.430 ;
        RECT 87.475 107.525 88.225 108.045 ;
        RECT 88.395 107.695 89.145 108.215 ;
        RECT 89.315 108.215 90.525 109.305 ;
        RECT 89.315 107.675 89.835 108.215 ;
        RECT 87.475 106.755 89.145 107.525 ;
        RECT 90.005 107.505 90.525 108.045 ;
        RECT 89.315 106.755 90.525 107.505 ;
        RECT 100.090 107.520 100.760 110.780 ;
        RECT 101.430 110.210 105.470 110.380 ;
        RECT 101.090 108.150 101.260 110.150 ;
        RECT 105.640 108.150 105.810 110.150 ;
        RECT 101.430 107.920 105.470 108.090 ;
        RECT 106.150 107.520 106.320 110.780 ;
        RECT 100.090 107.510 106.320 107.520 ;
        RECT 107.910 116.780 117.740 116.820 ;
        RECT 120.510 116.800 126.250 116.810 ;
        RECT 107.910 116.650 118.540 116.780 ;
        RECT 107.910 114.390 108.080 116.650 ;
        RECT 108.805 116.080 116.845 116.250 ;
        RECT 108.420 115.020 108.590 116.020 ;
        RECT 117.060 115.020 117.230 116.020 ;
        RECT 108.805 114.790 116.845 114.960 ;
        RECT 117.570 114.390 118.540 116.650 ;
        RECT 107.910 114.220 118.540 114.390 ;
        RECT 107.910 110.960 108.080 114.220 ;
        RECT 108.805 113.650 116.845 113.820 ;
        RECT 108.420 111.590 108.590 113.590 ;
        RECT 117.060 111.590 117.230 113.590 ;
        RECT 108.805 111.360 116.845 111.530 ;
        RECT 117.570 110.960 118.540 114.220 ;
        RECT 107.910 110.790 118.540 110.960 ;
        RECT 107.910 107.530 108.080 110.790 ;
        RECT 108.805 110.220 116.845 110.390 ;
        RECT 108.420 108.160 108.590 110.160 ;
        RECT 117.060 108.160 117.230 110.160 ;
        RECT 108.805 107.930 116.845 108.100 ;
        RECT 117.570 107.530 118.540 110.790 ;
        RECT 100.090 107.410 106.330 107.510 ;
        RECT 100.080 106.850 106.330 107.410 ;
        RECT 100.080 106.830 105.250 106.850 ;
        RECT 100.080 106.760 104.070 106.830 ;
        RECT 11.950 106.585 90.610 106.755 ;
        RECT 12.035 105.835 13.245 106.585 ;
        RECT 13.880 106.110 14.215 106.370 ;
        RECT 14.385 106.185 14.715 106.585 ;
        RECT 14.885 106.185 16.500 106.355 ;
        RECT 12.035 105.295 12.555 105.835 ;
        RECT 12.725 105.125 13.245 105.665 ;
        RECT 12.035 104.035 13.245 105.125 ;
        RECT 13.880 104.755 14.135 106.110 ;
        RECT 14.885 106.015 15.055 106.185 ;
        RECT 14.495 105.845 15.055 106.015 ;
        RECT 15.320 105.905 15.590 106.005 ;
        RECT 15.780 105.905 16.070 106.005 ;
        RECT 14.495 105.675 14.665 105.845 ;
        RECT 15.315 105.735 15.590 105.905 ;
        RECT 15.775 105.735 16.070 105.905 ;
        RECT 14.360 105.345 14.665 105.675 ;
        RECT 14.860 105.565 15.110 105.675 ;
        RECT 14.855 105.395 15.110 105.565 ;
        RECT 14.860 105.345 15.110 105.395 ;
        RECT 15.320 105.345 15.590 105.735 ;
        RECT 15.780 105.345 16.070 105.735 ;
        RECT 16.240 105.345 16.660 106.010 ;
        RECT 17.045 105.865 17.375 106.585 ;
        RECT 17.560 105.745 17.820 106.585 ;
        RECT 17.995 105.840 18.250 106.415 ;
        RECT 18.420 106.205 18.750 106.585 ;
        RECT 18.965 106.035 19.135 106.415 ;
        RECT 18.420 105.865 19.135 106.035 ;
        RECT 16.970 105.565 17.320 105.675 ;
        RECT 16.970 105.395 17.325 105.565 ;
        RECT 16.970 105.345 17.320 105.395 ;
        RECT 14.495 105.175 14.665 105.345 ;
        RECT 14.495 105.005 16.865 105.175 ;
        RECT 17.115 105.055 17.320 105.345 ;
        RECT 13.880 104.245 14.215 104.755 ;
        RECT 14.465 104.035 14.795 104.835 ;
        RECT 15.040 104.625 16.465 104.795 ;
        RECT 15.040 104.205 15.325 104.625 ;
        RECT 15.580 104.035 15.910 104.455 ;
        RECT 16.135 104.375 16.465 104.625 ;
        RECT 16.695 104.545 16.865 105.005 ;
        RECT 17.125 104.375 17.295 104.875 ;
        RECT 16.135 104.205 17.295 104.375 ;
        RECT 17.560 104.035 17.820 105.185 ;
        RECT 17.995 105.110 18.165 105.840 ;
        RECT 18.420 105.675 18.590 105.865 ;
        RECT 20.315 105.785 20.625 106.585 ;
        RECT 20.830 105.785 21.525 106.415 ;
        RECT 21.785 106.035 21.955 106.415 ;
        RECT 22.135 106.205 22.465 106.585 ;
        RECT 21.785 105.865 22.450 106.035 ;
        RECT 22.645 105.910 22.905 106.415 ;
        RECT 23.625 106.245 23.795 106.280 ;
        RECT 23.595 106.075 23.795 106.245 ;
        RECT 18.335 105.345 18.590 105.675 ;
        RECT 18.420 105.135 18.590 105.345 ;
        RECT 18.870 105.315 19.225 105.685 ;
        RECT 20.325 105.345 20.660 105.615 ;
        RECT 20.830 105.225 21.000 105.785 ;
        RECT 21.170 105.345 21.505 105.595 ;
        RECT 21.715 105.315 22.055 105.685 ;
        RECT 22.280 105.610 22.450 105.865 ;
        RECT 22.280 105.280 22.555 105.610 ;
        RECT 20.830 105.185 21.005 105.225 ;
        RECT 17.995 104.205 18.250 105.110 ;
        RECT 18.420 104.965 19.135 105.135 ;
        RECT 18.420 104.035 18.750 104.795 ;
        RECT 18.965 104.205 19.135 104.965 ;
        RECT 20.315 104.035 20.595 105.175 ;
        RECT 20.765 104.205 21.095 105.185 ;
        RECT 21.265 104.035 21.525 105.175 ;
        RECT 22.280 105.135 22.450 105.280 ;
        RECT 21.775 104.965 22.450 105.135 ;
        RECT 22.725 105.110 22.905 105.910 ;
        RECT 23.625 105.715 23.795 106.075 ;
        RECT 23.985 106.055 24.215 106.360 ;
        RECT 24.385 106.225 24.715 106.585 ;
        RECT 24.910 106.055 25.200 106.405 ;
        RECT 23.985 105.885 25.200 106.055 ;
        RECT 25.375 105.835 26.585 106.585 ;
        RECT 26.755 105.845 27.140 106.415 ;
        RECT 27.310 106.125 27.635 106.585 ;
        RECT 28.155 105.955 28.435 106.415 ;
        RECT 23.625 105.545 24.145 105.715 ;
        RECT 21.775 104.205 21.955 104.965 ;
        RECT 22.135 104.035 22.465 104.795 ;
        RECT 22.635 104.205 22.905 105.110 ;
        RECT 23.540 105.015 23.785 105.375 ;
        RECT 23.975 105.165 24.145 105.545 ;
        RECT 24.315 105.345 24.700 105.675 ;
        RECT 24.880 105.565 25.140 105.675 ;
        RECT 24.880 105.395 25.145 105.565 ;
        RECT 24.880 105.345 25.140 105.395 ;
        RECT 23.975 104.885 24.325 105.165 ;
        RECT 23.540 104.035 23.795 104.835 ;
        RECT 23.995 104.205 24.325 104.885 ;
        RECT 24.505 104.295 24.700 105.345 ;
        RECT 25.375 105.295 25.895 105.835 ;
        RECT 24.880 104.035 25.200 105.175 ;
        RECT 26.065 105.125 26.585 105.665 ;
        RECT 25.375 104.035 26.585 105.125 ;
        RECT 26.755 105.175 27.035 105.845 ;
        RECT 27.310 105.785 28.435 105.955 ;
        RECT 27.310 105.675 27.760 105.785 ;
        RECT 27.205 105.345 27.760 105.675 ;
        RECT 28.625 105.615 29.025 106.415 ;
        RECT 29.425 106.125 29.695 106.585 ;
        RECT 29.865 105.955 30.150 106.415 ;
        RECT 26.755 104.205 27.140 105.175 ;
        RECT 27.310 104.885 27.760 105.345 ;
        RECT 27.930 105.055 29.025 105.615 ;
        RECT 27.310 104.665 28.435 104.885 ;
        RECT 27.310 104.035 27.635 104.495 ;
        RECT 28.155 104.205 28.435 104.665 ;
        RECT 28.625 104.205 29.025 105.055 ;
        RECT 29.195 105.785 30.150 105.955 ;
        RECT 30.525 106.035 30.695 106.325 ;
        RECT 30.865 106.205 31.195 106.585 ;
        RECT 30.525 105.865 31.190 106.035 ;
        RECT 29.195 104.885 29.405 105.785 ;
        RECT 29.575 105.055 30.265 105.615 ;
        RECT 30.440 105.045 30.790 105.695 ;
        RECT 29.195 104.665 30.150 104.885 ;
        RECT 30.960 104.875 31.190 105.865 ;
        RECT 29.425 104.035 29.695 104.495 ;
        RECT 29.865 104.205 30.150 104.665 ;
        RECT 30.525 104.705 31.190 104.875 ;
        RECT 30.525 104.205 30.695 104.705 ;
        RECT 30.865 104.035 31.195 104.535 ;
        RECT 31.365 104.205 31.550 106.325 ;
        RECT 31.805 106.125 32.055 106.585 ;
        RECT 32.225 106.135 32.560 106.305 ;
        RECT 32.755 106.135 33.430 106.305 ;
        RECT 32.225 105.995 32.395 106.135 ;
        RECT 31.720 105.005 32.000 105.955 ;
        RECT 32.170 105.865 32.395 105.995 ;
        RECT 32.170 104.760 32.340 105.865 ;
        RECT 32.565 105.715 33.090 105.935 ;
        RECT 32.510 104.950 32.750 105.545 ;
        RECT 32.920 105.015 33.090 105.715 ;
        RECT 33.260 105.355 33.430 106.135 ;
        RECT 33.750 106.085 34.120 106.585 ;
        RECT 34.300 106.135 34.705 106.305 ;
        RECT 34.875 106.135 35.660 106.305 ;
        RECT 34.300 105.905 34.470 106.135 ;
        RECT 33.640 105.605 34.470 105.905 ;
        RECT 34.855 105.635 35.320 105.965 ;
        RECT 33.640 105.575 33.840 105.605 ;
        RECT 33.960 105.355 34.130 105.425 ;
        RECT 33.260 105.185 34.130 105.355 ;
        RECT 33.620 105.095 34.130 105.185 ;
        RECT 32.170 104.630 32.475 104.760 ;
        RECT 32.920 104.650 33.450 105.015 ;
        RECT 31.790 104.035 32.055 104.495 ;
        RECT 32.225 104.205 32.475 104.630 ;
        RECT 33.620 104.480 33.790 105.095 ;
        RECT 32.685 104.310 33.790 104.480 ;
        RECT 33.960 104.035 34.130 104.835 ;
        RECT 34.300 104.535 34.470 105.605 ;
        RECT 34.640 104.705 34.830 105.425 ;
        RECT 35.000 104.675 35.320 105.635 ;
        RECT 35.490 105.675 35.660 106.135 ;
        RECT 35.935 106.055 36.145 106.585 ;
        RECT 36.405 105.845 36.735 106.370 ;
        RECT 36.905 105.975 37.075 106.585 ;
        RECT 37.245 105.930 37.575 106.365 ;
        RECT 37.245 105.845 37.625 105.930 ;
        RECT 37.795 105.860 38.085 106.585 ;
        RECT 38.275 105.855 38.565 106.585 ;
        RECT 36.535 105.675 36.735 105.845 ;
        RECT 37.400 105.805 37.625 105.845 ;
        RECT 35.490 105.345 36.365 105.675 ;
        RECT 36.535 105.345 37.285 105.675 ;
        RECT 34.300 104.205 34.550 104.535 ;
        RECT 35.490 104.505 35.660 105.345 ;
        RECT 36.535 105.140 36.725 105.345 ;
        RECT 37.455 105.225 37.625 105.805 ;
        RECT 38.265 105.345 38.565 105.675 ;
        RECT 38.745 105.655 38.975 106.295 ;
        RECT 39.155 106.035 39.465 106.405 ;
        RECT 39.645 106.215 40.315 106.585 ;
        RECT 39.155 105.835 40.385 106.035 ;
        RECT 38.745 105.345 39.270 105.655 ;
        RECT 39.450 105.345 39.915 105.655 ;
        RECT 37.410 105.175 37.625 105.225 ;
        RECT 35.830 104.765 36.725 105.140 ;
        RECT 37.235 105.095 37.625 105.175 ;
        RECT 34.775 104.335 35.660 104.505 ;
        RECT 35.840 104.035 36.155 104.535 ;
        RECT 36.385 104.205 36.725 104.765 ;
        RECT 36.895 104.035 37.065 105.045 ;
        RECT 37.235 104.250 37.565 105.095 ;
        RECT 37.795 104.035 38.085 105.200 ;
        RECT 40.095 105.165 40.385 105.835 ;
        RECT 38.275 104.925 39.435 105.165 ;
        RECT 38.275 104.215 38.535 104.925 ;
        RECT 38.705 104.035 39.035 104.745 ;
        RECT 39.205 104.215 39.435 104.925 ;
        RECT 39.615 104.945 40.385 105.165 ;
        RECT 39.615 104.215 39.885 104.945 ;
        RECT 40.065 104.035 40.405 104.765 ;
        RECT 40.575 104.215 40.835 106.405 ;
        RECT 41.025 105.775 41.295 106.585 ;
        RECT 41.465 105.775 41.795 106.415 ;
        RECT 41.965 105.775 42.205 106.585 ;
        RECT 42.485 106.035 42.655 106.325 ;
        RECT 42.825 106.205 43.155 106.585 ;
        RECT 42.485 105.865 43.150 106.035 ;
        RECT 41.015 105.345 41.365 105.595 ;
        RECT 41.535 105.175 41.705 105.775 ;
        RECT 41.875 105.345 42.225 105.595 ;
        RECT 41.025 104.035 41.355 105.175 ;
        RECT 41.535 105.005 42.215 105.175 ;
        RECT 42.400 105.045 42.750 105.695 ;
        RECT 41.885 104.220 42.215 105.005 ;
        RECT 42.920 104.875 43.150 105.865 ;
        RECT 42.485 104.705 43.150 104.875 ;
        RECT 42.485 104.205 42.655 104.705 ;
        RECT 42.825 104.035 43.155 104.535 ;
        RECT 43.325 104.205 43.510 106.325 ;
        RECT 43.765 106.125 44.015 106.585 ;
        RECT 44.185 106.135 44.520 106.305 ;
        RECT 44.715 106.135 45.390 106.305 ;
        RECT 44.185 105.995 44.355 106.135 ;
        RECT 43.680 105.005 43.960 105.955 ;
        RECT 44.130 105.865 44.355 105.995 ;
        RECT 44.130 104.760 44.300 105.865 ;
        RECT 44.525 105.715 45.050 105.935 ;
        RECT 44.470 104.950 44.710 105.545 ;
        RECT 44.880 105.015 45.050 105.715 ;
        RECT 45.220 105.355 45.390 106.135 ;
        RECT 45.710 106.085 46.080 106.585 ;
        RECT 46.260 106.135 46.665 106.305 ;
        RECT 46.835 106.135 47.620 106.305 ;
        RECT 46.260 105.905 46.430 106.135 ;
        RECT 45.600 105.605 46.430 105.905 ;
        RECT 46.815 105.635 47.280 105.965 ;
        RECT 45.600 105.575 45.800 105.605 ;
        RECT 45.920 105.355 46.090 105.425 ;
        RECT 45.220 105.185 46.090 105.355 ;
        RECT 45.580 105.095 46.090 105.185 ;
        RECT 44.130 104.630 44.435 104.760 ;
        RECT 44.880 104.650 45.410 105.015 ;
        RECT 43.750 104.035 44.015 104.495 ;
        RECT 44.185 104.205 44.435 104.630 ;
        RECT 45.580 104.480 45.750 105.095 ;
        RECT 44.645 104.310 45.750 104.480 ;
        RECT 45.920 104.035 46.090 104.835 ;
        RECT 46.260 104.535 46.430 105.605 ;
        RECT 46.600 104.705 46.790 105.425 ;
        RECT 46.960 104.675 47.280 105.635 ;
        RECT 47.450 105.675 47.620 106.135 ;
        RECT 47.895 106.055 48.105 106.585 ;
        RECT 48.365 105.845 48.695 106.370 ;
        RECT 48.865 105.975 49.035 106.585 ;
        RECT 49.205 105.930 49.535 106.365 ;
        RECT 49.205 105.845 49.585 105.930 ;
        RECT 48.495 105.675 48.695 105.845 ;
        RECT 49.360 105.805 49.585 105.845 ;
        RECT 47.450 105.345 48.325 105.675 ;
        RECT 48.495 105.345 49.245 105.675 ;
        RECT 46.260 104.205 46.510 104.535 ;
        RECT 47.450 104.505 47.620 105.345 ;
        RECT 48.495 105.140 48.685 105.345 ;
        RECT 49.415 105.225 49.585 105.805 ;
        RECT 49.370 105.175 49.585 105.225 ;
        RECT 47.790 104.765 48.685 105.140 ;
        RECT 49.195 105.095 49.585 105.175 ;
        RECT 50.675 105.845 51.060 106.415 ;
        RECT 51.230 106.125 51.555 106.585 ;
        RECT 52.075 105.955 52.355 106.415 ;
        RECT 50.675 105.175 50.955 105.845 ;
        RECT 51.230 105.785 52.355 105.955 ;
        RECT 51.230 105.675 51.680 105.785 ;
        RECT 51.125 105.345 51.680 105.675 ;
        RECT 52.545 105.615 52.945 106.415 ;
        RECT 53.345 106.125 53.615 106.585 ;
        RECT 53.785 105.955 54.070 106.415 ;
        RECT 54.815 106.205 55.705 106.375 ;
        RECT 46.735 104.335 47.620 104.505 ;
        RECT 47.800 104.035 48.115 104.535 ;
        RECT 48.345 104.205 48.685 104.765 ;
        RECT 48.855 104.035 49.025 105.045 ;
        RECT 49.195 104.250 49.525 105.095 ;
        RECT 50.675 104.205 51.060 105.175 ;
        RECT 51.230 104.885 51.680 105.345 ;
        RECT 51.850 105.055 52.945 105.615 ;
        RECT 51.230 104.665 52.355 104.885 ;
        RECT 51.230 104.035 51.555 104.495 ;
        RECT 52.075 104.205 52.355 104.665 ;
        RECT 52.545 104.205 52.945 105.055 ;
        RECT 53.115 105.785 54.070 105.955 ;
        RECT 53.115 104.885 53.325 105.785 ;
        RECT 54.815 105.650 55.365 106.035 ;
        RECT 53.495 105.055 54.185 105.615 ;
        RECT 55.535 105.480 55.705 106.205 ;
        RECT 54.815 105.410 55.705 105.480 ;
        RECT 55.875 105.880 56.095 106.365 ;
        RECT 56.265 106.045 56.515 106.585 ;
        RECT 56.685 105.935 56.945 106.415 ;
        RECT 55.875 105.455 56.205 105.880 ;
        RECT 54.815 105.385 55.710 105.410 ;
        RECT 54.815 105.370 55.720 105.385 ;
        RECT 54.815 105.355 55.725 105.370 ;
        RECT 54.815 105.350 55.735 105.355 ;
        RECT 54.815 105.340 55.740 105.350 ;
        RECT 54.815 105.330 55.745 105.340 ;
        RECT 54.815 105.325 55.755 105.330 ;
        RECT 54.815 105.315 55.765 105.325 ;
        RECT 54.815 105.310 55.775 105.315 ;
        RECT 53.115 104.665 54.070 104.885 ;
        RECT 54.815 104.860 55.075 105.310 ;
        RECT 55.440 105.305 55.775 105.310 ;
        RECT 55.440 105.300 55.790 105.305 ;
        RECT 55.440 105.290 55.805 105.300 ;
        RECT 55.440 105.285 55.830 105.290 ;
        RECT 56.375 105.285 56.605 105.680 ;
        RECT 55.440 105.280 56.605 105.285 ;
        RECT 55.470 105.245 56.605 105.280 ;
        RECT 55.505 105.220 56.605 105.245 ;
        RECT 55.535 105.190 56.605 105.220 ;
        RECT 55.555 105.160 56.605 105.190 ;
        RECT 55.575 105.130 56.605 105.160 ;
        RECT 55.645 105.120 56.605 105.130 ;
        RECT 55.670 105.110 56.605 105.120 ;
        RECT 55.690 105.095 56.605 105.110 ;
        RECT 55.710 105.080 56.605 105.095 ;
        RECT 55.715 105.070 56.500 105.080 ;
        RECT 55.730 105.035 56.500 105.070 ;
        RECT 55.245 104.715 55.575 104.960 ;
        RECT 55.745 104.785 56.500 105.035 ;
        RECT 56.775 104.905 56.945 105.935 ;
        RECT 57.230 105.955 57.515 106.415 ;
        RECT 57.685 106.125 57.955 106.585 ;
        RECT 57.230 105.785 58.185 105.955 ;
        RECT 57.115 105.055 57.805 105.615 ;
        RECT 55.245 104.690 55.430 104.715 ;
        RECT 53.345 104.035 53.615 104.495 ;
        RECT 53.785 104.205 54.070 104.665 ;
        RECT 54.815 104.590 55.430 104.690 ;
        RECT 54.815 104.035 55.420 104.590 ;
        RECT 55.595 104.205 56.075 104.545 ;
        RECT 56.245 104.035 56.500 104.580 ;
        RECT 56.670 104.205 56.945 104.905 ;
        RECT 57.975 104.885 58.185 105.785 ;
        RECT 57.230 104.665 58.185 104.885 ;
        RECT 58.355 105.615 58.755 106.415 ;
        RECT 58.945 105.955 59.225 106.415 ;
        RECT 59.745 106.125 60.070 106.585 ;
        RECT 58.945 105.785 60.070 105.955 ;
        RECT 60.240 105.845 60.625 106.415 ;
        RECT 59.620 105.675 60.070 105.785 ;
        RECT 58.355 105.055 59.450 105.615 ;
        RECT 59.620 105.345 60.175 105.675 ;
        RECT 57.230 104.205 57.515 104.665 ;
        RECT 57.685 104.035 57.955 104.495 ;
        RECT 58.355 104.205 58.755 105.055 ;
        RECT 59.620 104.885 60.070 105.345 ;
        RECT 60.345 105.175 60.625 105.845 ;
        RECT 60.795 105.815 63.385 106.585 ;
        RECT 63.555 105.860 63.845 106.585 ;
        RECT 64.020 106.055 64.310 106.405 ;
        RECT 64.505 106.225 64.835 106.585 ;
        RECT 65.005 106.055 65.235 106.360 ;
        RECT 64.020 105.885 65.235 106.055 ;
        RECT 60.795 105.295 62.005 105.815 ;
        RECT 65.425 105.715 65.595 106.280 ;
        RECT 65.855 106.040 71.200 106.585 ;
        RECT 71.855 106.075 72.095 106.585 ;
        RECT 72.265 106.075 72.555 106.415 ;
        RECT 72.785 106.075 73.100 106.585 ;
        RECT 58.945 104.665 60.070 104.885 ;
        RECT 58.945 104.205 59.225 104.665 ;
        RECT 59.745 104.035 60.070 104.495 ;
        RECT 60.240 104.205 60.625 105.175 ;
        RECT 62.175 105.125 63.385 105.645 ;
        RECT 64.080 105.565 64.340 105.675 ;
        RECT 64.075 105.395 64.340 105.565 ;
        RECT 64.080 105.345 64.340 105.395 ;
        RECT 64.520 105.345 64.905 105.675 ;
        RECT 65.075 105.545 65.595 105.715 ;
        RECT 60.795 104.035 63.385 105.125 ;
        RECT 63.555 104.035 63.845 105.200 ;
        RECT 64.020 104.035 64.340 105.175 ;
        RECT 64.520 104.295 64.715 105.345 ;
        RECT 65.075 105.165 65.245 105.545 ;
        RECT 64.895 104.885 65.245 105.165 ;
        RECT 65.435 105.015 65.680 105.375 ;
        RECT 67.440 105.210 67.780 106.040 ;
        RECT 64.895 104.205 65.225 104.885 ;
        RECT 65.425 104.035 65.680 104.835 ;
        RECT 69.260 104.470 69.610 105.720 ;
        RECT 71.900 105.565 72.095 105.905 ;
        RECT 71.895 105.395 72.095 105.565 ;
        RECT 71.900 105.345 72.095 105.395 ;
        RECT 72.265 105.175 72.445 106.075 ;
        RECT 73.270 106.015 73.440 106.285 ;
        RECT 73.610 106.185 73.940 106.585 ;
        RECT 72.615 105.345 73.025 105.905 ;
        RECT 73.270 105.845 73.965 106.015 ;
        RECT 73.195 105.175 73.365 105.675 ;
        RECT 71.905 105.005 73.365 105.175 ;
        RECT 71.905 104.830 72.265 105.005 ;
        RECT 73.535 104.835 73.965 105.845 ;
        RECT 74.340 105.805 74.840 106.415 ;
        RECT 74.135 105.345 74.485 105.595 ;
        RECT 74.670 105.175 74.840 105.805 ;
        RECT 75.470 105.935 75.800 106.415 ;
        RECT 75.970 106.125 76.195 106.585 ;
        RECT 76.365 105.935 76.695 106.415 ;
        RECT 75.470 105.765 76.695 105.935 ;
        RECT 76.885 105.785 77.135 106.585 ;
        RECT 77.305 105.785 77.645 106.415 ;
        RECT 75.010 105.395 75.340 105.595 ;
        RECT 75.510 105.395 75.840 105.595 ;
        RECT 76.010 105.395 76.430 105.595 ;
        RECT 76.605 105.425 77.300 105.595 ;
        RECT 76.605 105.175 76.775 105.425 ;
        RECT 77.470 105.175 77.645 105.785 ;
        RECT 77.820 105.745 78.080 106.585 ;
        RECT 78.255 105.840 78.510 106.415 ;
        RECT 78.680 106.205 79.010 106.585 ;
        RECT 79.225 106.035 79.395 106.415 ;
        RECT 78.680 105.865 79.395 106.035 ;
        RECT 65.855 104.035 71.200 104.470 ;
        RECT 72.850 104.035 73.020 104.835 ;
        RECT 73.190 104.665 73.965 104.835 ;
        RECT 74.340 105.005 76.775 105.175 ;
        RECT 73.190 104.205 73.520 104.665 ;
        RECT 73.690 104.035 73.860 104.495 ;
        RECT 74.340 104.205 74.670 105.005 ;
        RECT 74.840 104.035 75.170 104.835 ;
        RECT 75.470 104.205 75.800 105.005 ;
        RECT 76.445 104.035 76.695 104.835 ;
        RECT 76.965 104.035 77.135 105.175 ;
        RECT 77.305 104.205 77.645 105.175 ;
        RECT 77.820 104.035 78.080 105.185 ;
        RECT 78.255 105.110 78.425 105.840 ;
        RECT 78.680 105.675 78.850 105.865 ;
        RECT 79.655 105.815 83.165 106.585 ;
        RECT 83.335 105.835 84.545 106.585 ;
        RECT 84.715 105.845 85.100 106.415 ;
        RECT 85.270 106.125 85.595 106.585 ;
        RECT 86.115 105.955 86.395 106.415 ;
        RECT 78.595 105.345 78.850 105.675 ;
        RECT 78.680 105.135 78.850 105.345 ;
        RECT 79.130 105.315 79.485 105.685 ;
        RECT 79.655 105.295 81.305 105.815 ;
        RECT 78.255 104.205 78.510 105.110 ;
        RECT 78.680 104.965 79.395 105.135 ;
        RECT 81.475 105.125 83.165 105.645 ;
        RECT 83.335 105.295 83.855 105.835 ;
        RECT 84.025 105.125 84.545 105.665 ;
        RECT 78.680 104.035 79.010 104.795 ;
        RECT 79.225 104.205 79.395 104.965 ;
        RECT 79.655 104.035 83.165 105.125 ;
        RECT 83.335 104.035 84.545 105.125 ;
        RECT 84.715 105.175 84.995 105.845 ;
        RECT 85.270 105.785 86.395 105.955 ;
        RECT 85.270 105.675 85.720 105.785 ;
        RECT 85.165 105.345 85.720 105.675 ;
        RECT 86.585 105.615 86.985 106.415 ;
        RECT 87.385 106.125 87.655 106.585 ;
        RECT 87.825 105.955 88.110 106.415 ;
        RECT 84.715 104.205 85.100 105.175 ;
        RECT 85.270 104.885 85.720 105.345 ;
        RECT 85.890 105.055 86.985 105.615 ;
        RECT 85.270 104.665 86.395 104.885 ;
        RECT 85.270 104.035 85.595 104.495 ;
        RECT 86.115 104.205 86.395 104.665 ;
        RECT 86.585 104.205 86.985 105.055 ;
        RECT 87.155 105.785 88.110 105.955 ;
        RECT 89.315 105.835 90.525 106.585 ;
        RECT 87.155 104.885 87.365 105.785 ;
        RECT 87.535 105.055 88.225 105.615 ;
        RECT 89.315 105.125 89.835 105.665 ;
        RECT 90.005 105.295 90.525 105.835 ;
        RECT 100.080 105.490 102.000 106.760 ;
        RECT 103.510 106.750 104.070 106.760 ;
        RECT 103.740 105.660 104.070 106.750 ;
        RECT 104.440 106.280 105.480 106.450 ;
        RECT 104.440 105.840 105.480 106.010 ;
        RECT 105.650 105.980 105.820 106.310 ;
        RECT 103.900 105.440 104.070 105.660 ;
        RECT 106.160 105.440 106.330 106.850 ;
        RECT 103.900 105.270 106.330 105.440 ;
        RECT 107.910 107.360 118.540 107.530 ;
        RECT 120.020 116.640 126.250 116.800 ;
        RECT 120.020 114.380 120.690 116.640 ;
        RECT 121.360 116.070 125.400 116.240 ;
        RECT 121.020 115.010 121.190 116.010 ;
        RECT 125.570 115.010 125.740 116.010 ;
        RECT 121.360 114.780 125.400 114.950 ;
        RECT 126.080 114.380 126.250 116.640 ;
        RECT 120.020 114.210 126.250 114.380 ;
        RECT 120.020 110.950 120.690 114.210 ;
        RECT 121.360 113.640 125.400 113.810 ;
        RECT 121.020 111.580 121.190 113.580 ;
        RECT 125.570 111.580 125.740 113.580 ;
        RECT 121.360 111.350 125.400 111.520 ;
        RECT 126.080 110.950 126.250 114.210 ;
        RECT 120.020 110.780 126.250 110.950 ;
        RECT 120.020 107.520 120.690 110.780 ;
        RECT 121.360 110.210 125.400 110.380 ;
        RECT 121.020 108.150 121.190 110.150 ;
        RECT 125.570 108.150 125.740 110.150 ;
        RECT 121.360 107.920 125.400 108.090 ;
        RECT 126.080 107.520 126.250 110.780 ;
        RECT 120.020 107.510 126.250 107.520 ;
        RECT 127.840 116.780 137.670 116.820 ;
        RECT 140.540 116.800 146.280 116.810 ;
        RECT 127.840 116.650 138.470 116.780 ;
        RECT 127.840 114.390 128.010 116.650 ;
        RECT 128.735 116.080 136.775 116.250 ;
        RECT 128.350 115.020 128.520 116.020 ;
        RECT 136.990 115.020 137.160 116.020 ;
        RECT 128.735 114.790 136.775 114.960 ;
        RECT 137.500 114.390 138.470 116.650 ;
        RECT 127.840 114.220 138.470 114.390 ;
        RECT 127.840 110.960 128.010 114.220 ;
        RECT 128.735 113.650 136.775 113.820 ;
        RECT 128.350 111.590 128.520 113.590 ;
        RECT 136.990 111.590 137.160 113.590 ;
        RECT 128.735 111.360 136.775 111.530 ;
        RECT 137.500 110.960 138.470 114.220 ;
        RECT 127.840 110.790 138.470 110.960 ;
        RECT 127.840 107.530 128.010 110.790 ;
        RECT 128.735 110.220 136.775 110.390 ;
        RECT 128.350 108.160 128.520 110.160 ;
        RECT 136.990 108.160 137.160 110.160 ;
        RECT 128.735 107.930 136.775 108.100 ;
        RECT 137.500 107.530 138.470 110.790 ;
        RECT 120.020 107.410 126.260 107.510 ;
        RECT 87.155 104.665 88.110 104.885 ;
        RECT 87.385 104.035 87.655 104.495 ;
        RECT 87.825 104.205 88.110 104.665 ;
        RECT 89.315 104.035 90.525 105.125 ;
        RECT 107.910 105.100 108.080 107.360 ;
        RECT 108.805 106.790 116.845 106.960 ;
        RECT 108.420 105.730 108.590 106.730 ;
        RECT 117.060 105.730 117.230 106.730 ;
        RECT 108.805 105.500 116.845 105.670 ;
        RECT 117.570 105.100 118.540 107.360 ;
        RECT 120.010 106.850 126.260 107.410 ;
        RECT 120.010 106.830 125.180 106.850 ;
        RECT 120.010 106.760 124.000 106.830 ;
        RECT 120.010 106.250 121.930 106.760 ;
        RECT 123.440 106.750 124.000 106.760 ;
        RECT 107.910 105.070 118.540 105.100 ;
        RECT 107.880 104.960 118.540 105.070 ;
        RECT 106.130 104.910 118.540 104.960 ;
        RECT 101.790 104.740 118.540 104.910 ;
        RECT 11.950 103.865 90.610 104.035 ;
        RECT 12.035 102.775 13.245 103.865 ;
        RECT 12.035 102.065 12.555 102.605 ;
        RECT 12.725 102.235 13.245 102.775 ;
        RECT 13.415 102.895 13.685 103.665 ;
        RECT 13.855 103.085 14.185 103.865 ;
        RECT 14.390 103.260 14.575 103.665 ;
        RECT 14.745 103.440 15.080 103.865 ;
        RECT 14.390 103.085 15.055 103.260 ;
        RECT 13.415 102.725 14.545 102.895 ;
        RECT 12.035 101.315 13.245 102.065 ;
        RECT 13.415 101.815 13.585 102.725 ;
        RECT 13.755 101.975 14.115 102.555 ;
        RECT 14.295 102.225 14.545 102.725 ;
        RECT 14.715 102.055 15.055 103.085 ;
        RECT 16.175 102.725 16.455 103.865 ;
        RECT 16.625 102.715 16.955 103.695 ;
        RECT 17.125 102.725 17.385 103.865 ;
        RECT 17.670 103.235 17.955 103.695 ;
        RECT 18.125 103.405 18.395 103.865 ;
        RECT 17.670 103.015 18.625 103.235 ;
        RECT 16.185 102.285 16.520 102.555 ;
        RECT 16.690 102.115 16.860 102.715 ;
        RECT 17.030 102.305 17.365 102.555 ;
        RECT 17.555 102.285 18.245 102.845 ;
        RECT 18.415 102.115 18.625 103.015 ;
        RECT 14.370 101.885 15.055 102.055 ;
        RECT 13.415 101.485 13.675 101.815 ;
        RECT 13.885 101.315 14.160 101.795 ;
        RECT 14.370 101.485 14.575 101.885 ;
        RECT 14.745 101.315 15.080 101.715 ;
        RECT 16.175 101.315 16.485 102.115 ;
        RECT 16.690 101.485 17.385 102.115 ;
        RECT 17.670 101.945 18.625 102.115 ;
        RECT 18.795 102.845 19.195 103.695 ;
        RECT 19.385 103.235 19.665 103.695 ;
        RECT 20.185 103.405 20.510 103.865 ;
        RECT 19.385 103.015 20.510 103.235 ;
        RECT 18.795 102.285 19.890 102.845 ;
        RECT 20.060 102.555 20.510 103.015 ;
        RECT 20.680 102.725 21.065 103.695 ;
        RECT 21.695 103.355 21.995 103.865 ;
        RECT 22.165 103.185 22.495 103.695 ;
        RECT 22.665 103.355 23.295 103.865 ;
        RECT 23.875 103.355 24.255 103.525 ;
        RECT 24.425 103.355 24.725 103.865 ;
        RECT 24.085 103.185 24.255 103.355 ;
        RECT 17.670 101.485 17.955 101.945 ;
        RECT 18.125 101.315 18.395 101.775 ;
        RECT 18.795 101.485 19.195 102.285 ;
        RECT 20.060 102.225 20.615 102.555 ;
        RECT 20.060 102.115 20.510 102.225 ;
        RECT 19.385 101.945 20.510 102.115 ;
        RECT 20.785 102.055 21.065 102.725 ;
        RECT 19.385 101.485 19.665 101.945 ;
        RECT 20.185 101.315 20.510 101.775 ;
        RECT 20.680 101.485 21.065 102.055 ;
        RECT 21.695 103.015 23.915 103.185 ;
        RECT 21.695 102.055 21.865 103.015 ;
        RECT 22.035 102.675 23.575 102.845 ;
        RECT 22.035 102.225 22.280 102.675 ;
        RECT 22.540 102.305 23.235 102.505 ;
        RECT 23.405 102.475 23.575 102.675 ;
        RECT 23.745 102.815 23.915 103.015 ;
        RECT 24.085 102.985 24.745 103.185 ;
        RECT 23.745 102.645 24.405 102.815 ;
        RECT 23.405 102.305 24.005 102.475 ;
        RECT 24.235 102.225 24.405 102.645 ;
        RECT 21.695 101.510 22.160 102.055 ;
        RECT 22.665 101.315 22.835 102.135 ;
        RECT 23.005 102.055 23.915 102.135 ;
        RECT 24.575 102.055 24.745 102.985 ;
        RECT 24.915 102.700 25.205 103.865 ;
        RECT 25.465 103.195 25.635 103.695 ;
        RECT 25.805 103.365 26.135 103.865 ;
        RECT 25.465 103.025 26.130 103.195 ;
        RECT 25.380 102.205 25.730 102.855 ;
        RECT 23.005 101.965 24.255 102.055 ;
        RECT 23.005 101.485 23.335 101.965 ;
        RECT 23.745 101.885 24.255 101.965 ;
        RECT 23.505 101.315 23.855 101.705 ;
        RECT 24.025 101.485 24.255 101.885 ;
        RECT 24.425 101.575 24.745 102.055 ;
        RECT 24.915 101.315 25.205 102.040 ;
        RECT 25.900 102.035 26.130 103.025 ;
        RECT 25.465 101.865 26.130 102.035 ;
        RECT 25.465 101.575 25.635 101.865 ;
        RECT 25.805 101.315 26.135 101.695 ;
        RECT 26.305 101.575 26.490 103.695 ;
        RECT 26.730 103.405 26.995 103.865 ;
        RECT 27.165 103.270 27.415 103.695 ;
        RECT 27.625 103.420 28.730 103.590 ;
        RECT 27.110 103.140 27.415 103.270 ;
        RECT 26.660 101.945 26.940 102.895 ;
        RECT 27.110 102.035 27.280 103.140 ;
        RECT 27.450 102.355 27.690 102.950 ;
        RECT 27.860 102.885 28.390 103.250 ;
        RECT 27.860 102.185 28.030 102.885 ;
        RECT 28.560 102.805 28.730 103.420 ;
        RECT 28.900 103.065 29.070 103.865 ;
        RECT 29.240 103.365 29.490 103.695 ;
        RECT 29.715 103.395 30.600 103.565 ;
        RECT 28.560 102.715 29.070 102.805 ;
        RECT 27.110 101.905 27.335 102.035 ;
        RECT 27.505 101.965 28.030 102.185 ;
        RECT 28.200 102.545 29.070 102.715 ;
        RECT 26.745 101.315 26.995 101.775 ;
        RECT 27.165 101.765 27.335 101.905 ;
        RECT 28.200 101.765 28.370 102.545 ;
        RECT 28.900 102.475 29.070 102.545 ;
        RECT 28.580 102.295 28.780 102.325 ;
        RECT 29.240 102.295 29.410 103.365 ;
        RECT 29.580 102.475 29.770 103.195 ;
        RECT 28.580 101.995 29.410 102.295 ;
        RECT 29.940 102.265 30.260 103.225 ;
        RECT 27.165 101.595 27.500 101.765 ;
        RECT 27.695 101.595 28.370 101.765 ;
        RECT 28.690 101.315 29.060 101.815 ;
        RECT 29.240 101.765 29.410 101.995 ;
        RECT 29.795 101.935 30.260 102.265 ;
        RECT 30.430 102.555 30.600 103.395 ;
        RECT 30.780 103.365 31.095 103.865 ;
        RECT 31.325 103.135 31.665 103.695 ;
        RECT 30.770 102.760 31.665 103.135 ;
        RECT 31.835 102.855 32.005 103.865 ;
        RECT 31.475 102.555 31.665 102.760 ;
        RECT 32.175 102.805 32.505 103.650 ;
        RECT 32.175 102.725 32.565 102.805 ;
        RECT 32.735 102.775 36.245 103.865 ;
        RECT 32.350 102.675 32.565 102.725 ;
        RECT 30.430 102.225 31.305 102.555 ;
        RECT 31.475 102.225 32.225 102.555 ;
        RECT 30.430 101.765 30.600 102.225 ;
        RECT 31.475 102.055 31.675 102.225 ;
        RECT 32.395 102.095 32.565 102.675 ;
        RECT 32.340 102.055 32.565 102.095 ;
        RECT 29.240 101.595 29.645 101.765 ;
        RECT 29.815 101.595 30.600 101.765 ;
        RECT 30.875 101.315 31.085 101.845 ;
        RECT 31.345 101.530 31.675 102.055 ;
        RECT 32.185 101.970 32.565 102.055 ;
        RECT 32.735 102.085 34.385 102.605 ;
        RECT 34.555 102.255 36.245 102.775 ;
        RECT 36.875 102.725 37.135 103.865 ;
        RECT 37.305 102.715 37.635 103.695 ;
        RECT 37.805 102.725 38.085 103.865 ;
        RECT 38.720 102.915 38.985 103.685 ;
        RECT 39.155 103.145 39.485 103.865 ;
        RECT 39.675 103.325 39.935 103.685 ;
        RECT 40.105 103.495 40.435 103.865 ;
        RECT 40.605 103.325 40.865 103.685 ;
        RECT 39.675 103.095 40.865 103.325 ;
        RECT 41.435 102.915 41.725 103.685 ;
        RECT 36.895 102.305 37.230 102.555 ;
        RECT 37.400 102.115 37.570 102.715 ;
        RECT 37.740 102.285 38.075 102.555 ;
        RECT 31.845 101.315 32.015 101.925 ;
        RECT 32.185 101.535 32.515 101.970 ;
        RECT 32.735 101.315 36.245 102.085 ;
        RECT 36.875 101.485 37.570 102.115 ;
        RECT 37.775 101.315 38.085 102.115 ;
        RECT 38.720 101.495 39.055 102.915 ;
        RECT 39.230 102.735 41.725 102.915 ;
        RECT 39.230 102.045 39.455 102.735 ;
        RECT 41.935 102.725 42.225 103.865 ;
        RECT 43.020 103.525 44.385 103.695 ;
        RECT 43.020 103.315 43.350 103.525 ;
        RECT 42.395 103.065 43.350 103.315 ;
        RECT 39.655 102.225 39.935 102.555 ;
        RECT 40.115 102.225 40.690 102.555 ;
        RECT 40.870 102.225 41.305 102.555 ;
        RECT 41.485 102.225 41.755 102.555 ;
        RECT 41.935 102.225 42.210 102.555 ;
        RECT 42.395 102.055 42.565 103.065 ;
        RECT 42.735 102.225 43.090 102.890 ;
        RECT 43.275 102.225 43.550 102.890 ;
        RECT 43.720 102.555 44.045 103.355 ;
        RECT 44.215 102.895 44.385 103.525 ;
        RECT 44.555 103.065 44.845 103.865 ;
        RECT 44.215 102.725 44.890 102.895 ;
        RECT 45.060 102.725 45.445 103.685 ;
        RECT 45.615 102.775 49.125 103.865 ;
        RECT 44.720 102.555 44.890 102.725 ;
        RECT 43.720 102.225 44.065 102.555 ;
        RECT 44.275 102.305 44.525 102.555 ;
        RECT 44.720 102.305 45.085 102.555 ;
        RECT 44.355 102.225 44.525 102.305 ;
        RECT 44.895 102.225 45.085 102.305 ;
        RECT 45.270 102.055 45.445 102.725 ;
        RECT 39.230 101.855 41.715 102.045 ;
        RECT 39.235 101.315 39.980 101.685 ;
        RECT 40.545 101.495 40.800 101.855 ;
        RECT 40.980 101.315 41.310 101.685 ;
        RECT 41.490 101.495 41.715 101.855 ;
        RECT 41.935 101.695 42.225 101.965 ;
        RECT 42.395 101.865 42.820 102.055 ;
        RECT 42.990 101.885 44.390 102.055 ;
        RECT 42.990 101.695 43.320 101.885 ;
        RECT 41.935 101.485 43.320 101.695 ;
        RECT 43.555 101.315 43.885 101.715 ;
        RECT 44.060 101.485 44.390 101.885 ;
        RECT 44.595 101.315 44.765 101.875 ;
        RECT 44.935 101.485 45.445 102.055 ;
        RECT 45.615 102.085 47.265 102.605 ;
        RECT 47.435 102.255 49.125 102.775 ;
        RECT 49.355 102.725 49.565 103.865 ;
        RECT 49.735 102.715 50.065 103.695 ;
        RECT 50.235 102.725 50.465 103.865 ;
        RECT 45.615 101.315 49.125 102.085 ;
        RECT 49.355 101.315 49.565 102.135 ;
        RECT 49.735 102.115 49.985 102.715 ;
        RECT 50.675 102.700 50.965 103.865 ;
        RECT 52.115 102.805 52.445 103.650 ;
        RECT 52.615 102.855 52.785 103.865 ;
        RECT 52.955 103.135 53.295 103.695 ;
        RECT 53.525 103.365 53.840 103.865 ;
        RECT 54.020 103.395 54.905 103.565 ;
        RECT 52.055 102.725 52.445 102.805 ;
        RECT 52.955 102.760 53.850 103.135 ;
        RECT 52.055 102.675 52.270 102.725 ;
        RECT 50.155 102.305 50.485 102.555 ;
        RECT 49.735 101.485 50.065 102.115 ;
        RECT 50.235 101.315 50.465 102.135 ;
        RECT 52.055 102.095 52.225 102.675 ;
        RECT 52.955 102.555 53.145 102.760 ;
        RECT 54.020 102.555 54.190 103.395 ;
        RECT 55.130 103.365 55.380 103.695 ;
        RECT 52.395 102.225 53.145 102.555 ;
        RECT 53.315 102.225 54.190 102.555 ;
        RECT 52.055 102.055 52.280 102.095 ;
        RECT 52.945 102.055 53.145 102.225 ;
        RECT 50.675 101.315 50.965 102.040 ;
        RECT 52.055 101.970 52.435 102.055 ;
        RECT 52.105 101.535 52.435 101.970 ;
        RECT 52.605 101.315 52.775 101.925 ;
        RECT 52.945 101.530 53.275 102.055 ;
        RECT 53.535 101.315 53.745 101.845 ;
        RECT 54.020 101.765 54.190 102.225 ;
        RECT 54.360 102.265 54.680 103.225 ;
        RECT 54.850 102.475 55.040 103.195 ;
        RECT 55.210 102.295 55.380 103.365 ;
        RECT 55.550 103.065 55.720 103.865 ;
        RECT 55.890 103.420 56.995 103.590 ;
        RECT 55.890 102.805 56.060 103.420 ;
        RECT 57.205 103.270 57.455 103.695 ;
        RECT 57.625 103.405 57.890 103.865 ;
        RECT 56.230 102.885 56.760 103.250 ;
        RECT 57.205 103.140 57.510 103.270 ;
        RECT 55.550 102.715 56.060 102.805 ;
        RECT 55.550 102.545 56.420 102.715 ;
        RECT 55.550 102.475 55.720 102.545 ;
        RECT 55.840 102.295 56.040 102.325 ;
        RECT 54.360 101.935 54.825 102.265 ;
        RECT 55.210 101.995 56.040 102.295 ;
        RECT 55.210 101.765 55.380 101.995 ;
        RECT 54.020 101.595 54.805 101.765 ;
        RECT 54.975 101.595 55.380 101.765 ;
        RECT 55.560 101.315 55.930 101.815 ;
        RECT 56.250 101.765 56.420 102.545 ;
        RECT 56.590 102.185 56.760 102.885 ;
        RECT 56.930 102.355 57.170 102.950 ;
        RECT 56.590 101.965 57.115 102.185 ;
        RECT 57.340 102.035 57.510 103.140 ;
        RECT 57.285 101.905 57.510 102.035 ;
        RECT 57.680 101.945 57.960 102.895 ;
        RECT 57.285 101.765 57.455 101.905 ;
        RECT 56.250 101.595 56.925 101.765 ;
        RECT 57.120 101.595 57.455 101.765 ;
        RECT 57.625 101.315 57.875 101.775 ;
        RECT 58.130 101.575 58.315 103.695 ;
        RECT 58.485 103.365 58.815 103.865 ;
        RECT 58.985 103.195 59.155 103.695 ;
        RECT 58.490 103.025 59.155 103.195 ;
        RECT 58.490 102.035 58.720 103.025 ;
        RECT 58.890 102.205 59.240 102.855 ;
        RECT 59.420 102.725 59.755 103.695 ;
        RECT 59.925 102.725 60.095 103.865 ;
        RECT 60.265 103.525 62.295 103.695 ;
        RECT 59.420 102.055 59.590 102.725 ;
        RECT 60.265 102.555 60.435 103.525 ;
        RECT 59.760 102.225 60.015 102.555 ;
        RECT 60.240 102.225 60.435 102.555 ;
        RECT 60.605 103.185 61.730 103.355 ;
        RECT 59.845 102.055 60.015 102.225 ;
        RECT 60.605 102.055 60.775 103.185 ;
        RECT 58.490 101.865 59.155 102.035 ;
        RECT 58.485 101.315 58.815 101.695 ;
        RECT 58.985 101.575 59.155 101.865 ;
        RECT 59.420 101.485 59.675 102.055 ;
        RECT 59.845 101.885 60.775 102.055 ;
        RECT 60.945 102.845 61.955 103.015 ;
        RECT 60.945 102.045 61.115 102.845 ;
        RECT 61.320 102.165 61.595 102.645 ;
        RECT 61.315 101.995 61.595 102.165 ;
        RECT 60.600 101.850 60.775 101.885 ;
        RECT 59.845 101.315 60.175 101.715 ;
        RECT 60.600 101.485 61.130 101.850 ;
        RECT 61.320 101.485 61.595 101.995 ;
        RECT 61.765 101.485 61.955 102.845 ;
        RECT 62.125 102.860 62.295 103.525 ;
        RECT 62.465 103.105 62.635 103.865 ;
        RECT 62.870 103.105 63.385 103.515 ;
        RECT 62.125 102.670 62.875 102.860 ;
        RECT 63.045 102.295 63.385 103.105 ;
        RECT 63.645 102.935 63.815 103.695 ;
        RECT 64.030 103.105 64.360 103.865 ;
        RECT 63.645 102.765 64.360 102.935 ;
        RECT 64.530 102.790 64.785 103.695 ;
        RECT 62.155 102.125 63.385 102.295 ;
        RECT 63.555 102.215 63.910 102.585 ;
        RECT 64.190 102.555 64.360 102.765 ;
        RECT 64.190 102.225 64.445 102.555 ;
        RECT 62.135 101.315 62.645 101.850 ;
        RECT 62.865 101.520 63.110 102.125 ;
        RECT 64.190 102.035 64.360 102.225 ;
        RECT 64.615 102.060 64.785 102.790 ;
        RECT 64.960 102.715 65.220 103.865 ;
        RECT 65.405 102.895 65.735 103.680 ;
        RECT 65.405 102.725 66.085 102.895 ;
        RECT 66.265 102.725 66.595 103.865 ;
        RECT 66.775 102.775 70.285 103.865 ;
        RECT 65.395 102.305 65.745 102.555 ;
        RECT 63.645 101.865 64.360 102.035 ;
        RECT 63.645 101.485 63.815 101.865 ;
        RECT 64.030 101.315 64.360 101.695 ;
        RECT 64.530 101.485 64.785 102.060 ;
        RECT 64.960 101.315 65.220 102.155 ;
        RECT 65.915 102.125 66.085 102.725 ;
        RECT 66.255 102.305 66.605 102.555 ;
        RECT 65.415 101.315 65.655 102.125 ;
        RECT 65.825 101.485 66.155 102.125 ;
        RECT 66.325 101.315 66.595 102.125 ;
        RECT 66.775 102.085 68.425 102.605 ;
        RECT 68.595 102.255 70.285 102.775 ;
        RECT 71.375 102.725 71.635 103.865 ;
        RECT 71.805 102.715 72.135 103.695 ;
        RECT 72.305 102.725 72.585 103.865 ;
        RECT 71.895 102.675 72.070 102.715 ;
        RECT 72.755 102.685 73.075 103.865 ;
        RECT 73.245 102.845 73.445 103.635 ;
        RECT 73.770 103.035 74.155 103.695 ;
        RECT 74.550 103.105 75.335 103.865 ;
        RECT 73.745 102.935 74.155 103.035 ;
        RECT 73.245 102.675 73.575 102.845 ;
        RECT 73.745 102.725 75.355 102.935 ;
        RECT 71.395 102.305 71.730 102.555 ;
        RECT 71.900 102.115 72.070 102.675 ;
        RECT 73.395 102.555 73.575 102.675 ;
        RECT 72.240 102.285 72.575 102.555 ;
        RECT 72.755 102.305 73.220 102.505 ;
        RECT 73.395 102.305 73.725 102.555 ;
        RECT 73.895 102.505 74.360 102.555 ;
        RECT 73.895 102.335 74.365 102.505 ;
        RECT 73.895 102.305 74.360 102.335 ;
        RECT 74.555 102.305 74.910 102.555 ;
        RECT 75.080 102.125 75.355 102.725 ;
        RECT 66.775 101.315 70.285 102.085 ;
        RECT 71.375 101.485 72.070 102.115 ;
        RECT 72.275 101.315 72.585 102.115 ;
        RECT 72.755 101.925 73.935 102.095 ;
        RECT 72.755 101.510 73.095 101.925 ;
        RECT 73.265 101.315 73.435 101.755 ;
        RECT 73.605 101.705 73.935 101.925 ;
        RECT 74.105 101.945 75.355 102.125 ;
        RECT 74.105 101.875 74.470 101.945 ;
        RECT 73.605 101.525 74.855 101.705 ;
        RECT 75.125 101.315 75.295 101.775 ;
        RECT 75.525 101.595 75.805 103.695 ;
        RECT 76.435 102.700 76.725 103.865 ;
        RECT 76.895 102.775 78.565 103.865 ;
        RECT 79.285 103.195 79.455 103.695 ;
        RECT 79.625 103.365 79.955 103.865 ;
        RECT 79.285 103.025 79.950 103.195 ;
        RECT 76.895 102.085 77.645 102.605 ;
        RECT 77.815 102.255 78.565 102.775 ;
        RECT 79.200 102.205 79.550 102.855 ;
        RECT 76.435 101.315 76.725 102.040 ;
        RECT 76.895 101.315 78.565 102.085 ;
        RECT 79.720 102.035 79.950 103.025 ;
        RECT 79.285 101.865 79.950 102.035 ;
        RECT 79.285 101.575 79.455 101.865 ;
        RECT 79.625 101.315 79.955 101.695 ;
        RECT 80.125 101.575 80.310 103.695 ;
        RECT 80.550 103.405 80.815 103.865 ;
        RECT 80.985 103.270 81.235 103.695 ;
        RECT 81.445 103.420 82.550 103.590 ;
        RECT 80.930 103.140 81.235 103.270 ;
        RECT 80.480 101.945 80.760 102.895 ;
        RECT 80.930 102.035 81.100 103.140 ;
        RECT 81.270 102.355 81.510 102.950 ;
        RECT 81.680 102.885 82.210 103.250 ;
        RECT 81.680 102.185 81.850 102.885 ;
        RECT 82.380 102.805 82.550 103.420 ;
        RECT 82.720 103.065 82.890 103.865 ;
        RECT 83.060 103.365 83.310 103.695 ;
        RECT 83.535 103.395 84.420 103.565 ;
        RECT 82.380 102.715 82.890 102.805 ;
        RECT 80.930 101.905 81.155 102.035 ;
        RECT 81.325 101.965 81.850 102.185 ;
        RECT 82.020 102.545 82.890 102.715 ;
        RECT 80.565 101.315 80.815 101.775 ;
        RECT 80.985 101.765 81.155 101.905 ;
        RECT 82.020 101.765 82.190 102.545 ;
        RECT 82.720 102.475 82.890 102.545 ;
        RECT 82.400 102.295 82.600 102.325 ;
        RECT 83.060 102.295 83.230 103.365 ;
        RECT 83.400 102.475 83.590 103.195 ;
        RECT 82.400 101.995 83.230 102.295 ;
        RECT 83.760 102.265 84.080 103.225 ;
        RECT 80.985 101.595 81.320 101.765 ;
        RECT 81.515 101.595 82.190 101.765 ;
        RECT 82.510 101.315 82.880 101.815 ;
        RECT 83.060 101.765 83.230 101.995 ;
        RECT 83.615 101.935 84.080 102.265 ;
        RECT 84.250 102.555 84.420 103.395 ;
        RECT 84.600 103.365 84.915 103.865 ;
        RECT 85.145 103.135 85.485 103.695 ;
        RECT 84.590 102.760 85.485 103.135 ;
        RECT 85.655 102.855 85.825 103.865 ;
        RECT 85.295 102.555 85.485 102.760 ;
        RECT 85.995 102.805 86.325 103.650 ;
        RECT 85.995 102.725 86.385 102.805 ;
        RECT 86.555 102.775 89.145 103.865 ;
        RECT 86.170 102.675 86.385 102.725 ;
        RECT 84.250 102.225 85.125 102.555 ;
        RECT 85.295 102.225 86.045 102.555 ;
        RECT 84.250 101.765 84.420 102.225 ;
        RECT 85.295 102.055 85.495 102.225 ;
        RECT 86.215 102.095 86.385 102.675 ;
        RECT 86.160 102.055 86.385 102.095 ;
        RECT 83.060 101.595 83.465 101.765 ;
        RECT 83.635 101.595 84.420 101.765 ;
        RECT 84.695 101.315 84.905 101.845 ;
        RECT 85.165 101.530 85.495 102.055 ;
        RECT 86.005 101.970 86.385 102.055 ;
        RECT 86.555 102.085 87.765 102.605 ;
        RECT 87.935 102.255 89.145 102.775 ;
        RECT 89.315 102.775 90.525 103.865 ;
        RECT 101.790 103.330 101.960 104.740 ;
        RECT 102.330 104.170 105.370 104.340 ;
        RECT 102.330 103.730 105.370 103.900 ;
        RECT 105.585 103.870 105.755 104.200 ;
        RECT 106.090 103.980 118.540 104.740 ;
        RECT 120.000 105.490 121.930 106.250 ;
        RECT 123.670 105.660 124.000 106.750 ;
        RECT 124.370 106.280 125.410 106.450 ;
        RECT 124.370 105.840 125.410 106.010 ;
        RECT 125.580 105.980 125.750 106.310 ;
        RECT 106.090 103.970 118.430 103.980 ;
        RECT 106.090 103.960 111.970 103.970 ;
        RECT 106.090 103.940 106.660 103.960 ;
        RECT 107.880 103.950 111.970 103.960 ;
        RECT 106.100 103.330 106.270 103.940 ;
        RECT 101.790 103.160 106.270 103.330 ;
        RECT 89.315 102.235 89.835 102.775 ;
        RECT 120.000 102.740 120.960 105.490 ;
        RECT 123.830 105.440 124.000 105.660 ;
        RECT 126.090 105.440 126.260 106.850 ;
        RECT 123.830 105.270 126.260 105.440 ;
        RECT 127.840 107.360 138.470 107.530 ;
        RECT 140.050 116.640 146.280 116.800 ;
        RECT 140.050 114.380 140.720 116.640 ;
        RECT 141.390 116.070 145.430 116.240 ;
        RECT 141.050 115.010 141.220 116.010 ;
        RECT 145.600 115.010 145.770 116.010 ;
        RECT 141.390 114.780 145.430 114.950 ;
        RECT 146.110 114.380 146.280 116.640 ;
        RECT 140.050 114.210 146.280 114.380 ;
        RECT 140.050 110.950 140.720 114.210 ;
        RECT 141.390 113.640 145.430 113.810 ;
        RECT 141.050 111.580 141.220 113.580 ;
        RECT 145.600 111.580 145.770 113.580 ;
        RECT 141.390 111.350 145.430 111.520 ;
        RECT 146.110 110.950 146.280 114.210 ;
        RECT 140.050 110.780 146.280 110.950 ;
        RECT 140.050 107.520 140.720 110.780 ;
        RECT 141.390 110.210 145.430 110.380 ;
        RECT 141.050 108.150 141.220 110.150 ;
        RECT 145.600 108.150 145.770 110.150 ;
        RECT 141.390 107.920 145.430 108.090 ;
        RECT 146.110 107.520 146.280 110.780 ;
        RECT 140.050 107.510 146.280 107.520 ;
        RECT 147.870 116.780 157.700 116.820 ;
        RECT 147.870 116.650 158.500 116.780 ;
        RECT 147.870 114.390 148.040 116.650 ;
        RECT 148.765 116.080 156.805 116.250 ;
        RECT 148.380 115.020 148.550 116.020 ;
        RECT 157.020 115.020 157.190 116.020 ;
        RECT 148.765 114.790 156.805 114.960 ;
        RECT 157.530 114.390 158.500 116.650 ;
        RECT 147.870 114.220 158.500 114.390 ;
        RECT 147.870 110.960 148.040 114.220 ;
        RECT 148.765 113.650 156.805 113.820 ;
        RECT 148.380 111.590 148.550 113.590 ;
        RECT 157.020 111.590 157.190 113.590 ;
        RECT 148.765 111.360 156.805 111.530 ;
        RECT 157.530 110.960 158.500 114.220 ;
        RECT 147.870 110.790 158.500 110.960 ;
        RECT 147.870 107.530 148.040 110.790 ;
        RECT 148.765 110.220 156.805 110.390 ;
        RECT 148.380 108.160 148.550 110.160 ;
        RECT 157.020 108.160 157.190 110.160 ;
        RECT 148.765 107.930 156.805 108.100 ;
        RECT 157.530 107.530 158.500 110.790 ;
        RECT 140.050 107.410 146.290 107.510 ;
        RECT 127.840 105.100 128.010 107.360 ;
        RECT 128.735 106.790 136.775 106.960 ;
        RECT 128.350 105.730 128.520 106.730 ;
        RECT 136.990 105.730 137.160 106.730 ;
        RECT 128.735 105.500 136.775 105.670 ;
        RECT 137.500 105.100 138.470 107.360 ;
        RECT 140.040 106.850 146.290 107.410 ;
        RECT 140.040 106.830 145.210 106.850 ;
        RECT 140.040 106.760 144.030 106.830 ;
        RECT 140.040 105.490 141.960 106.760 ;
        RECT 143.470 106.750 144.030 106.760 ;
        RECT 143.700 105.660 144.030 106.750 ;
        RECT 144.400 106.280 145.440 106.450 ;
        RECT 144.400 105.840 145.440 106.010 ;
        RECT 145.610 105.980 145.780 106.310 ;
        RECT 143.860 105.440 144.030 105.660 ;
        RECT 146.120 105.440 146.290 106.850 ;
        RECT 143.860 105.270 146.290 105.440 ;
        RECT 147.870 107.360 158.500 107.530 ;
        RECT 127.840 105.070 138.470 105.100 ;
        RECT 147.870 105.100 148.040 107.360 ;
        RECT 148.765 106.790 156.805 106.960 ;
        RECT 148.380 105.730 148.550 106.730 ;
        RECT 157.020 105.730 157.190 106.730 ;
        RECT 148.765 105.500 156.805 105.670 ;
        RECT 157.530 105.100 158.500 107.360 ;
        RECT 147.870 105.070 158.500 105.100 ;
        RECT 127.810 104.960 138.470 105.070 ;
        RECT 147.840 104.960 158.500 105.070 ;
        RECT 126.060 104.910 138.470 104.960 ;
        RECT 146.090 104.910 158.500 104.960 ;
        RECT 121.720 104.740 138.470 104.910 ;
        RECT 121.720 103.330 121.890 104.740 ;
        RECT 122.260 104.170 125.300 104.340 ;
        RECT 122.260 103.730 125.300 103.900 ;
        RECT 125.515 103.870 125.685 104.200 ;
        RECT 126.020 103.980 138.470 104.740 ;
        RECT 141.750 104.740 158.500 104.910 ;
        RECT 126.020 103.970 138.360 103.980 ;
        RECT 126.020 103.960 131.900 103.970 ;
        RECT 126.020 103.940 126.590 103.960 ;
        RECT 127.810 103.950 131.900 103.960 ;
        RECT 126.030 103.330 126.200 103.940 ;
        RECT 121.720 103.160 126.200 103.330 ;
        RECT 141.750 103.330 141.920 104.740 ;
        RECT 142.290 104.170 145.330 104.340 ;
        RECT 142.290 103.730 145.330 103.900 ;
        RECT 145.545 103.870 145.715 104.200 ;
        RECT 146.050 103.980 158.500 104.740 ;
        RECT 146.050 103.970 158.390 103.980 ;
        RECT 146.050 103.960 151.930 103.970 ;
        RECT 146.050 103.940 146.620 103.960 ;
        RECT 147.840 103.950 151.930 103.960 ;
        RECT 146.060 103.330 146.230 103.940 ;
        RECT 141.750 103.160 146.230 103.330 ;
        RECT 85.665 101.315 85.835 101.925 ;
        RECT 86.005 101.535 86.335 101.970 ;
        RECT 86.555 101.315 89.145 102.085 ;
        RECT 90.005 102.065 90.525 102.605 ;
        RECT 89.315 101.315 90.525 102.065 ;
        RECT 120.000 102.570 158.300 102.740 ;
        RECT 120.000 101.720 134.620 102.570 ;
        RECT 120.000 101.650 120.960 101.720 ;
        RECT 11.950 101.145 90.610 101.315 ;
        RECT 12.035 100.395 13.245 101.145 ;
        RECT 13.505 100.595 13.675 100.885 ;
        RECT 13.845 100.765 14.175 101.145 ;
        RECT 13.505 100.425 14.170 100.595 ;
        RECT 12.035 99.855 12.555 100.395 ;
        RECT 12.725 99.685 13.245 100.225 ;
        RECT 12.035 98.595 13.245 99.685 ;
        RECT 13.420 99.605 13.770 100.255 ;
        RECT 13.940 99.435 14.170 100.425 ;
        RECT 13.505 99.265 14.170 99.435 ;
        RECT 13.505 98.765 13.675 99.265 ;
        RECT 13.845 98.595 14.175 99.095 ;
        RECT 14.345 98.765 14.530 100.885 ;
        RECT 14.785 100.685 15.035 101.145 ;
        RECT 15.205 100.695 15.540 100.865 ;
        RECT 15.735 100.695 16.410 100.865 ;
        RECT 15.205 100.555 15.375 100.695 ;
        RECT 14.700 99.565 14.980 100.515 ;
        RECT 15.150 100.425 15.375 100.555 ;
        RECT 15.150 99.320 15.320 100.425 ;
        RECT 15.545 100.275 16.070 100.495 ;
        RECT 15.490 99.510 15.730 100.105 ;
        RECT 15.900 99.575 16.070 100.275 ;
        RECT 16.240 99.915 16.410 100.695 ;
        RECT 16.730 100.645 17.100 101.145 ;
        RECT 17.280 100.695 17.685 100.865 ;
        RECT 17.855 100.695 18.640 100.865 ;
        RECT 17.280 100.465 17.450 100.695 ;
        RECT 16.620 100.165 17.450 100.465 ;
        RECT 17.835 100.195 18.300 100.525 ;
        RECT 16.620 100.135 16.820 100.165 ;
        RECT 16.940 99.915 17.110 99.985 ;
        RECT 16.240 99.745 17.110 99.915 ;
        RECT 16.600 99.655 17.110 99.745 ;
        RECT 15.150 99.190 15.455 99.320 ;
        RECT 15.900 99.210 16.430 99.575 ;
        RECT 14.770 98.595 15.035 99.055 ;
        RECT 15.205 98.765 15.455 99.190 ;
        RECT 16.600 99.040 16.770 99.655 ;
        RECT 15.665 98.870 16.770 99.040 ;
        RECT 16.940 98.595 17.110 99.395 ;
        RECT 17.280 99.095 17.450 100.165 ;
        RECT 17.620 99.265 17.810 99.985 ;
        RECT 17.980 99.235 18.300 100.195 ;
        RECT 18.470 100.235 18.640 100.695 ;
        RECT 18.915 100.615 19.125 101.145 ;
        RECT 19.385 100.405 19.715 100.930 ;
        RECT 19.885 100.535 20.055 101.145 ;
        RECT 20.225 100.490 20.555 100.925 ;
        RECT 20.780 100.890 21.115 100.935 ;
        RECT 20.225 100.405 20.605 100.490 ;
        RECT 19.515 100.235 19.715 100.405 ;
        RECT 20.380 100.365 20.605 100.405 ;
        RECT 18.470 99.905 19.345 100.235 ;
        RECT 19.515 99.905 20.265 100.235 ;
        RECT 17.280 98.765 17.530 99.095 ;
        RECT 18.470 99.065 18.640 99.905 ;
        RECT 19.515 99.700 19.705 99.905 ;
        RECT 20.435 99.785 20.605 100.365 ;
        RECT 20.390 99.735 20.605 99.785 ;
        RECT 18.810 99.325 19.705 99.700 ;
        RECT 20.215 99.655 20.605 99.735 ;
        RECT 20.775 100.425 21.115 100.890 ;
        RECT 21.285 100.765 21.615 101.145 ;
        RECT 22.075 100.805 22.345 100.810 ;
        RECT 22.075 100.635 22.385 100.805 ;
        RECT 20.775 99.735 20.945 100.425 ;
        RECT 21.115 99.905 21.375 100.235 ;
        RECT 17.755 98.895 18.640 99.065 ;
        RECT 18.820 98.595 19.135 99.095 ;
        RECT 19.365 98.765 19.705 99.325 ;
        RECT 19.875 98.595 20.045 99.605 ;
        RECT 20.215 98.810 20.545 99.655 ;
        RECT 20.775 98.765 21.035 99.735 ;
        RECT 21.205 99.355 21.375 99.905 ;
        RECT 21.545 99.535 21.885 100.565 ;
        RECT 22.075 99.535 22.345 100.635 ;
        RECT 22.570 99.535 22.850 100.810 ;
        RECT 23.050 100.645 23.280 100.975 ;
        RECT 23.525 100.765 23.855 101.145 ;
        RECT 23.050 99.355 23.220 100.645 ;
        RECT 24.025 100.575 24.200 100.975 ;
        RECT 23.570 100.405 24.200 100.575 ;
        RECT 23.570 100.235 23.740 100.405 ;
        RECT 24.455 100.345 24.765 101.145 ;
        RECT 24.970 100.345 25.665 100.975 ;
        RECT 25.835 100.600 31.180 101.145 ;
        RECT 31.355 100.600 36.700 101.145 ;
        RECT 24.970 100.295 25.145 100.345 ;
        RECT 23.390 99.905 23.740 100.235 ;
        RECT 21.205 99.185 23.220 99.355 ;
        RECT 23.570 99.385 23.740 99.905 ;
        RECT 23.920 99.555 24.285 100.235 ;
        RECT 24.465 99.905 24.800 100.175 ;
        RECT 24.970 99.745 25.140 100.295 ;
        RECT 25.310 99.905 25.645 100.155 ;
        RECT 27.420 99.770 27.760 100.600 ;
        RECT 23.570 99.215 24.200 99.385 ;
        RECT 21.230 98.595 21.560 99.005 ;
        RECT 21.760 98.765 21.930 99.185 ;
        RECT 22.145 98.595 22.815 99.005 ;
        RECT 23.050 98.765 23.220 99.185 ;
        RECT 23.525 98.595 23.855 99.035 ;
        RECT 24.025 98.765 24.200 99.215 ;
        RECT 24.455 98.595 24.735 99.735 ;
        RECT 24.905 98.765 25.235 99.745 ;
        RECT 25.405 98.595 25.665 99.735 ;
        RECT 29.240 99.030 29.590 100.280 ;
        RECT 32.940 99.770 33.280 100.600 ;
        RECT 37.795 100.420 38.085 101.145 ;
        RECT 38.255 100.375 40.845 101.145 ;
        RECT 41.480 100.405 41.735 100.975 ;
        RECT 41.905 100.745 42.235 101.145 ;
        RECT 42.660 100.610 43.190 100.975 ;
        RECT 43.380 100.805 43.655 100.975 ;
        RECT 43.375 100.635 43.655 100.805 ;
        RECT 42.660 100.575 42.835 100.610 ;
        RECT 41.905 100.405 42.835 100.575 ;
        RECT 34.760 99.030 35.110 100.280 ;
        RECT 38.255 99.855 39.465 100.375 ;
        RECT 25.835 98.595 31.180 99.030 ;
        RECT 31.355 98.595 36.700 99.030 ;
        RECT 37.795 98.595 38.085 99.760 ;
        RECT 39.635 99.685 40.845 100.205 ;
        RECT 38.255 98.595 40.845 99.685 ;
        RECT 41.480 99.735 41.650 100.405 ;
        RECT 41.905 100.235 42.075 100.405 ;
        RECT 41.820 99.905 42.075 100.235 ;
        RECT 42.300 99.905 42.495 100.235 ;
        RECT 41.480 98.765 41.815 99.735 ;
        RECT 41.985 98.595 42.155 99.735 ;
        RECT 42.325 98.935 42.495 99.905 ;
        RECT 42.665 99.275 42.835 100.405 ;
        RECT 43.005 99.615 43.175 100.415 ;
        RECT 43.380 99.815 43.655 100.635 ;
        RECT 43.825 99.615 44.015 100.975 ;
        RECT 44.195 100.610 44.705 101.145 ;
        RECT 44.925 100.335 45.170 100.940 ;
        RECT 45.705 100.595 45.875 100.885 ;
        RECT 46.045 100.765 46.375 101.145 ;
        RECT 45.705 100.425 46.370 100.595 ;
        RECT 44.215 100.165 45.445 100.335 ;
        RECT 43.005 99.445 44.015 99.615 ;
        RECT 44.185 99.600 44.935 99.790 ;
        RECT 42.665 99.105 43.790 99.275 ;
        RECT 44.185 98.935 44.355 99.600 ;
        RECT 45.105 99.355 45.445 100.165 ;
        RECT 45.620 99.605 45.970 100.255 ;
        RECT 46.140 99.435 46.370 100.425 ;
        RECT 42.325 98.765 44.355 98.935 ;
        RECT 44.525 98.595 44.695 99.355 ;
        RECT 44.930 98.945 45.445 99.355 ;
        RECT 45.705 99.265 46.370 99.435 ;
        RECT 45.705 98.765 45.875 99.265 ;
        RECT 46.045 98.595 46.375 99.095 ;
        RECT 46.545 98.765 46.730 100.885 ;
        RECT 46.985 100.685 47.235 101.145 ;
        RECT 47.405 100.695 47.740 100.865 ;
        RECT 47.935 100.695 48.610 100.865 ;
        RECT 47.405 100.555 47.575 100.695 ;
        RECT 46.900 99.565 47.180 100.515 ;
        RECT 47.350 100.425 47.575 100.555 ;
        RECT 47.350 99.320 47.520 100.425 ;
        RECT 47.745 100.275 48.270 100.495 ;
        RECT 47.690 99.510 47.930 100.105 ;
        RECT 48.100 99.575 48.270 100.275 ;
        RECT 48.440 99.915 48.610 100.695 ;
        RECT 48.930 100.645 49.300 101.145 ;
        RECT 49.480 100.695 49.885 100.865 ;
        RECT 50.055 100.695 50.840 100.865 ;
        RECT 49.480 100.465 49.650 100.695 ;
        RECT 48.820 100.165 49.650 100.465 ;
        RECT 50.035 100.195 50.500 100.525 ;
        RECT 48.820 100.135 49.020 100.165 ;
        RECT 49.140 99.915 49.310 99.985 ;
        RECT 48.440 99.745 49.310 99.915 ;
        RECT 48.800 99.655 49.310 99.745 ;
        RECT 47.350 99.190 47.655 99.320 ;
        RECT 48.100 99.210 48.630 99.575 ;
        RECT 46.970 98.595 47.235 99.055 ;
        RECT 47.405 98.765 47.655 99.190 ;
        RECT 48.800 99.040 48.970 99.655 ;
        RECT 47.865 98.870 48.970 99.040 ;
        RECT 49.140 98.595 49.310 99.395 ;
        RECT 49.480 99.095 49.650 100.165 ;
        RECT 49.820 99.265 50.010 99.985 ;
        RECT 50.180 99.235 50.500 100.195 ;
        RECT 50.670 100.235 50.840 100.695 ;
        RECT 51.115 100.615 51.325 101.145 ;
        RECT 51.585 100.405 51.915 100.930 ;
        RECT 52.085 100.535 52.255 101.145 ;
        RECT 52.425 100.490 52.755 100.925 ;
        RECT 53.160 100.665 53.330 101.145 ;
        RECT 53.500 100.495 53.830 100.965 ;
        RECT 54.000 100.665 54.170 101.145 ;
        RECT 54.340 100.495 54.670 100.965 ;
        RECT 52.425 100.405 52.805 100.490 ;
        RECT 51.715 100.235 51.915 100.405 ;
        RECT 52.580 100.365 52.805 100.405 ;
        RECT 50.670 99.905 51.545 100.235 ;
        RECT 51.715 99.905 52.465 100.235 ;
        RECT 49.480 98.765 49.730 99.095 ;
        RECT 50.670 99.065 50.840 99.905 ;
        RECT 51.715 99.700 51.905 99.905 ;
        RECT 52.635 99.785 52.805 100.365 ;
        RECT 52.590 99.735 52.805 99.785 ;
        RECT 51.010 99.325 51.905 99.700 ;
        RECT 52.415 99.655 52.805 99.735 ;
        RECT 52.975 100.325 54.670 100.495 ;
        RECT 54.880 100.405 55.050 101.145 ;
        RECT 55.265 100.405 55.595 100.940 ;
        RECT 55.765 100.635 56.005 101.145 ;
        RECT 56.285 100.595 56.455 100.885 ;
        RECT 56.625 100.765 56.955 101.145 ;
        RECT 52.975 99.735 53.320 100.325 ;
        RECT 53.490 99.985 54.700 100.155 ;
        RECT 54.495 99.735 54.700 99.985 ;
        RECT 54.870 99.905 55.245 100.235 ;
        RECT 55.415 99.735 55.595 100.405 ;
        RECT 55.765 99.905 56.020 100.465 ;
        RECT 56.285 100.425 56.950 100.595 ;
        RECT 49.955 98.895 50.840 99.065 ;
        RECT 51.020 98.595 51.335 99.095 ;
        RECT 51.565 98.765 51.905 99.325 ;
        RECT 52.075 98.595 52.245 99.605 ;
        RECT 52.415 98.810 52.745 99.655 ;
        RECT 52.975 99.565 53.830 99.735 ;
        RECT 54.495 99.565 55.955 99.735 ;
        RECT 56.200 99.605 56.550 100.255 ;
        RECT 53.500 99.395 53.830 99.565 ;
        RECT 53.160 98.595 53.330 99.395 ;
        RECT 53.500 99.225 54.670 99.395 ;
        RECT 53.500 98.765 53.830 99.225 ;
        RECT 54.000 98.595 54.170 99.055 ;
        RECT 54.340 98.765 54.670 99.225 ;
        RECT 54.880 98.595 55.050 99.395 ;
        RECT 55.595 98.765 55.955 99.565 ;
        RECT 56.720 99.435 56.950 100.425 ;
        RECT 56.285 99.265 56.950 99.435 ;
        RECT 56.285 98.765 56.455 99.265 ;
        RECT 56.625 98.595 56.955 99.095 ;
        RECT 57.125 98.765 57.310 100.885 ;
        RECT 57.565 100.685 57.815 101.145 ;
        RECT 57.985 100.695 58.320 100.865 ;
        RECT 58.515 100.695 59.190 100.865 ;
        RECT 57.985 100.555 58.155 100.695 ;
        RECT 57.480 99.565 57.760 100.515 ;
        RECT 57.930 100.425 58.155 100.555 ;
        RECT 57.930 99.320 58.100 100.425 ;
        RECT 58.325 100.275 58.850 100.495 ;
        RECT 58.270 99.510 58.510 100.105 ;
        RECT 58.680 99.575 58.850 100.275 ;
        RECT 59.020 99.915 59.190 100.695 ;
        RECT 59.510 100.645 59.880 101.145 ;
        RECT 60.060 100.695 60.465 100.865 ;
        RECT 60.635 100.695 61.420 100.865 ;
        RECT 60.060 100.465 60.230 100.695 ;
        RECT 59.400 100.165 60.230 100.465 ;
        RECT 60.615 100.195 61.080 100.525 ;
        RECT 59.400 100.135 59.600 100.165 ;
        RECT 59.720 99.915 59.890 99.985 ;
        RECT 59.020 99.745 59.890 99.915 ;
        RECT 59.380 99.655 59.890 99.745 ;
        RECT 57.930 99.190 58.235 99.320 ;
        RECT 58.680 99.210 59.210 99.575 ;
        RECT 57.550 98.595 57.815 99.055 ;
        RECT 57.985 98.765 58.235 99.190 ;
        RECT 59.380 99.040 59.550 99.655 ;
        RECT 58.445 98.870 59.550 99.040 ;
        RECT 59.720 98.595 59.890 99.395 ;
        RECT 60.060 99.095 60.230 100.165 ;
        RECT 60.400 99.265 60.590 99.985 ;
        RECT 60.760 99.235 61.080 100.195 ;
        RECT 61.250 100.235 61.420 100.695 ;
        RECT 61.695 100.615 61.905 101.145 ;
        RECT 62.165 100.405 62.495 100.930 ;
        RECT 62.665 100.535 62.835 101.145 ;
        RECT 63.005 100.490 63.335 100.925 ;
        RECT 63.005 100.405 63.385 100.490 ;
        RECT 63.555 100.420 63.845 101.145 ;
        RECT 62.295 100.235 62.495 100.405 ;
        RECT 63.160 100.365 63.385 100.405 ;
        RECT 61.250 99.905 62.125 100.235 ;
        RECT 62.295 99.905 63.045 100.235 ;
        RECT 60.060 98.765 60.310 99.095 ;
        RECT 61.250 99.065 61.420 99.905 ;
        RECT 62.295 99.700 62.485 99.905 ;
        RECT 63.215 99.785 63.385 100.365 ;
        RECT 63.170 99.735 63.385 99.785 ;
        RECT 64.020 100.405 64.275 100.975 ;
        RECT 64.445 100.745 64.775 101.145 ;
        RECT 65.200 100.610 65.730 100.975 ;
        RECT 65.200 100.575 65.375 100.610 ;
        RECT 64.445 100.405 65.375 100.575 ;
        RECT 61.590 99.325 62.485 99.700 ;
        RECT 62.995 99.655 63.385 99.735 ;
        RECT 60.535 98.895 61.420 99.065 ;
        RECT 61.600 98.595 61.915 99.095 ;
        RECT 62.145 98.765 62.485 99.325 ;
        RECT 62.655 98.595 62.825 99.605 ;
        RECT 62.995 98.810 63.325 99.655 ;
        RECT 63.555 98.595 63.845 99.760 ;
        RECT 64.020 99.735 64.190 100.405 ;
        RECT 64.445 100.235 64.615 100.405 ;
        RECT 64.360 99.905 64.615 100.235 ;
        RECT 64.840 99.905 65.035 100.235 ;
        RECT 64.020 98.765 64.355 99.735 ;
        RECT 64.525 98.595 64.695 99.735 ;
        RECT 64.865 98.935 65.035 99.905 ;
        RECT 65.205 99.275 65.375 100.405 ;
        RECT 65.545 99.615 65.715 100.415 ;
        RECT 65.920 100.125 66.195 100.975 ;
        RECT 65.915 99.955 66.195 100.125 ;
        RECT 65.920 99.815 66.195 99.955 ;
        RECT 66.365 99.615 66.555 100.975 ;
        RECT 66.735 100.610 67.245 101.145 ;
        RECT 67.465 100.335 67.710 100.940 ;
        RECT 68.155 100.375 69.825 101.145 ;
        RECT 70.455 100.405 70.945 100.975 ;
        RECT 71.115 100.575 71.345 100.975 ;
        RECT 71.515 100.745 71.935 101.145 ;
        RECT 72.105 100.575 72.275 100.975 ;
        RECT 71.115 100.405 72.275 100.575 ;
        RECT 72.445 100.405 72.895 101.145 ;
        RECT 73.065 100.405 73.505 100.965 ;
        RECT 73.725 100.675 74.015 101.145 ;
        RECT 74.185 100.505 74.515 100.975 ;
        RECT 74.685 100.675 74.855 101.145 ;
        RECT 75.025 100.505 75.355 100.975 ;
        RECT 74.185 100.495 75.355 100.505 ;
        RECT 66.755 100.165 67.985 100.335 ;
        RECT 65.545 99.445 66.555 99.615 ;
        RECT 66.725 99.600 67.475 99.790 ;
        RECT 65.205 99.105 66.330 99.275 ;
        RECT 66.725 98.935 66.895 99.600 ;
        RECT 67.645 99.355 67.985 100.165 ;
        RECT 68.155 99.855 68.905 100.375 ;
        RECT 69.075 99.685 69.825 100.205 ;
        RECT 64.865 98.765 66.895 98.935 ;
        RECT 67.065 98.595 67.235 99.355 ;
        RECT 67.470 98.945 67.985 99.355 ;
        RECT 68.155 98.595 69.825 99.685 ;
        RECT 70.455 99.735 70.625 100.405 ;
        RECT 70.795 99.905 71.200 100.235 ;
        RECT 70.455 99.565 71.225 99.735 ;
        RECT 70.465 98.595 70.795 99.395 ;
        RECT 70.975 98.935 71.225 99.565 ;
        RECT 71.415 99.105 71.665 100.235 ;
        RECT 71.865 99.905 72.110 100.235 ;
        RECT 72.295 99.955 72.685 100.235 ;
        RECT 71.865 99.105 72.065 99.905 ;
        RECT 72.855 99.785 73.025 100.235 ;
        RECT 72.235 99.615 73.025 99.785 ;
        RECT 72.235 98.935 72.405 99.615 ;
        RECT 70.975 98.765 72.405 98.935 ;
        RECT 72.575 98.595 72.890 99.445 ;
        RECT 73.195 99.395 73.505 100.405 ;
        RECT 73.755 100.325 75.355 100.495 ;
        RECT 75.525 100.325 75.800 101.145 ;
        RECT 75.980 100.470 76.255 100.815 ;
        RECT 76.445 100.745 76.825 101.145 ;
        RECT 76.995 100.575 77.165 100.925 ;
        RECT 77.335 100.745 77.665 101.145 ;
        RECT 77.835 100.575 78.090 100.925 ;
        RECT 78.295 100.635 78.535 101.145 ;
        RECT 78.705 100.635 78.995 100.975 ;
        RECT 79.225 100.635 79.540 101.145 ;
        RECT 73.755 99.785 73.970 100.325 ;
        RECT 74.140 99.955 74.910 100.155 ;
        RECT 75.080 99.955 75.800 100.155 ;
        RECT 73.755 99.565 74.515 99.785 ;
        RECT 73.065 98.765 73.505 99.395 ;
        RECT 73.715 98.935 74.015 99.395 ;
        RECT 74.185 99.105 74.515 99.565 ;
        RECT 74.685 99.565 75.800 99.775 ;
        RECT 74.685 98.935 74.855 99.565 ;
        RECT 73.715 98.765 74.855 98.935 ;
        RECT 75.025 98.595 75.355 99.395 ;
        RECT 75.525 98.765 75.800 99.565 ;
        RECT 75.980 99.735 76.150 100.470 ;
        RECT 76.425 100.405 78.090 100.575 ;
        RECT 76.425 100.235 76.595 100.405 ;
        RECT 76.320 99.905 76.595 100.235 ;
        RECT 76.765 99.905 77.590 100.235 ;
        RECT 77.760 99.905 78.105 100.235 ;
        RECT 78.340 100.125 78.535 100.465 ;
        RECT 78.335 99.955 78.535 100.125 ;
        RECT 78.340 99.905 78.535 99.955 ;
        RECT 76.425 99.735 76.595 99.905 ;
        RECT 75.980 98.765 76.255 99.735 ;
        RECT 76.425 99.565 77.085 99.735 ;
        RECT 77.395 99.615 77.590 99.905 ;
        RECT 78.705 99.735 78.885 100.635 ;
        RECT 79.710 100.575 79.880 100.845 ;
        RECT 80.050 100.745 80.380 101.145 ;
        RECT 79.055 99.905 79.465 100.465 ;
        RECT 79.710 100.405 80.405 100.575 ;
        RECT 79.635 99.735 79.805 100.235 ;
        RECT 76.915 99.445 77.085 99.565 ;
        RECT 77.760 99.445 78.085 99.735 ;
        RECT 76.465 98.595 76.745 99.395 ;
        RECT 76.915 99.275 78.085 99.445 ;
        RECT 78.345 99.565 79.805 99.735 ;
        RECT 78.345 99.390 78.705 99.565 ;
        RECT 79.975 99.395 80.405 100.405 ;
        RECT 76.915 98.815 78.105 99.105 ;
        RECT 79.290 98.595 79.460 99.395 ;
        RECT 79.630 99.225 80.405 99.395 ;
        RECT 81.040 100.405 81.295 100.975 ;
        RECT 81.465 100.745 81.795 101.145 ;
        RECT 82.220 100.610 82.750 100.975 ;
        RECT 82.940 100.805 83.215 100.975 ;
        RECT 82.935 100.635 83.215 100.805 ;
        RECT 82.220 100.575 82.395 100.610 ;
        RECT 81.465 100.405 82.395 100.575 ;
        RECT 81.040 99.735 81.210 100.405 ;
        RECT 81.465 100.235 81.635 100.405 ;
        RECT 81.380 99.905 81.635 100.235 ;
        RECT 81.860 99.905 82.055 100.235 ;
        RECT 79.630 98.765 79.960 99.225 ;
        RECT 80.130 98.595 80.300 99.055 ;
        RECT 81.040 98.765 81.375 99.735 ;
        RECT 81.545 98.595 81.715 99.735 ;
        RECT 81.885 98.935 82.055 99.905 ;
        RECT 82.225 99.275 82.395 100.405 ;
        RECT 82.565 99.615 82.735 100.415 ;
        RECT 82.940 99.815 83.215 100.635 ;
        RECT 83.385 99.615 83.575 100.975 ;
        RECT 83.755 100.610 84.265 101.145 ;
        RECT 84.485 100.335 84.730 100.940 ;
        RECT 85.175 100.375 88.685 101.145 ;
        RECT 89.315 100.395 90.525 101.145 ;
        RECT 100.030 100.395 112.740 101.005 ;
        RECT 83.775 100.165 85.005 100.335 ;
        RECT 82.565 99.445 83.575 99.615 ;
        RECT 83.745 99.600 84.495 99.790 ;
        RECT 82.225 99.105 83.350 99.275 ;
        RECT 83.745 98.935 83.915 99.600 ;
        RECT 84.665 99.355 85.005 100.165 ;
        RECT 85.175 99.855 86.825 100.375 ;
        RECT 86.995 99.685 88.685 100.205 ;
        RECT 81.885 98.765 83.915 98.935 ;
        RECT 84.085 98.595 84.255 99.355 ;
        RECT 84.490 98.945 85.005 99.355 ;
        RECT 85.175 98.595 88.685 99.685 ;
        RECT 89.315 99.685 89.835 100.225 ;
        RECT 90.005 99.855 90.525 100.395 ;
        RECT 99.980 100.195 112.790 100.395 ;
        RECT 89.315 98.595 90.525 99.685 ;
        RECT 11.950 98.425 90.610 98.595 ;
        RECT 12.035 97.335 13.245 98.425 ;
        RECT 13.415 97.335 16.925 98.425 ;
        RECT 12.035 96.625 12.555 97.165 ;
        RECT 12.725 96.795 13.245 97.335 ;
        RECT 13.415 96.645 15.065 97.165 ;
        RECT 15.235 96.815 16.925 97.335 ;
        RECT 17.100 97.285 17.420 98.425 ;
        RECT 17.600 97.115 17.795 98.165 ;
        RECT 17.975 97.575 18.305 98.255 ;
        RECT 18.505 97.625 18.760 98.425 ;
        RECT 17.975 97.295 18.325 97.575 ;
        RECT 17.160 97.065 17.420 97.115 ;
        RECT 17.155 96.895 17.420 97.065 ;
        RECT 17.160 96.785 17.420 96.895 ;
        RECT 17.600 96.785 17.985 97.115 ;
        RECT 18.155 96.915 18.325 97.295 ;
        RECT 18.515 97.085 18.760 97.445 ;
        RECT 18.935 97.285 19.320 98.255 ;
        RECT 19.490 97.965 19.815 98.425 ;
        RECT 20.335 97.795 20.615 98.255 ;
        RECT 19.490 97.575 20.615 97.795 ;
        RECT 18.155 96.745 18.675 96.915 ;
        RECT 12.035 95.875 13.245 96.625 ;
        RECT 13.415 95.875 16.925 96.645 ;
        RECT 17.100 96.405 18.315 96.575 ;
        RECT 17.100 96.055 17.390 96.405 ;
        RECT 17.585 95.875 17.915 96.235 ;
        RECT 18.085 96.100 18.315 96.405 ;
        RECT 18.505 96.180 18.675 96.745 ;
        RECT 18.935 96.615 19.215 97.285 ;
        RECT 19.490 97.115 19.940 97.575 ;
        RECT 20.805 97.405 21.205 98.255 ;
        RECT 21.605 97.965 21.875 98.425 ;
        RECT 22.045 97.795 22.330 98.255 ;
        RECT 19.385 96.785 19.940 97.115 ;
        RECT 20.110 96.845 21.205 97.405 ;
        RECT 19.490 96.675 19.940 96.785 ;
        RECT 18.935 96.045 19.320 96.615 ;
        RECT 19.490 96.505 20.615 96.675 ;
        RECT 19.490 95.875 19.815 96.335 ;
        RECT 20.335 96.045 20.615 96.505 ;
        RECT 20.805 96.045 21.205 96.845 ;
        RECT 21.375 97.575 22.330 97.795 ;
        RECT 21.375 96.675 21.585 97.575 ;
        RECT 21.755 96.845 22.445 97.405 ;
        RECT 22.615 97.335 24.285 98.425 ;
        RECT 21.375 96.505 22.330 96.675 ;
        RECT 21.605 95.875 21.875 96.335 ;
        RECT 22.045 96.045 22.330 96.505 ;
        RECT 22.615 96.645 23.365 97.165 ;
        RECT 23.535 96.815 24.285 97.335 ;
        RECT 24.915 97.260 25.205 98.425 ;
        RECT 25.375 97.990 30.720 98.425 ;
        RECT 22.615 95.875 24.285 96.645 ;
        RECT 24.915 95.875 25.205 96.600 ;
        RECT 26.960 96.420 27.300 97.250 ;
        RECT 28.780 96.740 29.130 97.990 ;
        RECT 30.895 97.335 32.565 98.425 ;
        RECT 32.825 97.755 32.995 98.255 ;
        RECT 33.165 97.925 33.495 98.425 ;
        RECT 32.825 97.585 33.490 97.755 ;
        RECT 30.895 96.645 31.645 97.165 ;
        RECT 31.815 96.815 32.565 97.335 ;
        RECT 32.740 96.765 33.090 97.415 ;
        RECT 25.375 95.875 30.720 96.420 ;
        RECT 30.895 95.875 32.565 96.645 ;
        RECT 33.260 96.595 33.490 97.585 ;
        RECT 32.825 96.425 33.490 96.595 ;
        RECT 32.825 96.135 32.995 96.425 ;
        RECT 33.165 95.875 33.495 96.255 ;
        RECT 33.665 96.135 33.850 98.255 ;
        RECT 34.090 97.965 34.355 98.425 ;
        RECT 34.525 97.830 34.775 98.255 ;
        RECT 34.985 97.980 36.090 98.150 ;
        RECT 34.470 97.700 34.775 97.830 ;
        RECT 34.020 96.505 34.300 97.455 ;
        RECT 34.470 96.595 34.640 97.700 ;
        RECT 34.810 96.915 35.050 97.510 ;
        RECT 35.220 97.445 35.750 97.810 ;
        RECT 35.220 96.745 35.390 97.445 ;
        RECT 35.920 97.365 36.090 97.980 ;
        RECT 36.260 97.625 36.430 98.425 ;
        RECT 36.600 97.925 36.850 98.255 ;
        RECT 37.075 97.955 37.960 98.125 ;
        RECT 35.920 97.275 36.430 97.365 ;
        RECT 34.470 96.465 34.695 96.595 ;
        RECT 34.865 96.525 35.390 96.745 ;
        RECT 35.560 97.105 36.430 97.275 ;
        RECT 34.105 95.875 34.355 96.335 ;
        RECT 34.525 96.325 34.695 96.465 ;
        RECT 35.560 96.325 35.730 97.105 ;
        RECT 36.260 97.035 36.430 97.105 ;
        RECT 35.940 96.855 36.140 96.885 ;
        RECT 36.600 96.855 36.770 97.925 ;
        RECT 36.940 97.035 37.130 97.755 ;
        RECT 35.940 96.555 36.770 96.855 ;
        RECT 37.300 96.825 37.620 97.785 ;
        RECT 34.525 96.155 34.860 96.325 ;
        RECT 35.055 96.155 35.730 96.325 ;
        RECT 36.050 95.875 36.420 96.375 ;
        RECT 36.600 96.325 36.770 96.555 ;
        RECT 37.155 96.495 37.620 96.825 ;
        RECT 37.790 97.115 37.960 97.955 ;
        RECT 38.140 97.925 38.455 98.425 ;
        RECT 38.685 97.695 39.025 98.255 ;
        RECT 38.130 97.320 39.025 97.695 ;
        RECT 39.195 97.415 39.365 98.425 ;
        RECT 38.835 97.115 39.025 97.320 ;
        RECT 39.535 97.365 39.865 98.210 ;
        RECT 39.535 97.285 39.925 97.365 ;
        RECT 39.710 97.235 39.925 97.285 ;
        RECT 37.790 96.785 38.665 97.115 ;
        RECT 38.835 96.785 39.585 97.115 ;
        RECT 37.790 96.325 37.960 96.785 ;
        RECT 38.835 96.615 39.035 96.785 ;
        RECT 39.755 96.655 39.925 97.235 ;
        RECT 39.700 96.615 39.925 96.655 ;
        RECT 36.600 96.155 37.005 96.325 ;
        RECT 37.175 96.155 37.960 96.325 ;
        RECT 38.235 95.875 38.445 96.405 ;
        RECT 38.705 96.090 39.035 96.615 ;
        RECT 39.545 96.530 39.925 96.615 ;
        RECT 40.095 97.285 40.480 98.255 ;
        RECT 40.650 97.965 40.975 98.425 ;
        RECT 41.495 97.795 41.775 98.255 ;
        RECT 40.650 97.575 41.775 97.795 ;
        RECT 40.095 96.615 40.375 97.285 ;
        RECT 40.650 97.115 41.100 97.575 ;
        RECT 41.965 97.405 42.365 98.255 ;
        RECT 42.765 97.965 43.035 98.425 ;
        RECT 43.205 97.795 43.490 98.255 ;
        RECT 40.545 96.785 41.100 97.115 ;
        RECT 41.270 96.845 42.365 97.405 ;
        RECT 40.650 96.675 41.100 96.785 ;
        RECT 39.205 95.875 39.375 96.485 ;
        RECT 39.545 96.095 39.875 96.530 ;
        RECT 40.095 96.045 40.480 96.615 ;
        RECT 40.650 96.505 41.775 96.675 ;
        RECT 40.650 95.875 40.975 96.335 ;
        RECT 41.495 96.045 41.775 96.505 ;
        RECT 41.965 96.045 42.365 96.845 ;
        RECT 42.535 97.575 43.490 97.795 ;
        RECT 42.535 96.675 42.745 97.575 ;
        RECT 42.915 96.845 43.605 97.405 ;
        RECT 43.775 97.335 46.365 98.425 ;
        RECT 42.535 96.505 43.490 96.675 ;
        RECT 42.765 95.875 43.035 96.335 ;
        RECT 43.205 96.045 43.490 96.505 ;
        RECT 43.775 96.645 44.985 97.165 ;
        RECT 45.155 96.815 46.365 97.335 ;
        RECT 46.540 97.285 46.875 98.255 ;
        RECT 47.045 97.285 47.215 98.425 ;
        RECT 47.385 98.085 49.415 98.255 ;
        RECT 43.775 95.875 46.365 96.645 ;
        RECT 46.540 96.615 46.710 97.285 ;
        RECT 47.385 97.115 47.555 98.085 ;
        RECT 46.880 96.785 47.135 97.115 ;
        RECT 47.360 96.785 47.555 97.115 ;
        RECT 47.725 97.745 48.850 97.915 ;
        RECT 46.965 96.615 47.135 96.785 ;
        RECT 47.725 96.615 47.895 97.745 ;
        RECT 46.540 96.045 46.795 96.615 ;
        RECT 46.965 96.445 47.895 96.615 ;
        RECT 48.065 97.405 49.075 97.575 ;
        RECT 48.065 96.605 48.235 97.405 ;
        RECT 48.440 96.725 48.715 97.205 ;
        RECT 48.435 96.555 48.715 96.725 ;
        RECT 47.720 96.410 47.895 96.445 ;
        RECT 46.965 95.875 47.295 96.275 ;
        RECT 47.720 96.045 48.250 96.410 ;
        RECT 48.440 96.045 48.715 96.555 ;
        RECT 48.885 96.045 49.075 97.405 ;
        RECT 49.245 97.420 49.415 98.085 ;
        RECT 49.585 97.665 49.755 98.425 ;
        RECT 49.990 97.665 50.505 98.075 ;
        RECT 49.245 97.230 49.995 97.420 ;
        RECT 50.165 96.855 50.505 97.665 ;
        RECT 50.675 97.260 50.965 98.425 ;
        RECT 51.140 97.285 51.475 98.255 ;
        RECT 51.645 97.285 51.815 98.425 ;
        RECT 51.985 98.085 54.015 98.255 ;
        RECT 49.275 96.685 50.505 96.855 ;
        RECT 49.255 95.875 49.765 96.410 ;
        RECT 49.985 96.080 50.230 96.685 ;
        RECT 51.140 96.615 51.310 97.285 ;
        RECT 51.985 97.115 52.155 98.085 ;
        RECT 51.480 96.785 51.735 97.115 ;
        RECT 51.960 96.785 52.155 97.115 ;
        RECT 52.325 97.745 53.450 97.915 ;
        RECT 51.565 96.615 51.735 96.785 ;
        RECT 52.325 96.615 52.495 97.745 ;
        RECT 50.675 95.875 50.965 96.600 ;
        RECT 51.140 96.045 51.395 96.615 ;
        RECT 51.565 96.445 52.495 96.615 ;
        RECT 52.665 97.405 53.675 97.575 ;
        RECT 52.665 96.605 52.835 97.405 ;
        RECT 53.040 97.065 53.315 97.205 ;
        RECT 53.035 96.895 53.315 97.065 ;
        RECT 52.320 96.410 52.495 96.445 ;
        RECT 51.565 95.875 51.895 96.275 ;
        RECT 52.320 96.045 52.850 96.410 ;
        RECT 53.040 96.045 53.315 96.895 ;
        RECT 53.485 96.045 53.675 97.405 ;
        RECT 53.845 97.420 54.015 98.085 ;
        RECT 54.185 97.665 54.355 98.425 ;
        RECT 54.590 97.665 55.105 98.075 ;
        RECT 53.845 97.230 54.595 97.420 ;
        RECT 54.765 96.855 55.105 97.665 ;
        RECT 55.275 97.335 58.785 98.425 ;
        RECT 58.955 97.335 60.165 98.425 ;
        RECT 60.450 97.795 60.735 98.255 ;
        RECT 60.905 97.965 61.175 98.425 ;
        RECT 60.450 97.575 61.405 97.795 ;
        RECT 53.875 96.685 55.105 96.855 ;
        RECT 53.855 95.875 54.365 96.410 ;
        RECT 54.585 96.080 54.830 96.685 ;
        RECT 55.275 96.645 56.925 97.165 ;
        RECT 57.095 96.815 58.785 97.335 ;
        RECT 55.275 95.875 58.785 96.645 ;
        RECT 58.955 96.625 59.475 97.165 ;
        RECT 59.645 96.795 60.165 97.335 ;
        RECT 60.335 96.845 61.025 97.405 ;
        RECT 61.195 96.675 61.405 97.575 ;
        RECT 58.955 95.875 60.165 96.625 ;
        RECT 60.450 96.505 61.405 96.675 ;
        RECT 61.575 97.405 61.975 98.255 ;
        RECT 62.165 97.795 62.445 98.255 ;
        RECT 62.965 97.965 63.290 98.425 ;
        RECT 62.165 97.575 63.290 97.795 ;
        RECT 61.575 96.845 62.670 97.405 ;
        RECT 62.840 97.115 63.290 97.575 ;
        RECT 63.460 97.285 63.845 98.255 ;
        RECT 64.015 97.335 65.685 98.425 ;
        RECT 60.450 96.045 60.735 96.505 ;
        RECT 60.905 95.875 61.175 96.335 ;
        RECT 61.575 96.045 61.975 96.845 ;
        RECT 62.840 96.785 63.395 97.115 ;
        RECT 62.840 96.675 63.290 96.785 ;
        RECT 62.165 96.505 63.290 96.675 ;
        RECT 63.565 96.615 63.845 97.285 ;
        RECT 62.165 96.045 62.445 96.505 ;
        RECT 62.965 95.875 63.290 96.335 ;
        RECT 63.460 96.045 63.845 96.615 ;
        RECT 64.015 96.645 64.765 97.165 ;
        RECT 64.935 96.815 65.685 97.335 ;
        RECT 65.855 97.555 66.130 98.255 ;
        RECT 66.300 97.880 66.555 98.425 ;
        RECT 66.725 97.915 67.205 98.255 ;
        RECT 67.380 97.870 67.985 98.425 ;
        RECT 67.370 97.770 67.985 97.870 ;
        RECT 67.370 97.745 67.555 97.770 ;
        RECT 64.015 95.875 65.685 96.645 ;
        RECT 65.855 96.525 66.025 97.555 ;
        RECT 66.300 97.425 67.055 97.675 ;
        RECT 67.225 97.500 67.555 97.745 ;
        RECT 66.300 97.390 67.070 97.425 ;
        RECT 66.300 97.380 67.085 97.390 ;
        RECT 66.195 97.365 67.090 97.380 ;
        RECT 66.195 97.350 67.110 97.365 ;
        RECT 66.195 97.340 67.130 97.350 ;
        RECT 66.195 97.330 67.155 97.340 ;
        RECT 66.195 97.300 67.225 97.330 ;
        RECT 66.195 97.270 67.245 97.300 ;
        RECT 66.195 97.240 67.265 97.270 ;
        RECT 66.195 97.215 67.295 97.240 ;
        RECT 66.195 97.180 67.330 97.215 ;
        RECT 66.195 97.175 67.360 97.180 ;
        RECT 66.195 96.780 66.425 97.175 ;
        RECT 66.970 97.170 67.360 97.175 ;
        RECT 66.995 97.160 67.360 97.170 ;
        RECT 67.010 97.155 67.360 97.160 ;
        RECT 67.025 97.150 67.360 97.155 ;
        RECT 67.725 97.150 67.985 97.600 ;
        RECT 68.165 97.455 68.495 98.240 ;
        RECT 68.165 97.285 68.845 97.455 ;
        RECT 69.025 97.285 69.355 98.425 ;
        RECT 69.535 97.335 72.125 98.425 ;
        RECT 72.755 97.915 73.945 98.205 ;
        RECT 67.025 97.145 67.985 97.150 ;
        RECT 67.035 97.135 67.985 97.145 ;
        RECT 67.045 97.130 67.985 97.135 ;
        RECT 67.055 97.120 67.985 97.130 ;
        RECT 67.060 97.110 67.985 97.120 ;
        RECT 67.065 97.105 67.985 97.110 ;
        RECT 67.075 97.090 67.985 97.105 ;
        RECT 67.080 97.075 67.985 97.090 ;
        RECT 67.090 97.050 67.985 97.075 ;
        RECT 66.595 96.580 66.925 97.005 ;
        RECT 65.855 96.045 66.115 96.525 ;
        RECT 66.285 95.875 66.535 96.415 ;
        RECT 66.705 96.095 66.925 96.580 ;
        RECT 67.095 96.980 67.985 97.050 ;
        RECT 67.095 96.255 67.265 96.980 ;
        RECT 68.155 96.865 68.505 97.115 ;
        RECT 67.435 96.425 67.985 96.810 ;
        RECT 68.675 96.685 68.845 97.285 ;
        RECT 69.015 96.865 69.365 97.115 ;
        RECT 67.095 96.085 67.985 96.255 ;
        RECT 68.175 95.875 68.415 96.685 ;
        RECT 68.585 96.045 68.915 96.685 ;
        RECT 69.085 95.875 69.355 96.685 ;
        RECT 69.535 96.645 70.745 97.165 ;
        RECT 70.915 96.815 72.125 97.335 ;
        RECT 72.775 97.575 73.945 97.745 ;
        RECT 74.115 97.625 74.395 98.425 ;
        RECT 72.775 97.285 73.100 97.575 ;
        RECT 73.775 97.455 73.945 97.575 ;
        RECT 73.270 97.115 73.465 97.405 ;
        RECT 73.775 97.285 74.435 97.455 ;
        RECT 74.605 97.285 74.880 98.255 ;
        RECT 75.055 97.335 76.265 98.425 ;
        RECT 74.265 97.115 74.435 97.285 ;
        RECT 72.755 96.785 73.100 97.115 ;
        RECT 73.270 96.785 74.095 97.115 ;
        RECT 74.265 96.785 74.540 97.115 ;
        RECT 69.535 95.875 72.125 96.645 ;
        RECT 74.265 96.615 74.435 96.785 ;
        RECT 72.770 96.445 74.435 96.615 ;
        RECT 74.710 96.550 74.880 97.285 ;
        RECT 72.770 96.095 73.025 96.445 ;
        RECT 73.195 95.875 73.525 96.275 ;
        RECT 73.695 96.095 73.865 96.445 ;
        RECT 74.035 95.875 74.415 96.275 ;
        RECT 74.605 96.205 74.880 96.550 ;
        RECT 75.055 96.625 75.575 97.165 ;
        RECT 75.745 96.795 76.265 97.335 ;
        RECT 76.435 97.260 76.725 98.425 ;
        RECT 77.815 97.665 78.330 98.075 ;
        RECT 78.565 97.665 78.735 98.425 ;
        RECT 78.905 98.085 80.935 98.255 ;
        RECT 77.815 96.855 78.155 97.665 ;
        RECT 78.905 97.420 79.075 98.085 ;
        RECT 79.470 97.745 80.595 97.915 ;
        RECT 78.325 97.230 79.075 97.420 ;
        RECT 79.245 97.405 80.255 97.575 ;
        RECT 77.815 96.685 79.045 96.855 ;
        RECT 75.055 95.875 76.265 96.625 ;
        RECT 76.435 95.875 76.725 96.600 ;
        RECT 78.090 96.080 78.335 96.685 ;
        RECT 78.555 95.875 79.065 96.410 ;
        RECT 79.245 96.045 79.435 97.405 ;
        RECT 79.605 96.385 79.880 97.205 ;
        RECT 80.085 96.605 80.255 97.405 ;
        RECT 80.425 96.615 80.595 97.745 ;
        RECT 80.765 97.115 80.935 98.085 ;
        RECT 81.105 97.285 81.275 98.425 ;
        RECT 81.445 97.285 81.780 98.255 ;
        RECT 81.955 97.990 87.300 98.425 ;
        RECT 80.765 96.785 80.960 97.115 ;
        RECT 81.185 96.785 81.440 97.115 ;
        RECT 81.185 96.615 81.355 96.785 ;
        RECT 81.610 96.615 81.780 97.285 ;
        RECT 80.425 96.445 81.355 96.615 ;
        RECT 80.425 96.410 80.600 96.445 ;
        RECT 79.605 96.215 79.885 96.385 ;
        RECT 79.605 96.045 79.880 96.215 ;
        RECT 80.070 96.045 80.600 96.410 ;
        RECT 81.025 95.875 81.355 96.275 ;
        RECT 81.525 96.045 81.780 96.615 ;
        RECT 83.540 96.420 83.880 97.250 ;
        RECT 85.360 96.740 85.710 97.990 ;
        RECT 87.475 97.335 89.145 98.425 ;
        RECT 87.475 96.645 88.225 97.165 ;
        RECT 88.395 96.815 89.145 97.335 ;
        RECT 89.315 97.335 90.525 98.425 ;
        RECT 89.315 96.795 89.835 97.335 ;
        RECT 81.955 95.875 87.300 96.420 ;
        RECT 87.475 95.875 89.145 96.645 ;
        RECT 90.005 96.625 90.525 97.165 ;
        RECT 89.315 95.875 90.525 96.625 ;
        RECT 11.950 95.705 90.610 95.875 ;
        RECT 12.035 94.955 13.245 95.705 ;
        RECT 13.415 94.955 14.625 95.705 ;
        RECT 14.800 94.965 15.055 95.535 ;
        RECT 15.225 95.305 15.555 95.705 ;
        RECT 15.980 95.170 16.510 95.535 ;
        RECT 15.980 95.135 16.155 95.170 ;
        RECT 15.225 94.965 16.155 95.135 ;
        RECT 12.035 94.415 12.555 94.955 ;
        RECT 12.725 94.245 13.245 94.785 ;
        RECT 13.415 94.415 13.935 94.955 ;
        RECT 14.105 94.245 14.625 94.785 ;
        RECT 12.035 93.155 13.245 94.245 ;
        RECT 13.415 93.155 14.625 94.245 ;
        RECT 14.800 94.295 14.970 94.965 ;
        RECT 15.225 94.795 15.395 94.965 ;
        RECT 15.140 94.465 15.395 94.795 ;
        RECT 15.620 94.465 15.815 94.795 ;
        RECT 14.800 93.325 15.135 94.295 ;
        RECT 15.305 93.155 15.475 94.295 ;
        RECT 15.645 93.495 15.815 94.465 ;
        RECT 15.985 93.835 16.155 94.965 ;
        RECT 16.325 94.175 16.495 94.975 ;
        RECT 16.700 94.685 16.975 95.535 ;
        RECT 16.695 94.515 16.975 94.685 ;
        RECT 16.700 94.375 16.975 94.515 ;
        RECT 17.145 94.175 17.335 95.535 ;
        RECT 17.515 95.170 18.025 95.705 ;
        RECT 18.245 94.895 18.490 95.500 ;
        RECT 19.415 95.135 19.670 95.485 ;
        RECT 19.840 95.305 20.170 95.705 ;
        RECT 20.340 95.135 20.510 95.485 ;
        RECT 20.680 95.305 21.060 95.705 ;
        RECT 19.415 94.965 21.080 95.135 ;
        RECT 21.250 95.030 21.525 95.375 ;
        RECT 17.535 94.725 18.765 94.895 ;
        RECT 20.910 94.795 21.080 94.965 ;
        RECT 16.325 94.005 17.335 94.175 ;
        RECT 17.505 94.160 18.255 94.350 ;
        RECT 15.985 93.665 17.110 93.835 ;
        RECT 17.505 93.495 17.675 94.160 ;
        RECT 18.425 93.915 18.765 94.725 ;
        RECT 19.395 94.465 19.745 94.795 ;
        RECT 19.915 94.465 20.740 94.795 ;
        RECT 20.910 94.465 21.185 94.795 ;
        RECT 15.645 93.325 17.675 93.495 ;
        RECT 17.845 93.155 18.015 93.915 ;
        RECT 18.250 93.505 18.765 93.915 ;
        RECT 19.415 94.005 19.745 94.295 ;
        RECT 19.915 94.175 20.140 94.465 ;
        RECT 20.910 94.295 21.080 94.465 ;
        RECT 21.355 94.295 21.525 95.030 ;
        RECT 21.695 94.875 21.985 95.705 ;
        RECT 22.155 94.935 24.745 95.705 ;
        RECT 25.005 95.155 25.175 95.445 ;
        RECT 25.345 95.325 25.675 95.705 ;
        RECT 25.005 94.985 25.670 95.155 ;
        RECT 22.155 94.415 23.365 94.935 ;
        RECT 20.410 94.125 21.080 94.295 ;
        RECT 20.410 94.005 20.580 94.125 ;
        RECT 19.415 93.835 20.580 94.005 ;
        RECT 19.395 93.375 20.590 93.665 ;
        RECT 20.760 93.155 21.040 93.955 ;
        RECT 21.250 93.325 21.525 94.295 ;
        RECT 21.695 93.155 21.985 94.360 ;
        RECT 23.535 94.245 24.745 94.765 ;
        RECT 22.155 93.155 24.745 94.245 ;
        RECT 24.920 94.165 25.270 94.815 ;
        RECT 25.440 93.995 25.670 94.985 ;
        RECT 25.005 93.825 25.670 93.995 ;
        RECT 25.005 93.325 25.175 93.825 ;
        RECT 25.345 93.155 25.675 93.655 ;
        RECT 25.845 93.325 26.030 95.445 ;
        RECT 26.285 95.245 26.535 95.705 ;
        RECT 26.705 95.255 27.040 95.425 ;
        RECT 27.235 95.255 27.910 95.425 ;
        RECT 26.705 95.115 26.875 95.255 ;
        RECT 26.200 94.125 26.480 95.075 ;
        RECT 26.650 94.985 26.875 95.115 ;
        RECT 26.650 93.880 26.820 94.985 ;
        RECT 27.045 94.835 27.570 95.055 ;
        RECT 26.990 94.070 27.230 94.665 ;
        RECT 27.400 94.135 27.570 94.835 ;
        RECT 27.740 94.475 27.910 95.255 ;
        RECT 28.230 95.205 28.600 95.705 ;
        RECT 28.780 95.255 29.185 95.425 ;
        RECT 29.355 95.255 30.140 95.425 ;
        RECT 28.780 95.025 28.950 95.255 ;
        RECT 28.120 94.725 28.950 95.025 ;
        RECT 29.335 94.755 29.800 95.085 ;
        RECT 28.120 94.695 28.320 94.725 ;
        RECT 28.440 94.475 28.610 94.545 ;
        RECT 27.740 94.305 28.610 94.475 ;
        RECT 28.100 94.215 28.610 94.305 ;
        RECT 26.650 93.750 26.955 93.880 ;
        RECT 27.400 93.770 27.930 94.135 ;
        RECT 26.270 93.155 26.535 93.615 ;
        RECT 26.705 93.325 26.955 93.750 ;
        RECT 28.100 93.600 28.270 94.215 ;
        RECT 27.165 93.430 28.270 93.600 ;
        RECT 28.440 93.155 28.610 93.955 ;
        RECT 28.780 93.655 28.950 94.725 ;
        RECT 29.120 93.825 29.310 94.545 ;
        RECT 29.480 93.795 29.800 94.755 ;
        RECT 29.970 94.795 30.140 95.255 ;
        RECT 30.415 95.175 30.625 95.705 ;
        RECT 30.885 94.965 31.215 95.490 ;
        RECT 31.385 95.095 31.555 95.705 ;
        RECT 31.725 95.050 32.055 95.485 ;
        RECT 32.225 95.190 32.395 95.705 ;
        RECT 31.725 94.965 32.105 95.050 ;
        RECT 31.015 94.795 31.215 94.965 ;
        RECT 31.880 94.925 32.105 94.965 ;
        RECT 29.970 94.465 30.845 94.795 ;
        RECT 31.015 94.465 31.765 94.795 ;
        RECT 28.780 93.325 29.030 93.655 ;
        RECT 29.970 93.625 30.140 94.465 ;
        RECT 31.015 94.260 31.205 94.465 ;
        RECT 31.935 94.345 32.105 94.925 ;
        RECT 31.890 94.295 32.105 94.345 ;
        RECT 30.310 93.885 31.205 94.260 ;
        RECT 31.715 94.215 32.105 94.295 ;
        RECT 33.660 94.965 33.915 95.535 ;
        RECT 34.085 95.305 34.415 95.705 ;
        RECT 34.840 95.170 35.370 95.535 ;
        RECT 35.560 95.365 35.835 95.535 ;
        RECT 35.555 95.195 35.835 95.365 ;
        RECT 34.840 95.135 35.015 95.170 ;
        RECT 34.085 94.965 35.015 95.135 ;
        RECT 33.660 94.295 33.830 94.965 ;
        RECT 34.085 94.795 34.255 94.965 ;
        RECT 34.000 94.465 34.255 94.795 ;
        RECT 34.480 94.465 34.675 94.795 ;
        RECT 29.255 93.455 30.140 93.625 ;
        RECT 30.320 93.155 30.635 93.655 ;
        RECT 30.865 93.325 31.205 93.885 ;
        RECT 31.375 93.155 31.545 94.165 ;
        RECT 31.715 93.370 32.045 94.215 ;
        RECT 32.215 93.155 32.385 94.070 ;
        RECT 33.660 93.325 33.995 94.295 ;
        RECT 34.165 93.155 34.335 94.295 ;
        RECT 34.505 93.495 34.675 94.465 ;
        RECT 34.845 93.835 35.015 94.965 ;
        RECT 35.185 94.175 35.355 94.975 ;
        RECT 35.560 94.375 35.835 95.195 ;
        RECT 36.005 94.175 36.195 95.535 ;
        RECT 36.375 95.170 36.885 95.705 ;
        RECT 37.105 94.895 37.350 95.500 ;
        RECT 37.795 94.980 38.085 95.705 ;
        RECT 38.720 94.965 38.975 95.535 ;
        RECT 39.145 95.305 39.475 95.705 ;
        RECT 39.900 95.170 40.430 95.535 ;
        RECT 39.900 95.135 40.075 95.170 ;
        RECT 39.145 94.965 40.075 95.135 ;
        RECT 36.395 94.725 37.625 94.895 ;
        RECT 35.185 94.005 36.195 94.175 ;
        RECT 36.365 94.160 37.115 94.350 ;
        RECT 34.845 93.665 35.970 93.835 ;
        RECT 36.365 93.495 36.535 94.160 ;
        RECT 37.285 93.915 37.625 94.725 ;
        RECT 34.505 93.325 36.535 93.495 ;
        RECT 36.705 93.155 36.875 93.915 ;
        RECT 37.110 93.505 37.625 93.915 ;
        RECT 37.795 93.155 38.085 94.320 ;
        RECT 38.720 94.295 38.890 94.965 ;
        RECT 39.145 94.795 39.315 94.965 ;
        RECT 39.060 94.465 39.315 94.795 ;
        RECT 39.540 94.465 39.735 94.795 ;
        RECT 38.720 93.325 39.055 94.295 ;
        RECT 39.225 93.155 39.395 94.295 ;
        RECT 39.565 93.495 39.735 94.465 ;
        RECT 39.905 93.835 40.075 94.965 ;
        RECT 40.245 94.175 40.415 94.975 ;
        RECT 40.620 94.685 40.895 95.535 ;
        RECT 40.615 94.515 40.895 94.685 ;
        RECT 40.620 94.375 40.895 94.515 ;
        RECT 41.065 94.175 41.255 95.535 ;
        RECT 41.435 95.170 41.945 95.705 ;
        RECT 42.165 94.895 42.410 95.500 ;
        RECT 42.855 95.325 43.745 95.495 ;
        RECT 41.455 94.725 42.685 94.895 ;
        RECT 42.855 94.770 43.405 95.155 ;
        RECT 40.245 94.005 41.255 94.175 ;
        RECT 41.425 94.160 42.175 94.350 ;
        RECT 39.905 93.665 41.030 93.835 ;
        RECT 41.425 93.495 41.595 94.160 ;
        RECT 42.345 93.915 42.685 94.725 ;
        RECT 43.575 94.600 43.745 95.325 ;
        RECT 42.855 94.530 43.745 94.600 ;
        RECT 43.915 95.000 44.135 95.485 ;
        RECT 44.305 95.165 44.555 95.705 ;
        RECT 44.725 95.055 44.985 95.535 ;
        RECT 45.155 95.160 50.500 95.705 ;
        RECT 43.915 94.575 44.245 95.000 ;
        RECT 42.855 94.505 43.750 94.530 ;
        RECT 42.855 94.490 43.760 94.505 ;
        RECT 42.855 94.475 43.765 94.490 ;
        RECT 42.855 94.470 43.775 94.475 ;
        RECT 42.855 94.460 43.780 94.470 ;
        RECT 42.855 94.450 43.785 94.460 ;
        RECT 42.855 94.445 43.795 94.450 ;
        RECT 42.855 94.435 43.805 94.445 ;
        RECT 42.855 94.430 43.815 94.435 ;
        RECT 42.855 93.980 43.115 94.430 ;
        RECT 43.480 94.425 43.815 94.430 ;
        RECT 43.480 94.420 43.830 94.425 ;
        RECT 43.480 94.410 43.845 94.420 ;
        RECT 43.480 94.405 43.870 94.410 ;
        RECT 44.415 94.405 44.645 94.800 ;
        RECT 43.480 94.400 44.645 94.405 ;
        RECT 43.510 94.365 44.645 94.400 ;
        RECT 43.545 94.340 44.645 94.365 ;
        RECT 43.575 94.310 44.645 94.340 ;
        RECT 43.595 94.280 44.645 94.310 ;
        RECT 43.615 94.250 44.645 94.280 ;
        RECT 43.685 94.240 44.645 94.250 ;
        RECT 43.710 94.230 44.645 94.240 ;
        RECT 43.730 94.215 44.645 94.230 ;
        RECT 43.750 94.200 44.645 94.215 ;
        RECT 43.755 94.190 44.540 94.200 ;
        RECT 43.770 94.155 44.540 94.190 ;
        RECT 39.565 93.325 41.595 93.495 ;
        RECT 41.765 93.155 41.935 93.915 ;
        RECT 42.170 93.505 42.685 93.915 ;
        RECT 43.285 93.835 43.615 94.080 ;
        RECT 43.785 93.905 44.540 94.155 ;
        RECT 44.815 94.025 44.985 95.055 ;
        RECT 46.740 94.330 47.080 95.160 ;
        RECT 50.675 94.935 53.265 95.705 ;
        RECT 53.945 95.050 54.275 95.485 ;
        RECT 54.445 95.095 54.615 95.705 ;
        RECT 53.895 94.965 54.275 95.050 ;
        RECT 54.785 94.965 55.115 95.490 ;
        RECT 55.375 95.175 55.585 95.705 ;
        RECT 55.860 95.255 56.645 95.425 ;
        RECT 56.815 95.255 57.220 95.425 ;
        RECT 43.285 93.810 43.470 93.835 ;
        RECT 42.855 93.710 43.470 93.810 ;
        RECT 42.855 93.155 43.460 93.710 ;
        RECT 43.635 93.325 44.115 93.665 ;
        RECT 44.285 93.155 44.540 93.700 ;
        RECT 44.710 93.325 44.985 94.025 ;
        RECT 48.560 93.590 48.910 94.840 ;
        RECT 50.675 94.415 51.885 94.935 ;
        RECT 53.895 94.925 54.120 94.965 ;
        RECT 52.055 94.245 53.265 94.765 ;
        RECT 45.155 93.155 50.500 93.590 ;
        RECT 50.675 93.155 53.265 94.245 ;
        RECT 53.895 94.345 54.065 94.925 ;
        RECT 54.785 94.795 54.985 94.965 ;
        RECT 55.860 94.795 56.030 95.255 ;
        RECT 54.235 94.465 54.985 94.795 ;
        RECT 55.155 94.465 56.030 94.795 ;
        RECT 53.895 94.295 54.110 94.345 ;
        RECT 53.895 94.215 54.285 94.295 ;
        RECT 53.955 93.370 54.285 94.215 ;
        RECT 54.795 94.260 54.985 94.465 ;
        RECT 54.455 93.155 54.625 94.165 ;
        RECT 54.795 93.885 55.690 94.260 ;
        RECT 54.795 93.325 55.135 93.885 ;
        RECT 55.365 93.155 55.680 93.655 ;
        RECT 55.860 93.625 56.030 94.465 ;
        RECT 56.200 94.755 56.665 95.085 ;
        RECT 57.050 95.025 57.220 95.255 ;
        RECT 57.400 95.205 57.770 95.705 ;
        RECT 58.090 95.255 58.765 95.425 ;
        RECT 58.960 95.255 59.295 95.425 ;
        RECT 56.200 93.795 56.520 94.755 ;
        RECT 57.050 94.725 57.880 95.025 ;
        RECT 56.690 93.825 56.880 94.545 ;
        RECT 57.050 93.655 57.220 94.725 ;
        RECT 57.680 94.695 57.880 94.725 ;
        RECT 57.390 94.475 57.560 94.545 ;
        RECT 58.090 94.475 58.260 95.255 ;
        RECT 59.125 95.115 59.295 95.255 ;
        RECT 59.465 95.245 59.715 95.705 ;
        RECT 57.390 94.305 58.260 94.475 ;
        RECT 58.430 94.835 58.955 95.055 ;
        RECT 59.125 94.985 59.350 95.115 ;
        RECT 57.390 94.215 57.900 94.305 ;
        RECT 55.860 93.455 56.745 93.625 ;
        RECT 56.970 93.325 57.220 93.655 ;
        RECT 57.390 93.155 57.560 93.955 ;
        RECT 57.730 93.600 57.900 94.215 ;
        RECT 58.430 94.135 58.600 94.835 ;
        RECT 58.070 93.770 58.600 94.135 ;
        RECT 58.770 94.070 59.010 94.665 ;
        RECT 59.180 93.880 59.350 94.985 ;
        RECT 59.520 94.125 59.800 95.075 ;
        RECT 59.045 93.750 59.350 93.880 ;
        RECT 57.730 93.430 58.835 93.600 ;
        RECT 59.045 93.325 59.295 93.750 ;
        RECT 59.465 93.155 59.730 93.615 ;
        RECT 59.970 93.325 60.155 95.445 ;
        RECT 60.325 95.325 60.655 95.705 ;
        RECT 60.825 95.155 60.995 95.445 ;
        RECT 60.330 94.985 60.995 95.155 ;
        RECT 60.330 93.995 60.560 94.985 ;
        RECT 61.255 94.935 62.925 95.705 ;
        RECT 63.555 94.980 63.845 95.705 ;
        RECT 64.015 95.205 64.275 95.535 ;
        RECT 64.445 95.345 64.775 95.705 ;
        RECT 65.030 95.325 66.330 95.535 ;
        RECT 64.015 95.195 64.245 95.205 ;
        RECT 60.730 94.165 61.080 94.815 ;
        RECT 61.255 94.415 62.005 94.935 ;
        RECT 62.175 94.245 62.925 94.765 ;
        RECT 60.330 93.825 60.995 93.995 ;
        RECT 60.325 93.155 60.655 93.655 ;
        RECT 60.825 93.325 60.995 93.825 ;
        RECT 61.255 93.155 62.925 94.245 ;
        RECT 63.555 93.155 63.845 94.320 ;
        RECT 64.015 94.005 64.185 95.195 ;
        RECT 65.030 95.175 65.200 95.325 ;
        RECT 64.445 95.050 65.200 95.175 ;
        RECT 64.355 95.005 65.200 95.050 ;
        RECT 64.355 94.885 64.625 95.005 ;
        RECT 64.355 94.310 64.525 94.885 ;
        RECT 64.755 94.445 65.165 94.750 ;
        RECT 65.455 94.715 65.665 95.115 ;
        RECT 65.335 94.505 65.665 94.715 ;
        RECT 65.910 94.715 66.130 95.115 ;
        RECT 66.605 94.940 67.060 95.705 ;
        RECT 65.910 94.505 66.385 94.715 ;
        RECT 66.575 94.515 67.065 94.715 ;
        RECT 64.355 94.275 64.555 94.310 ;
        RECT 65.885 94.275 67.060 94.335 ;
        RECT 64.355 94.165 67.060 94.275 ;
        RECT 64.415 94.105 66.215 94.165 ;
        RECT 65.885 94.075 66.215 94.105 ;
        RECT 64.015 93.325 64.275 94.005 ;
        RECT 64.445 93.155 64.695 93.935 ;
        RECT 64.945 93.905 65.780 93.915 ;
        RECT 66.370 93.905 66.555 93.995 ;
        RECT 64.945 93.705 66.555 93.905 ;
        RECT 64.945 93.325 65.195 93.705 ;
        RECT 66.325 93.665 66.555 93.705 ;
        RECT 66.805 93.545 67.060 94.165 ;
        RECT 65.365 93.155 65.720 93.535 ;
        RECT 66.725 93.325 67.060 93.545 ;
        RECT 67.700 94.105 68.035 95.525 ;
        RECT 68.215 95.335 68.960 95.705 ;
        RECT 69.525 95.165 69.780 95.525 ;
        RECT 69.960 95.335 70.290 95.705 ;
        RECT 70.470 95.165 70.695 95.525 ;
        RECT 68.210 94.975 70.695 95.165 ;
        RECT 68.210 94.285 68.435 94.975 ;
        RECT 70.915 94.935 72.585 95.705 ;
        RECT 72.770 95.135 73.025 95.485 ;
        RECT 73.195 95.305 73.525 95.705 ;
        RECT 73.695 95.135 73.865 95.485 ;
        RECT 74.035 95.305 74.415 95.705 ;
        RECT 72.770 94.965 74.435 95.135 ;
        RECT 74.605 95.030 74.880 95.375 ;
        RECT 75.220 95.195 75.460 95.705 ;
        RECT 75.640 95.195 75.920 95.525 ;
        RECT 76.150 95.195 76.365 95.705 ;
        RECT 68.635 94.465 68.915 94.795 ;
        RECT 69.095 94.465 69.670 94.795 ;
        RECT 69.850 94.465 70.285 94.795 ;
        RECT 70.465 94.465 70.735 94.795 ;
        RECT 70.915 94.415 71.665 94.935 ;
        RECT 74.265 94.795 74.435 94.965 ;
        RECT 68.210 94.105 70.705 94.285 ;
        RECT 71.835 94.245 72.585 94.765 ;
        RECT 72.755 94.465 73.100 94.795 ;
        RECT 73.270 94.465 74.095 94.795 ;
        RECT 74.265 94.465 74.540 94.795 ;
        RECT 67.700 93.335 67.965 94.105 ;
        RECT 68.135 93.155 68.465 93.875 ;
        RECT 68.655 93.695 69.845 93.925 ;
        RECT 68.655 93.335 68.915 93.695 ;
        RECT 69.085 93.155 69.415 93.525 ;
        RECT 69.585 93.335 69.845 93.695 ;
        RECT 70.415 93.335 70.705 94.105 ;
        RECT 70.915 93.155 72.585 94.245 ;
        RECT 72.775 94.005 73.100 94.295 ;
        RECT 73.270 94.175 73.465 94.465 ;
        RECT 74.265 94.295 74.435 94.465 ;
        RECT 74.710 94.295 74.880 95.030 ;
        RECT 75.115 94.465 75.470 95.025 ;
        RECT 75.640 94.295 75.810 95.195 ;
        RECT 75.980 94.465 76.245 95.025 ;
        RECT 76.535 94.965 77.150 95.535 ;
        RECT 76.495 94.295 76.665 94.795 ;
        RECT 73.775 94.125 74.435 94.295 ;
        RECT 73.775 94.005 73.945 94.125 ;
        RECT 72.775 93.835 73.945 94.005 ;
        RECT 72.755 93.375 73.945 93.665 ;
        RECT 74.115 93.155 74.395 93.955 ;
        RECT 74.605 93.325 74.880 94.295 ;
        RECT 75.240 94.125 76.665 94.295 ;
        RECT 75.240 93.950 75.630 94.125 ;
        RECT 76.115 93.155 76.445 93.955 ;
        RECT 76.835 93.945 77.150 94.965 ;
        RECT 78.280 94.940 78.735 95.705 ;
        RECT 79.010 95.325 80.310 95.535 ;
        RECT 80.565 95.345 80.895 95.705 ;
        RECT 80.140 95.175 80.310 95.325 ;
        RECT 81.065 95.205 81.325 95.535 ;
        RECT 81.095 95.195 81.325 95.205 ;
        RECT 79.210 94.715 79.430 95.115 ;
        RECT 78.275 94.515 78.765 94.715 ;
        RECT 78.955 94.505 79.430 94.715 ;
        RECT 79.675 94.715 79.885 95.115 ;
        RECT 80.140 95.050 80.895 95.175 ;
        RECT 80.140 95.005 80.985 95.050 ;
        RECT 80.715 94.885 80.985 95.005 ;
        RECT 79.675 94.505 80.005 94.715 ;
        RECT 80.175 94.445 80.585 94.750 ;
        RECT 76.615 93.325 77.150 93.945 ;
        RECT 78.280 94.275 79.455 94.335 ;
        RECT 80.815 94.310 80.985 94.885 ;
        RECT 80.785 94.275 80.985 94.310 ;
        RECT 78.280 94.165 80.985 94.275 ;
        RECT 78.280 93.545 78.535 94.165 ;
        RECT 79.125 94.105 80.925 94.165 ;
        RECT 79.125 94.075 79.455 94.105 ;
        RECT 81.155 94.005 81.325 95.195 ;
        RECT 81.495 95.160 86.840 95.705 ;
        RECT 83.080 94.330 83.420 95.160 ;
        RECT 87.015 94.935 88.685 95.705 ;
        RECT 89.315 94.955 90.525 95.705 ;
        RECT 78.785 93.905 78.970 93.995 ;
        RECT 79.560 93.905 80.395 93.915 ;
        RECT 78.785 93.705 80.395 93.905 ;
        RECT 78.785 93.665 79.015 93.705 ;
        RECT 78.280 93.325 78.615 93.545 ;
        RECT 79.620 93.155 79.975 93.535 ;
        RECT 80.145 93.325 80.395 93.705 ;
        RECT 80.645 93.155 80.895 93.935 ;
        RECT 81.065 93.325 81.325 94.005 ;
        RECT 84.900 93.590 85.250 94.840 ;
        RECT 87.015 94.415 87.765 94.935 ;
        RECT 87.935 94.245 88.685 94.765 ;
        RECT 81.495 93.155 86.840 93.590 ;
        RECT 87.015 93.155 88.685 94.245 ;
        RECT 89.315 94.245 89.835 94.785 ;
        RECT 90.005 94.415 90.525 94.955 ;
        RECT 89.315 93.155 90.525 94.245 ;
        RECT 11.950 92.985 90.610 93.155 ;
        RECT 99.980 93.085 100.150 100.195 ;
        RECT 100.550 93.815 100.720 99.855 ;
        RECT 100.990 93.815 101.160 99.855 ;
        RECT 100.690 93.430 101.020 93.600 ;
        RECT 101.560 93.085 101.730 100.195 ;
        RECT 102.130 93.815 102.300 99.855 ;
        RECT 102.570 93.815 102.740 99.855 ;
        RECT 102.270 93.430 102.600 93.600 ;
        RECT 103.140 93.085 103.310 100.195 ;
        RECT 103.710 93.815 103.880 99.855 ;
        RECT 104.150 93.815 104.320 99.855 ;
        RECT 103.850 93.430 104.180 93.600 ;
        RECT 104.720 93.085 104.890 100.195 ;
        RECT 105.290 93.815 105.460 99.855 ;
        RECT 105.730 93.815 105.900 99.855 ;
        RECT 105.430 93.430 105.760 93.600 ;
        RECT 106.300 93.085 106.470 100.195 ;
        RECT 106.870 93.815 107.040 99.855 ;
        RECT 107.310 93.815 107.480 99.855 ;
        RECT 107.010 93.430 107.340 93.600 ;
        RECT 107.880 93.085 108.050 100.195 ;
        RECT 108.450 93.815 108.620 99.855 ;
        RECT 108.890 93.815 109.060 99.855 ;
        RECT 108.590 93.430 108.920 93.600 ;
        RECT 109.460 93.085 109.630 100.195 ;
        RECT 110.030 93.815 110.200 99.855 ;
        RECT 110.470 93.815 110.640 99.855 ;
        RECT 110.170 93.430 110.500 93.600 ;
        RECT 111.040 93.085 111.210 100.195 ;
        RECT 111.610 93.815 111.780 99.855 ;
        RECT 112.050 93.815 112.220 99.855 ;
        RECT 111.750 93.430 112.080 93.600 ;
        RECT 112.620 93.085 112.790 100.195 ;
        RECT 134.450 96.750 134.620 101.720 ;
        RECT 135.100 99.930 135.450 102.090 ;
        RECT 135.100 97.230 135.450 99.390 ;
        RECT 135.930 96.750 136.100 102.570 ;
        RECT 136.580 99.930 136.930 102.090 ;
        RECT 136.580 97.230 136.930 99.390 ;
        RECT 137.410 96.750 137.580 102.570 ;
        RECT 138.060 99.930 138.410 102.090 ;
        RECT 138.060 97.230 138.410 99.390 ;
        RECT 138.890 96.750 139.060 102.570 ;
        RECT 139.540 99.930 139.890 102.090 ;
        RECT 139.540 97.230 139.890 99.390 ;
        RECT 140.370 96.750 140.540 102.570 ;
        RECT 141.020 99.930 141.370 102.090 ;
        RECT 141.020 97.230 141.370 99.390 ;
        RECT 141.850 96.750 142.020 102.570 ;
        RECT 142.500 99.930 142.850 102.090 ;
        RECT 142.500 97.230 142.850 99.390 ;
        RECT 143.330 96.750 143.500 102.570 ;
        RECT 143.980 99.930 144.330 102.090 ;
        RECT 143.980 97.230 144.330 99.390 ;
        RECT 144.810 96.750 144.980 102.570 ;
        RECT 145.460 99.930 145.810 102.090 ;
        RECT 145.460 97.230 145.810 99.390 ;
        RECT 146.290 96.750 146.460 102.570 ;
        RECT 146.940 99.930 147.290 102.090 ;
        RECT 146.940 97.230 147.290 99.390 ;
        RECT 147.770 96.750 147.940 102.570 ;
        RECT 148.420 99.930 148.770 102.090 ;
        RECT 148.420 97.230 148.770 99.390 ;
        RECT 149.250 96.750 149.420 102.570 ;
        RECT 149.900 99.930 150.250 102.090 ;
        RECT 149.900 97.230 150.250 99.390 ;
        RECT 150.730 96.750 150.900 102.570 ;
        RECT 151.380 99.930 151.730 102.090 ;
        RECT 151.380 97.230 151.730 99.390 ;
        RECT 152.210 96.750 152.380 102.570 ;
        RECT 152.860 99.930 153.210 102.090 ;
        RECT 152.860 97.230 153.210 99.390 ;
        RECT 153.690 96.750 153.860 102.570 ;
        RECT 154.340 99.930 154.690 102.090 ;
        RECT 154.340 97.230 154.690 99.390 ;
        RECT 155.170 96.750 155.340 102.570 ;
        RECT 155.820 99.930 156.170 102.090 ;
        RECT 155.820 97.230 156.170 99.390 ;
        RECT 156.650 96.750 156.820 102.570 ;
        RECT 157.300 99.930 157.650 102.090 ;
        RECT 157.300 97.230 157.650 99.390 ;
        RECT 158.130 96.750 158.300 102.570 ;
        RECT 134.450 96.580 158.300 96.750 ;
        RECT 12.035 91.895 13.245 92.985 ;
        RECT 13.505 92.315 13.675 92.815 ;
        RECT 13.845 92.485 14.175 92.985 ;
        RECT 13.505 92.145 14.170 92.315 ;
        RECT 12.035 91.185 12.555 91.725 ;
        RECT 12.725 91.355 13.245 91.895 ;
        RECT 13.420 91.325 13.770 91.975 ;
        RECT 12.035 90.435 13.245 91.185 ;
        RECT 13.940 91.155 14.170 92.145 ;
        RECT 13.505 90.985 14.170 91.155 ;
        RECT 13.505 90.695 13.675 90.985 ;
        RECT 13.845 90.435 14.175 90.815 ;
        RECT 14.345 90.695 14.530 92.815 ;
        RECT 14.770 92.525 15.035 92.985 ;
        RECT 15.205 92.390 15.455 92.815 ;
        RECT 15.665 92.540 16.770 92.710 ;
        RECT 15.150 92.260 15.455 92.390 ;
        RECT 14.700 91.065 14.980 92.015 ;
        RECT 15.150 91.155 15.320 92.260 ;
        RECT 15.490 91.475 15.730 92.070 ;
        RECT 15.900 92.005 16.430 92.370 ;
        RECT 15.900 91.305 16.070 92.005 ;
        RECT 16.600 91.925 16.770 92.540 ;
        RECT 16.940 92.185 17.110 92.985 ;
        RECT 17.280 92.485 17.530 92.815 ;
        RECT 17.755 92.515 18.640 92.685 ;
        RECT 16.600 91.835 17.110 91.925 ;
        RECT 15.150 91.025 15.375 91.155 ;
        RECT 15.545 91.085 16.070 91.305 ;
        RECT 16.240 91.665 17.110 91.835 ;
        RECT 14.785 90.435 15.035 90.895 ;
        RECT 15.205 90.885 15.375 91.025 ;
        RECT 16.240 90.885 16.410 91.665 ;
        RECT 16.940 91.595 17.110 91.665 ;
        RECT 16.620 91.415 16.820 91.445 ;
        RECT 17.280 91.415 17.450 92.485 ;
        RECT 17.620 91.595 17.810 92.315 ;
        RECT 16.620 91.115 17.450 91.415 ;
        RECT 17.980 91.385 18.300 92.345 ;
        RECT 15.205 90.715 15.540 90.885 ;
        RECT 15.735 90.715 16.410 90.885 ;
        RECT 16.730 90.435 17.100 90.935 ;
        RECT 17.280 90.885 17.450 91.115 ;
        RECT 17.835 91.055 18.300 91.385 ;
        RECT 18.470 91.675 18.640 92.515 ;
        RECT 18.820 92.485 19.135 92.985 ;
        RECT 19.365 92.255 19.705 92.815 ;
        RECT 18.810 91.880 19.705 92.255 ;
        RECT 19.875 91.975 20.045 92.985 ;
        RECT 19.515 91.675 19.705 91.880 ;
        RECT 20.215 91.925 20.545 92.770 ;
        RECT 20.715 92.070 20.885 92.985 ;
        RECT 22.155 92.430 22.760 92.985 ;
        RECT 22.935 92.475 23.415 92.815 ;
        RECT 23.585 92.440 23.840 92.985 ;
        RECT 22.155 92.330 22.770 92.430 ;
        RECT 22.585 92.305 22.770 92.330 ;
        RECT 20.215 91.845 20.605 91.925 ;
        RECT 20.390 91.795 20.605 91.845 ;
        RECT 18.470 91.345 19.345 91.675 ;
        RECT 19.515 91.345 20.265 91.675 ;
        RECT 18.470 90.885 18.640 91.345 ;
        RECT 19.515 91.175 19.715 91.345 ;
        RECT 20.435 91.215 20.605 91.795 ;
        RECT 22.155 91.710 22.415 92.160 ;
        RECT 22.585 92.060 22.915 92.305 ;
        RECT 23.085 91.985 23.840 92.235 ;
        RECT 24.010 92.115 24.285 92.815 ;
        RECT 23.070 91.950 23.840 91.985 ;
        RECT 23.055 91.940 23.840 91.950 ;
        RECT 23.050 91.925 23.945 91.940 ;
        RECT 23.030 91.910 23.945 91.925 ;
        RECT 23.010 91.900 23.945 91.910 ;
        RECT 22.985 91.890 23.945 91.900 ;
        RECT 22.915 91.860 23.945 91.890 ;
        RECT 22.895 91.830 23.945 91.860 ;
        RECT 22.875 91.800 23.945 91.830 ;
        RECT 22.845 91.775 23.945 91.800 ;
        RECT 22.810 91.740 23.945 91.775 ;
        RECT 22.780 91.735 23.945 91.740 ;
        RECT 22.780 91.730 23.170 91.735 ;
        RECT 22.780 91.720 23.145 91.730 ;
        RECT 22.780 91.715 23.130 91.720 ;
        RECT 22.780 91.710 23.115 91.715 ;
        RECT 22.155 91.705 23.115 91.710 ;
        RECT 22.155 91.695 23.105 91.705 ;
        RECT 22.155 91.690 23.095 91.695 ;
        RECT 22.155 91.680 23.085 91.690 ;
        RECT 22.155 91.670 23.080 91.680 ;
        RECT 22.155 91.665 23.075 91.670 ;
        RECT 22.155 91.650 23.065 91.665 ;
        RECT 22.155 91.635 23.060 91.650 ;
        RECT 22.155 91.610 23.050 91.635 ;
        RECT 22.155 91.540 23.045 91.610 ;
        RECT 20.380 91.175 20.605 91.215 ;
        RECT 17.280 90.715 17.685 90.885 ;
        RECT 17.855 90.715 18.640 90.885 ;
        RECT 18.915 90.435 19.125 90.965 ;
        RECT 19.385 90.650 19.715 91.175 ;
        RECT 20.225 91.090 20.605 91.175 ;
        RECT 19.885 90.435 20.055 91.045 ;
        RECT 20.225 90.655 20.555 91.090 ;
        RECT 22.155 90.985 22.705 91.370 ;
        RECT 20.725 90.435 20.895 90.950 ;
        RECT 22.875 90.815 23.045 91.540 ;
        RECT 22.155 90.645 23.045 90.815 ;
        RECT 23.215 91.140 23.545 91.565 ;
        RECT 23.715 91.340 23.945 91.735 ;
        RECT 23.215 90.655 23.435 91.140 ;
        RECT 24.115 91.085 24.285 92.115 ;
        RECT 24.915 91.820 25.205 92.985 ;
        RECT 25.840 91.845 26.175 92.815 ;
        RECT 26.345 91.845 26.515 92.985 ;
        RECT 26.685 92.645 28.715 92.815 ;
        RECT 25.840 91.175 26.010 91.845 ;
        RECT 26.685 91.675 26.855 92.645 ;
        RECT 26.180 91.345 26.435 91.675 ;
        RECT 26.660 91.345 26.855 91.675 ;
        RECT 27.025 92.305 28.150 92.475 ;
        RECT 26.265 91.175 26.435 91.345 ;
        RECT 27.025 91.175 27.195 92.305 ;
        RECT 23.605 90.435 23.855 90.975 ;
        RECT 24.025 90.605 24.285 91.085 ;
        RECT 24.915 90.435 25.205 91.160 ;
        RECT 25.840 90.605 26.095 91.175 ;
        RECT 26.265 91.005 27.195 91.175 ;
        RECT 27.365 91.965 28.375 92.135 ;
        RECT 27.365 91.165 27.535 91.965 ;
        RECT 27.740 91.285 28.015 91.765 ;
        RECT 27.735 91.115 28.015 91.285 ;
        RECT 27.020 90.970 27.195 91.005 ;
        RECT 26.265 90.435 26.595 90.835 ;
        RECT 27.020 90.605 27.550 90.970 ;
        RECT 27.740 90.605 28.015 91.115 ;
        RECT 28.185 90.605 28.375 91.965 ;
        RECT 28.545 91.980 28.715 92.645 ;
        RECT 28.885 92.225 29.055 92.985 ;
        RECT 29.290 92.225 29.805 92.635 ;
        RECT 29.975 92.550 35.320 92.985 ;
        RECT 28.545 91.790 29.295 91.980 ;
        RECT 29.465 91.415 29.805 92.225 ;
        RECT 28.575 91.245 29.805 91.415 ;
        RECT 28.555 90.435 29.065 90.970 ;
        RECT 29.285 90.640 29.530 91.245 ;
        RECT 31.560 90.980 31.900 91.810 ;
        RECT 33.380 91.300 33.730 92.550 ;
        RECT 35.495 91.895 39.005 92.985 ;
        RECT 39.290 92.355 39.575 92.815 ;
        RECT 39.745 92.525 40.015 92.985 ;
        RECT 39.290 92.135 40.245 92.355 ;
        RECT 35.495 91.205 37.145 91.725 ;
        RECT 37.315 91.375 39.005 91.895 ;
        RECT 39.175 91.405 39.865 91.965 ;
        RECT 40.035 91.235 40.245 92.135 ;
        RECT 29.975 90.435 35.320 90.980 ;
        RECT 35.495 90.435 39.005 91.205 ;
        RECT 39.290 91.065 40.245 91.235 ;
        RECT 40.415 91.965 40.815 92.815 ;
        RECT 41.005 92.355 41.285 92.815 ;
        RECT 41.805 92.525 42.130 92.985 ;
        RECT 41.005 92.135 42.130 92.355 ;
        RECT 40.415 91.405 41.510 91.965 ;
        RECT 41.680 91.675 42.130 92.135 ;
        RECT 42.300 91.845 42.685 92.815 ;
        RECT 42.855 91.895 44.525 92.985 ;
        RECT 45.155 91.910 45.495 92.985 ;
        RECT 45.680 92.475 47.730 92.765 ;
        RECT 39.290 90.605 39.575 91.065 ;
        RECT 39.745 90.435 40.015 90.895 ;
        RECT 40.415 90.605 40.815 91.405 ;
        RECT 41.680 91.345 42.235 91.675 ;
        RECT 41.680 91.235 42.130 91.345 ;
        RECT 41.005 91.065 42.130 91.235 ;
        RECT 42.405 91.175 42.685 91.845 ;
        RECT 41.005 90.605 41.285 91.065 ;
        RECT 41.805 90.435 42.130 90.895 ;
        RECT 42.300 90.605 42.685 91.175 ;
        RECT 42.855 91.205 43.605 91.725 ;
        RECT 43.775 91.375 44.525 91.895 ;
        RECT 45.665 91.675 45.905 92.270 ;
        RECT 46.100 92.135 47.730 92.305 ;
        RECT 47.900 92.185 48.180 92.985 ;
        RECT 46.100 91.845 46.420 92.135 ;
        RECT 47.560 92.015 47.730 92.135 ;
        RECT 42.855 90.435 44.525 91.205 ;
        RECT 45.155 91.105 45.495 91.675 ;
        RECT 45.665 91.345 46.320 91.675 ;
        RECT 46.590 91.345 47.330 91.965 ;
        RECT 47.560 91.845 48.220 92.015 ;
        RECT 48.390 91.845 48.665 92.815 ;
        RECT 48.835 91.895 50.505 92.985 ;
        RECT 48.050 91.675 48.220 91.845 ;
        RECT 47.500 91.345 47.880 91.675 ;
        RECT 48.050 91.345 48.325 91.675 ;
        RECT 45.155 90.435 45.495 90.935 ;
        RECT 45.665 90.655 45.910 91.345 ;
        RECT 48.050 91.175 48.220 91.345 ;
        RECT 46.635 91.005 48.220 91.175 ;
        RECT 48.495 91.110 48.665 91.845 ;
        RECT 46.105 90.435 46.435 90.935 ;
        RECT 46.635 90.655 46.805 91.005 ;
        RECT 46.980 90.435 47.310 90.835 ;
        RECT 47.480 90.655 47.650 91.005 ;
        RECT 47.820 90.435 48.200 90.835 ;
        RECT 48.390 90.765 48.665 91.110 ;
        RECT 48.835 91.205 49.585 91.725 ;
        RECT 49.755 91.375 50.505 91.895 ;
        RECT 50.675 91.820 50.965 92.985 ;
        RECT 51.135 92.550 56.480 92.985 ;
        RECT 56.655 92.550 62.000 92.985 ;
        RECT 48.835 90.435 50.505 91.205 ;
        RECT 50.675 90.435 50.965 91.160 ;
        RECT 52.720 90.980 53.060 91.810 ;
        RECT 54.540 91.300 54.890 92.550 ;
        RECT 58.240 90.980 58.580 91.810 ;
        RECT 60.060 91.300 60.410 92.550 ;
        RECT 62.175 91.895 65.685 92.985 ;
        RECT 65.960 92.185 66.215 92.985 ;
        RECT 66.385 92.015 66.715 92.815 ;
        RECT 66.885 92.185 67.055 92.985 ;
        RECT 67.225 92.015 67.555 92.815 ;
        RECT 62.175 91.205 63.825 91.725 ;
        RECT 63.995 91.375 65.685 91.895 ;
        RECT 65.855 91.845 67.555 92.015 ;
        RECT 67.725 91.845 67.985 92.985 ;
        RECT 68.155 91.895 69.825 92.985 ;
        RECT 69.995 92.430 70.600 92.985 ;
        RECT 70.775 92.475 71.255 92.815 ;
        RECT 71.425 92.440 71.680 92.985 ;
        RECT 69.995 92.330 70.610 92.430 ;
        RECT 70.425 92.305 70.610 92.330 ;
        RECT 65.855 91.255 66.135 91.845 ;
        RECT 66.305 91.425 67.055 91.675 ;
        RECT 67.225 91.425 67.985 91.675 ;
        RECT 51.135 90.435 56.480 90.980 ;
        RECT 56.655 90.435 62.000 90.980 ;
        RECT 62.175 90.435 65.685 91.205 ;
        RECT 65.855 91.005 66.715 91.255 ;
        RECT 66.885 91.065 67.985 91.235 ;
        RECT 65.965 90.815 66.295 90.835 ;
        RECT 66.885 90.815 67.135 91.065 ;
        RECT 65.965 90.605 67.135 90.815 ;
        RECT 67.305 90.435 67.475 90.895 ;
        RECT 67.645 90.605 67.985 91.065 ;
        RECT 68.155 91.205 68.905 91.725 ;
        RECT 69.075 91.375 69.825 91.895 ;
        RECT 69.995 91.710 70.255 92.160 ;
        RECT 70.425 92.060 70.755 92.305 ;
        RECT 70.925 91.985 71.680 92.235 ;
        RECT 71.850 92.115 72.125 92.815 ;
        RECT 70.910 91.950 71.680 91.985 ;
        RECT 70.895 91.940 71.680 91.950 ;
        RECT 70.890 91.925 71.785 91.940 ;
        RECT 70.870 91.910 71.785 91.925 ;
        RECT 70.850 91.900 71.785 91.910 ;
        RECT 70.825 91.890 71.785 91.900 ;
        RECT 70.755 91.860 71.785 91.890 ;
        RECT 70.735 91.830 71.785 91.860 ;
        RECT 70.715 91.800 71.785 91.830 ;
        RECT 70.685 91.775 71.785 91.800 ;
        RECT 70.650 91.740 71.785 91.775 ;
        RECT 70.620 91.735 71.785 91.740 ;
        RECT 70.620 91.730 71.010 91.735 ;
        RECT 70.620 91.720 70.985 91.730 ;
        RECT 70.620 91.715 70.970 91.720 ;
        RECT 70.620 91.710 70.955 91.715 ;
        RECT 69.995 91.705 70.955 91.710 ;
        RECT 69.995 91.695 70.945 91.705 ;
        RECT 69.995 91.690 70.935 91.695 ;
        RECT 69.995 91.680 70.925 91.690 ;
        RECT 69.995 91.670 70.920 91.680 ;
        RECT 69.995 91.665 70.915 91.670 ;
        RECT 69.995 91.650 70.905 91.665 ;
        RECT 69.995 91.635 70.900 91.650 ;
        RECT 69.995 91.610 70.890 91.635 ;
        RECT 69.995 91.540 70.885 91.610 ;
        RECT 68.155 90.435 69.825 91.205 ;
        RECT 69.995 90.985 70.545 91.370 ;
        RECT 70.715 90.815 70.885 91.540 ;
        RECT 69.995 90.645 70.885 90.815 ;
        RECT 71.055 91.140 71.385 91.565 ;
        RECT 71.555 91.340 71.785 91.735 ;
        RECT 71.055 90.655 71.275 91.140 ;
        RECT 71.955 91.085 72.125 92.115 ;
        RECT 72.295 91.895 75.805 92.985 ;
        RECT 71.445 90.435 71.695 90.975 ;
        RECT 71.865 90.605 72.125 91.085 ;
        RECT 72.295 91.205 73.945 91.725 ;
        RECT 74.115 91.375 75.805 91.895 ;
        RECT 76.435 91.820 76.725 92.985 ;
        RECT 76.900 92.015 77.175 92.815 ;
        RECT 77.345 92.185 77.675 92.985 ;
        RECT 77.845 92.645 78.985 92.815 ;
        RECT 77.845 92.015 78.015 92.645 ;
        RECT 76.900 91.805 78.015 92.015 ;
        RECT 78.185 92.015 78.515 92.475 ;
        RECT 78.685 92.185 78.985 92.645 ;
        RECT 78.185 91.965 78.945 92.015 ;
        RECT 78.185 91.795 78.965 91.965 ;
        RECT 79.255 91.845 79.465 92.985 ;
        RECT 79.635 91.835 79.965 92.815 ;
        RECT 80.135 91.845 80.365 92.985 ;
        RECT 80.575 91.895 84.085 92.985 ;
        RECT 84.255 91.895 85.465 92.985 ;
        RECT 76.900 91.425 77.620 91.625 ;
        RECT 77.790 91.425 78.560 91.625 ;
        RECT 78.730 91.255 78.945 91.795 ;
        RECT 72.295 90.435 75.805 91.205 ;
        RECT 76.435 90.435 76.725 91.160 ;
        RECT 76.900 90.435 77.175 91.255 ;
        RECT 77.345 91.085 78.945 91.255 ;
        RECT 77.345 91.075 78.515 91.085 ;
        RECT 77.345 90.605 77.675 91.075 ;
        RECT 77.845 90.435 78.015 90.905 ;
        RECT 78.185 90.605 78.515 91.075 ;
        RECT 78.685 90.435 78.975 90.905 ;
        RECT 79.255 90.435 79.465 91.255 ;
        RECT 79.635 91.235 79.885 91.835 ;
        RECT 80.055 91.425 80.385 91.675 ;
        RECT 79.635 90.605 79.965 91.235 ;
        RECT 80.135 90.435 80.365 91.255 ;
        RECT 80.575 91.205 82.225 91.725 ;
        RECT 82.395 91.375 84.085 91.895 ;
        RECT 80.575 90.435 84.085 91.205 ;
        RECT 84.255 91.185 84.775 91.725 ;
        RECT 84.945 91.355 85.465 91.895 ;
        RECT 85.635 91.845 86.020 92.815 ;
        RECT 86.190 92.525 86.515 92.985 ;
        RECT 87.035 92.355 87.315 92.815 ;
        RECT 86.190 92.135 87.315 92.355 ;
        RECT 84.255 90.435 85.465 91.185 ;
        RECT 85.635 91.175 85.915 91.845 ;
        RECT 86.190 91.675 86.640 92.135 ;
        RECT 87.505 91.965 87.905 92.815 ;
        RECT 88.305 92.525 88.575 92.985 ;
        RECT 88.745 92.355 89.030 92.815 ;
        RECT 86.085 91.345 86.640 91.675 ;
        RECT 86.810 91.405 87.905 91.965 ;
        RECT 86.190 91.235 86.640 91.345 ;
        RECT 85.635 90.605 86.020 91.175 ;
        RECT 86.190 91.065 87.315 91.235 ;
        RECT 86.190 90.435 86.515 90.895 ;
        RECT 87.035 90.605 87.315 91.065 ;
        RECT 87.505 90.605 87.905 91.405 ;
        RECT 88.075 92.135 89.030 92.355 ;
        RECT 88.075 91.235 88.285 92.135 ;
        RECT 88.455 91.405 89.145 91.965 ;
        RECT 89.315 91.895 90.525 92.985 ;
        RECT 99.980 92.915 112.790 93.085 ;
        RECT 117.630 93.120 130.430 93.230 ;
        RECT 117.630 92.430 130.440 93.120 ;
        RECT 117.590 92.260 130.440 92.430 ;
        RECT 89.315 91.355 89.835 91.895 ;
        RECT 88.075 91.065 89.030 91.235 ;
        RECT 90.005 91.185 90.525 91.725 ;
        RECT 88.305 90.435 88.575 90.895 ;
        RECT 88.745 90.605 89.030 91.065 ;
        RECT 89.315 90.435 90.525 91.185 ;
        RECT 99.990 91.675 112.800 91.845 ;
        RECT 11.950 90.265 90.610 90.435 ;
        RECT 12.035 89.515 13.245 90.265 ;
        RECT 12.035 88.975 12.555 89.515 ;
        RECT 13.415 89.495 15.085 90.265 ;
        RECT 15.720 89.590 15.995 89.935 ;
        RECT 16.185 89.865 16.565 90.265 ;
        RECT 16.735 89.695 16.905 90.045 ;
        RECT 17.075 89.865 17.405 90.265 ;
        RECT 17.575 89.695 17.830 90.045 ;
        RECT 12.725 88.805 13.245 89.345 ;
        RECT 13.415 88.975 14.165 89.495 ;
        RECT 14.335 88.805 15.085 89.325 ;
        RECT 12.035 87.715 13.245 88.805 ;
        RECT 13.415 87.715 15.085 88.805 ;
        RECT 15.720 88.855 15.890 89.590 ;
        RECT 16.165 89.525 17.830 89.695 ;
        RECT 18.105 89.715 18.275 90.005 ;
        RECT 18.445 89.885 18.775 90.265 ;
        RECT 18.105 89.545 18.770 89.715 ;
        RECT 16.165 89.355 16.335 89.525 ;
        RECT 16.060 89.025 16.335 89.355 ;
        RECT 16.505 89.025 17.330 89.355 ;
        RECT 17.500 89.025 17.845 89.355 ;
        RECT 16.165 88.855 16.335 89.025 ;
        RECT 15.720 87.885 15.995 88.855 ;
        RECT 16.165 88.685 16.825 88.855 ;
        RECT 17.135 88.735 17.330 89.025 ;
        RECT 16.655 88.565 16.825 88.685 ;
        RECT 17.500 88.565 17.825 88.855 ;
        RECT 18.020 88.725 18.370 89.375 ;
        RECT 16.205 87.715 16.485 88.515 ;
        RECT 16.655 88.395 17.825 88.565 ;
        RECT 18.540 88.555 18.770 89.545 ;
        RECT 18.105 88.385 18.770 88.555 ;
        RECT 16.655 87.935 17.845 88.225 ;
        RECT 18.105 87.885 18.275 88.385 ;
        RECT 18.445 87.715 18.775 88.215 ;
        RECT 18.945 87.885 19.130 90.005 ;
        RECT 19.385 89.805 19.635 90.265 ;
        RECT 19.805 89.815 20.140 89.985 ;
        RECT 20.335 89.815 21.010 89.985 ;
        RECT 19.805 89.675 19.975 89.815 ;
        RECT 19.300 88.685 19.580 89.635 ;
        RECT 19.750 89.545 19.975 89.675 ;
        RECT 19.750 88.440 19.920 89.545 ;
        RECT 20.145 89.395 20.670 89.615 ;
        RECT 20.090 88.630 20.330 89.225 ;
        RECT 20.500 88.695 20.670 89.395 ;
        RECT 20.840 89.035 21.010 89.815 ;
        RECT 21.330 89.765 21.700 90.265 ;
        RECT 21.880 89.815 22.285 89.985 ;
        RECT 22.455 89.815 23.240 89.985 ;
        RECT 21.880 89.585 22.050 89.815 ;
        RECT 21.220 89.285 22.050 89.585 ;
        RECT 22.435 89.315 22.900 89.645 ;
        RECT 21.220 89.255 21.420 89.285 ;
        RECT 21.540 89.035 21.710 89.105 ;
        RECT 20.840 88.865 21.710 89.035 ;
        RECT 21.200 88.775 21.710 88.865 ;
        RECT 19.750 88.310 20.055 88.440 ;
        RECT 20.500 88.330 21.030 88.695 ;
        RECT 19.370 87.715 19.635 88.175 ;
        RECT 19.805 87.885 20.055 88.310 ;
        RECT 21.200 88.160 21.370 88.775 ;
        RECT 20.265 87.990 21.370 88.160 ;
        RECT 21.540 87.715 21.710 88.515 ;
        RECT 21.880 88.215 22.050 89.285 ;
        RECT 22.220 88.385 22.410 89.105 ;
        RECT 22.580 88.355 22.900 89.315 ;
        RECT 23.070 89.355 23.240 89.815 ;
        RECT 23.515 89.735 23.725 90.265 ;
        RECT 23.985 89.525 24.315 90.050 ;
        RECT 24.485 89.655 24.655 90.265 ;
        RECT 24.825 89.610 25.155 90.045 ;
        RECT 25.375 89.885 26.265 90.055 ;
        RECT 24.825 89.525 25.205 89.610 ;
        RECT 24.115 89.355 24.315 89.525 ;
        RECT 24.980 89.485 25.205 89.525 ;
        RECT 23.070 89.025 23.945 89.355 ;
        RECT 24.115 89.025 24.865 89.355 ;
        RECT 21.880 87.885 22.130 88.215 ;
        RECT 23.070 88.185 23.240 89.025 ;
        RECT 24.115 88.820 24.305 89.025 ;
        RECT 25.035 88.905 25.205 89.485 ;
        RECT 25.375 89.330 25.925 89.715 ;
        RECT 26.095 89.160 26.265 89.885 ;
        RECT 24.990 88.855 25.205 88.905 ;
        RECT 23.410 88.445 24.305 88.820 ;
        RECT 24.815 88.775 25.205 88.855 ;
        RECT 25.375 89.090 26.265 89.160 ;
        RECT 26.435 89.560 26.655 90.045 ;
        RECT 26.825 89.725 27.075 90.265 ;
        RECT 27.245 89.615 27.505 90.095 ;
        RECT 26.435 89.135 26.765 89.560 ;
        RECT 25.375 89.065 26.270 89.090 ;
        RECT 25.375 89.050 26.280 89.065 ;
        RECT 25.375 89.035 26.285 89.050 ;
        RECT 25.375 89.030 26.295 89.035 ;
        RECT 25.375 89.020 26.300 89.030 ;
        RECT 25.375 89.010 26.305 89.020 ;
        RECT 25.375 89.005 26.315 89.010 ;
        RECT 25.375 88.995 26.325 89.005 ;
        RECT 25.375 88.990 26.335 88.995 ;
        RECT 22.355 88.015 23.240 88.185 ;
        RECT 23.420 87.715 23.735 88.215 ;
        RECT 23.965 87.885 24.305 88.445 ;
        RECT 24.475 87.715 24.645 88.725 ;
        RECT 24.815 87.930 25.145 88.775 ;
        RECT 25.375 88.540 25.635 88.990 ;
        RECT 26.000 88.985 26.335 88.990 ;
        RECT 26.000 88.980 26.350 88.985 ;
        RECT 26.000 88.970 26.365 88.980 ;
        RECT 26.000 88.965 26.390 88.970 ;
        RECT 26.935 88.965 27.165 89.360 ;
        RECT 26.000 88.960 27.165 88.965 ;
        RECT 26.030 88.925 27.165 88.960 ;
        RECT 26.065 88.900 27.165 88.925 ;
        RECT 26.095 88.870 27.165 88.900 ;
        RECT 26.115 88.840 27.165 88.870 ;
        RECT 26.135 88.810 27.165 88.840 ;
        RECT 26.205 88.800 27.165 88.810 ;
        RECT 26.230 88.790 27.165 88.800 ;
        RECT 26.250 88.775 27.165 88.790 ;
        RECT 26.270 88.760 27.165 88.775 ;
        RECT 26.275 88.750 27.060 88.760 ;
        RECT 26.290 88.715 27.060 88.750 ;
        RECT 25.805 88.395 26.135 88.640 ;
        RECT 26.305 88.465 27.060 88.715 ;
        RECT 27.335 88.585 27.505 89.615 ;
        RECT 27.675 89.495 30.265 90.265 ;
        RECT 30.525 89.715 30.695 90.005 ;
        RECT 30.865 89.885 31.195 90.265 ;
        RECT 30.525 89.545 31.190 89.715 ;
        RECT 27.675 88.975 28.885 89.495 ;
        RECT 29.055 88.805 30.265 89.325 ;
        RECT 25.805 88.370 25.990 88.395 ;
        RECT 25.375 88.270 25.990 88.370 ;
        RECT 25.375 87.715 25.980 88.270 ;
        RECT 26.155 87.885 26.635 88.225 ;
        RECT 26.805 87.715 27.060 88.260 ;
        RECT 27.230 87.885 27.505 88.585 ;
        RECT 27.675 87.715 30.265 88.805 ;
        RECT 30.440 88.725 30.790 89.375 ;
        RECT 30.960 88.555 31.190 89.545 ;
        RECT 30.525 88.385 31.190 88.555 ;
        RECT 30.525 87.885 30.695 88.385 ;
        RECT 30.865 87.715 31.195 88.215 ;
        RECT 31.365 87.885 31.550 90.005 ;
        RECT 31.805 89.805 32.055 90.265 ;
        RECT 32.225 89.815 32.560 89.985 ;
        RECT 32.755 89.815 33.430 89.985 ;
        RECT 32.225 89.675 32.395 89.815 ;
        RECT 31.720 88.685 32.000 89.635 ;
        RECT 32.170 89.545 32.395 89.675 ;
        RECT 32.170 88.440 32.340 89.545 ;
        RECT 32.565 89.395 33.090 89.615 ;
        RECT 32.510 88.630 32.750 89.225 ;
        RECT 32.920 88.695 33.090 89.395 ;
        RECT 33.260 89.035 33.430 89.815 ;
        RECT 33.750 89.765 34.120 90.265 ;
        RECT 34.300 89.815 34.705 89.985 ;
        RECT 34.875 89.815 35.660 89.985 ;
        RECT 34.300 89.585 34.470 89.815 ;
        RECT 33.640 89.285 34.470 89.585 ;
        RECT 34.855 89.315 35.320 89.645 ;
        RECT 33.640 89.255 33.840 89.285 ;
        RECT 33.960 89.035 34.130 89.105 ;
        RECT 33.260 88.865 34.130 89.035 ;
        RECT 33.620 88.775 34.130 88.865 ;
        RECT 32.170 88.310 32.475 88.440 ;
        RECT 32.920 88.330 33.450 88.695 ;
        RECT 31.790 87.715 32.055 88.175 ;
        RECT 32.225 87.885 32.475 88.310 ;
        RECT 33.620 88.160 33.790 88.775 ;
        RECT 32.685 87.990 33.790 88.160 ;
        RECT 33.960 87.715 34.130 88.515 ;
        RECT 34.300 88.215 34.470 89.285 ;
        RECT 34.640 88.385 34.830 89.105 ;
        RECT 35.000 88.355 35.320 89.315 ;
        RECT 35.490 89.355 35.660 89.815 ;
        RECT 35.935 89.735 36.145 90.265 ;
        RECT 36.405 89.525 36.735 90.050 ;
        RECT 36.905 89.655 37.075 90.265 ;
        RECT 37.245 89.610 37.575 90.045 ;
        RECT 37.245 89.525 37.625 89.610 ;
        RECT 37.795 89.540 38.085 90.265 ;
        RECT 36.535 89.355 36.735 89.525 ;
        RECT 37.400 89.485 37.625 89.525 ;
        RECT 35.490 89.025 36.365 89.355 ;
        RECT 36.535 89.025 37.285 89.355 ;
        RECT 34.300 87.885 34.550 88.215 ;
        RECT 35.490 88.185 35.660 89.025 ;
        RECT 36.535 88.820 36.725 89.025 ;
        RECT 37.455 88.905 37.625 89.485 ;
        RECT 37.410 88.855 37.625 88.905 ;
        RECT 38.260 89.525 38.515 90.095 ;
        RECT 38.685 89.865 39.015 90.265 ;
        RECT 39.440 89.730 39.970 90.095 ;
        RECT 40.160 89.925 40.435 90.095 ;
        RECT 40.155 89.755 40.435 89.925 ;
        RECT 39.440 89.695 39.615 89.730 ;
        RECT 38.685 89.525 39.615 89.695 ;
        RECT 35.830 88.445 36.725 88.820 ;
        RECT 37.235 88.775 37.625 88.855 ;
        RECT 34.775 88.015 35.660 88.185 ;
        RECT 35.840 87.715 36.155 88.215 ;
        RECT 36.385 87.885 36.725 88.445 ;
        RECT 36.895 87.715 37.065 88.725 ;
        RECT 37.235 87.930 37.565 88.775 ;
        RECT 37.795 87.715 38.085 88.880 ;
        RECT 38.260 88.855 38.430 89.525 ;
        RECT 38.685 89.355 38.855 89.525 ;
        RECT 38.600 89.025 38.855 89.355 ;
        RECT 39.080 89.025 39.275 89.355 ;
        RECT 38.260 87.885 38.595 88.855 ;
        RECT 38.765 87.715 38.935 88.855 ;
        RECT 39.105 88.055 39.275 89.025 ;
        RECT 39.445 88.395 39.615 89.525 ;
        RECT 39.785 88.735 39.955 89.535 ;
        RECT 40.160 88.935 40.435 89.755 ;
        RECT 40.605 88.735 40.795 90.095 ;
        RECT 40.975 89.730 41.485 90.265 ;
        RECT 41.705 89.455 41.950 90.060 ;
        RECT 42.395 89.495 44.065 90.265 ;
        RECT 40.995 89.285 42.225 89.455 ;
        RECT 39.785 88.565 40.795 88.735 ;
        RECT 40.965 88.720 41.715 88.910 ;
        RECT 39.445 88.225 40.570 88.395 ;
        RECT 40.965 88.055 41.135 88.720 ;
        RECT 41.885 88.475 42.225 89.285 ;
        RECT 42.395 88.975 43.145 89.495 ;
        RECT 44.235 89.465 44.575 90.095 ;
        RECT 44.745 89.465 44.995 90.265 ;
        RECT 45.185 89.615 45.515 90.095 ;
        RECT 45.685 89.805 45.910 90.265 ;
        RECT 46.080 89.615 46.410 90.095 ;
        RECT 43.315 88.805 44.065 89.325 ;
        RECT 39.105 87.885 41.135 88.055 ;
        RECT 41.305 87.715 41.475 88.475 ;
        RECT 41.710 88.065 42.225 88.475 ;
        RECT 42.395 87.715 44.065 88.805 ;
        RECT 44.235 88.855 44.410 89.465 ;
        RECT 45.185 89.445 46.410 89.615 ;
        RECT 47.040 89.485 47.540 90.095 ;
        RECT 47.915 89.615 48.175 90.095 ;
        RECT 48.345 89.805 48.675 90.265 ;
        RECT 48.865 89.625 49.065 90.045 ;
        RECT 44.580 89.105 45.275 89.275 ;
        RECT 45.105 88.855 45.275 89.105 ;
        RECT 45.450 89.075 45.870 89.275 ;
        RECT 46.040 89.075 46.370 89.275 ;
        RECT 46.540 89.075 46.870 89.275 ;
        RECT 47.040 88.855 47.210 89.485 ;
        RECT 47.395 89.025 47.745 89.275 ;
        RECT 44.235 87.885 44.575 88.855 ;
        RECT 44.745 87.715 44.915 88.855 ;
        RECT 45.105 88.685 47.540 88.855 ;
        RECT 45.185 87.715 45.435 88.515 ;
        RECT 46.080 87.885 46.410 88.685 ;
        RECT 46.710 87.715 47.040 88.515 ;
        RECT 47.210 87.885 47.540 88.685 ;
        RECT 47.915 88.585 48.085 89.615 ;
        RECT 48.255 88.925 48.485 89.355 ;
        RECT 48.655 89.105 49.065 89.625 ;
        RECT 49.235 89.780 50.025 90.045 ;
        RECT 49.235 88.925 49.490 89.780 ;
        RECT 50.205 89.445 50.535 89.865 ;
        RECT 50.705 89.445 50.965 90.265 ;
        RECT 51.155 89.575 51.395 90.095 ;
        RECT 51.565 89.770 51.960 90.265 ;
        RECT 52.525 89.935 52.695 90.080 ;
        RECT 52.320 89.740 52.695 89.935 ;
        RECT 50.205 89.355 50.455 89.445 ;
        RECT 49.660 89.105 50.455 89.355 ;
        RECT 48.255 88.755 50.045 88.925 ;
        RECT 47.915 87.885 48.190 88.585 ;
        RECT 48.360 88.460 49.075 88.755 ;
        RECT 49.295 88.395 49.625 88.585 ;
        RECT 48.400 87.715 48.615 88.260 ;
        RECT 48.785 87.885 49.260 88.225 ;
        RECT 49.430 88.220 49.625 88.395 ;
        RECT 49.795 88.390 50.045 88.755 ;
        RECT 49.430 87.715 50.045 88.220 ;
        RECT 50.285 87.885 50.455 89.105 ;
        RECT 50.625 88.395 50.965 89.275 ;
        RECT 51.155 88.770 51.330 89.575 ;
        RECT 52.320 89.405 52.490 89.740 ;
        RECT 52.975 89.695 53.215 90.070 ;
        RECT 53.385 89.760 53.720 90.265 ;
        RECT 52.975 89.545 53.195 89.695 ;
        RECT 51.505 89.045 52.490 89.405 ;
        RECT 52.660 89.215 53.195 89.545 ;
        RECT 51.505 89.025 52.790 89.045 ;
        RECT 51.930 88.875 52.790 89.025 ;
        RECT 50.705 87.715 50.965 88.225 ;
        RECT 51.155 87.985 51.460 88.770 ;
        RECT 51.635 88.395 52.330 88.705 ;
        RECT 51.640 87.715 52.325 88.185 ;
        RECT 52.505 87.930 52.790 88.875 ;
        RECT 52.960 88.565 53.195 89.215 ;
        RECT 53.365 88.735 53.665 89.585 ;
        RECT 53.895 89.495 55.565 90.265 ;
        RECT 55.825 89.715 55.995 90.005 ;
        RECT 56.165 89.885 56.495 90.265 ;
        RECT 55.825 89.545 56.490 89.715 ;
        RECT 53.895 88.975 54.645 89.495 ;
        RECT 54.815 88.805 55.565 89.325 ;
        RECT 52.960 88.335 53.635 88.565 ;
        RECT 52.965 87.715 53.295 88.165 ;
        RECT 53.465 87.905 53.635 88.335 ;
        RECT 53.895 87.715 55.565 88.805 ;
        RECT 55.740 88.725 56.090 89.375 ;
        RECT 56.260 88.555 56.490 89.545 ;
        RECT 55.825 88.385 56.490 88.555 ;
        RECT 55.825 87.885 55.995 88.385 ;
        RECT 56.165 87.715 56.495 88.215 ;
        RECT 56.665 87.885 56.850 90.005 ;
        RECT 57.105 89.805 57.355 90.265 ;
        RECT 57.525 89.815 57.860 89.985 ;
        RECT 58.055 89.815 58.730 89.985 ;
        RECT 57.525 89.675 57.695 89.815 ;
        RECT 57.020 88.685 57.300 89.635 ;
        RECT 57.470 89.545 57.695 89.675 ;
        RECT 57.470 88.440 57.640 89.545 ;
        RECT 57.865 89.395 58.390 89.615 ;
        RECT 57.810 88.630 58.050 89.225 ;
        RECT 58.220 88.695 58.390 89.395 ;
        RECT 58.560 89.035 58.730 89.815 ;
        RECT 59.050 89.765 59.420 90.265 ;
        RECT 59.600 89.815 60.005 89.985 ;
        RECT 60.175 89.815 60.960 89.985 ;
        RECT 59.600 89.585 59.770 89.815 ;
        RECT 58.940 89.285 59.770 89.585 ;
        RECT 60.155 89.315 60.620 89.645 ;
        RECT 58.940 89.255 59.140 89.285 ;
        RECT 59.260 89.035 59.430 89.105 ;
        RECT 58.560 88.865 59.430 89.035 ;
        RECT 58.920 88.775 59.430 88.865 ;
        RECT 57.470 88.310 57.775 88.440 ;
        RECT 58.220 88.330 58.750 88.695 ;
        RECT 57.090 87.715 57.355 88.175 ;
        RECT 57.525 87.885 57.775 88.310 ;
        RECT 58.920 88.160 59.090 88.775 ;
        RECT 57.985 87.990 59.090 88.160 ;
        RECT 59.260 87.715 59.430 88.515 ;
        RECT 59.600 88.215 59.770 89.285 ;
        RECT 59.940 88.385 60.130 89.105 ;
        RECT 60.300 88.355 60.620 89.315 ;
        RECT 60.790 89.355 60.960 89.815 ;
        RECT 61.235 89.735 61.445 90.265 ;
        RECT 61.705 89.525 62.035 90.050 ;
        RECT 62.205 89.655 62.375 90.265 ;
        RECT 62.545 89.610 62.875 90.045 ;
        RECT 62.545 89.525 62.925 89.610 ;
        RECT 63.555 89.540 63.845 90.265 ;
        RECT 64.020 89.790 64.355 90.050 ;
        RECT 64.525 89.865 64.855 90.265 ;
        RECT 65.025 89.865 66.640 90.035 ;
        RECT 61.835 89.355 62.035 89.525 ;
        RECT 62.700 89.485 62.925 89.525 ;
        RECT 60.790 89.025 61.665 89.355 ;
        RECT 61.835 89.025 62.585 89.355 ;
        RECT 59.600 87.885 59.850 88.215 ;
        RECT 60.790 88.185 60.960 89.025 ;
        RECT 61.835 88.820 62.025 89.025 ;
        RECT 62.755 88.905 62.925 89.485 ;
        RECT 62.710 88.855 62.925 88.905 ;
        RECT 61.130 88.445 62.025 88.820 ;
        RECT 62.535 88.775 62.925 88.855 ;
        RECT 60.075 88.015 60.960 88.185 ;
        RECT 61.140 87.715 61.455 88.215 ;
        RECT 61.685 87.885 62.025 88.445 ;
        RECT 62.195 87.715 62.365 88.725 ;
        RECT 62.535 87.930 62.865 88.775 ;
        RECT 63.555 87.715 63.845 88.880 ;
        RECT 64.020 88.435 64.275 89.790 ;
        RECT 65.025 89.695 65.195 89.865 ;
        RECT 64.635 89.525 65.195 89.695 ;
        RECT 64.635 89.355 64.805 89.525 ;
        RECT 64.500 89.025 64.805 89.355 ;
        RECT 65.000 89.245 65.250 89.355 ;
        RECT 65.460 89.245 65.730 89.685 ;
        RECT 65.920 89.585 66.210 89.685 ;
        RECT 65.915 89.415 66.210 89.585 ;
        RECT 64.995 89.075 65.250 89.245 ;
        RECT 65.455 89.075 65.730 89.245 ;
        RECT 65.000 89.025 65.250 89.075 ;
        RECT 65.460 89.025 65.730 89.075 ;
        RECT 65.920 89.025 66.210 89.415 ;
        RECT 66.380 89.025 66.800 89.690 ;
        RECT 67.185 89.545 67.515 90.265 ;
        RECT 68.620 89.760 68.955 90.265 ;
        RECT 69.125 89.695 69.365 90.070 ;
        RECT 69.645 89.935 69.815 90.080 ;
        RECT 69.645 89.740 70.020 89.935 ;
        RECT 70.380 89.770 70.775 90.265 ;
        RECT 67.110 89.245 67.460 89.355 ;
        RECT 67.110 89.075 67.465 89.245 ;
        RECT 67.110 89.025 67.460 89.075 ;
        RECT 64.635 88.855 64.805 89.025 ;
        RECT 64.635 88.685 67.005 88.855 ;
        RECT 67.255 88.735 67.460 89.025 ;
        RECT 68.675 88.735 68.975 89.585 ;
        RECT 69.145 89.545 69.365 89.695 ;
        RECT 69.145 89.215 69.680 89.545 ;
        RECT 69.850 89.405 70.020 89.740 ;
        RECT 70.945 89.575 71.185 90.095 ;
        RECT 64.020 87.925 64.355 88.435 ;
        RECT 64.605 87.715 64.935 88.515 ;
        RECT 65.180 88.305 66.605 88.475 ;
        RECT 65.180 87.885 65.465 88.305 ;
        RECT 65.720 87.715 66.050 88.135 ;
        RECT 66.275 88.055 66.605 88.305 ;
        RECT 66.835 88.225 67.005 88.685 ;
        RECT 69.145 88.565 69.380 89.215 ;
        RECT 69.850 89.045 70.835 89.405 ;
        RECT 67.265 88.055 67.435 88.555 ;
        RECT 66.275 87.885 67.435 88.055 ;
        RECT 68.705 88.335 69.380 88.565 ;
        RECT 69.550 89.025 70.835 89.045 ;
        RECT 69.550 88.875 70.410 89.025 ;
        RECT 68.705 87.905 68.875 88.335 ;
        RECT 69.045 87.715 69.375 88.165 ;
        RECT 69.550 87.930 69.835 88.875 ;
        RECT 71.010 88.770 71.185 89.575 ;
        RECT 71.380 89.735 71.670 90.085 ;
        RECT 71.865 89.905 72.195 90.265 ;
        RECT 72.365 89.735 72.595 90.040 ;
        RECT 71.380 89.565 72.595 89.735 ;
        RECT 72.785 89.925 72.955 89.960 ;
        RECT 72.785 89.755 72.985 89.925 ;
        RECT 72.785 89.395 72.955 89.755 ;
        RECT 71.440 89.245 71.700 89.355 ;
        RECT 71.435 89.075 71.700 89.245 ;
        RECT 71.440 89.025 71.700 89.075 ;
        RECT 71.880 89.025 72.265 89.355 ;
        RECT 72.435 89.225 72.955 89.395 ;
        RECT 73.215 89.495 75.805 90.265 ;
        RECT 76.440 89.500 76.895 90.265 ;
        RECT 77.170 89.885 78.470 90.095 ;
        RECT 78.725 89.905 79.055 90.265 ;
        RECT 78.300 89.735 78.470 89.885 ;
        RECT 79.225 89.765 79.485 90.095 ;
        RECT 70.010 88.395 70.705 88.705 ;
        RECT 70.015 87.715 70.700 88.185 ;
        RECT 70.880 87.985 71.185 88.770 ;
        RECT 71.380 87.715 71.700 88.855 ;
        RECT 71.880 87.975 72.075 89.025 ;
        RECT 72.435 88.845 72.605 89.225 ;
        RECT 72.255 88.565 72.605 88.845 ;
        RECT 72.795 88.695 73.040 89.055 ;
        RECT 73.215 88.975 74.425 89.495 ;
        RECT 74.595 88.805 75.805 89.325 ;
        RECT 77.370 89.275 77.590 89.675 ;
        RECT 76.435 89.075 76.925 89.275 ;
        RECT 77.115 89.065 77.590 89.275 ;
        RECT 77.835 89.275 78.045 89.675 ;
        RECT 78.300 89.610 79.055 89.735 ;
        RECT 78.300 89.565 79.145 89.610 ;
        RECT 78.875 89.445 79.145 89.565 ;
        RECT 77.835 89.065 78.165 89.275 ;
        RECT 78.335 89.005 78.745 89.310 ;
        RECT 72.255 87.885 72.585 88.565 ;
        RECT 72.785 87.715 73.040 88.515 ;
        RECT 73.215 87.715 75.805 88.805 ;
        RECT 76.440 88.835 77.615 88.895 ;
        RECT 78.975 88.870 79.145 89.445 ;
        RECT 78.945 88.835 79.145 88.870 ;
        RECT 76.440 88.725 79.145 88.835 ;
        RECT 76.440 88.105 76.695 88.725 ;
        RECT 77.285 88.665 79.085 88.725 ;
        RECT 77.285 88.635 77.615 88.665 ;
        RECT 79.315 88.565 79.485 89.765 ;
        RECT 80.205 89.715 80.375 90.005 ;
        RECT 80.545 89.885 80.875 90.265 ;
        RECT 80.205 89.545 80.870 89.715 ;
        RECT 80.120 88.725 80.470 89.375 ;
        RECT 76.945 88.465 77.130 88.555 ;
        RECT 77.720 88.465 78.555 88.475 ;
        RECT 76.945 88.265 78.555 88.465 ;
        RECT 76.945 88.225 77.175 88.265 ;
        RECT 76.440 87.885 76.775 88.105 ;
        RECT 77.780 87.715 78.135 88.095 ;
        RECT 78.305 87.885 78.555 88.265 ;
        RECT 78.805 87.715 79.055 88.495 ;
        RECT 79.225 87.885 79.485 88.565 ;
        RECT 80.640 88.555 80.870 89.545 ;
        RECT 80.205 88.385 80.870 88.555 ;
        RECT 80.205 87.885 80.375 88.385 ;
        RECT 80.545 87.715 80.875 88.215 ;
        RECT 81.045 87.885 81.230 90.005 ;
        RECT 81.485 89.805 81.735 90.265 ;
        RECT 81.905 89.815 82.240 89.985 ;
        RECT 82.435 89.815 83.110 89.985 ;
        RECT 81.905 89.675 82.075 89.815 ;
        RECT 81.400 88.685 81.680 89.635 ;
        RECT 81.850 89.545 82.075 89.675 ;
        RECT 81.850 88.440 82.020 89.545 ;
        RECT 82.245 89.395 82.770 89.615 ;
        RECT 82.190 88.630 82.430 89.225 ;
        RECT 82.600 88.695 82.770 89.395 ;
        RECT 82.940 89.035 83.110 89.815 ;
        RECT 83.430 89.765 83.800 90.265 ;
        RECT 83.980 89.815 84.385 89.985 ;
        RECT 84.555 89.815 85.340 89.985 ;
        RECT 83.980 89.585 84.150 89.815 ;
        RECT 83.320 89.285 84.150 89.585 ;
        RECT 84.535 89.315 85.000 89.645 ;
        RECT 83.320 89.255 83.520 89.285 ;
        RECT 83.640 89.035 83.810 89.105 ;
        RECT 82.940 88.865 83.810 89.035 ;
        RECT 83.300 88.775 83.810 88.865 ;
        RECT 81.850 88.310 82.155 88.440 ;
        RECT 82.600 88.330 83.130 88.695 ;
        RECT 81.470 87.715 81.735 88.175 ;
        RECT 81.905 87.885 82.155 88.310 ;
        RECT 83.300 88.160 83.470 88.775 ;
        RECT 82.365 87.990 83.470 88.160 ;
        RECT 83.640 87.715 83.810 88.515 ;
        RECT 83.980 88.215 84.150 89.285 ;
        RECT 84.320 88.385 84.510 89.105 ;
        RECT 84.680 88.355 85.000 89.315 ;
        RECT 85.170 89.355 85.340 89.815 ;
        RECT 85.615 89.735 85.825 90.265 ;
        RECT 86.085 89.525 86.415 90.050 ;
        RECT 86.585 89.655 86.755 90.265 ;
        RECT 86.925 89.610 87.255 90.045 ;
        RECT 87.565 89.715 87.735 90.095 ;
        RECT 87.950 89.885 88.280 90.265 ;
        RECT 86.925 89.525 87.305 89.610 ;
        RECT 87.565 89.545 88.280 89.715 ;
        RECT 86.215 89.355 86.415 89.525 ;
        RECT 87.080 89.485 87.305 89.525 ;
        RECT 85.170 89.025 86.045 89.355 ;
        RECT 86.215 89.025 86.965 89.355 ;
        RECT 83.980 87.885 84.230 88.215 ;
        RECT 85.170 88.185 85.340 89.025 ;
        RECT 86.215 88.820 86.405 89.025 ;
        RECT 87.135 88.905 87.305 89.485 ;
        RECT 87.475 88.995 87.830 89.365 ;
        RECT 88.110 89.355 88.280 89.545 ;
        RECT 88.450 89.520 88.705 90.095 ;
        RECT 88.110 89.025 88.365 89.355 ;
        RECT 87.090 88.855 87.305 88.905 ;
        RECT 85.510 88.445 86.405 88.820 ;
        RECT 86.915 88.775 87.305 88.855 ;
        RECT 88.110 88.815 88.280 89.025 ;
        RECT 84.455 88.015 85.340 88.185 ;
        RECT 85.520 87.715 85.835 88.215 ;
        RECT 86.065 87.885 86.405 88.445 ;
        RECT 86.575 87.715 86.745 88.725 ;
        RECT 86.915 87.930 87.245 88.775 ;
        RECT 87.565 88.645 88.280 88.815 ;
        RECT 88.535 88.790 88.705 89.520 ;
        RECT 88.880 89.425 89.140 90.265 ;
        RECT 89.315 89.515 90.525 90.265 ;
        RECT 87.565 87.885 87.735 88.645 ;
        RECT 87.950 87.715 88.280 88.475 ;
        RECT 88.450 87.885 88.705 88.790 ;
        RECT 88.880 87.715 89.140 88.865 ;
        RECT 89.315 88.805 89.835 89.345 ;
        RECT 90.005 88.975 90.525 89.515 ;
        RECT 89.315 87.715 90.525 88.805 ;
        RECT 99.990 88.605 100.160 91.675 ;
        RECT 100.700 91.165 101.030 91.335 ;
        RECT 100.560 88.955 100.730 90.995 ;
        RECT 101.000 88.955 101.170 90.995 ;
        RECT 101.570 88.605 101.740 91.675 ;
        RECT 102.280 91.165 102.610 91.335 ;
        RECT 102.140 88.955 102.310 90.995 ;
        RECT 102.580 88.955 102.750 90.995 ;
        RECT 103.150 88.605 103.320 91.675 ;
        RECT 103.860 91.165 104.190 91.335 ;
        RECT 103.720 88.955 103.890 90.995 ;
        RECT 104.160 88.955 104.330 90.995 ;
        RECT 104.730 88.605 104.900 91.675 ;
        RECT 105.440 91.165 105.770 91.335 ;
        RECT 105.300 88.955 105.470 90.995 ;
        RECT 105.740 88.955 105.910 90.995 ;
        RECT 106.310 88.605 106.480 91.675 ;
        RECT 107.020 91.165 107.350 91.335 ;
        RECT 106.880 88.955 107.050 90.995 ;
        RECT 107.320 88.955 107.490 90.995 ;
        RECT 107.890 88.605 108.060 91.675 ;
        RECT 108.600 91.165 108.930 91.335 ;
        RECT 108.460 88.955 108.630 90.995 ;
        RECT 108.900 88.955 109.070 90.995 ;
        RECT 109.470 88.605 109.640 91.675 ;
        RECT 110.180 91.165 110.510 91.335 ;
        RECT 110.040 88.955 110.210 90.995 ;
        RECT 110.480 88.955 110.650 90.995 ;
        RECT 111.050 88.605 111.220 91.675 ;
        RECT 111.760 91.165 112.090 91.335 ;
        RECT 111.620 88.955 111.790 90.995 ;
        RECT 112.060 88.955 112.230 90.995 ;
        RECT 112.630 88.605 112.800 91.675 ;
        RECT 99.990 88.415 112.800 88.605 ;
        RECT 100.070 87.785 112.760 88.415 ;
        RECT 11.950 87.545 90.610 87.715 ;
        RECT 99.990 87.615 113.480 87.785 ;
        RECT 12.035 86.455 13.245 87.545 ;
        RECT 13.415 86.455 16.925 87.545 ;
        RECT 17.095 86.455 18.305 87.545 ;
        RECT 12.035 85.745 12.555 86.285 ;
        RECT 12.725 85.915 13.245 86.455 ;
        RECT 13.415 85.765 15.065 86.285 ;
        RECT 15.235 85.935 16.925 86.455 ;
        RECT 12.035 84.995 13.245 85.745 ;
        RECT 13.415 84.995 16.925 85.765 ;
        RECT 17.095 85.745 17.615 86.285 ;
        RECT 17.785 85.915 18.305 86.455 ;
        RECT 18.660 86.575 19.050 86.750 ;
        RECT 19.535 86.745 19.865 87.545 ;
        RECT 20.035 86.755 20.570 87.375 ;
        RECT 18.660 86.405 20.085 86.575 ;
        RECT 17.095 84.995 18.305 85.745 ;
        RECT 18.535 85.675 18.890 86.235 ;
        RECT 19.060 85.505 19.230 86.405 ;
        RECT 19.400 85.675 19.665 86.235 ;
        RECT 19.915 85.905 20.085 86.405 ;
        RECT 20.255 85.735 20.570 86.755 ;
        RECT 18.640 84.995 18.880 85.505 ;
        RECT 19.060 85.175 19.340 85.505 ;
        RECT 19.570 84.995 19.785 85.505 ;
        RECT 19.955 85.165 20.570 85.735 ;
        RECT 20.775 86.825 21.235 87.375 ;
        RECT 21.425 86.825 21.755 87.545 ;
        RECT 20.775 85.455 21.025 86.825 ;
        RECT 21.955 86.655 22.255 87.205 ;
        RECT 22.425 86.875 22.705 87.545 ;
        RECT 21.315 86.485 22.255 86.655 ;
        RECT 21.315 86.235 21.485 86.485 ;
        RECT 22.625 86.235 22.890 86.595 ;
        RECT 23.575 86.405 23.805 87.545 ;
        RECT 23.975 86.395 24.305 87.375 ;
        RECT 24.475 86.405 24.685 87.545 ;
        RECT 21.195 85.905 21.485 86.235 ;
        RECT 21.655 85.985 21.995 86.235 ;
        RECT 22.215 85.985 22.890 86.235 ;
        RECT 23.555 85.985 23.885 86.235 ;
        RECT 21.315 85.815 21.485 85.905 ;
        RECT 21.315 85.625 22.705 85.815 ;
        RECT 20.775 85.165 21.335 85.455 ;
        RECT 21.505 84.995 21.755 85.455 ;
        RECT 22.375 85.265 22.705 85.625 ;
        RECT 23.575 84.995 23.805 85.815 ;
        RECT 24.055 85.795 24.305 86.395 ;
        RECT 24.915 86.380 25.205 87.545 ;
        RECT 26.385 86.875 26.555 87.375 ;
        RECT 26.725 87.045 27.055 87.545 ;
        RECT 26.385 86.705 27.050 86.875 ;
        RECT 26.300 85.885 26.650 86.535 ;
        RECT 23.975 85.165 24.305 85.795 ;
        RECT 24.475 84.995 24.685 85.815 ;
        RECT 24.915 84.995 25.205 85.720 ;
        RECT 26.820 85.715 27.050 86.705 ;
        RECT 26.385 85.545 27.050 85.715 ;
        RECT 26.385 85.255 26.555 85.545 ;
        RECT 26.725 84.995 27.055 85.375 ;
        RECT 27.225 85.255 27.410 87.375 ;
        RECT 27.650 87.085 27.915 87.545 ;
        RECT 28.085 86.950 28.335 87.375 ;
        RECT 28.545 87.100 29.650 87.270 ;
        RECT 28.030 86.820 28.335 86.950 ;
        RECT 27.580 85.625 27.860 86.575 ;
        RECT 28.030 85.715 28.200 86.820 ;
        RECT 28.370 86.035 28.610 86.630 ;
        RECT 28.780 86.565 29.310 86.930 ;
        RECT 28.780 85.865 28.950 86.565 ;
        RECT 29.480 86.485 29.650 87.100 ;
        RECT 29.820 86.745 29.990 87.545 ;
        RECT 30.160 87.045 30.410 87.375 ;
        RECT 30.635 87.075 31.520 87.245 ;
        RECT 29.480 86.395 29.990 86.485 ;
        RECT 28.030 85.585 28.255 85.715 ;
        RECT 28.425 85.645 28.950 85.865 ;
        RECT 29.120 86.225 29.990 86.395 ;
        RECT 27.665 84.995 27.915 85.455 ;
        RECT 28.085 85.445 28.255 85.585 ;
        RECT 29.120 85.445 29.290 86.225 ;
        RECT 29.820 86.155 29.990 86.225 ;
        RECT 29.500 85.975 29.700 86.005 ;
        RECT 30.160 85.975 30.330 87.045 ;
        RECT 30.500 86.155 30.690 86.875 ;
        RECT 29.500 85.675 30.330 85.975 ;
        RECT 30.860 85.945 31.180 86.905 ;
        RECT 28.085 85.275 28.420 85.445 ;
        RECT 28.615 85.275 29.290 85.445 ;
        RECT 29.610 84.995 29.980 85.495 ;
        RECT 30.160 85.445 30.330 85.675 ;
        RECT 30.715 85.615 31.180 85.945 ;
        RECT 31.350 86.235 31.520 87.075 ;
        RECT 31.700 87.045 32.015 87.545 ;
        RECT 32.245 86.815 32.585 87.375 ;
        RECT 31.690 86.440 32.585 86.815 ;
        RECT 32.755 86.535 32.925 87.545 ;
        RECT 32.395 86.235 32.585 86.440 ;
        RECT 33.095 86.485 33.425 87.330 ;
        RECT 33.595 86.630 33.765 87.545 ;
        RECT 33.095 86.405 33.485 86.485 ;
        RECT 34.115 86.455 37.625 87.545 ;
        RECT 33.270 86.355 33.485 86.405 ;
        RECT 31.350 85.905 32.225 86.235 ;
        RECT 32.395 85.905 33.145 86.235 ;
        RECT 31.350 85.445 31.520 85.905 ;
        RECT 32.395 85.735 32.595 85.905 ;
        RECT 33.315 85.775 33.485 86.355 ;
        RECT 33.260 85.735 33.485 85.775 ;
        RECT 30.160 85.275 30.565 85.445 ;
        RECT 30.735 85.275 31.520 85.445 ;
        RECT 31.795 84.995 32.005 85.525 ;
        RECT 32.265 85.210 32.595 85.735 ;
        RECT 33.105 85.650 33.485 85.735 ;
        RECT 34.115 85.765 35.765 86.285 ;
        RECT 35.935 85.935 37.625 86.455 ;
        RECT 38.715 86.405 39.100 87.375 ;
        RECT 39.270 87.085 39.595 87.545 ;
        RECT 40.115 86.915 40.395 87.375 ;
        RECT 39.270 86.695 40.395 86.915 ;
        RECT 32.765 84.995 32.935 85.605 ;
        RECT 33.105 85.215 33.435 85.650 ;
        RECT 33.605 84.995 33.775 85.510 ;
        RECT 34.115 84.995 37.625 85.765 ;
        RECT 38.715 85.735 38.995 86.405 ;
        RECT 39.270 86.235 39.720 86.695 ;
        RECT 40.585 86.525 40.985 87.375 ;
        RECT 41.385 87.085 41.655 87.545 ;
        RECT 41.825 86.915 42.110 87.375 ;
        RECT 42.395 87.035 42.655 87.545 ;
        RECT 39.165 85.905 39.720 86.235 ;
        RECT 39.890 85.965 40.985 86.525 ;
        RECT 39.270 85.795 39.720 85.905 ;
        RECT 38.715 85.165 39.100 85.735 ;
        RECT 39.270 85.625 40.395 85.795 ;
        RECT 39.270 84.995 39.595 85.455 ;
        RECT 40.115 85.165 40.395 85.625 ;
        RECT 40.585 85.165 40.985 85.965 ;
        RECT 41.155 86.695 42.110 86.915 ;
        RECT 41.155 85.795 41.365 86.695 ;
        RECT 41.535 85.965 42.225 86.525 ;
        RECT 42.395 85.985 42.735 86.865 ;
        RECT 42.905 86.155 43.075 87.375 ;
        RECT 43.315 87.040 43.930 87.545 ;
        RECT 43.315 86.505 43.565 86.870 ;
        RECT 43.735 86.865 43.930 87.040 ;
        RECT 44.100 87.035 44.575 87.375 ;
        RECT 44.745 87.000 44.960 87.545 ;
        RECT 43.735 86.675 44.065 86.865 ;
        RECT 44.285 86.505 45.000 86.800 ;
        RECT 45.170 86.675 45.445 87.375 ;
        RECT 43.315 86.335 45.105 86.505 ;
        RECT 42.905 85.905 43.700 86.155 ;
        RECT 42.905 85.815 43.155 85.905 ;
        RECT 41.155 85.625 42.110 85.795 ;
        RECT 41.385 84.995 41.655 85.455 ;
        RECT 41.825 85.165 42.110 85.625 ;
        RECT 42.395 84.995 42.655 85.815 ;
        RECT 42.825 85.395 43.155 85.815 ;
        RECT 43.870 85.480 44.125 86.335 ;
        RECT 43.335 85.215 44.125 85.480 ;
        RECT 44.295 85.635 44.705 86.155 ;
        RECT 44.875 85.905 45.105 86.335 ;
        RECT 45.275 85.645 45.445 86.675 ;
        RECT 44.295 85.215 44.495 85.635 ;
        RECT 44.685 84.995 45.015 85.455 ;
        RECT 45.185 85.165 45.445 85.645 ;
        RECT 46.555 86.490 46.860 87.275 ;
        RECT 47.040 87.075 47.725 87.545 ;
        RECT 47.035 86.555 47.730 86.865 ;
        RECT 46.555 85.685 46.730 86.490 ;
        RECT 47.905 86.385 48.190 87.330 ;
        RECT 48.365 87.095 48.695 87.545 ;
        RECT 48.865 86.925 49.035 87.355 ;
        RECT 47.330 86.235 48.190 86.385 ;
        RECT 46.905 86.215 48.190 86.235 ;
        RECT 48.360 86.695 49.035 86.925 ;
        RECT 46.905 85.855 47.890 86.215 ;
        RECT 48.360 86.045 48.595 86.695 ;
        RECT 46.555 85.165 46.795 85.685 ;
        RECT 47.720 85.520 47.890 85.855 ;
        RECT 48.060 85.715 48.595 86.045 ;
        RECT 48.375 85.565 48.595 85.715 ;
        RECT 48.765 85.675 49.065 86.525 ;
        RECT 49.295 86.455 50.505 87.545 ;
        RECT 49.295 85.745 49.815 86.285 ;
        RECT 49.985 85.915 50.505 86.455 ;
        RECT 50.675 86.380 50.965 87.545 ;
        RECT 51.140 86.405 51.475 87.375 ;
        RECT 51.645 86.405 51.815 87.545 ;
        RECT 51.985 87.205 54.015 87.375 ;
        RECT 46.965 84.995 47.360 85.490 ;
        RECT 47.720 85.325 48.095 85.520 ;
        RECT 47.925 85.180 48.095 85.325 ;
        RECT 48.375 85.190 48.615 85.565 ;
        RECT 48.785 84.995 49.120 85.500 ;
        RECT 49.295 84.995 50.505 85.745 ;
        RECT 51.140 85.735 51.310 86.405 ;
        RECT 51.985 86.235 52.155 87.205 ;
        RECT 51.480 85.905 51.735 86.235 ;
        RECT 51.960 85.905 52.155 86.235 ;
        RECT 52.325 86.865 53.450 87.035 ;
        RECT 51.565 85.735 51.735 85.905 ;
        RECT 52.325 85.735 52.495 86.865 ;
        RECT 50.675 84.995 50.965 85.720 ;
        RECT 51.140 85.165 51.395 85.735 ;
        RECT 51.565 85.565 52.495 85.735 ;
        RECT 52.665 86.525 53.675 86.695 ;
        RECT 52.665 85.725 52.835 86.525 ;
        RECT 52.320 85.530 52.495 85.565 ;
        RECT 51.565 84.995 51.895 85.395 ;
        RECT 52.320 85.165 52.850 85.530 ;
        RECT 53.040 85.505 53.315 86.325 ;
        RECT 53.035 85.335 53.315 85.505 ;
        RECT 53.040 85.165 53.315 85.335 ;
        RECT 53.485 85.165 53.675 86.525 ;
        RECT 53.845 86.540 54.015 87.205 ;
        RECT 54.185 86.785 54.355 87.545 ;
        RECT 54.590 86.785 55.105 87.195 ;
        RECT 53.845 86.350 54.595 86.540 ;
        RECT 54.765 85.975 55.105 86.785 ;
        RECT 55.825 86.875 55.995 87.375 ;
        RECT 56.165 87.045 56.495 87.545 ;
        RECT 55.825 86.705 56.490 86.875 ;
        RECT 53.875 85.805 55.105 85.975 ;
        RECT 55.740 85.885 56.090 86.535 ;
        RECT 53.855 84.995 54.365 85.530 ;
        RECT 54.585 85.200 54.830 85.805 ;
        RECT 56.260 85.715 56.490 86.705 ;
        RECT 55.825 85.545 56.490 85.715 ;
        RECT 55.825 85.255 55.995 85.545 ;
        RECT 56.165 84.995 56.495 85.375 ;
        RECT 56.665 85.255 56.850 87.375 ;
        RECT 57.090 87.085 57.355 87.545 ;
        RECT 57.525 86.950 57.775 87.375 ;
        RECT 57.985 87.100 59.090 87.270 ;
        RECT 57.470 86.820 57.775 86.950 ;
        RECT 57.020 85.625 57.300 86.575 ;
        RECT 57.470 85.715 57.640 86.820 ;
        RECT 57.810 86.035 58.050 86.630 ;
        RECT 58.220 86.565 58.750 86.930 ;
        RECT 58.220 85.865 58.390 86.565 ;
        RECT 58.920 86.485 59.090 87.100 ;
        RECT 59.260 86.745 59.430 87.545 ;
        RECT 59.600 87.045 59.850 87.375 ;
        RECT 60.075 87.075 60.960 87.245 ;
        RECT 58.920 86.395 59.430 86.485 ;
        RECT 57.470 85.585 57.695 85.715 ;
        RECT 57.865 85.645 58.390 85.865 ;
        RECT 58.560 86.225 59.430 86.395 ;
        RECT 57.105 84.995 57.355 85.455 ;
        RECT 57.525 85.445 57.695 85.585 ;
        RECT 58.560 85.445 58.730 86.225 ;
        RECT 59.260 86.155 59.430 86.225 ;
        RECT 58.940 85.975 59.140 86.005 ;
        RECT 59.600 85.975 59.770 87.045 ;
        RECT 59.940 86.155 60.130 86.875 ;
        RECT 58.940 85.675 59.770 85.975 ;
        RECT 60.300 85.945 60.620 86.905 ;
        RECT 57.525 85.275 57.860 85.445 ;
        RECT 58.055 85.275 58.730 85.445 ;
        RECT 59.050 84.995 59.420 85.495 ;
        RECT 59.600 85.445 59.770 85.675 ;
        RECT 60.155 85.615 60.620 85.945 ;
        RECT 60.790 86.235 60.960 87.075 ;
        RECT 61.140 87.045 61.455 87.545 ;
        RECT 61.685 86.815 62.025 87.375 ;
        RECT 61.130 86.440 62.025 86.815 ;
        RECT 62.195 86.535 62.365 87.545 ;
        RECT 61.835 86.235 62.025 86.440 ;
        RECT 62.535 86.485 62.865 87.330 ;
        RECT 63.100 86.595 63.365 87.365 ;
        RECT 63.535 86.825 63.865 87.545 ;
        RECT 64.055 87.005 64.315 87.365 ;
        RECT 64.485 87.175 64.815 87.545 ;
        RECT 64.985 87.005 65.245 87.365 ;
        RECT 64.055 86.775 65.245 87.005 ;
        RECT 65.815 86.595 66.105 87.365 ;
        RECT 62.535 86.405 62.925 86.485 ;
        RECT 62.710 86.355 62.925 86.405 ;
        RECT 60.790 85.905 61.665 86.235 ;
        RECT 61.835 85.905 62.585 86.235 ;
        RECT 60.790 85.445 60.960 85.905 ;
        RECT 61.835 85.735 62.035 85.905 ;
        RECT 62.755 85.775 62.925 86.355 ;
        RECT 62.700 85.735 62.925 85.775 ;
        RECT 59.600 85.275 60.005 85.445 ;
        RECT 60.175 85.275 60.960 85.445 ;
        RECT 61.235 84.995 61.445 85.525 ;
        RECT 61.705 85.210 62.035 85.735 ;
        RECT 62.545 85.650 62.925 85.735 ;
        RECT 62.205 84.995 62.375 85.605 ;
        RECT 62.545 85.215 62.875 85.650 ;
        RECT 63.100 85.175 63.435 86.595 ;
        RECT 63.610 86.415 66.105 86.595 ;
        RECT 66.350 86.755 66.885 87.375 ;
        RECT 63.610 85.725 63.835 86.415 ;
        RECT 64.035 85.905 64.315 86.235 ;
        RECT 64.495 85.905 65.070 86.235 ;
        RECT 65.250 85.905 65.685 86.235 ;
        RECT 65.865 85.905 66.135 86.235 ;
        RECT 66.350 85.735 66.665 86.755 ;
        RECT 67.055 86.745 67.385 87.545 ;
        RECT 67.870 86.575 68.260 86.750 ;
        RECT 66.835 86.405 68.260 86.575 ;
        RECT 68.615 86.405 68.875 87.545 ;
        RECT 66.835 85.905 67.005 86.405 ;
        RECT 63.610 85.535 66.095 85.725 ;
        RECT 63.615 84.995 64.360 85.365 ;
        RECT 64.925 85.175 65.180 85.535 ;
        RECT 65.360 84.995 65.690 85.365 ;
        RECT 65.870 85.175 66.095 85.535 ;
        RECT 66.350 85.165 66.965 85.735 ;
        RECT 67.255 85.675 67.520 86.235 ;
        RECT 67.690 85.505 67.860 86.405 ;
        RECT 69.045 86.395 69.375 87.375 ;
        RECT 69.545 86.405 69.825 87.545 ;
        RECT 69.995 86.455 71.205 87.545 ;
        RECT 68.030 85.675 68.385 86.235 ;
        RECT 68.635 85.985 68.970 86.235 ;
        RECT 69.140 85.795 69.310 86.395 ;
        RECT 69.480 85.965 69.815 86.235 ;
        RECT 67.135 84.995 67.350 85.505 ;
        RECT 67.580 85.175 67.860 85.505 ;
        RECT 68.040 84.995 68.280 85.505 ;
        RECT 68.615 85.165 69.310 85.795 ;
        RECT 69.515 84.995 69.825 85.795 ;
        RECT 69.995 85.745 70.515 86.285 ;
        RECT 70.685 85.915 71.205 86.455 ;
        RECT 71.380 86.405 71.700 87.545 ;
        RECT 71.880 86.235 72.075 87.285 ;
        RECT 72.255 86.695 72.585 87.375 ;
        RECT 72.785 86.745 73.040 87.545 ;
        RECT 72.255 86.415 72.605 86.695 ;
        RECT 74.320 86.575 74.710 86.750 ;
        RECT 75.195 86.745 75.525 87.545 ;
        RECT 75.695 86.755 76.230 87.375 ;
        RECT 71.440 86.185 71.700 86.235 ;
        RECT 71.435 86.015 71.700 86.185 ;
        RECT 71.440 85.905 71.700 86.015 ;
        RECT 71.880 85.905 72.265 86.235 ;
        RECT 72.435 86.035 72.605 86.415 ;
        RECT 72.795 86.205 73.040 86.565 ;
        RECT 74.320 86.405 75.745 86.575 ;
        RECT 72.435 85.865 72.955 86.035 ;
        RECT 69.995 84.995 71.205 85.745 ;
        RECT 71.380 85.525 72.595 85.695 ;
        RECT 71.380 85.175 71.670 85.525 ;
        RECT 71.865 84.995 72.195 85.355 ;
        RECT 72.365 85.220 72.595 85.525 ;
        RECT 72.785 85.505 72.955 85.865 ;
        RECT 74.195 85.675 74.550 86.235 ;
        RECT 74.720 85.505 74.890 86.405 ;
        RECT 75.060 85.675 75.325 86.235 ;
        RECT 75.575 85.905 75.745 86.405 ;
        RECT 75.915 85.735 76.230 86.755 ;
        RECT 76.435 86.380 76.725 87.545 ;
        RECT 77.050 86.535 77.350 87.375 ;
        RECT 77.545 86.705 77.795 87.545 ;
        RECT 78.385 86.955 79.190 87.375 ;
        RECT 77.965 86.785 79.530 86.955 ;
        RECT 77.965 86.535 78.135 86.785 ;
        RECT 77.050 86.365 78.135 86.535 ;
        RECT 76.895 85.905 77.225 86.195 ;
        RECT 77.395 85.735 77.565 86.365 ;
        RECT 78.305 86.235 78.625 86.615 ;
        RECT 78.815 86.525 79.190 86.615 ;
        RECT 78.795 86.355 79.190 86.525 ;
        RECT 79.360 86.535 79.530 86.785 ;
        RECT 79.700 86.705 80.030 87.545 ;
        RECT 80.200 86.785 80.865 87.375 ;
        RECT 79.360 86.365 80.280 86.535 ;
        RECT 77.735 85.985 78.065 86.195 ;
        RECT 78.245 85.985 78.625 86.235 ;
        RECT 78.815 86.195 79.190 86.355 ;
        RECT 80.110 86.195 80.280 86.365 ;
        RECT 78.815 85.985 79.300 86.195 ;
        RECT 79.490 85.985 79.940 86.195 ;
        RECT 80.110 85.985 80.445 86.195 ;
        RECT 80.615 85.815 80.865 86.785 ;
        RECT 72.785 85.335 72.985 85.505 ;
        RECT 72.785 85.300 72.955 85.335 ;
        RECT 74.300 84.995 74.540 85.505 ;
        RECT 74.720 85.175 75.000 85.505 ;
        RECT 75.230 84.995 75.445 85.505 ;
        RECT 75.615 85.165 76.230 85.735 ;
        RECT 76.435 84.995 76.725 85.720 ;
        RECT 77.055 85.555 77.565 85.735 ;
        RECT 77.970 85.645 79.670 85.815 ;
        RECT 77.970 85.555 78.355 85.645 ;
        RECT 77.055 85.165 77.385 85.555 ;
        RECT 77.555 85.215 78.740 85.385 ;
        RECT 79.000 84.995 79.170 85.465 ;
        RECT 79.340 85.180 79.670 85.645 ;
        RECT 79.840 84.995 80.010 85.815 ;
        RECT 80.180 85.175 80.865 85.815 ;
        RECT 81.960 86.405 82.295 87.375 ;
        RECT 82.465 86.405 82.635 87.545 ;
        RECT 82.805 87.205 84.835 87.375 ;
        RECT 81.960 85.735 82.130 86.405 ;
        RECT 82.805 86.235 82.975 87.205 ;
        RECT 82.300 85.905 82.555 86.235 ;
        RECT 82.780 85.905 82.975 86.235 ;
        RECT 83.145 86.865 84.270 87.035 ;
        RECT 82.385 85.735 82.555 85.905 ;
        RECT 83.145 85.735 83.315 86.865 ;
        RECT 81.960 85.165 82.215 85.735 ;
        RECT 82.385 85.565 83.315 85.735 ;
        RECT 83.485 86.525 84.495 86.695 ;
        RECT 83.485 85.725 83.655 86.525 ;
        RECT 83.860 86.185 84.135 86.325 ;
        RECT 83.855 86.015 84.135 86.185 ;
        RECT 83.140 85.530 83.315 85.565 ;
        RECT 82.385 84.995 82.715 85.395 ;
        RECT 83.140 85.165 83.670 85.530 ;
        RECT 83.860 85.165 84.135 86.015 ;
        RECT 84.305 85.165 84.495 86.525 ;
        RECT 84.665 86.540 84.835 87.205 ;
        RECT 85.005 86.785 85.175 87.545 ;
        RECT 85.410 86.785 85.925 87.195 ;
        RECT 84.665 86.350 85.415 86.540 ;
        RECT 85.585 85.975 85.925 86.785 ;
        RECT 86.185 86.615 86.355 87.375 ;
        RECT 86.535 86.785 86.865 87.545 ;
        RECT 86.185 86.445 86.850 86.615 ;
        RECT 87.035 86.470 87.305 87.375 ;
        RECT 86.680 86.300 86.850 86.445 ;
        RECT 84.695 85.805 85.925 85.975 ;
        RECT 86.115 85.895 86.445 86.265 ;
        RECT 86.680 85.970 86.965 86.300 ;
        RECT 84.675 84.995 85.185 85.530 ;
        RECT 85.405 85.200 85.650 85.805 ;
        RECT 86.680 85.715 86.850 85.970 ;
        RECT 86.185 85.545 86.850 85.715 ;
        RECT 87.135 85.670 87.305 86.470 ;
        RECT 87.475 86.455 89.145 87.545 ;
        RECT 86.185 85.165 86.355 85.545 ;
        RECT 86.535 84.995 86.865 85.375 ;
        RECT 87.045 85.165 87.305 85.670 ;
        RECT 87.475 85.765 88.225 86.285 ;
        RECT 88.395 85.935 89.145 86.455 ;
        RECT 89.315 86.455 90.525 87.545 ;
        RECT 89.315 85.915 89.835 86.455 ;
        RECT 87.475 84.995 89.145 85.765 ;
        RECT 90.005 85.745 90.525 86.285 ;
        RECT 89.315 84.995 90.525 85.745 ;
        RECT 11.950 84.825 90.610 84.995 ;
        RECT 12.035 84.075 13.245 84.825 ;
        RECT 13.415 84.280 18.760 84.825 ;
        RECT 18.935 84.280 24.280 84.825 ;
        RECT 12.035 83.535 12.555 84.075 ;
        RECT 12.725 83.365 13.245 83.905 ;
        RECT 15.000 83.450 15.340 84.280 ;
        RECT 12.035 82.275 13.245 83.365 ;
        RECT 16.820 82.710 17.170 83.960 ;
        RECT 20.520 83.450 20.860 84.280 ;
        RECT 24.455 84.055 26.125 84.825 ;
        RECT 26.760 84.085 27.015 84.655 ;
        RECT 27.185 84.425 27.515 84.825 ;
        RECT 27.940 84.290 28.470 84.655 ;
        RECT 27.940 84.255 28.115 84.290 ;
        RECT 27.185 84.085 28.115 84.255 ;
        RECT 22.340 82.710 22.690 83.960 ;
        RECT 24.455 83.535 25.205 84.055 ;
        RECT 25.375 83.365 26.125 83.885 ;
        RECT 13.415 82.275 18.760 82.710 ;
        RECT 18.935 82.275 24.280 82.710 ;
        RECT 24.455 82.275 26.125 83.365 ;
        RECT 26.760 83.415 26.930 84.085 ;
        RECT 27.185 83.915 27.355 84.085 ;
        RECT 27.100 83.585 27.355 83.915 ;
        RECT 27.580 83.585 27.775 83.915 ;
        RECT 26.760 82.445 27.095 83.415 ;
        RECT 27.265 82.275 27.435 83.415 ;
        RECT 27.605 82.615 27.775 83.585 ;
        RECT 27.945 82.955 28.115 84.085 ;
        RECT 28.285 83.295 28.455 84.095 ;
        RECT 28.660 83.805 28.935 84.655 ;
        RECT 28.655 83.635 28.935 83.805 ;
        RECT 28.660 83.495 28.935 83.635 ;
        RECT 29.105 83.295 29.295 84.655 ;
        RECT 29.475 84.290 29.985 84.825 ;
        RECT 30.205 84.015 30.450 84.620 ;
        RECT 30.895 84.280 36.240 84.825 ;
        RECT 29.495 83.845 30.725 84.015 ;
        RECT 28.285 83.125 29.295 83.295 ;
        RECT 29.465 83.280 30.215 83.470 ;
        RECT 27.945 82.785 29.070 82.955 ;
        RECT 29.465 82.615 29.635 83.280 ;
        RECT 30.385 83.035 30.725 83.845 ;
        RECT 32.480 83.450 32.820 84.280 ;
        RECT 36.415 84.075 37.625 84.825 ;
        RECT 37.795 84.100 38.085 84.825 ;
        RECT 38.345 84.275 38.515 84.565 ;
        RECT 38.685 84.445 39.015 84.825 ;
        RECT 38.345 84.105 39.010 84.275 ;
        RECT 27.605 82.445 29.635 82.615 ;
        RECT 29.805 82.275 29.975 83.035 ;
        RECT 30.210 82.625 30.725 83.035 ;
        RECT 34.300 82.710 34.650 83.960 ;
        RECT 36.415 83.535 36.935 84.075 ;
        RECT 37.105 83.365 37.625 83.905 ;
        RECT 30.895 82.275 36.240 82.710 ;
        RECT 36.415 82.275 37.625 83.365 ;
        RECT 37.795 82.275 38.085 83.440 ;
        RECT 38.260 83.285 38.610 83.935 ;
        RECT 38.780 83.115 39.010 84.105 ;
        RECT 38.345 82.945 39.010 83.115 ;
        RECT 38.345 82.445 38.515 82.945 ;
        RECT 38.685 82.275 39.015 82.775 ;
        RECT 39.185 82.445 39.370 84.565 ;
        RECT 39.625 84.365 39.875 84.825 ;
        RECT 40.045 84.375 40.380 84.545 ;
        RECT 40.575 84.375 41.250 84.545 ;
        RECT 40.045 84.235 40.215 84.375 ;
        RECT 39.540 83.245 39.820 84.195 ;
        RECT 39.990 84.105 40.215 84.235 ;
        RECT 39.990 83.000 40.160 84.105 ;
        RECT 40.385 83.955 40.910 84.175 ;
        RECT 40.330 83.190 40.570 83.785 ;
        RECT 40.740 83.255 40.910 83.955 ;
        RECT 41.080 83.595 41.250 84.375 ;
        RECT 41.570 84.325 41.940 84.825 ;
        RECT 42.120 84.375 42.525 84.545 ;
        RECT 42.695 84.375 43.480 84.545 ;
        RECT 42.120 84.145 42.290 84.375 ;
        RECT 41.460 83.845 42.290 84.145 ;
        RECT 42.675 83.875 43.140 84.205 ;
        RECT 41.460 83.815 41.660 83.845 ;
        RECT 41.780 83.595 41.950 83.665 ;
        RECT 41.080 83.425 41.950 83.595 ;
        RECT 41.440 83.335 41.950 83.425 ;
        RECT 39.990 82.870 40.295 83.000 ;
        RECT 40.740 82.890 41.270 83.255 ;
        RECT 39.610 82.275 39.875 82.735 ;
        RECT 40.045 82.445 40.295 82.870 ;
        RECT 41.440 82.720 41.610 83.335 ;
        RECT 40.505 82.550 41.610 82.720 ;
        RECT 41.780 82.275 41.950 83.075 ;
        RECT 42.120 82.775 42.290 83.845 ;
        RECT 42.460 82.945 42.650 83.665 ;
        RECT 42.820 82.915 43.140 83.875 ;
        RECT 43.310 83.915 43.480 84.375 ;
        RECT 43.755 84.295 43.965 84.825 ;
        RECT 44.225 84.085 44.555 84.610 ;
        RECT 44.725 84.215 44.895 84.825 ;
        RECT 45.065 84.170 45.395 84.605 ;
        RECT 45.065 84.085 45.445 84.170 ;
        RECT 44.355 83.915 44.555 84.085 ;
        RECT 45.220 84.045 45.445 84.085 ;
        RECT 43.310 83.585 44.185 83.915 ;
        RECT 44.355 83.585 45.105 83.915 ;
        RECT 42.120 82.445 42.370 82.775 ;
        RECT 43.310 82.745 43.480 83.585 ;
        RECT 44.355 83.380 44.545 83.585 ;
        RECT 45.275 83.465 45.445 84.045 ;
        RECT 45.230 83.415 45.445 83.465 ;
        RECT 43.650 83.005 44.545 83.380 ;
        RECT 45.055 83.335 45.445 83.415 ;
        RECT 45.615 84.150 45.885 84.495 ;
        RECT 46.075 84.425 46.455 84.825 ;
        RECT 46.625 84.255 46.795 84.605 ;
        RECT 46.965 84.425 47.295 84.825 ;
        RECT 47.495 84.255 47.665 84.605 ;
        RECT 47.865 84.325 48.195 84.825 ;
        RECT 45.615 83.415 45.785 84.150 ;
        RECT 46.055 84.085 47.665 84.255 ;
        RECT 48.925 84.275 49.095 84.565 ;
        RECT 49.265 84.445 49.595 84.825 ;
        RECT 46.055 83.915 46.225 84.085 ;
        RECT 45.955 83.585 46.225 83.915 ;
        RECT 46.395 83.585 46.800 83.915 ;
        RECT 46.055 83.415 46.225 83.585 ;
        RECT 42.595 82.575 43.480 82.745 ;
        RECT 43.660 82.275 43.975 82.775 ;
        RECT 44.205 82.445 44.545 83.005 ;
        RECT 44.715 82.275 44.885 83.285 ;
        RECT 45.055 82.490 45.385 83.335 ;
        RECT 45.615 82.445 45.885 83.415 ;
        RECT 46.055 83.245 46.780 83.415 ;
        RECT 46.970 83.295 47.680 83.915 ;
        RECT 47.850 83.585 48.200 84.155 ;
        RECT 48.925 84.105 49.590 84.275 ;
        RECT 46.610 83.125 46.780 83.245 ;
        RECT 47.880 83.125 48.200 83.415 ;
        RECT 48.840 83.285 49.190 83.935 ;
        RECT 46.095 82.275 46.375 83.075 ;
        RECT 46.610 82.955 48.200 83.125 ;
        RECT 49.360 83.115 49.590 84.105 ;
        RECT 48.925 82.945 49.590 83.115 ;
        RECT 46.545 82.495 48.200 82.785 ;
        RECT 48.925 82.445 49.095 82.945 ;
        RECT 49.265 82.275 49.595 82.775 ;
        RECT 49.765 82.445 49.950 84.565 ;
        RECT 50.205 84.365 50.455 84.825 ;
        RECT 50.625 84.375 50.960 84.545 ;
        RECT 51.155 84.375 51.830 84.545 ;
        RECT 50.625 84.235 50.795 84.375 ;
        RECT 50.120 83.245 50.400 84.195 ;
        RECT 50.570 84.105 50.795 84.235 ;
        RECT 50.570 83.000 50.740 84.105 ;
        RECT 50.965 83.955 51.490 84.175 ;
        RECT 50.910 83.190 51.150 83.785 ;
        RECT 51.320 83.255 51.490 83.955 ;
        RECT 51.660 83.595 51.830 84.375 ;
        RECT 52.150 84.325 52.520 84.825 ;
        RECT 52.700 84.375 53.105 84.545 ;
        RECT 53.275 84.375 54.060 84.545 ;
        RECT 52.700 84.145 52.870 84.375 ;
        RECT 52.040 83.845 52.870 84.145 ;
        RECT 53.255 83.875 53.720 84.205 ;
        RECT 52.040 83.815 52.240 83.845 ;
        RECT 52.360 83.595 52.530 83.665 ;
        RECT 51.660 83.425 52.530 83.595 ;
        RECT 52.020 83.335 52.530 83.425 ;
        RECT 50.570 82.870 50.875 83.000 ;
        RECT 51.320 82.890 51.850 83.255 ;
        RECT 50.190 82.275 50.455 82.735 ;
        RECT 50.625 82.445 50.875 82.870 ;
        RECT 52.020 82.720 52.190 83.335 ;
        RECT 51.085 82.550 52.190 82.720 ;
        RECT 52.360 82.275 52.530 83.075 ;
        RECT 52.700 82.775 52.870 83.845 ;
        RECT 53.040 82.945 53.230 83.665 ;
        RECT 53.400 82.915 53.720 83.875 ;
        RECT 53.890 83.915 54.060 84.375 ;
        RECT 54.335 84.295 54.545 84.825 ;
        RECT 54.805 84.085 55.135 84.610 ;
        RECT 55.305 84.215 55.475 84.825 ;
        RECT 55.645 84.170 55.975 84.605 ;
        RECT 55.645 84.085 56.025 84.170 ;
        RECT 54.935 83.915 55.135 84.085 ;
        RECT 55.800 84.045 56.025 84.085 ;
        RECT 53.890 83.585 54.765 83.915 ;
        RECT 54.935 83.585 55.685 83.915 ;
        RECT 52.700 82.445 52.950 82.775 ;
        RECT 53.890 82.745 54.060 83.585 ;
        RECT 54.935 83.380 55.125 83.585 ;
        RECT 55.855 83.465 56.025 84.045 ;
        RECT 55.810 83.415 56.025 83.465 ;
        RECT 54.230 83.005 55.125 83.380 ;
        RECT 55.635 83.335 56.025 83.415 ;
        RECT 56.195 84.085 56.580 84.655 ;
        RECT 56.750 84.365 57.075 84.825 ;
        RECT 57.595 84.195 57.875 84.655 ;
        RECT 56.195 83.415 56.475 84.085 ;
        RECT 56.750 84.025 57.875 84.195 ;
        RECT 56.750 83.915 57.200 84.025 ;
        RECT 56.645 83.585 57.200 83.915 ;
        RECT 58.065 83.855 58.465 84.655 ;
        RECT 58.865 84.365 59.135 84.825 ;
        RECT 59.305 84.195 59.590 84.655 ;
        RECT 53.175 82.575 54.060 82.745 ;
        RECT 54.240 82.275 54.555 82.775 ;
        RECT 54.785 82.445 55.125 83.005 ;
        RECT 55.295 82.275 55.465 83.285 ;
        RECT 55.635 82.490 55.965 83.335 ;
        RECT 56.195 82.445 56.580 83.415 ;
        RECT 56.750 83.125 57.200 83.585 ;
        RECT 57.370 83.295 58.465 83.855 ;
        RECT 56.750 82.905 57.875 83.125 ;
        RECT 56.750 82.275 57.075 82.735 ;
        RECT 57.595 82.445 57.875 82.905 ;
        RECT 58.065 82.445 58.465 83.295 ;
        RECT 58.635 84.025 59.590 84.195 ;
        RECT 59.875 84.055 63.385 84.825 ;
        RECT 63.555 84.100 63.845 84.825 ;
        RECT 58.635 83.125 58.845 84.025 ;
        RECT 59.015 83.295 59.705 83.855 ;
        RECT 59.875 83.535 61.525 84.055 ;
        RECT 64.935 84.005 65.195 84.825 ;
        RECT 65.365 84.005 65.695 84.425 ;
        RECT 65.875 84.340 66.665 84.605 ;
        RECT 65.445 83.915 65.695 84.005 ;
        RECT 61.695 83.365 63.385 83.885 ;
        RECT 58.635 82.905 59.590 83.125 ;
        RECT 58.865 82.275 59.135 82.735 ;
        RECT 59.305 82.445 59.590 82.905 ;
        RECT 59.875 82.275 63.385 83.365 ;
        RECT 63.555 82.275 63.845 83.440 ;
        RECT 64.935 82.955 65.275 83.835 ;
        RECT 65.445 83.665 66.240 83.915 ;
        RECT 64.935 82.275 65.195 82.785 ;
        RECT 65.445 82.445 65.615 83.665 ;
        RECT 66.410 83.485 66.665 84.340 ;
        RECT 66.835 84.185 67.035 84.605 ;
        RECT 67.225 84.365 67.555 84.825 ;
        RECT 66.835 83.665 67.245 84.185 ;
        RECT 67.725 84.175 67.985 84.655 ;
        RECT 67.415 83.485 67.645 83.915 ;
        RECT 65.855 83.315 67.645 83.485 ;
        RECT 65.855 82.950 66.105 83.315 ;
        RECT 66.275 82.955 66.605 83.145 ;
        RECT 66.825 83.020 67.540 83.315 ;
        RECT 67.815 83.145 67.985 84.175 ;
        RECT 66.275 82.780 66.470 82.955 ;
        RECT 65.855 82.275 66.470 82.780 ;
        RECT 66.640 82.445 67.115 82.785 ;
        RECT 67.285 82.275 67.500 82.820 ;
        RECT 67.710 82.445 67.985 83.145 ;
        RECT 68.175 84.135 68.415 84.655 ;
        RECT 68.585 84.330 68.980 84.825 ;
        RECT 69.545 84.495 69.715 84.640 ;
        RECT 69.340 84.300 69.715 84.495 ;
        RECT 68.175 83.330 68.350 84.135 ;
        RECT 69.340 83.965 69.510 84.300 ;
        RECT 69.995 84.255 70.235 84.630 ;
        RECT 70.405 84.320 70.740 84.825 ;
        RECT 69.995 84.105 70.215 84.255 ;
        RECT 68.525 83.605 69.510 83.965 ;
        RECT 69.680 83.775 70.215 84.105 ;
        RECT 68.525 83.585 69.810 83.605 ;
        RECT 68.950 83.435 69.810 83.585 ;
        RECT 68.175 82.545 68.480 83.330 ;
        RECT 68.655 82.955 69.350 83.265 ;
        RECT 68.660 82.275 69.345 82.745 ;
        RECT 69.525 82.490 69.810 83.435 ;
        RECT 69.980 83.125 70.215 83.775 ;
        RECT 70.385 83.295 70.685 84.145 ;
        RECT 70.915 84.055 73.505 84.825 ;
        RECT 73.675 84.175 73.935 84.655 ;
        RECT 74.105 84.285 74.355 84.825 ;
        RECT 70.915 83.535 72.125 84.055 ;
        RECT 72.295 83.365 73.505 83.885 ;
        RECT 69.980 82.895 70.655 83.125 ;
        RECT 69.985 82.275 70.315 82.725 ;
        RECT 70.485 82.465 70.655 82.895 ;
        RECT 70.915 82.275 73.505 83.365 ;
        RECT 73.675 83.145 73.845 84.175 ;
        RECT 74.525 84.120 74.745 84.605 ;
        RECT 74.015 83.525 74.245 83.920 ;
        RECT 74.415 83.695 74.745 84.120 ;
        RECT 74.915 84.445 75.805 84.615 ;
        RECT 74.915 83.720 75.085 84.445 ;
        RECT 75.975 84.280 81.320 84.825 ;
        RECT 75.255 83.890 75.805 84.275 ;
        RECT 74.915 83.650 75.805 83.720 ;
        RECT 74.910 83.625 75.805 83.650 ;
        RECT 74.900 83.610 75.805 83.625 ;
        RECT 74.895 83.595 75.805 83.610 ;
        RECT 74.885 83.590 75.805 83.595 ;
        RECT 74.880 83.580 75.805 83.590 ;
        RECT 74.875 83.570 75.805 83.580 ;
        RECT 74.865 83.565 75.805 83.570 ;
        RECT 74.855 83.555 75.805 83.565 ;
        RECT 74.845 83.550 75.805 83.555 ;
        RECT 74.845 83.545 75.180 83.550 ;
        RECT 74.830 83.540 75.180 83.545 ;
        RECT 74.815 83.530 75.180 83.540 ;
        RECT 74.790 83.525 75.180 83.530 ;
        RECT 74.015 83.520 75.180 83.525 ;
        RECT 74.015 83.485 75.150 83.520 ;
        RECT 74.015 83.460 75.115 83.485 ;
        RECT 74.015 83.430 75.085 83.460 ;
        RECT 74.015 83.400 75.065 83.430 ;
        RECT 74.015 83.370 75.045 83.400 ;
        RECT 74.015 83.360 74.975 83.370 ;
        RECT 74.015 83.350 74.950 83.360 ;
        RECT 74.015 83.335 74.930 83.350 ;
        RECT 74.015 83.320 74.910 83.335 ;
        RECT 74.120 83.310 74.905 83.320 ;
        RECT 74.120 83.275 74.890 83.310 ;
        RECT 73.675 82.445 73.950 83.145 ;
        RECT 74.120 83.025 74.875 83.275 ;
        RECT 75.045 82.955 75.375 83.200 ;
        RECT 75.545 83.100 75.805 83.550 ;
        RECT 77.560 83.450 77.900 84.280 ;
        RECT 81.495 84.055 84.085 84.825 ;
        RECT 84.345 84.275 84.515 84.655 ;
        RECT 84.695 84.445 85.025 84.825 ;
        RECT 84.345 84.105 85.010 84.275 ;
        RECT 85.205 84.150 85.465 84.655 ;
        RECT 75.190 82.930 75.375 82.955 ;
        RECT 75.190 82.830 75.805 82.930 ;
        RECT 74.120 82.275 74.375 82.820 ;
        RECT 74.545 82.445 75.025 82.785 ;
        RECT 75.200 82.275 75.805 82.830 ;
        RECT 79.380 82.710 79.730 83.960 ;
        RECT 81.495 83.535 82.705 84.055 ;
        RECT 82.875 83.365 84.085 83.885 ;
        RECT 84.275 83.555 84.605 83.925 ;
        RECT 84.840 83.850 85.010 84.105 ;
        RECT 84.840 83.520 85.125 83.850 ;
        RECT 84.840 83.375 85.010 83.520 ;
        RECT 75.975 82.275 81.320 82.710 ;
        RECT 81.495 82.275 84.085 83.365 ;
        RECT 84.345 83.205 85.010 83.375 ;
        RECT 85.295 83.350 85.465 84.150 ;
        RECT 84.345 82.445 84.515 83.205 ;
        RECT 84.695 82.275 85.025 83.035 ;
        RECT 85.195 82.445 85.465 83.350 ;
        RECT 85.635 84.085 86.020 84.655 ;
        RECT 86.190 84.365 86.515 84.825 ;
        RECT 87.035 84.195 87.315 84.655 ;
        RECT 85.635 83.415 85.915 84.085 ;
        RECT 86.190 84.025 87.315 84.195 ;
        RECT 86.190 83.915 86.640 84.025 ;
        RECT 86.085 83.585 86.640 83.915 ;
        RECT 87.505 83.855 87.905 84.655 ;
        RECT 88.305 84.365 88.575 84.825 ;
        RECT 88.745 84.195 89.030 84.655 ;
        RECT 85.635 82.445 86.020 83.415 ;
        RECT 86.190 83.125 86.640 83.585 ;
        RECT 86.810 83.295 87.905 83.855 ;
        RECT 86.190 82.905 87.315 83.125 ;
        RECT 86.190 82.275 86.515 82.735 ;
        RECT 87.035 82.445 87.315 82.905 ;
        RECT 87.505 82.445 87.905 83.295 ;
        RECT 88.075 84.025 89.030 84.195 ;
        RECT 89.315 84.075 90.525 84.825 ;
        RECT 88.075 83.125 88.285 84.025 ;
        RECT 88.455 83.295 89.145 83.855 ;
        RECT 89.315 83.365 89.835 83.905 ;
        RECT 90.005 83.535 90.525 84.075 ;
        RECT 88.075 82.905 89.030 83.125 ;
        RECT 88.305 82.275 88.575 82.735 ;
        RECT 88.745 82.445 89.030 82.905 ;
        RECT 89.315 82.275 90.525 83.365 ;
        RECT 11.950 82.105 90.610 82.275 ;
        RECT 12.035 81.015 13.245 82.105 ;
        RECT 13.415 81.015 15.085 82.105 ;
        RECT 12.035 80.305 12.555 80.845 ;
        RECT 12.725 80.475 13.245 81.015 ;
        RECT 13.415 80.325 14.165 80.845 ;
        RECT 14.335 80.495 15.085 81.015 ;
        RECT 15.715 81.385 16.175 81.935 ;
        RECT 16.365 81.385 16.695 82.105 ;
        RECT 12.035 79.555 13.245 80.305 ;
        RECT 13.415 79.555 15.085 80.325 ;
        RECT 15.715 80.015 15.965 81.385 ;
        RECT 16.895 81.215 17.195 81.765 ;
        RECT 17.365 81.435 17.645 82.105 ;
        RECT 16.255 81.045 17.195 81.215 ;
        RECT 16.255 80.795 16.425 81.045 ;
        RECT 17.565 80.795 17.830 81.155 ;
        RECT 18.015 80.965 18.275 82.105 ;
        RECT 18.445 80.955 18.775 81.935 ;
        RECT 18.945 80.965 19.225 82.105 ;
        RECT 19.405 81.135 19.735 81.920 ;
        RECT 19.405 80.965 20.085 81.135 ;
        RECT 20.265 80.965 20.595 82.105 ;
        RECT 21.695 80.965 21.955 82.105 ;
        RECT 22.195 81.595 23.810 81.925 ;
        RECT 18.535 80.915 18.710 80.955 ;
        RECT 16.135 80.465 16.425 80.795 ;
        RECT 16.595 80.545 16.935 80.795 ;
        RECT 17.155 80.545 17.830 80.795 ;
        RECT 18.035 80.545 18.370 80.795 ;
        RECT 16.255 80.375 16.425 80.465 ;
        RECT 16.255 80.185 17.645 80.375 ;
        RECT 18.540 80.355 18.710 80.915 ;
        RECT 18.880 80.525 19.215 80.795 ;
        RECT 19.395 80.545 19.745 80.795 ;
        RECT 19.915 80.365 20.085 80.965 ;
        RECT 22.205 80.795 22.375 81.355 ;
        RECT 22.635 81.255 23.810 81.425 ;
        RECT 23.980 81.305 24.260 82.105 ;
        RECT 22.635 80.965 22.965 81.255 ;
        RECT 23.640 81.135 23.810 81.255 ;
        RECT 23.135 80.795 23.380 81.085 ;
        RECT 23.640 80.965 24.300 81.135 ;
        RECT 24.470 80.965 24.745 81.935 ;
        RECT 24.130 80.795 24.300 80.965 ;
        RECT 20.255 80.545 20.605 80.795 ;
        RECT 21.700 80.545 22.035 80.795 ;
        RECT 22.205 80.465 22.920 80.795 ;
        RECT 23.135 80.465 23.960 80.795 ;
        RECT 24.130 80.465 24.405 80.795 ;
        RECT 22.205 80.375 22.455 80.465 ;
        RECT 15.715 79.725 16.275 80.015 ;
        RECT 16.445 79.555 16.695 80.015 ;
        RECT 17.315 79.825 17.645 80.185 ;
        RECT 18.015 79.725 18.710 80.355 ;
        RECT 18.915 79.555 19.225 80.355 ;
        RECT 19.415 79.555 19.655 80.365 ;
        RECT 19.825 79.725 20.155 80.365 ;
        RECT 20.325 79.555 20.595 80.365 ;
        RECT 21.695 79.555 21.955 80.375 ;
        RECT 22.125 79.955 22.455 80.375 ;
        RECT 24.130 80.295 24.300 80.465 ;
        RECT 22.635 80.125 24.300 80.295 ;
        RECT 24.575 80.230 24.745 80.965 ;
        RECT 24.915 80.940 25.205 82.105 ;
        RECT 25.375 81.015 26.585 82.105 ;
        RECT 25.375 80.305 25.895 80.845 ;
        RECT 26.065 80.475 26.585 81.015 ;
        RECT 26.760 80.965 27.095 81.935 ;
        RECT 27.265 80.965 27.435 82.105 ;
        RECT 27.605 81.765 29.635 81.935 ;
        RECT 22.635 79.725 22.895 80.125 ;
        RECT 23.065 79.555 23.395 79.955 ;
        RECT 23.565 79.775 23.735 80.125 ;
        RECT 23.905 79.555 24.280 79.955 ;
        RECT 24.470 79.885 24.745 80.230 ;
        RECT 24.915 79.555 25.205 80.280 ;
        RECT 25.375 79.555 26.585 80.305 ;
        RECT 26.760 80.295 26.930 80.965 ;
        RECT 27.605 80.795 27.775 81.765 ;
        RECT 27.100 80.465 27.355 80.795 ;
        RECT 27.580 80.465 27.775 80.795 ;
        RECT 27.945 81.425 29.070 81.595 ;
        RECT 27.185 80.295 27.355 80.465 ;
        RECT 27.945 80.295 28.115 81.425 ;
        RECT 26.760 79.725 27.015 80.295 ;
        RECT 27.185 80.125 28.115 80.295 ;
        RECT 28.285 81.085 29.295 81.255 ;
        RECT 28.285 80.285 28.455 81.085 ;
        RECT 28.660 80.745 28.935 80.885 ;
        RECT 28.655 80.575 28.935 80.745 ;
        RECT 27.940 80.090 28.115 80.125 ;
        RECT 27.185 79.555 27.515 79.955 ;
        RECT 27.940 79.725 28.470 80.090 ;
        RECT 28.660 79.725 28.935 80.575 ;
        RECT 29.105 79.725 29.295 81.085 ;
        RECT 29.465 81.100 29.635 81.765 ;
        RECT 29.805 81.345 29.975 82.105 ;
        RECT 30.210 81.345 30.725 81.755 ;
        RECT 30.895 81.670 36.240 82.105 ;
        RECT 29.465 80.910 30.215 81.100 ;
        RECT 30.385 80.535 30.725 81.345 ;
        RECT 29.495 80.365 30.725 80.535 ;
        RECT 29.475 79.555 29.985 80.090 ;
        RECT 30.205 79.760 30.450 80.365 ;
        RECT 32.480 80.100 32.820 80.930 ;
        RECT 34.300 80.420 34.650 81.670 ;
        RECT 37.335 81.345 37.850 81.755 ;
        RECT 38.085 81.345 38.255 82.105 ;
        RECT 38.425 81.765 40.455 81.935 ;
        RECT 37.335 80.535 37.675 81.345 ;
        RECT 38.425 81.100 38.595 81.765 ;
        RECT 38.990 81.425 40.115 81.595 ;
        RECT 37.845 80.910 38.595 81.100 ;
        RECT 38.765 81.085 39.775 81.255 ;
        RECT 37.335 80.365 38.565 80.535 ;
        RECT 30.895 79.555 36.240 80.100 ;
        RECT 37.610 79.760 37.855 80.365 ;
        RECT 38.075 79.555 38.585 80.090 ;
        RECT 38.765 79.725 38.955 81.085 ;
        RECT 39.125 80.065 39.400 80.885 ;
        RECT 39.605 80.285 39.775 81.085 ;
        RECT 39.945 80.295 40.115 81.425 ;
        RECT 40.285 80.795 40.455 81.765 ;
        RECT 40.625 80.965 40.795 82.105 ;
        RECT 40.965 80.965 41.300 81.935 ;
        RECT 41.475 81.015 43.145 82.105 ;
        RECT 40.285 80.465 40.480 80.795 ;
        RECT 40.705 80.465 40.960 80.795 ;
        RECT 40.705 80.295 40.875 80.465 ;
        RECT 41.130 80.295 41.300 80.965 ;
        RECT 39.945 80.125 40.875 80.295 ;
        RECT 39.945 80.090 40.120 80.125 ;
        RECT 39.125 79.895 39.405 80.065 ;
        RECT 39.125 79.725 39.400 79.895 ;
        RECT 39.590 79.725 40.120 80.090 ;
        RECT 40.545 79.555 40.875 79.955 ;
        RECT 41.045 79.725 41.300 80.295 ;
        RECT 41.475 80.325 42.225 80.845 ;
        RECT 42.395 80.495 43.145 81.015 ;
        RECT 43.315 80.965 43.700 81.935 ;
        RECT 43.870 81.645 44.195 82.105 ;
        RECT 44.715 81.475 44.995 81.935 ;
        RECT 43.870 81.255 44.995 81.475 ;
        RECT 41.475 79.555 43.145 80.325 ;
        RECT 43.315 80.295 43.595 80.965 ;
        RECT 43.870 80.795 44.320 81.255 ;
        RECT 45.185 81.085 45.585 81.935 ;
        RECT 45.985 81.645 46.255 82.105 ;
        RECT 46.425 81.475 46.710 81.935 ;
        RECT 43.765 80.465 44.320 80.795 ;
        RECT 44.490 80.525 45.585 81.085 ;
        RECT 43.870 80.355 44.320 80.465 ;
        RECT 43.315 79.725 43.700 80.295 ;
        RECT 43.870 80.185 44.995 80.355 ;
        RECT 43.870 79.555 44.195 80.015 ;
        RECT 44.715 79.725 44.995 80.185 ;
        RECT 45.185 79.725 45.585 80.525 ;
        RECT 45.755 81.255 46.710 81.475 ;
        RECT 47.110 81.475 47.395 81.935 ;
        RECT 47.565 81.645 47.835 82.105 ;
        RECT 47.110 81.255 48.065 81.475 ;
        RECT 45.755 80.355 45.965 81.255 ;
        RECT 46.135 80.525 46.825 81.085 ;
        RECT 46.995 80.525 47.685 81.085 ;
        RECT 47.855 80.355 48.065 81.255 ;
        RECT 45.755 80.185 46.710 80.355 ;
        RECT 45.985 79.555 46.255 80.015 ;
        RECT 46.425 79.725 46.710 80.185 ;
        RECT 47.110 80.185 48.065 80.355 ;
        RECT 48.235 81.085 48.635 81.935 ;
        RECT 48.825 81.475 49.105 81.935 ;
        RECT 49.625 81.645 49.950 82.105 ;
        RECT 48.825 81.255 49.950 81.475 ;
        RECT 48.235 80.525 49.330 81.085 ;
        RECT 49.500 80.795 49.950 81.255 ;
        RECT 50.120 80.965 50.505 81.935 ;
        RECT 47.110 79.725 47.395 80.185 ;
        RECT 47.565 79.555 47.835 80.015 ;
        RECT 48.235 79.725 48.635 80.525 ;
        RECT 49.500 80.465 50.055 80.795 ;
        RECT 49.500 80.355 49.950 80.465 ;
        RECT 48.825 80.185 49.950 80.355 ;
        RECT 50.225 80.295 50.505 80.965 ;
        RECT 50.675 80.940 50.965 82.105 ;
        RECT 51.135 81.235 51.410 81.935 ;
        RECT 51.580 81.560 51.835 82.105 ;
        RECT 52.005 81.595 52.485 81.935 ;
        RECT 52.660 81.550 53.265 82.105 ;
        RECT 52.650 81.450 53.265 81.550 ;
        RECT 52.650 81.425 52.835 81.450 ;
        RECT 48.825 79.725 49.105 80.185 ;
        RECT 49.625 79.555 49.950 80.015 ;
        RECT 50.120 79.725 50.505 80.295 ;
        RECT 50.675 79.555 50.965 80.280 ;
        RECT 51.135 80.205 51.305 81.235 ;
        RECT 51.580 81.105 52.335 81.355 ;
        RECT 52.505 81.180 52.835 81.425 ;
        RECT 51.580 81.070 52.350 81.105 ;
        RECT 51.580 81.060 52.365 81.070 ;
        RECT 51.475 81.045 52.370 81.060 ;
        RECT 51.475 81.030 52.390 81.045 ;
        RECT 51.475 81.020 52.410 81.030 ;
        RECT 51.475 81.010 52.435 81.020 ;
        RECT 51.475 80.980 52.505 81.010 ;
        RECT 51.475 80.950 52.525 80.980 ;
        RECT 51.475 80.920 52.545 80.950 ;
        RECT 51.475 80.895 52.575 80.920 ;
        RECT 51.475 80.860 52.610 80.895 ;
        RECT 51.475 80.855 52.640 80.860 ;
        RECT 51.475 80.460 51.705 80.855 ;
        RECT 52.250 80.850 52.640 80.855 ;
        RECT 52.275 80.840 52.640 80.850 ;
        RECT 52.290 80.835 52.640 80.840 ;
        RECT 52.305 80.830 52.640 80.835 ;
        RECT 53.005 80.830 53.265 81.280 ;
        RECT 52.305 80.825 53.265 80.830 ;
        RECT 52.315 80.815 53.265 80.825 ;
        RECT 52.325 80.810 53.265 80.815 ;
        RECT 52.335 80.800 53.265 80.810 ;
        RECT 52.340 80.790 53.265 80.800 ;
        RECT 52.345 80.785 53.265 80.790 ;
        RECT 52.355 80.770 53.265 80.785 ;
        RECT 52.360 80.755 53.265 80.770 ;
        RECT 52.370 80.730 53.265 80.755 ;
        RECT 51.875 80.260 52.205 80.685 ;
        RECT 51.135 79.725 51.395 80.205 ;
        RECT 51.565 79.555 51.815 80.095 ;
        RECT 51.985 79.775 52.205 80.260 ;
        RECT 52.375 80.660 53.265 80.730 ;
        RECT 53.440 80.965 53.775 81.935 ;
        RECT 53.945 80.965 54.115 82.105 ;
        RECT 54.285 81.765 56.315 81.935 ;
        RECT 52.375 79.935 52.545 80.660 ;
        RECT 52.715 80.105 53.265 80.490 ;
        RECT 53.440 80.295 53.610 80.965 ;
        RECT 54.285 80.795 54.455 81.765 ;
        RECT 53.780 80.465 54.035 80.795 ;
        RECT 54.260 80.465 54.455 80.795 ;
        RECT 54.625 81.425 55.750 81.595 ;
        RECT 53.865 80.295 54.035 80.465 ;
        RECT 54.625 80.295 54.795 81.425 ;
        RECT 52.375 79.765 53.265 79.935 ;
        RECT 53.440 79.725 53.695 80.295 ;
        RECT 53.865 80.125 54.795 80.295 ;
        RECT 54.965 81.085 55.975 81.255 ;
        RECT 54.965 80.285 55.135 81.085 ;
        RECT 54.620 80.090 54.795 80.125 ;
        RECT 53.865 79.555 54.195 79.955 ;
        RECT 54.620 79.725 55.150 80.090 ;
        RECT 55.340 80.065 55.615 80.885 ;
        RECT 55.335 79.895 55.615 80.065 ;
        RECT 55.340 79.725 55.615 79.895 ;
        RECT 55.785 79.725 55.975 81.085 ;
        RECT 56.145 81.100 56.315 81.765 ;
        RECT 56.485 81.345 56.655 82.105 ;
        RECT 56.890 81.345 57.405 81.755 ;
        RECT 57.575 81.670 62.920 82.105 ;
        RECT 56.145 80.910 56.895 81.100 ;
        RECT 57.065 80.535 57.405 81.345 ;
        RECT 56.175 80.365 57.405 80.535 ;
        RECT 56.155 79.555 56.665 80.090 ;
        RECT 56.885 79.760 57.130 80.365 ;
        RECT 59.160 80.100 59.500 80.930 ;
        RECT 60.980 80.420 61.330 81.670 ;
        RECT 63.210 81.475 63.495 81.935 ;
        RECT 63.665 81.645 63.935 82.105 ;
        RECT 63.210 81.255 64.165 81.475 ;
        RECT 63.095 80.525 63.785 81.085 ;
        RECT 63.955 80.355 64.165 81.255 ;
        RECT 63.210 80.185 64.165 80.355 ;
        RECT 64.335 81.085 64.735 81.935 ;
        RECT 64.925 81.475 65.205 81.935 ;
        RECT 65.725 81.645 66.050 82.105 ;
        RECT 64.925 81.255 66.050 81.475 ;
        RECT 64.335 80.525 65.430 81.085 ;
        RECT 65.600 80.795 66.050 81.255 ;
        RECT 66.220 80.965 66.605 81.935 ;
        RECT 66.775 81.550 67.380 82.105 ;
        RECT 67.555 81.595 68.035 81.935 ;
        RECT 68.205 81.560 68.460 82.105 ;
        RECT 66.775 81.450 67.390 81.550 ;
        RECT 67.205 81.425 67.390 81.450 ;
        RECT 57.575 79.555 62.920 80.100 ;
        RECT 63.210 79.725 63.495 80.185 ;
        RECT 63.665 79.555 63.935 80.015 ;
        RECT 64.335 79.725 64.735 80.525 ;
        RECT 65.600 80.465 66.155 80.795 ;
        RECT 65.600 80.355 66.050 80.465 ;
        RECT 64.925 80.185 66.050 80.355 ;
        RECT 66.325 80.295 66.605 80.965 ;
        RECT 66.775 80.830 67.035 81.280 ;
        RECT 67.205 81.180 67.535 81.425 ;
        RECT 67.705 81.105 68.460 81.355 ;
        RECT 68.630 81.235 68.905 81.935 ;
        RECT 67.690 81.070 68.460 81.105 ;
        RECT 67.675 81.060 68.460 81.070 ;
        RECT 67.670 81.045 68.565 81.060 ;
        RECT 67.650 81.030 68.565 81.045 ;
        RECT 67.630 81.020 68.565 81.030 ;
        RECT 67.605 81.010 68.565 81.020 ;
        RECT 67.535 80.980 68.565 81.010 ;
        RECT 67.515 80.950 68.565 80.980 ;
        RECT 67.495 80.920 68.565 80.950 ;
        RECT 67.465 80.895 68.565 80.920 ;
        RECT 67.430 80.860 68.565 80.895 ;
        RECT 67.400 80.855 68.565 80.860 ;
        RECT 67.400 80.850 67.790 80.855 ;
        RECT 67.400 80.840 67.765 80.850 ;
        RECT 67.400 80.835 67.750 80.840 ;
        RECT 67.400 80.830 67.735 80.835 ;
        RECT 66.775 80.825 67.735 80.830 ;
        RECT 66.775 80.815 67.725 80.825 ;
        RECT 66.775 80.810 67.715 80.815 ;
        RECT 66.775 80.800 67.705 80.810 ;
        RECT 66.775 80.790 67.700 80.800 ;
        RECT 66.775 80.785 67.695 80.790 ;
        RECT 66.775 80.770 67.685 80.785 ;
        RECT 66.775 80.755 67.680 80.770 ;
        RECT 66.775 80.730 67.670 80.755 ;
        RECT 66.775 80.660 67.665 80.730 ;
        RECT 64.925 79.725 65.205 80.185 ;
        RECT 65.725 79.555 66.050 80.015 ;
        RECT 66.220 79.725 66.605 80.295 ;
        RECT 66.775 80.105 67.325 80.490 ;
        RECT 67.495 79.935 67.665 80.660 ;
        RECT 66.775 79.765 67.665 79.935 ;
        RECT 67.835 80.260 68.165 80.685 ;
        RECT 68.335 80.460 68.565 80.855 ;
        RECT 67.835 79.775 68.055 80.260 ;
        RECT 68.735 80.205 68.905 81.235 ;
        RECT 69.075 81.015 71.665 82.105 ;
        RECT 68.225 79.555 68.475 80.095 ;
        RECT 68.645 79.725 68.905 80.205 ;
        RECT 69.075 80.325 70.285 80.845 ;
        RECT 70.455 80.495 71.665 81.015 ;
        RECT 72.450 81.095 72.750 81.935 ;
        RECT 72.945 81.265 73.195 82.105 ;
        RECT 73.785 81.515 74.590 81.935 ;
        RECT 73.365 81.345 74.930 81.515 ;
        RECT 73.365 81.095 73.535 81.345 ;
        RECT 72.450 80.925 73.535 81.095 ;
        RECT 72.295 80.465 72.625 80.755 ;
        RECT 69.075 79.555 71.665 80.325 ;
        RECT 72.795 80.295 72.965 80.925 ;
        RECT 73.705 80.795 74.025 81.175 ;
        RECT 73.135 80.545 73.465 80.755 ;
        RECT 73.645 80.545 74.025 80.795 ;
        RECT 74.215 80.755 74.590 81.175 ;
        RECT 74.760 81.095 74.930 81.345 ;
        RECT 75.100 81.265 75.430 82.105 ;
        RECT 75.600 81.345 76.265 81.935 ;
        RECT 74.760 80.925 75.680 81.095 ;
        RECT 75.510 80.755 75.680 80.925 ;
        RECT 74.215 80.745 74.700 80.755 ;
        RECT 74.195 80.575 74.700 80.745 ;
        RECT 74.215 80.545 74.700 80.575 ;
        RECT 74.890 80.545 75.340 80.755 ;
        RECT 75.510 80.545 75.845 80.755 ;
        RECT 76.015 80.375 76.265 81.345 ;
        RECT 76.435 80.940 76.725 82.105 ;
        RECT 76.900 81.715 77.235 81.935 ;
        RECT 78.240 81.725 78.595 82.105 ;
        RECT 76.900 81.095 77.155 81.715 ;
        RECT 77.405 81.555 77.635 81.595 ;
        RECT 78.765 81.555 79.015 81.935 ;
        RECT 77.405 81.355 79.015 81.555 ;
        RECT 77.405 81.265 77.590 81.355 ;
        RECT 78.180 81.345 79.015 81.355 ;
        RECT 79.265 81.325 79.515 82.105 ;
        RECT 79.685 81.255 79.945 81.935 ;
        RECT 80.205 81.435 80.375 81.935 ;
        RECT 80.545 81.605 80.875 82.105 ;
        RECT 80.205 81.265 80.870 81.435 ;
        RECT 77.745 81.155 78.075 81.185 ;
        RECT 77.745 81.095 79.545 81.155 ;
        RECT 76.900 80.985 79.605 81.095 ;
        RECT 76.900 80.925 78.075 80.985 ;
        RECT 79.405 80.950 79.605 80.985 ;
        RECT 76.895 80.545 77.385 80.745 ;
        RECT 77.575 80.545 78.050 80.755 ;
        RECT 72.455 80.115 72.965 80.295 ;
        RECT 73.370 80.205 75.070 80.375 ;
        RECT 73.370 80.115 73.755 80.205 ;
        RECT 72.455 79.725 72.785 80.115 ;
        RECT 72.955 79.775 74.140 79.945 ;
        RECT 74.400 79.555 74.570 80.025 ;
        RECT 74.740 79.740 75.070 80.205 ;
        RECT 75.240 79.555 75.410 80.375 ;
        RECT 75.580 79.735 76.265 80.375 ;
        RECT 76.435 79.555 76.725 80.280 ;
        RECT 76.900 79.555 77.355 80.320 ;
        RECT 77.830 80.145 78.050 80.545 ;
        RECT 78.295 80.545 78.625 80.755 ;
        RECT 78.295 80.145 78.505 80.545 ;
        RECT 78.795 80.510 79.205 80.815 ;
        RECT 79.435 80.375 79.605 80.950 ;
        RECT 79.335 80.255 79.605 80.375 ;
        RECT 78.760 80.210 79.605 80.255 ;
        RECT 78.760 80.085 79.515 80.210 ;
        RECT 78.760 79.935 78.930 80.085 ;
        RECT 79.775 80.065 79.945 81.255 ;
        RECT 80.120 80.445 80.470 81.095 ;
        RECT 80.640 80.275 80.870 81.265 ;
        RECT 79.715 80.055 79.945 80.065 ;
        RECT 77.630 79.725 78.930 79.935 ;
        RECT 79.185 79.555 79.515 79.915 ;
        RECT 79.685 79.725 79.945 80.055 ;
        RECT 80.205 80.105 80.870 80.275 ;
        RECT 80.205 79.815 80.375 80.105 ;
        RECT 80.545 79.555 80.875 79.935 ;
        RECT 81.045 79.815 81.230 81.935 ;
        RECT 81.470 81.645 81.735 82.105 ;
        RECT 81.905 81.510 82.155 81.935 ;
        RECT 82.365 81.660 83.470 81.830 ;
        RECT 81.850 81.380 82.155 81.510 ;
        RECT 81.400 80.185 81.680 81.135 ;
        RECT 81.850 80.275 82.020 81.380 ;
        RECT 82.190 80.595 82.430 81.190 ;
        RECT 82.600 81.125 83.130 81.490 ;
        RECT 82.600 80.425 82.770 81.125 ;
        RECT 83.300 81.045 83.470 81.660 ;
        RECT 83.640 81.305 83.810 82.105 ;
        RECT 83.980 81.605 84.230 81.935 ;
        RECT 84.455 81.635 85.340 81.805 ;
        RECT 83.300 80.955 83.810 81.045 ;
        RECT 81.850 80.145 82.075 80.275 ;
        RECT 82.245 80.205 82.770 80.425 ;
        RECT 82.940 80.785 83.810 80.955 ;
        RECT 81.485 79.555 81.735 80.015 ;
        RECT 81.905 80.005 82.075 80.145 ;
        RECT 82.940 80.005 83.110 80.785 ;
        RECT 83.640 80.715 83.810 80.785 ;
        RECT 83.320 80.535 83.520 80.565 ;
        RECT 83.980 80.535 84.150 81.605 ;
        RECT 84.320 80.715 84.510 81.435 ;
        RECT 83.320 80.235 84.150 80.535 ;
        RECT 84.680 80.505 85.000 81.465 ;
        RECT 81.905 79.835 82.240 80.005 ;
        RECT 82.435 79.835 83.110 80.005 ;
        RECT 83.430 79.555 83.800 80.055 ;
        RECT 83.980 80.005 84.150 80.235 ;
        RECT 84.535 80.175 85.000 80.505 ;
        RECT 85.170 80.795 85.340 81.635 ;
        RECT 85.520 81.605 85.835 82.105 ;
        RECT 86.065 81.375 86.405 81.935 ;
        RECT 85.510 81.000 86.405 81.375 ;
        RECT 86.575 81.095 86.745 82.105 ;
        RECT 86.215 80.795 86.405 81.000 ;
        RECT 86.915 81.045 87.245 81.890 ;
        RECT 87.565 81.175 87.735 81.935 ;
        RECT 87.950 81.345 88.280 82.105 ;
        RECT 86.915 80.965 87.305 81.045 ;
        RECT 87.565 81.005 88.280 81.175 ;
        RECT 88.450 81.030 88.705 81.935 ;
        RECT 87.090 80.915 87.305 80.965 ;
        RECT 85.170 80.465 86.045 80.795 ;
        RECT 86.215 80.465 86.965 80.795 ;
        RECT 85.170 80.005 85.340 80.465 ;
        RECT 86.215 80.295 86.415 80.465 ;
        RECT 87.135 80.335 87.305 80.915 ;
        RECT 87.475 80.455 87.830 80.825 ;
        RECT 88.110 80.795 88.280 81.005 ;
        RECT 88.110 80.465 88.365 80.795 ;
        RECT 87.080 80.295 87.305 80.335 ;
        RECT 83.980 79.835 84.385 80.005 ;
        RECT 84.555 79.835 85.340 80.005 ;
        RECT 85.615 79.555 85.825 80.085 ;
        RECT 86.085 79.770 86.415 80.295 ;
        RECT 86.925 80.210 87.305 80.295 ;
        RECT 88.110 80.275 88.280 80.465 ;
        RECT 88.535 80.300 88.705 81.030 ;
        RECT 88.880 80.955 89.140 82.105 ;
        RECT 89.315 81.015 90.525 82.105 ;
        RECT 99.990 81.095 100.160 87.615 ;
        RECT 100.640 84.975 100.990 87.135 ;
        RECT 100.640 81.575 100.990 83.735 ;
        RECT 101.470 81.095 101.640 87.615 ;
        RECT 102.120 84.975 102.470 87.135 ;
        RECT 102.120 81.575 102.470 83.735 ;
        RECT 102.950 81.095 103.120 87.615 ;
        RECT 103.600 84.975 103.950 87.135 ;
        RECT 103.600 81.575 103.950 83.735 ;
        RECT 104.430 81.095 104.600 87.615 ;
        RECT 105.080 84.975 105.430 87.135 ;
        RECT 105.080 81.575 105.430 83.735 ;
        RECT 105.910 81.095 106.080 87.615 ;
        RECT 106.560 84.975 106.910 87.135 ;
        RECT 106.560 81.575 106.910 83.735 ;
        RECT 107.390 81.095 107.560 87.615 ;
        RECT 108.040 84.975 108.390 87.135 ;
        RECT 108.040 81.575 108.390 83.735 ;
        RECT 108.870 81.095 109.040 87.615 ;
        RECT 109.520 84.975 109.870 87.135 ;
        RECT 109.520 81.575 109.870 83.735 ;
        RECT 110.350 81.095 110.520 87.615 ;
        RECT 111.000 84.975 111.350 87.135 ;
        RECT 111.000 81.575 111.350 83.735 ;
        RECT 111.830 81.095 112.000 87.615 ;
        RECT 112.480 84.975 112.830 87.135 ;
        RECT 112.480 81.575 112.830 83.735 ;
        RECT 113.310 81.095 113.480 87.615 ;
        RECT 117.590 82.770 117.760 92.260 ;
        RECT 118.390 91.750 119.390 91.920 ;
        RECT 118.160 83.495 118.330 91.535 ;
        RECT 119.450 83.495 119.620 91.535 ;
        RECT 118.390 83.110 119.390 83.280 ;
        RECT 120.020 82.770 120.190 92.260 ;
        RECT 120.820 91.750 122.820 91.920 ;
        RECT 120.590 83.495 120.760 91.535 ;
        RECT 122.880 83.495 123.050 91.535 ;
        RECT 120.820 83.110 122.820 83.280 ;
        RECT 123.450 82.770 123.620 92.260 ;
        RECT 124.250 91.750 126.250 91.920 ;
        RECT 124.020 83.495 124.190 91.535 ;
        RECT 126.310 83.495 126.480 91.535 ;
        RECT 124.250 83.110 126.250 83.280 ;
        RECT 126.880 82.770 127.050 92.260 ;
        RECT 127.680 91.750 128.680 91.920 ;
        RECT 127.450 83.495 127.620 91.535 ;
        RECT 128.740 83.495 128.910 91.535 ;
        RECT 129.310 86.660 130.440 92.260 ;
        RECT 127.680 83.110 128.680 83.280 ;
        RECT 129.310 82.770 130.460 86.660 ;
        RECT 134.410 84.640 139.730 85.560 ;
        RECT 134.410 84.540 136.170 84.640 ;
        RECT 117.590 82.600 130.460 82.770 ;
        RECT 129.340 82.570 130.460 82.600 ;
        RECT 89.315 80.475 89.835 81.015 ;
        RECT 99.990 80.925 113.480 81.095 ;
        RECT 129.450 81.350 130.450 82.570 ;
        RECT 126.900 81.010 129.140 81.020 ;
        RECT 86.585 79.555 86.755 80.165 ;
        RECT 86.925 79.775 87.255 80.210 ;
        RECT 87.565 80.105 88.280 80.275 ;
        RECT 87.565 79.725 87.735 80.105 ;
        RECT 87.950 79.555 88.280 79.935 ;
        RECT 88.450 79.725 88.705 80.300 ;
        RECT 88.880 79.555 89.140 80.395 ;
        RECT 90.005 80.305 90.525 80.845 ;
        RECT 89.315 79.555 90.525 80.305 ;
        RECT 11.950 79.385 90.610 79.555 ;
        RECT 12.035 78.635 13.245 79.385 ;
        RECT 14.425 78.835 14.595 79.125 ;
        RECT 14.765 79.005 15.095 79.385 ;
        RECT 14.425 78.665 15.090 78.835 ;
        RECT 12.035 78.095 12.555 78.635 ;
        RECT 12.725 77.925 13.245 78.465 ;
        RECT 12.035 76.835 13.245 77.925 ;
        RECT 14.340 77.845 14.690 78.495 ;
        RECT 14.860 77.675 15.090 78.665 ;
        RECT 14.425 77.505 15.090 77.675 ;
        RECT 14.425 77.005 14.595 77.505 ;
        RECT 14.765 76.835 15.095 77.335 ;
        RECT 15.265 77.005 15.450 79.125 ;
        RECT 15.705 78.925 15.955 79.385 ;
        RECT 16.125 78.935 16.460 79.105 ;
        RECT 16.655 78.935 17.330 79.105 ;
        RECT 16.125 78.795 16.295 78.935 ;
        RECT 15.620 77.805 15.900 78.755 ;
        RECT 16.070 78.665 16.295 78.795 ;
        RECT 16.070 77.560 16.240 78.665 ;
        RECT 16.465 78.515 16.990 78.735 ;
        RECT 16.410 77.750 16.650 78.345 ;
        RECT 16.820 77.815 16.990 78.515 ;
        RECT 17.160 78.155 17.330 78.935 ;
        RECT 17.650 78.885 18.020 79.385 ;
        RECT 18.200 78.935 18.605 79.105 ;
        RECT 18.775 78.935 19.560 79.105 ;
        RECT 18.200 78.705 18.370 78.935 ;
        RECT 17.540 78.405 18.370 78.705 ;
        RECT 18.755 78.435 19.220 78.765 ;
        RECT 17.540 78.375 17.740 78.405 ;
        RECT 17.860 78.155 18.030 78.225 ;
        RECT 17.160 77.985 18.030 78.155 ;
        RECT 17.520 77.895 18.030 77.985 ;
        RECT 16.070 77.430 16.375 77.560 ;
        RECT 16.820 77.450 17.350 77.815 ;
        RECT 15.690 76.835 15.955 77.295 ;
        RECT 16.125 77.005 16.375 77.430 ;
        RECT 17.520 77.280 17.690 77.895 ;
        RECT 16.585 77.110 17.690 77.280 ;
        RECT 17.860 76.835 18.030 77.635 ;
        RECT 18.200 77.335 18.370 78.405 ;
        RECT 18.540 77.505 18.730 78.225 ;
        RECT 18.900 77.475 19.220 78.435 ;
        RECT 19.390 78.475 19.560 78.935 ;
        RECT 19.835 78.855 20.045 79.385 ;
        RECT 20.305 78.645 20.635 79.170 ;
        RECT 20.805 78.775 20.975 79.385 ;
        RECT 21.145 78.730 21.475 79.165 ;
        RECT 21.145 78.645 21.525 78.730 ;
        RECT 20.435 78.475 20.635 78.645 ;
        RECT 21.300 78.605 21.525 78.645 ;
        RECT 19.390 78.145 20.265 78.475 ;
        RECT 20.435 78.145 21.185 78.475 ;
        RECT 18.200 77.005 18.450 77.335 ;
        RECT 19.390 77.305 19.560 78.145 ;
        RECT 20.435 77.940 20.625 78.145 ;
        RECT 21.355 78.025 21.525 78.605 ;
        RECT 21.695 78.615 23.365 79.385 ;
        RECT 21.695 78.095 22.445 78.615 ;
        RECT 23.535 78.565 23.795 79.385 ;
        RECT 23.965 78.565 24.295 78.985 ;
        RECT 24.475 78.815 24.735 79.215 ;
        RECT 24.905 78.985 25.235 79.385 ;
        RECT 25.405 78.815 25.575 79.165 ;
        RECT 25.745 78.985 26.120 79.385 ;
        RECT 24.475 78.645 26.140 78.815 ;
        RECT 26.310 78.710 26.585 79.055 ;
        RECT 24.045 78.475 24.295 78.565 ;
        RECT 25.970 78.475 26.140 78.645 ;
        RECT 21.310 77.975 21.525 78.025 ;
        RECT 19.730 77.565 20.625 77.940 ;
        RECT 21.135 77.895 21.525 77.975 ;
        RECT 22.615 77.925 23.365 78.445 ;
        RECT 23.540 78.145 23.875 78.395 ;
        RECT 24.045 78.145 24.760 78.475 ;
        RECT 24.975 78.145 25.800 78.475 ;
        RECT 25.970 78.145 26.245 78.475 ;
        RECT 18.675 77.135 19.560 77.305 ;
        RECT 19.740 76.835 20.055 77.335 ;
        RECT 20.285 77.005 20.625 77.565 ;
        RECT 20.795 76.835 20.965 77.845 ;
        RECT 21.135 77.050 21.465 77.895 ;
        RECT 21.695 76.835 23.365 77.925 ;
        RECT 23.535 76.835 23.795 77.975 ;
        RECT 24.045 77.585 24.215 78.145 ;
        RECT 24.475 77.685 24.805 77.975 ;
        RECT 24.975 77.855 25.220 78.145 ;
        RECT 25.970 77.975 26.140 78.145 ;
        RECT 26.415 77.975 26.585 78.710 ;
        RECT 27.305 78.835 27.475 79.125 ;
        RECT 27.645 79.005 27.975 79.385 ;
        RECT 27.305 78.665 27.970 78.835 ;
        RECT 25.480 77.805 26.140 77.975 ;
        RECT 25.480 77.685 25.650 77.805 ;
        RECT 24.475 77.515 25.650 77.685 ;
        RECT 24.035 77.015 25.650 77.345 ;
        RECT 25.820 76.835 26.100 77.635 ;
        RECT 26.310 77.005 26.585 77.975 ;
        RECT 27.220 77.845 27.570 78.495 ;
        RECT 27.740 77.675 27.970 78.665 ;
        RECT 27.305 77.505 27.970 77.675 ;
        RECT 27.305 77.005 27.475 77.505 ;
        RECT 27.645 76.835 27.975 77.335 ;
        RECT 28.145 77.005 28.330 79.125 ;
        RECT 28.585 78.925 28.835 79.385 ;
        RECT 29.005 78.935 29.340 79.105 ;
        RECT 29.535 78.935 30.210 79.105 ;
        RECT 29.005 78.795 29.175 78.935 ;
        RECT 28.500 77.805 28.780 78.755 ;
        RECT 28.950 78.665 29.175 78.795 ;
        RECT 28.950 77.560 29.120 78.665 ;
        RECT 29.345 78.515 29.870 78.735 ;
        RECT 29.290 77.750 29.530 78.345 ;
        RECT 29.700 77.815 29.870 78.515 ;
        RECT 30.040 78.155 30.210 78.935 ;
        RECT 30.530 78.885 30.900 79.385 ;
        RECT 31.080 78.935 31.485 79.105 ;
        RECT 31.655 78.935 32.440 79.105 ;
        RECT 31.080 78.705 31.250 78.935 ;
        RECT 30.420 78.405 31.250 78.705 ;
        RECT 31.635 78.435 32.100 78.765 ;
        RECT 30.420 78.375 30.620 78.405 ;
        RECT 30.740 78.155 30.910 78.225 ;
        RECT 30.040 77.985 30.910 78.155 ;
        RECT 30.400 77.895 30.910 77.985 ;
        RECT 28.950 77.430 29.255 77.560 ;
        RECT 29.700 77.450 30.230 77.815 ;
        RECT 28.570 76.835 28.835 77.295 ;
        RECT 29.005 77.005 29.255 77.430 ;
        RECT 30.400 77.280 30.570 77.895 ;
        RECT 29.465 77.110 30.570 77.280 ;
        RECT 30.740 76.835 30.910 77.635 ;
        RECT 31.080 77.335 31.250 78.405 ;
        RECT 31.420 77.505 31.610 78.225 ;
        RECT 31.780 77.475 32.100 78.435 ;
        RECT 32.270 78.475 32.440 78.935 ;
        RECT 32.715 78.855 32.925 79.385 ;
        RECT 33.185 78.645 33.515 79.170 ;
        RECT 33.685 78.775 33.855 79.385 ;
        RECT 34.025 78.730 34.355 79.165 ;
        RECT 34.525 78.870 34.695 79.385 ;
        RECT 34.025 78.645 34.405 78.730 ;
        RECT 33.315 78.475 33.515 78.645 ;
        RECT 34.180 78.605 34.405 78.645 ;
        RECT 32.270 78.145 33.145 78.475 ;
        RECT 33.315 78.145 34.065 78.475 ;
        RECT 31.080 77.005 31.330 77.335 ;
        RECT 32.270 77.305 32.440 78.145 ;
        RECT 33.315 77.940 33.505 78.145 ;
        RECT 34.235 78.025 34.405 78.605 ;
        RECT 35.035 78.615 37.625 79.385 ;
        RECT 37.795 78.660 38.085 79.385 ;
        RECT 38.345 78.835 38.515 79.125 ;
        RECT 38.685 79.005 39.015 79.385 ;
        RECT 38.345 78.665 39.010 78.835 ;
        RECT 35.035 78.095 36.245 78.615 ;
        RECT 34.190 77.975 34.405 78.025 ;
        RECT 32.610 77.565 33.505 77.940 ;
        RECT 34.015 77.895 34.405 77.975 ;
        RECT 36.415 77.925 37.625 78.445 ;
        RECT 31.555 77.135 32.440 77.305 ;
        RECT 32.620 76.835 32.935 77.335 ;
        RECT 33.165 77.005 33.505 77.565 ;
        RECT 33.675 76.835 33.845 77.845 ;
        RECT 34.015 77.050 34.345 77.895 ;
        RECT 34.515 76.835 34.685 77.750 ;
        RECT 35.035 76.835 37.625 77.925 ;
        RECT 37.795 76.835 38.085 78.000 ;
        RECT 38.260 77.845 38.610 78.495 ;
        RECT 38.780 77.675 39.010 78.665 ;
        RECT 38.345 77.505 39.010 77.675 ;
        RECT 38.345 77.005 38.515 77.505 ;
        RECT 38.685 76.835 39.015 77.335 ;
        RECT 39.185 77.005 39.370 79.125 ;
        RECT 39.625 78.925 39.875 79.385 ;
        RECT 40.045 78.935 40.380 79.105 ;
        RECT 40.575 78.935 41.250 79.105 ;
        RECT 40.045 78.795 40.215 78.935 ;
        RECT 39.540 77.805 39.820 78.755 ;
        RECT 39.990 78.665 40.215 78.795 ;
        RECT 39.990 77.560 40.160 78.665 ;
        RECT 40.385 78.515 40.910 78.735 ;
        RECT 40.330 77.750 40.570 78.345 ;
        RECT 40.740 77.815 40.910 78.515 ;
        RECT 41.080 78.155 41.250 78.935 ;
        RECT 41.570 78.885 41.940 79.385 ;
        RECT 42.120 78.935 42.525 79.105 ;
        RECT 42.695 78.935 43.480 79.105 ;
        RECT 42.120 78.705 42.290 78.935 ;
        RECT 41.460 78.405 42.290 78.705 ;
        RECT 42.675 78.435 43.140 78.765 ;
        RECT 41.460 78.375 41.660 78.405 ;
        RECT 41.780 78.155 41.950 78.225 ;
        RECT 41.080 77.985 41.950 78.155 ;
        RECT 41.440 77.895 41.950 77.985 ;
        RECT 39.990 77.430 40.295 77.560 ;
        RECT 40.740 77.450 41.270 77.815 ;
        RECT 39.610 76.835 39.875 77.295 ;
        RECT 40.045 77.005 40.295 77.430 ;
        RECT 41.440 77.280 41.610 77.895 ;
        RECT 40.505 77.110 41.610 77.280 ;
        RECT 41.780 76.835 41.950 77.635 ;
        RECT 42.120 77.335 42.290 78.405 ;
        RECT 42.460 77.505 42.650 78.225 ;
        RECT 42.820 77.475 43.140 78.435 ;
        RECT 43.310 78.475 43.480 78.935 ;
        RECT 43.755 78.855 43.965 79.385 ;
        RECT 44.225 78.645 44.555 79.170 ;
        RECT 44.725 78.775 44.895 79.385 ;
        RECT 45.065 78.730 45.395 79.165 ;
        RECT 46.125 78.730 46.455 79.165 ;
        RECT 46.625 78.775 46.795 79.385 ;
        RECT 45.065 78.645 45.445 78.730 ;
        RECT 44.355 78.475 44.555 78.645 ;
        RECT 45.220 78.605 45.445 78.645 ;
        RECT 43.310 78.145 44.185 78.475 ;
        RECT 44.355 78.145 45.105 78.475 ;
        RECT 42.120 77.005 42.370 77.335 ;
        RECT 43.310 77.305 43.480 78.145 ;
        RECT 44.355 77.940 44.545 78.145 ;
        RECT 45.275 78.025 45.445 78.605 ;
        RECT 45.230 77.975 45.445 78.025 ;
        RECT 43.650 77.565 44.545 77.940 ;
        RECT 45.055 77.895 45.445 77.975 ;
        RECT 46.075 78.645 46.455 78.730 ;
        RECT 46.965 78.645 47.295 79.170 ;
        RECT 47.555 78.855 47.765 79.385 ;
        RECT 48.040 78.935 48.825 79.105 ;
        RECT 48.995 78.935 49.400 79.105 ;
        RECT 46.075 78.605 46.300 78.645 ;
        RECT 46.075 78.025 46.245 78.605 ;
        RECT 46.965 78.475 47.165 78.645 ;
        RECT 48.040 78.475 48.210 78.935 ;
        RECT 46.415 78.145 47.165 78.475 ;
        RECT 47.335 78.145 48.210 78.475 ;
        RECT 46.075 77.975 46.290 78.025 ;
        RECT 46.075 77.895 46.465 77.975 ;
        RECT 42.595 77.135 43.480 77.305 ;
        RECT 43.660 76.835 43.975 77.335 ;
        RECT 44.205 77.005 44.545 77.565 ;
        RECT 44.715 76.835 44.885 77.845 ;
        RECT 45.055 77.050 45.385 77.895 ;
        RECT 46.135 77.050 46.465 77.895 ;
        RECT 46.975 77.940 47.165 78.145 ;
        RECT 46.635 76.835 46.805 77.845 ;
        RECT 46.975 77.565 47.870 77.940 ;
        RECT 46.975 77.005 47.315 77.565 ;
        RECT 47.545 76.835 47.860 77.335 ;
        RECT 48.040 77.305 48.210 78.145 ;
        RECT 48.380 78.435 48.845 78.765 ;
        RECT 49.230 78.705 49.400 78.935 ;
        RECT 49.580 78.885 49.950 79.385 ;
        RECT 50.270 78.935 50.945 79.105 ;
        RECT 51.140 78.935 51.475 79.105 ;
        RECT 48.380 77.475 48.700 78.435 ;
        RECT 49.230 78.405 50.060 78.705 ;
        RECT 48.870 77.505 49.060 78.225 ;
        RECT 49.230 77.335 49.400 78.405 ;
        RECT 49.860 78.375 50.060 78.405 ;
        RECT 49.570 78.155 49.740 78.225 ;
        RECT 50.270 78.155 50.440 78.935 ;
        RECT 51.305 78.795 51.475 78.935 ;
        RECT 51.645 78.925 51.895 79.385 ;
        RECT 49.570 77.985 50.440 78.155 ;
        RECT 50.610 78.515 51.135 78.735 ;
        RECT 51.305 78.665 51.530 78.795 ;
        RECT 49.570 77.895 50.080 77.985 ;
        RECT 48.040 77.135 48.925 77.305 ;
        RECT 49.150 77.005 49.400 77.335 ;
        RECT 49.570 76.835 49.740 77.635 ;
        RECT 49.910 77.280 50.080 77.895 ;
        RECT 50.610 77.815 50.780 78.515 ;
        RECT 50.250 77.450 50.780 77.815 ;
        RECT 50.950 77.750 51.190 78.345 ;
        RECT 51.360 77.560 51.530 78.665 ;
        RECT 51.700 77.805 51.980 78.755 ;
        RECT 51.225 77.430 51.530 77.560 ;
        RECT 49.910 77.110 51.015 77.280 ;
        RECT 51.225 77.005 51.475 77.430 ;
        RECT 51.645 76.835 51.910 77.295 ;
        RECT 52.150 77.005 52.335 79.125 ;
        RECT 52.505 79.005 52.835 79.385 ;
        RECT 53.005 78.835 53.175 79.125 ;
        RECT 52.510 78.665 53.175 78.835 ;
        RECT 52.510 77.675 52.740 78.665 ;
        RECT 53.435 78.615 56.025 79.385 ;
        RECT 56.245 78.730 56.575 79.165 ;
        RECT 56.745 78.775 56.915 79.385 ;
        RECT 56.195 78.645 56.575 78.730 ;
        RECT 57.085 78.645 57.415 79.170 ;
        RECT 57.675 78.855 57.885 79.385 ;
        RECT 58.160 78.935 58.945 79.105 ;
        RECT 59.115 78.935 59.520 79.105 ;
        RECT 52.910 77.845 53.260 78.495 ;
        RECT 53.435 78.095 54.645 78.615 ;
        RECT 56.195 78.605 56.420 78.645 ;
        RECT 54.815 77.925 56.025 78.445 ;
        RECT 52.510 77.505 53.175 77.675 ;
        RECT 52.505 76.835 52.835 77.335 ;
        RECT 53.005 77.005 53.175 77.505 ;
        RECT 53.435 76.835 56.025 77.925 ;
        RECT 56.195 78.025 56.365 78.605 ;
        RECT 57.085 78.475 57.285 78.645 ;
        RECT 58.160 78.475 58.330 78.935 ;
        RECT 56.535 78.145 57.285 78.475 ;
        RECT 57.455 78.145 58.330 78.475 ;
        RECT 56.195 77.975 56.410 78.025 ;
        RECT 56.195 77.895 56.585 77.975 ;
        RECT 56.255 77.050 56.585 77.895 ;
        RECT 57.095 77.940 57.285 78.145 ;
        RECT 56.755 76.835 56.925 77.845 ;
        RECT 57.095 77.565 57.990 77.940 ;
        RECT 57.095 77.005 57.435 77.565 ;
        RECT 57.665 76.835 57.980 77.335 ;
        RECT 58.160 77.305 58.330 78.145 ;
        RECT 58.500 78.435 58.965 78.765 ;
        RECT 59.350 78.705 59.520 78.935 ;
        RECT 59.700 78.885 60.070 79.385 ;
        RECT 60.390 78.935 61.065 79.105 ;
        RECT 61.260 78.935 61.595 79.105 ;
        RECT 58.500 77.475 58.820 78.435 ;
        RECT 59.350 78.405 60.180 78.705 ;
        RECT 58.990 77.505 59.180 78.225 ;
        RECT 59.350 77.335 59.520 78.405 ;
        RECT 59.980 78.375 60.180 78.405 ;
        RECT 59.690 78.155 59.860 78.225 ;
        RECT 60.390 78.155 60.560 78.935 ;
        RECT 61.425 78.795 61.595 78.935 ;
        RECT 61.765 78.925 62.015 79.385 ;
        RECT 59.690 77.985 60.560 78.155 ;
        RECT 60.730 78.515 61.255 78.735 ;
        RECT 61.425 78.665 61.650 78.795 ;
        RECT 59.690 77.895 60.200 77.985 ;
        RECT 58.160 77.135 59.045 77.305 ;
        RECT 59.270 77.005 59.520 77.335 ;
        RECT 59.690 76.835 59.860 77.635 ;
        RECT 60.030 77.280 60.200 77.895 ;
        RECT 60.730 77.815 60.900 78.515 ;
        RECT 60.370 77.450 60.900 77.815 ;
        RECT 61.070 77.750 61.310 78.345 ;
        RECT 61.480 77.560 61.650 78.665 ;
        RECT 61.820 77.805 62.100 78.755 ;
        RECT 61.345 77.430 61.650 77.560 ;
        RECT 60.030 77.110 61.135 77.280 ;
        RECT 61.345 77.005 61.595 77.430 ;
        RECT 61.765 76.835 62.030 77.295 ;
        RECT 62.270 77.005 62.455 79.125 ;
        RECT 62.625 79.005 62.955 79.385 ;
        RECT 63.125 78.835 63.295 79.125 ;
        RECT 62.630 78.665 63.295 78.835 ;
        RECT 62.630 77.675 62.860 78.665 ;
        RECT 63.555 78.660 63.845 79.385 ;
        RECT 64.015 78.645 64.455 79.205 ;
        RECT 64.625 78.645 65.075 79.385 ;
        RECT 65.245 78.815 65.415 79.215 ;
        RECT 65.585 78.985 66.005 79.385 ;
        RECT 66.175 78.815 66.405 79.215 ;
        RECT 65.245 78.645 66.405 78.815 ;
        RECT 66.575 78.645 67.065 79.215 ;
        RECT 63.030 77.845 63.380 78.495 ;
        RECT 62.630 77.505 63.295 77.675 ;
        RECT 62.625 76.835 62.955 77.335 ;
        RECT 63.125 77.005 63.295 77.505 ;
        RECT 63.555 76.835 63.845 78.000 ;
        RECT 64.015 77.635 64.325 78.645 ;
        RECT 64.495 78.025 64.665 78.475 ;
        RECT 64.835 78.195 65.225 78.475 ;
        RECT 65.410 78.145 65.655 78.475 ;
        RECT 64.495 77.855 65.285 78.025 ;
        RECT 64.015 77.005 64.455 77.635 ;
        RECT 64.630 76.835 64.945 77.685 ;
        RECT 65.115 77.175 65.285 77.855 ;
        RECT 65.455 77.345 65.655 78.145 ;
        RECT 65.855 77.345 66.105 78.475 ;
        RECT 66.320 78.145 66.725 78.475 ;
        RECT 66.895 77.975 67.065 78.645 ;
        RECT 66.295 77.805 67.065 77.975 ;
        RECT 67.245 78.660 67.575 79.170 ;
        RECT 67.745 78.985 68.075 79.385 ;
        RECT 69.125 78.815 69.455 79.155 ;
        RECT 69.625 78.985 69.955 79.385 ;
        RECT 67.245 78.025 67.435 78.660 ;
        RECT 67.745 78.645 70.110 78.815 ;
        RECT 71.395 78.655 71.685 79.385 ;
        RECT 67.745 78.475 67.915 78.645 ;
        RECT 67.605 78.145 67.915 78.475 ;
        RECT 68.085 78.145 68.390 78.475 ;
        RECT 67.245 77.895 67.465 78.025 ;
        RECT 66.295 77.175 66.545 77.805 ;
        RECT 65.115 77.005 66.545 77.175 ;
        RECT 66.725 76.835 67.055 77.635 ;
        RECT 67.245 77.045 67.575 77.895 ;
        RECT 67.745 76.835 67.995 77.975 ;
        RECT 68.175 77.815 68.390 78.145 ;
        RECT 68.565 77.815 68.850 78.475 ;
        RECT 69.045 77.815 69.310 78.475 ;
        RECT 69.525 77.815 69.770 78.475 ;
        RECT 69.940 77.645 70.110 78.645 ;
        RECT 71.385 78.145 71.685 78.475 ;
        RECT 71.865 78.455 72.095 79.095 ;
        RECT 72.275 78.835 72.585 79.205 ;
        RECT 72.765 79.015 73.435 79.385 ;
        RECT 72.275 78.635 73.505 78.835 ;
        RECT 71.865 78.145 72.390 78.455 ;
        RECT 72.570 78.145 73.035 78.455 ;
        RECT 73.215 77.965 73.505 78.635 ;
        RECT 68.185 77.475 69.475 77.645 ;
        RECT 68.185 77.055 68.435 77.475 ;
        RECT 68.665 76.835 68.995 77.305 ;
        RECT 69.225 77.055 69.475 77.475 ;
        RECT 69.655 77.475 70.110 77.645 ;
        RECT 71.395 77.725 72.555 77.965 ;
        RECT 69.655 77.045 69.985 77.475 ;
        RECT 71.395 77.015 71.655 77.725 ;
        RECT 71.825 76.835 72.155 77.545 ;
        RECT 72.325 77.015 72.555 77.725 ;
        RECT 72.735 77.745 73.505 77.965 ;
        RECT 72.735 77.015 73.005 77.745 ;
        RECT 73.185 76.835 73.525 77.565 ;
        RECT 73.695 77.015 73.955 79.205 ;
        RECT 74.155 78.655 74.445 79.385 ;
        RECT 74.145 78.145 74.445 78.475 ;
        RECT 74.625 78.455 74.855 79.095 ;
        RECT 75.035 78.835 75.345 79.205 ;
        RECT 75.525 79.015 76.195 79.385 ;
        RECT 75.035 78.635 76.265 78.835 ;
        RECT 74.625 78.145 75.150 78.455 ;
        RECT 75.330 78.145 75.795 78.455 ;
        RECT 75.975 77.965 76.265 78.635 ;
        RECT 74.155 77.725 75.315 77.965 ;
        RECT 74.155 77.015 74.415 77.725 ;
        RECT 74.585 76.835 74.915 77.545 ;
        RECT 75.085 77.015 75.315 77.725 ;
        RECT 75.495 77.745 76.265 77.965 ;
        RECT 75.495 77.015 75.765 77.745 ;
        RECT 75.945 76.835 76.285 77.565 ;
        RECT 76.455 77.015 76.715 79.205 ;
        RECT 76.895 78.615 80.405 79.385 ;
        RECT 80.575 78.635 81.785 79.385 ;
        RECT 81.960 78.645 82.215 79.215 ;
        RECT 82.385 78.985 82.715 79.385 ;
        RECT 83.140 78.850 83.670 79.215 ;
        RECT 83.860 79.045 84.135 79.215 ;
        RECT 83.855 78.875 84.135 79.045 ;
        RECT 83.140 78.815 83.315 78.850 ;
        RECT 82.385 78.645 83.315 78.815 ;
        RECT 76.895 78.095 78.545 78.615 ;
        RECT 78.715 77.925 80.405 78.445 ;
        RECT 80.575 78.095 81.095 78.635 ;
        RECT 81.265 77.925 81.785 78.465 ;
        RECT 76.895 76.835 80.405 77.925 ;
        RECT 80.575 76.835 81.785 77.925 ;
        RECT 81.960 77.975 82.130 78.645 ;
        RECT 82.385 78.475 82.555 78.645 ;
        RECT 82.300 78.145 82.555 78.475 ;
        RECT 82.780 78.145 82.975 78.475 ;
        RECT 81.960 77.005 82.295 77.975 ;
        RECT 82.465 76.835 82.635 77.975 ;
        RECT 82.805 77.175 82.975 78.145 ;
        RECT 83.145 77.515 83.315 78.645 ;
        RECT 83.485 77.855 83.655 78.655 ;
        RECT 83.860 78.055 84.135 78.875 ;
        RECT 84.305 77.855 84.495 79.215 ;
        RECT 84.675 78.850 85.185 79.385 ;
        RECT 85.405 78.575 85.650 79.180 ;
        RECT 86.185 78.835 86.355 79.215 ;
        RECT 86.535 79.005 86.865 79.385 ;
        RECT 86.185 78.665 86.850 78.835 ;
        RECT 87.045 78.710 87.305 79.215 ;
        RECT 84.695 78.405 85.925 78.575 ;
        RECT 83.485 77.685 84.495 77.855 ;
        RECT 84.665 77.840 85.415 78.030 ;
        RECT 83.145 77.345 84.270 77.515 ;
        RECT 84.665 77.175 84.835 77.840 ;
        RECT 85.585 77.595 85.925 78.405 ;
        RECT 86.115 78.115 86.445 78.485 ;
        RECT 86.680 78.410 86.850 78.665 ;
        RECT 86.680 78.080 86.965 78.410 ;
        RECT 86.680 77.935 86.850 78.080 ;
        RECT 82.805 77.005 84.835 77.175 ;
        RECT 85.005 76.835 85.175 77.595 ;
        RECT 85.410 77.185 85.925 77.595 ;
        RECT 86.185 77.765 86.850 77.935 ;
        RECT 87.135 77.910 87.305 78.710 ;
        RECT 87.475 78.615 89.145 79.385 ;
        RECT 89.315 78.635 90.525 79.385 ;
        RECT 87.475 78.095 88.225 78.615 ;
        RECT 88.395 77.925 89.145 78.445 ;
        RECT 86.185 77.005 86.355 77.765 ;
        RECT 86.535 76.835 86.865 77.595 ;
        RECT 87.035 77.005 87.305 77.910 ;
        RECT 87.475 76.835 89.145 77.925 ;
        RECT 89.315 77.925 89.835 78.465 ;
        RECT 90.005 78.095 90.525 78.635 ;
        RECT 89.315 76.835 90.525 77.925 ;
        RECT 11.950 76.665 90.610 76.835 ;
        RECT 12.035 75.575 13.245 76.665 ;
        RECT 13.415 75.575 15.085 76.665 ;
        RECT 12.035 74.865 12.555 75.405 ;
        RECT 12.725 75.035 13.245 75.575 ;
        RECT 13.415 74.885 14.165 75.405 ;
        RECT 14.335 75.055 15.085 75.575 ;
        RECT 15.290 75.875 15.825 76.495 ;
        RECT 12.035 74.115 13.245 74.865 ;
        RECT 13.415 74.115 15.085 74.885 ;
        RECT 15.290 74.855 15.605 75.875 ;
        RECT 15.995 75.865 16.325 76.665 ;
        RECT 18.015 76.155 18.275 76.665 ;
        RECT 16.810 75.695 17.200 75.870 ;
        RECT 15.775 75.525 17.200 75.695 ;
        RECT 15.775 75.025 15.945 75.525 ;
        RECT 15.290 74.285 15.905 74.855 ;
        RECT 16.195 74.795 16.460 75.355 ;
        RECT 16.630 74.625 16.800 75.525 ;
        RECT 16.970 74.795 17.325 75.355 ;
        RECT 18.015 75.105 18.355 75.985 ;
        RECT 18.525 75.275 18.695 76.495 ;
        RECT 18.935 76.160 19.550 76.665 ;
        RECT 18.935 75.625 19.185 75.990 ;
        RECT 19.355 75.985 19.550 76.160 ;
        RECT 19.720 76.155 20.195 76.495 ;
        RECT 20.365 76.120 20.580 76.665 ;
        RECT 19.355 75.795 19.685 75.985 ;
        RECT 19.905 75.625 20.620 75.920 ;
        RECT 20.790 75.795 21.065 76.495 ;
        RECT 18.935 75.455 20.725 75.625 ;
        RECT 18.525 75.025 19.320 75.275 ;
        RECT 18.525 74.935 18.775 75.025 ;
        RECT 16.075 74.115 16.290 74.625 ;
        RECT 16.520 74.295 16.800 74.625 ;
        RECT 16.980 74.115 17.220 74.625 ;
        RECT 18.015 74.115 18.275 74.935 ;
        RECT 18.445 74.515 18.775 74.935 ;
        RECT 19.490 74.600 19.745 75.455 ;
        RECT 18.955 74.335 19.745 74.600 ;
        RECT 19.915 74.755 20.325 75.275 ;
        RECT 20.495 75.025 20.725 75.455 ;
        RECT 20.895 74.765 21.065 75.795 ;
        RECT 21.695 75.525 21.955 76.665 ;
        RECT 22.195 76.155 23.810 76.485 ;
        RECT 22.205 75.355 22.375 75.915 ;
        RECT 22.635 75.815 23.810 75.985 ;
        RECT 23.980 75.865 24.260 76.665 ;
        RECT 22.635 75.525 22.965 75.815 ;
        RECT 23.640 75.695 23.810 75.815 ;
        RECT 23.135 75.355 23.380 75.645 ;
        RECT 23.640 75.525 24.300 75.695 ;
        RECT 24.470 75.525 24.745 76.495 ;
        RECT 24.130 75.355 24.300 75.525 ;
        RECT 21.700 75.105 22.035 75.355 ;
        RECT 22.205 75.025 22.920 75.355 ;
        RECT 23.135 75.025 23.960 75.355 ;
        RECT 24.130 75.025 24.405 75.355 ;
        RECT 22.205 74.935 22.455 75.025 ;
        RECT 19.915 74.335 20.115 74.755 ;
        RECT 20.305 74.115 20.635 74.575 ;
        RECT 20.805 74.285 21.065 74.765 ;
        RECT 21.695 74.115 21.955 74.935 ;
        RECT 22.125 74.515 22.455 74.935 ;
        RECT 24.130 74.855 24.300 75.025 ;
        RECT 22.635 74.685 24.300 74.855 ;
        RECT 24.575 74.790 24.745 75.525 ;
        RECT 24.915 75.500 25.205 76.665 ;
        RECT 25.375 75.575 27.045 76.665 ;
        RECT 27.765 75.995 27.935 76.495 ;
        RECT 28.105 76.165 28.435 76.665 ;
        RECT 27.765 75.825 28.430 75.995 ;
        RECT 25.375 74.885 26.125 75.405 ;
        RECT 26.295 75.055 27.045 75.575 ;
        RECT 27.680 75.005 28.030 75.655 ;
        RECT 22.635 74.285 22.895 74.685 ;
        RECT 23.065 74.115 23.395 74.515 ;
        RECT 23.565 74.335 23.735 74.685 ;
        RECT 23.905 74.115 24.280 74.515 ;
        RECT 24.470 74.445 24.745 74.790 ;
        RECT 24.915 74.115 25.205 74.840 ;
        RECT 25.375 74.115 27.045 74.885 ;
        RECT 28.200 74.835 28.430 75.825 ;
        RECT 27.765 74.665 28.430 74.835 ;
        RECT 27.765 74.375 27.935 74.665 ;
        RECT 28.105 74.115 28.435 74.495 ;
        RECT 28.605 74.375 28.790 76.495 ;
        RECT 29.030 76.205 29.295 76.665 ;
        RECT 29.465 76.070 29.715 76.495 ;
        RECT 29.925 76.220 31.030 76.390 ;
        RECT 29.410 75.940 29.715 76.070 ;
        RECT 28.960 74.745 29.240 75.695 ;
        RECT 29.410 74.835 29.580 75.940 ;
        RECT 29.750 75.155 29.990 75.750 ;
        RECT 30.160 75.685 30.690 76.050 ;
        RECT 30.160 74.985 30.330 75.685 ;
        RECT 30.860 75.605 31.030 76.220 ;
        RECT 31.200 75.865 31.370 76.665 ;
        RECT 31.540 76.165 31.790 76.495 ;
        RECT 32.015 76.195 32.900 76.365 ;
        RECT 30.860 75.515 31.370 75.605 ;
        RECT 29.410 74.705 29.635 74.835 ;
        RECT 29.805 74.765 30.330 74.985 ;
        RECT 30.500 75.345 31.370 75.515 ;
        RECT 29.045 74.115 29.295 74.575 ;
        RECT 29.465 74.565 29.635 74.705 ;
        RECT 30.500 74.565 30.670 75.345 ;
        RECT 31.200 75.275 31.370 75.345 ;
        RECT 30.880 75.095 31.080 75.125 ;
        RECT 31.540 75.095 31.710 76.165 ;
        RECT 31.880 75.275 32.070 75.995 ;
        RECT 30.880 74.795 31.710 75.095 ;
        RECT 32.240 75.065 32.560 76.025 ;
        RECT 29.465 74.395 29.800 74.565 ;
        RECT 29.995 74.395 30.670 74.565 ;
        RECT 30.990 74.115 31.360 74.615 ;
        RECT 31.540 74.565 31.710 74.795 ;
        RECT 32.095 74.735 32.560 75.065 ;
        RECT 32.730 75.355 32.900 76.195 ;
        RECT 33.080 76.165 33.395 76.665 ;
        RECT 33.625 75.935 33.965 76.495 ;
        RECT 33.070 75.560 33.965 75.935 ;
        RECT 34.135 75.655 34.305 76.665 ;
        RECT 33.775 75.355 33.965 75.560 ;
        RECT 34.475 75.605 34.805 76.450 ;
        RECT 34.975 75.750 35.145 76.665 ;
        RECT 34.475 75.525 34.865 75.605 ;
        RECT 35.495 75.575 39.005 76.665 ;
        RECT 34.650 75.475 34.865 75.525 ;
        RECT 32.730 75.025 33.605 75.355 ;
        RECT 33.775 75.025 34.525 75.355 ;
        RECT 32.730 74.565 32.900 75.025 ;
        RECT 33.775 74.855 33.975 75.025 ;
        RECT 34.695 74.895 34.865 75.475 ;
        RECT 34.640 74.855 34.865 74.895 ;
        RECT 31.540 74.395 31.945 74.565 ;
        RECT 32.115 74.395 32.900 74.565 ;
        RECT 33.175 74.115 33.385 74.645 ;
        RECT 33.645 74.330 33.975 74.855 ;
        RECT 34.485 74.770 34.865 74.855 ;
        RECT 35.495 74.885 37.145 75.405 ;
        RECT 37.315 75.055 39.005 75.575 ;
        RECT 39.245 75.660 39.500 76.465 ;
        RECT 39.670 75.830 39.930 76.665 ;
        RECT 40.100 75.660 40.360 76.465 ;
        RECT 40.530 75.830 40.785 76.665 ;
        RECT 39.245 75.490 40.845 75.660 ;
        RECT 39.175 75.095 40.395 75.320 ;
        RECT 40.565 74.925 40.845 75.490 ;
        RECT 34.145 74.115 34.315 74.725 ;
        RECT 34.485 74.335 34.815 74.770 ;
        RECT 34.985 74.115 35.155 74.630 ;
        RECT 35.495 74.115 39.005 74.885 ;
        RECT 40.115 74.755 40.845 74.925 ;
        RECT 41.020 75.525 41.355 76.495 ;
        RECT 41.525 75.525 41.695 76.665 ;
        RECT 41.865 76.325 43.895 76.495 ;
        RECT 41.020 74.855 41.190 75.525 ;
        RECT 41.865 75.355 42.035 76.325 ;
        RECT 41.360 75.025 41.615 75.355 ;
        RECT 41.840 75.025 42.035 75.355 ;
        RECT 42.205 75.985 43.330 76.155 ;
        RECT 41.445 74.855 41.615 75.025 ;
        RECT 42.205 74.855 42.375 75.985 ;
        RECT 39.650 74.115 39.945 74.640 ;
        RECT 40.115 74.310 40.340 74.755 ;
        RECT 40.510 74.115 40.840 74.585 ;
        RECT 41.020 74.285 41.275 74.855 ;
        RECT 41.445 74.685 42.375 74.855 ;
        RECT 42.545 75.645 43.555 75.815 ;
        RECT 42.545 74.845 42.715 75.645 ;
        RECT 42.200 74.650 42.375 74.685 ;
        RECT 41.445 74.115 41.775 74.515 ;
        RECT 42.200 74.285 42.730 74.650 ;
        RECT 42.920 74.625 43.195 75.445 ;
        RECT 42.915 74.455 43.195 74.625 ;
        RECT 42.920 74.285 43.195 74.455 ;
        RECT 43.365 74.285 43.555 75.645 ;
        RECT 43.725 75.660 43.895 76.325 ;
        RECT 44.065 75.905 44.235 76.665 ;
        RECT 44.470 75.905 44.985 76.315 ;
        RECT 43.725 75.470 44.475 75.660 ;
        RECT 44.645 75.095 44.985 75.905 ;
        RECT 43.755 74.925 44.985 75.095 ;
        RECT 45.160 75.525 45.495 76.495 ;
        RECT 45.665 75.525 45.835 76.665 ;
        RECT 46.005 76.325 48.035 76.495 ;
        RECT 43.735 74.115 44.245 74.650 ;
        RECT 44.465 74.320 44.710 74.925 ;
        RECT 45.160 74.855 45.330 75.525 ;
        RECT 46.005 75.355 46.175 76.325 ;
        RECT 45.500 75.025 45.755 75.355 ;
        RECT 45.980 75.025 46.175 75.355 ;
        RECT 46.345 75.985 47.470 76.155 ;
        RECT 45.585 74.855 45.755 75.025 ;
        RECT 46.345 74.855 46.515 75.985 ;
        RECT 45.160 74.285 45.415 74.855 ;
        RECT 45.585 74.685 46.515 74.855 ;
        RECT 46.685 75.645 47.695 75.815 ;
        RECT 46.685 74.845 46.855 75.645 ;
        RECT 46.340 74.650 46.515 74.685 ;
        RECT 45.585 74.115 45.915 74.515 ;
        RECT 46.340 74.285 46.870 74.650 ;
        RECT 47.060 74.625 47.335 75.445 ;
        RECT 47.055 74.455 47.335 74.625 ;
        RECT 47.060 74.285 47.335 74.455 ;
        RECT 47.505 74.285 47.695 75.645 ;
        RECT 47.865 75.660 48.035 76.325 ;
        RECT 48.205 75.905 48.375 76.665 ;
        RECT 48.610 75.905 49.125 76.315 ;
        RECT 47.865 75.470 48.615 75.660 ;
        RECT 48.785 75.095 49.125 75.905 ;
        RECT 49.295 75.575 50.505 76.665 ;
        RECT 47.895 74.925 49.125 75.095 ;
        RECT 47.875 74.115 48.385 74.650 ;
        RECT 48.605 74.320 48.850 74.925 ;
        RECT 49.295 74.865 49.815 75.405 ;
        RECT 49.985 75.035 50.505 75.575 ;
        RECT 50.675 75.500 50.965 76.665 ;
        RECT 51.140 75.525 51.475 76.495 ;
        RECT 51.645 75.525 51.815 76.665 ;
        RECT 51.985 76.325 54.015 76.495 ;
        RECT 49.295 74.115 50.505 74.865 ;
        RECT 51.140 74.855 51.310 75.525 ;
        RECT 51.985 75.355 52.155 76.325 ;
        RECT 51.480 75.025 51.735 75.355 ;
        RECT 51.960 75.025 52.155 75.355 ;
        RECT 52.325 75.985 53.450 76.155 ;
        RECT 51.565 74.855 51.735 75.025 ;
        RECT 52.325 74.855 52.495 75.985 ;
        RECT 50.675 74.115 50.965 74.840 ;
        RECT 51.140 74.285 51.395 74.855 ;
        RECT 51.565 74.685 52.495 74.855 ;
        RECT 52.665 75.645 53.675 75.815 ;
        RECT 52.665 74.845 52.835 75.645 ;
        RECT 52.320 74.650 52.495 74.685 ;
        RECT 51.565 74.115 51.895 74.515 ;
        RECT 52.320 74.285 52.850 74.650 ;
        RECT 53.040 74.625 53.315 75.445 ;
        RECT 53.035 74.455 53.315 74.625 ;
        RECT 53.040 74.285 53.315 74.455 ;
        RECT 53.485 74.285 53.675 75.645 ;
        RECT 53.845 75.660 54.015 76.325 ;
        RECT 54.185 75.905 54.355 76.665 ;
        RECT 54.590 75.905 55.105 76.315 ;
        RECT 53.845 75.470 54.595 75.660 ;
        RECT 54.765 75.095 55.105 75.905 ;
        RECT 55.795 75.605 56.125 76.450 ;
        RECT 56.295 75.655 56.465 76.665 ;
        RECT 56.635 75.935 56.975 76.495 ;
        RECT 57.205 76.165 57.520 76.665 ;
        RECT 57.700 76.195 58.585 76.365 ;
        RECT 53.875 74.925 55.105 75.095 ;
        RECT 55.735 75.525 56.125 75.605 ;
        RECT 56.635 75.560 57.530 75.935 ;
        RECT 55.735 75.475 55.950 75.525 ;
        RECT 53.855 74.115 54.365 74.650 ;
        RECT 54.585 74.320 54.830 74.925 ;
        RECT 55.735 74.895 55.905 75.475 ;
        RECT 56.635 75.355 56.825 75.560 ;
        RECT 57.700 75.355 57.870 76.195 ;
        RECT 58.810 76.165 59.060 76.495 ;
        RECT 56.075 75.025 56.825 75.355 ;
        RECT 56.995 75.025 57.870 75.355 ;
        RECT 55.735 74.855 55.960 74.895 ;
        RECT 56.625 74.855 56.825 75.025 ;
        RECT 55.735 74.770 56.115 74.855 ;
        RECT 55.785 74.335 56.115 74.770 ;
        RECT 56.285 74.115 56.455 74.725 ;
        RECT 56.625 74.330 56.955 74.855 ;
        RECT 57.215 74.115 57.425 74.645 ;
        RECT 57.700 74.565 57.870 75.025 ;
        RECT 58.040 75.065 58.360 76.025 ;
        RECT 58.530 75.275 58.720 75.995 ;
        RECT 58.890 75.095 59.060 76.165 ;
        RECT 59.230 75.865 59.400 76.665 ;
        RECT 59.570 76.220 60.675 76.390 ;
        RECT 59.570 75.605 59.740 76.220 ;
        RECT 60.885 76.070 61.135 76.495 ;
        RECT 61.305 76.205 61.570 76.665 ;
        RECT 59.910 75.685 60.440 76.050 ;
        RECT 60.885 75.940 61.190 76.070 ;
        RECT 59.230 75.515 59.740 75.605 ;
        RECT 59.230 75.345 60.100 75.515 ;
        RECT 59.230 75.275 59.400 75.345 ;
        RECT 59.520 75.095 59.720 75.125 ;
        RECT 58.040 74.735 58.505 75.065 ;
        RECT 58.890 74.795 59.720 75.095 ;
        RECT 58.890 74.565 59.060 74.795 ;
        RECT 57.700 74.395 58.485 74.565 ;
        RECT 58.655 74.395 59.060 74.565 ;
        RECT 59.240 74.115 59.610 74.615 ;
        RECT 59.930 74.565 60.100 75.345 ;
        RECT 60.270 74.985 60.440 75.685 ;
        RECT 60.610 75.155 60.850 75.750 ;
        RECT 60.270 74.765 60.795 74.985 ;
        RECT 61.020 74.835 61.190 75.940 ;
        RECT 60.965 74.705 61.190 74.835 ;
        RECT 61.360 74.745 61.640 75.695 ;
        RECT 60.965 74.565 61.135 74.705 ;
        RECT 59.930 74.395 60.605 74.565 ;
        RECT 60.800 74.395 61.135 74.565 ;
        RECT 61.305 74.115 61.555 74.575 ;
        RECT 61.810 74.375 61.995 76.495 ;
        RECT 62.165 76.165 62.495 76.665 ;
        RECT 62.665 75.995 62.835 76.495 ;
        RECT 62.170 75.825 62.835 75.995 ;
        RECT 63.210 76.035 63.495 76.495 ;
        RECT 63.665 76.205 63.935 76.665 ;
        RECT 62.170 74.835 62.400 75.825 ;
        RECT 63.210 75.815 64.165 76.035 ;
        RECT 62.570 75.005 62.920 75.655 ;
        RECT 63.095 75.085 63.785 75.645 ;
        RECT 63.955 74.915 64.165 75.815 ;
        RECT 62.170 74.665 62.835 74.835 ;
        RECT 62.165 74.115 62.495 74.495 ;
        RECT 62.665 74.375 62.835 74.665 ;
        RECT 63.210 74.745 64.165 74.915 ;
        RECT 64.335 75.645 64.735 76.495 ;
        RECT 64.925 76.035 65.205 76.495 ;
        RECT 65.725 76.205 66.050 76.665 ;
        RECT 64.925 75.815 66.050 76.035 ;
        RECT 64.335 75.085 65.430 75.645 ;
        RECT 65.600 75.355 66.050 75.815 ;
        RECT 66.220 75.525 66.605 76.495 ;
        RECT 63.210 74.285 63.495 74.745 ;
        RECT 63.665 74.115 63.935 74.575 ;
        RECT 64.335 74.285 64.735 75.085 ;
        RECT 65.600 75.025 66.155 75.355 ;
        RECT 65.600 74.915 66.050 75.025 ;
        RECT 64.925 74.745 66.050 74.915 ;
        RECT 66.325 74.855 66.605 75.525 ;
        RECT 64.925 74.285 65.205 74.745 ;
        RECT 65.725 74.115 66.050 74.575 ;
        RECT 66.220 74.285 66.605 74.855 ;
        RECT 66.775 74.395 67.055 76.495 ;
        RECT 67.245 75.905 68.030 76.665 ;
        RECT 68.425 75.835 68.810 76.495 ;
        RECT 68.425 75.735 68.835 75.835 ;
        RECT 67.225 75.525 68.835 75.735 ;
        RECT 69.135 75.645 69.335 76.435 ;
        RECT 67.225 74.925 67.500 75.525 ;
        RECT 69.005 75.475 69.335 75.645 ;
        RECT 69.505 75.485 69.825 76.665 ;
        RECT 70.195 75.995 70.475 76.665 ;
        RECT 70.645 75.775 70.945 76.325 ;
        RECT 71.145 75.945 71.475 76.665 ;
        RECT 71.665 75.945 72.125 76.495 ;
        RECT 69.005 75.355 69.185 75.475 ;
        RECT 67.670 75.105 68.025 75.355 ;
        RECT 68.220 75.305 68.685 75.355 ;
        RECT 68.215 75.135 68.685 75.305 ;
        RECT 68.220 75.105 68.685 75.135 ;
        RECT 68.855 75.105 69.185 75.355 ;
        RECT 70.010 75.355 70.275 75.715 ;
        RECT 70.645 75.605 71.585 75.775 ;
        RECT 71.415 75.355 71.585 75.605 ;
        RECT 69.360 75.105 69.825 75.305 ;
        RECT 70.010 75.105 70.685 75.355 ;
        RECT 70.905 75.105 71.245 75.355 ;
        RECT 71.415 75.025 71.705 75.355 ;
        RECT 71.415 74.935 71.585 75.025 ;
        RECT 67.225 74.745 68.475 74.925 ;
        RECT 68.110 74.675 68.475 74.745 ;
        RECT 68.645 74.725 69.825 74.895 ;
        RECT 67.285 74.115 67.455 74.575 ;
        RECT 68.645 74.505 68.975 74.725 ;
        RECT 67.725 74.325 68.975 74.505 ;
        RECT 69.145 74.115 69.315 74.555 ;
        RECT 69.485 74.310 69.825 74.725 ;
        RECT 70.195 74.745 71.585 74.935 ;
        RECT 70.195 74.385 70.525 74.745 ;
        RECT 71.875 74.575 72.125 75.945 ;
        RECT 72.295 75.525 72.555 76.665 ;
        RECT 72.725 75.515 73.055 76.495 ;
        RECT 73.225 75.525 73.505 76.665 ;
        RECT 74.225 75.735 74.395 76.495 ;
        RECT 74.610 75.905 74.940 76.665 ;
        RECT 74.225 75.565 74.940 75.735 ;
        RECT 75.110 75.590 75.365 76.495 ;
        RECT 72.315 75.105 72.650 75.355 ;
        RECT 72.820 74.915 72.990 75.515 ;
        RECT 73.160 75.085 73.495 75.355 ;
        RECT 74.135 75.015 74.490 75.385 ;
        RECT 74.770 75.355 74.940 75.565 ;
        RECT 74.770 75.025 75.025 75.355 ;
        RECT 71.145 74.115 71.395 74.575 ;
        RECT 71.565 74.285 72.125 74.575 ;
        RECT 72.295 74.285 72.990 74.915 ;
        RECT 73.195 74.115 73.505 74.915 ;
        RECT 74.770 74.835 74.940 75.025 ;
        RECT 75.195 74.860 75.365 75.590 ;
        RECT 75.540 75.515 75.800 76.665 ;
        RECT 76.435 75.500 76.725 76.665 ;
        RECT 76.895 75.575 79.485 76.665 ;
        RECT 80.205 75.995 80.375 76.495 ;
        RECT 80.545 76.165 80.875 76.665 ;
        RECT 80.205 75.825 80.870 75.995 ;
        RECT 74.225 74.665 74.940 74.835 ;
        RECT 74.225 74.285 74.395 74.665 ;
        RECT 74.610 74.115 74.940 74.495 ;
        RECT 75.110 74.285 75.365 74.860 ;
        RECT 75.540 74.115 75.800 74.955 ;
        RECT 76.895 74.885 78.105 75.405 ;
        RECT 78.275 75.055 79.485 75.575 ;
        RECT 80.120 75.005 80.470 75.655 ;
        RECT 76.435 74.115 76.725 74.840 ;
        RECT 76.895 74.115 79.485 74.885 ;
        RECT 80.640 74.835 80.870 75.825 ;
        RECT 80.205 74.665 80.870 74.835 ;
        RECT 80.205 74.375 80.375 74.665 ;
        RECT 80.545 74.115 80.875 74.495 ;
        RECT 81.045 74.375 81.230 76.495 ;
        RECT 81.470 76.205 81.735 76.665 ;
        RECT 81.905 76.070 82.155 76.495 ;
        RECT 82.365 76.220 83.470 76.390 ;
        RECT 81.850 75.940 82.155 76.070 ;
        RECT 81.400 74.745 81.680 75.695 ;
        RECT 81.850 74.835 82.020 75.940 ;
        RECT 82.190 75.155 82.430 75.750 ;
        RECT 82.600 75.685 83.130 76.050 ;
        RECT 82.600 74.985 82.770 75.685 ;
        RECT 83.300 75.605 83.470 76.220 ;
        RECT 83.640 75.865 83.810 76.665 ;
        RECT 83.980 76.165 84.230 76.495 ;
        RECT 84.455 76.195 85.340 76.365 ;
        RECT 83.300 75.515 83.810 75.605 ;
        RECT 81.850 74.705 82.075 74.835 ;
        RECT 82.245 74.765 82.770 74.985 ;
        RECT 82.940 75.345 83.810 75.515 ;
        RECT 81.485 74.115 81.735 74.575 ;
        RECT 81.905 74.565 82.075 74.705 ;
        RECT 82.940 74.565 83.110 75.345 ;
        RECT 83.640 75.275 83.810 75.345 ;
        RECT 83.320 75.095 83.520 75.125 ;
        RECT 83.980 75.095 84.150 76.165 ;
        RECT 84.320 75.275 84.510 75.995 ;
        RECT 83.320 74.795 84.150 75.095 ;
        RECT 84.680 75.065 85.000 76.025 ;
        RECT 81.905 74.395 82.240 74.565 ;
        RECT 82.435 74.395 83.110 74.565 ;
        RECT 83.430 74.115 83.800 74.615 ;
        RECT 83.980 74.565 84.150 74.795 ;
        RECT 84.535 74.735 85.000 75.065 ;
        RECT 85.170 75.355 85.340 76.195 ;
        RECT 85.520 76.165 85.835 76.665 ;
        RECT 86.065 75.935 86.405 76.495 ;
        RECT 85.510 75.560 86.405 75.935 ;
        RECT 86.575 75.655 86.745 76.665 ;
        RECT 86.215 75.355 86.405 75.560 ;
        RECT 86.915 75.605 87.245 76.450 ;
        RECT 87.565 75.735 87.735 76.495 ;
        RECT 87.950 75.905 88.280 76.665 ;
        RECT 86.915 75.525 87.305 75.605 ;
        RECT 87.565 75.565 88.280 75.735 ;
        RECT 88.450 75.590 88.705 76.495 ;
        RECT 87.090 75.475 87.305 75.525 ;
        RECT 85.170 75.025 86.045 75.355 ;
        RECT 86.215 75.025 86.965 75.355 ;
        RECT 85.170 74.565 85.340 75.025 ;
        RECT 86.215 74.855 86.415 75.025 ;
        RECT 87.135 74.895 87.305 75.475 ;
        RECT 87.475 75.015 87.830 75.385 ;
        RECT 88.110 75.355 88.280 75.565 ;
        RECT 88.110 75.025 88.365 75.355 ;
        RECT 87.080 74.855 87.305 74.895 ;
        RECT 83.980 74.395 84.385 74.565 ;
        RECT 84.555 74.395 85.340 74.565 ;
        RECT 85.615 74.115 85.825 74.645 ;
        RECT 86.085 74.330 86.415 74.855 ;
        RECT 86.925 74.770 87.305 74.855 ;
        RECT 88.110 74.835 88.280 75.025 ;
        RECT 88.535 74.860 88.705 75.590 ;
        RECT 88.880 75.515 89.140 76.665 ;
        RECT 89.315 75.575 90.525 76.665 ;
        RECT 89.315 75.035 89.835 75.575 ;
        RECT 86.585 74.115 86.755 74.725 ;
        RECT 86.925 74.335 87.255 74.770 ;
        RECT 87.565 74.665 88.280 74.835 ;
        RECT 87.565 74.285 87.735 74.665 ;
        RECT 87.950 74.115 88.280 74.495 ;
        RECT 88.450 74.285 88.705 74.860 ;
        RECT 88.880 74.115 89.140 74.955 ;
        RECT 90.005 74.865 90.525 75.405 ;
        RECT 99.990 75.105 100.160 80.925 ;
        RECT 100.640 78.285 100.990 80.445 ;
        RECT 100.640 75.585 100.990 77.745 ;
        RECT 101.470 75.105 101.640 80.925 ;
        RECT 102.120 78.285 102.470 80.445 ;
        RECT 102.120 75.585 102.470 77.745 ;
        RECT 102.950 75.105 103.120 80.925 ;
        RECT 103.600 78.285 103.950 80.445 ;
        RECT 103.600 75.585 103.950 77.745 ;
        RECT 104.430 75.105 104.600 80.925 ;
        RECT 105.080 78.285 105.430 80.445 ;
        RECT 105.080 75.585 105.430 77.745 ;
        RECT 105.910 75.105 106.080 80.925 ;
        RECT 106.560 78.285 106.910 80.445 ;
        RECT 106.560 75.585 106.910 77.745 ;
        RECT 107.390 75.105 107.560 80.925 ;
        RECT 108.040 78.285 108.390 80.445 ;
        RECT 108.040 75.585 108.390 77.745 ;
        RECT 108.870 75.105 109.040 80.925 ;
        RECT 109.520 78.285 109.870 80.445 ;
        RECT 109.520 75.585 109.870 77.745 ;
        RECT 110.350 75.105 110.520 80.925 ;
        RECT 117.600 80.850 129.140 81.010 ;
        RECT 117.600 80.840 127.560 80.850 ;
        RECT 117.600 75.450 117.770 80.840 ;
        RECT 118.400 80.330 119.400 80.500 ;
        RECT 118.170 76.120 118.340 80.160 ;
        RECT 119.460 76.120 119.630 80.160 ;
        RECT 118.400 75.780 119.400 75.950 ;
        RECT 120.030 75.450 120.200 80.840 ;
        RECT 120.830 80.330 122.830 80.500 ;
        RECT 120.600 76.120 120.770 80.160 ;
        RECT 122.890 76.120 123.060 80.160 ;
        RECT 120.830 75.780 122.830 75.950 ;
        RECT 123.460 75.450 123.630 80.840 ;
        RECT 124.260 80.330 126.260 80.500 ;
        RECT 124.030 76.120 124.200 80.160 ;
        RECT 126.320 76.120 126.490 80.160 ;
        RECT 126.890 79.940 127.560 80.840 ;
        RECT 128.100 80.340 128.430 80.510 ;
        RECT 126.890 78.760 127.580 79.940 ;
        RECT 127.960 79.130 128.130 80.170 ;
        RECT 128.400 79.130 128.570 80.170 ;
        RECT 128.970 78.760 129.140 80.850 ;
        RECT 129.450 80.960 130.470 81.350 ;
        RECT 129.450 80.820 131.250 80.960 ;
        RECT 126.890 78.590 129.140 78.760 ;
        RECT 129.500 80.790 131.250 80.820 ;
        RECT 129.500 80.780 130.470 80.790 ;
        RECT 126.890 78.430 128.750 78.590 ;
        RECT 126.890 78.200 127.660 78.430 ;
        RECT 126.890 76.690 127.650 78.200 ;
        RECT 124.260 75.780 126.260 75.950 ;
        RECT 126.890 75.450 128.920 76.690 ;
        RECT 129.500 76.650 129.670 80.780 ;
        RECT 130.210 80.275 130.540 80.445 ;
        RECT 130.070 77.020 130.240 80.060 ;
        RECT 130.510 77.020 130.680 80.060 ;
        RECT 131.080 76.650 131.250 80.790 ;
        RECT 134.420 79.150 134.590 84.540 ;
        RECT 135.130 84.130 135.460 84.300 ;
        RECT 134.990 79.875 135.160 83.915 ;
        RECT 135.430 79.875 135.600 83.915 ;
        RECT 135.130 79.490 135.460 79.660 ;
        RECT 136.000 79.150 136.170 84.540 ;
        RECT 139.540 84.540 139.730 84.640 ;
        RECT 137.210 84.130 137.540 84.300 ;
        RECT 138.170 84.130 138.500 84.300 ;
        RECT 136.570 79.875 136.740 83.915 ;
        RECT 137.050 79.875 137.220 83.915 ;
        RECT 137.530 79.875 137.700 83.915 ;
        RECT 138.010 79.875 138.180 83.915 ;
        RECT 138.490 79.875 138.660 83.915 ;
        RECT 138.970 79.875 139.140 83.915 ;
        RECT 136.730 79.490 137.060 79.660 ;
        RECT 137.690 79.490 138.020 79.660 ;
        RECT 138.650 79.490 138.980 79.660 ;
        RECT 139.540 79.150 139.710 84.540 ;
        RECT 134.420 78.980 139.710 79.150 ;
        RECT 129.500 76.480 131.250 76.650 ;
        RECT 134.410 78.090 139.700 78.260 ;
        RECT 134.410 75.690 134.580 78.090 ;
        RECT 135.120 77.580 135.450 77.750 ;
        RECT 134.980 76.370 135.150 77.410 ;
        RECT 135.420 76.370 135.590 77.410 ;
        RECT 135.120 76.030 135.450 76.200 ;
        RECT 135.990 75.690 136.160 78.090 ;
        RECT 137.200 77.580 137.530 77.750 ;
        RECT 138.160 77.580 138.490 77.750 ;
        RECT 136.560 76.370 136.730 77.410 ;
        RECT 137.040 76.370 137.210 77.410 ;
        RECT 137.520 76.370 137.690 77.410 ;
        RECT 138.000 76.370 138.170 77.410 ;
        RECT 138.480 76.370 138.650 77.410 ;
        RECT 138.960 76.370 139.130 77.410 ;
        RECT 136.720 76.030 137.050 76.200 ;
        RECT 137.680 76.030 138.010 76.200 ;
        RECT 138.640 76.030 138.970 76.200 ;
        RECT 139.530 75.690 139.700 78.090 ;
        RECT 134.410 75.520 139.700 75.690 ;
        RECT 117.600 75.270 128.920 75.450 ;
        RECT 99.990 74.935 110.520 75.105 ;
        RECT 89.315 74.115 90.525 74.865 ;
        RECT 117.610 74.780 128.920 75.270 ;
        RECT 127.000 74.770 128.920 74.780 ;
        RECT 134.420 74.690 139.700 75.520 ;
        RECT 11.950 73.945 90.610 74.115 ;
        RECT 12.035 73.195 13.245 73.945 ;
        RECT 13.880 73.205 14.135 73.775 ;
        RECT 14.305 73.545 14.635 73.945 ;
        RECT 15.060 73.410 15.590 73.775 ;
        RECT 15.060 73.375 15.235 73.410 ;
        RECT 14.305 73.205 15.235 73.375 ;
        RECT 12.035 72.655 12.555 73.195 ;
        RECT 12.725 72.485 13.245 73.025 ;
        RECT 12.035 71.395 13.245 72.485 ;
        RECT 13.880 72.535 14.050 73.205 ;
        RECT 14.305 73.035 14.475 73.205 ;
        RECT 14.220 72.705 14.475 73.035 ;
        RECT 14.700 72.705 14.895 73.035 ;
        RECT 13.880 71.565 14.215 72.535 ;
        RECT 14.385 71.395 14.555 72.535 ;
        RECT 14.725 71.735 14.895 72.705 ;
        RECT 15.065 72.075 15.235 73.205 ;
        RECT 15.405 72.415 15.575 73.215 ;
        RECT 15.780 72.925 16.055 73.775 ;
        RECT 15.775 72.755 16.055 72.925 ;
        RECT 15.780 72.615 16.055 72.755 ;
        RECT 16.225 72.415 16.415 73.775 ;
        RECT 16.595 73.410 17.105 73.945 ;
        RECT 17.325 73.135 17.570 73.740 ;
        RECT 18.020 73.205 18.275 73.775 ;
        RECT 18.445 73.545 18.775 73.945 ;
        RECT 19.200 73.410 19.730 73.775 ;
        RECT 19.200 73.375 19.375 73.410 ;
        RECT 18.445 73.205 19.375 73.375 ;
        RECT 16.615 72.965 17.845 73.135 ;
        RECT 15.405 72.245 16.415 72.415 ;
        RECT 16.585 72.400 17.335 72.590 ;
        RECT 15.065 71.905 16.190 72.075 ;
        RECT 16.585 71.735 16.755 72.400 ;
        RECT 17.505 72.155 17.845 72.965 ;
        RECT 14.725 71.565 16.755 71.735 ;
        RECT 16.925 71.395 17.095 72.155 ;
        RECT 17.330 71.745 17.845 72.155 ;
        RECT 18.020 72.535 18.190 73.205 ;
        RECT 18.445 73.035 18.615 73.205 ;
        RECT 18.360 72.705 18.615 73.035 ;
        RECT 18.840 72.705 19.035 73.035 ;
        RECT 18.020 71.565 18.355 72.535 ;
        RECT 18.525 71.395 18.695 72.535 ;
        RECT 18.865 71.735 19.035 72.705 ;
        RECT 19.205 72.075 19.375 73.205 ;
        RECT 19.545 72.415 19.715 73.215 ;
        RECT 19.920 72.925 20.195 73.775 ;
        RECT 19.915 72.755 20.195 72.925 ;
        RECT 19.920 72.615 20.195 72.755 ;
        RECT 20.365 72.415 20.555 73.775 ;
        RECT 20.735 73.410 21.245 73.945 ;
        RECT 21.465 73.135 21.710 73.740 ;
        RECT 23.350 73.135 23.595 73.740 ;
        RECT 23.815 73.410 24.325 73.945 ;
        RECT 20.755 72.965 21.985 73.135 ;
        RECT 19.545 72.245 20.555 72.415 ;
        RECT 20.725 72.400 21.475 72.590 ;
        RECT 19.205 71.905 20.330 72.075 ;
        RECT 20.725 71.735 20.895 72.400 ;
        RECT 21.645 72.155 21.985 72.965 ;
        RECT 18.865 71.565 20.895 71.735 ;
        RECT 21.065 71.395 21.235 72.155 ;
        RECT 21.470 71.745 21.985 72.155 ;
        RECT 23.075 72.965 24.305 73.135 ;
        RECT 23.075 72.155 23.415 72.965 ;
        RECT 23.585 72.400 24.335 72.590 ;
        RECT 23.075 71.745 23.590 72.155 ;
        RECT 23.825 71.395 23.995 72.155 ;
        RECT 24.165 71.735 24.335 72.400 ;
        RECT 24.505 72.415 24.695 73.775 ;
        RECT 24.865 73.605 25.140 73.775 ;
        RECT 24.865 73.435 25.145 73.605 ;
        RECT 24.865 72.615 25.140 73.435 ;
        RECT 25.330 73.410 25.860 73.775 ;
        RECT 26.285 73.545 26.615 73.945 ;
        RECT 25.685 73.375 25.860 73.410 ;
        RECT 25.345 72.415 25.515 73.215 ;
        RECT 24.505 72.245 25.515 72.415 ;
        RECT 25.685 73.205 26.615 73.375 ;
        RECT 26.785 73.205 27.040 73.775 ;
        RECT 27.275 73.485 27.520 73.945 ;
        RECT 25.685 72.075 25.855 73.205 ;
        RECT 26.445 73.035 26.615 73.205 ;
        RECT 24.730 71.905 25.855 72.075 ;
        RECT 26.025 72.705 26.220 73.035 ;
        RECT 26.445 72.705 26.700 73.035 ;
        RECT 26.025 71.735 26.195 72.705 ;
        RECT 26.870 72.535 27.040 73.205 ;
        RECT 27.215 72.705 27.530 73.315 ;
        RECT 27.700 72.955 27.950 73.765 ;
        RECT 28.120 73.420 28.380 73.945 ;
        RECT 28.550 73.295 28.810 73.750 ;
        RECT 28.980 73.465 29.240 73.945 ;
        RECT 29.410 73.295 29.670 73.750 ;
        RECT 29.840 73.465 30.100 73.945 ;
        RECT 30.270 73.295 30.530 73.750 ;
        RECT 30.700 73.465 30.960 73.945 ;
        RECT 31.130 73.295 31.390 73.750 ;
        RECT 31.560 73.465 31.860 73.945 ;
        RECT 32.275 73.400 37.620 73.945 ;
        RECT 28.550 73.125 31.860 73.295 ;
        RECT 27.700 72.705 30.720 72.955 ;
        RECT 24.165 71.565 26.195 71.735 ;
        RECT 26.365 71.395 26.535 72.535 ;
        RECT 26.705 71.565 27.040 72.535 ;
        RECT 27.225 71.395 27.520 72.505 ;
        RECT 27.700 71.570 27.950 72.705 ;
        RECT 30.890 72.535 31.860 73.125 ;
        RECT 33.860 72.570 34.200 73.400 ;
        RECT 37.795 73.220 38.085 73.945 ;
        RECT 39.235 73.485 39.480 73.945 ;
        RECT 28.120 71.395 28.380 72.505 ;
        RECT 28.550 72.295 31.860 72.535 ;
        RECT 28.550 71.570 28.810 72.295 ;
        RECT 28.980 71.395 29.240 72.125 ;
        RECT 29.410 71.570 29.670 72.295 ;
        RECT 29.840 71.395 30.100 72.125 ;
        RECT 30.270 71.570 30.530 72.295 ;
        RECT 30.700 71.395 30.960 72.125 ;
        RECT 31.130 71.570 31.390 72.295 ;
        RECT 31.560 71.395 31.855 72.125 ;
        RECT 35.680 71.830 36.030 73.080 ;
        RECT 39.175 72.705 39.490 73.315 ;
        RECT 39.660 72.955 39.910 73.765 ;
        RECT 40.080 73.420 40.340 73.945 ;
        RECT 40.510 73.295 40.770 73.750 ;
        RECT 40.940 73.465 41.200 73.945 ;
        RECT 41.370 73.295 41.630 73.750 ;
        RECT 41.800 73.465 42.060 73.945 ;
        RECT 42.230 73.295 42.490 73.750 ;
        RECT 42.660 73.465 42.920 73.945 ;
        RECT 43.090 73.295 43.350 73.750 ;
        RECT 43.520 73.465 43.820 73.945 ;
        RECT 40.510 73.125 43.820 73.295 ;
        RECT 39.660 72.705 42.680 72.955 ;
        RECT 32.275 71.395 37.620 71.830 ;
        RECT 37.795 71.395 38.085 72.560 ;
        RECT 39.185 71.395 39.480 72.505 ;
        RECT 39.660 71.570 39.910 72.705 ;
        RECT 42.850 72.535 43.820 73.125 ;
        RECT 44.235 73.175 46.825 73.945 ;
        RECT 47.085 73.395 47.255 73.685 ;
        RECT 47.425 73.565 47.755 73.945 ;
        RECT 47.085 73.225 47.750 73.395 ;
        RECT 44.235 72.655 45.445 73.175 ;
        RECT 40.080 71.395 40.340 72.505 ;
        RECT 40.510 72.295 43.820 72.535 ;
        RECT 45.615 72.485 46.825 73.005 ;
        RECT 40.510 71.570 40.770 72.295 ;
        RECT 40.940 71.395 41.200 72.125 ;
        RECT 41.370 71.570 41.630 72.295 ;
        RECT 41.800 71.395 42.060 72.125 ;
        RECT 42.230 71.570 42.490 72.295 ;
        RECT 42.660 71.395 42.920 72.125 ;
        RECT 43.090 71.570 43.350 72.295 ;
        RECT 43.520 71.395 43.815 72.125 ;
        RECT 44.235 71.395 46.825 72.485 ;
        RECT 47.000 72.405 47.350 73.055 ;
        RECT 47.520 72.235 47.750 73.225 ;
        RECT 47.085 72.065 47.750 72.235 ;
        RECT 47.085 71.565 47.255 72.065 ;
        RECT 47.425 71.395 47.755 71.895 ;
        RECT 47.925 71.565 48.110 73.685 ;
        RECT 48.365 73.485 48.615 73.945 ;
        RECT 48.785 73.495 49.120 73.665 ;
        RECT 49.315 73.495 49.990 73.665 ;
        RECT 48.785 73.355 48.955 73.495 ;
        RECT 48.280 72.365 48.560 73.315 ;
        RECT 48.730 73.225 48.955 73.355 ;
        RECT 48.730 72.120 48.900 73.225 ;
        RECT 49.125 73.075 49.650 73.295 ;
        RECT 49.070 72.310 49.310 72.905 ;
        RECT 49.480 72.375 49.650 73.075 ;
        RECT 49.820 72.715 49.990 73.495 ;
        RECT 50.310 73.445 50.680 73.945 ;
        RECT 50.860 73.495 51.265 73.665 ;
        RECT 51.435 73.495 52.220 73.665 ;
        RECT 50.860 73.265 51.030 73.495 ;
        RECT 50.200 72.965 51.030 73.265 ;
        RECT 51.415 72.995 51.880 73.325 ;
        RECT 50.200 72.935 50.400 72.965 ;
        RECT 50.520 72.715 50.690 72.785 ;
        RECT 49.820 72.545 50.690 72.715 ;
        RECT 50.180 72.455 50.690 72.545 ;
        RECT 48.730 71.990 49.035 72.120 ;
        RECT 49.480 72.010 50.010 72.375 ;
        RECT 48.350 71.395 48.615 71.855 ;
        RECT 48.785 71.565 49.035 71.990 ;
        RECT 50.180 71.840 50.350 72.455 ;
        RECT 49.245 71.670 50.350 71.840 ;
        RECT 50.520 71.395 50.690 72.195 ;
        RECT 50.860 71.895 51.030 72.965 ;
        RECT 51.200 72.065 51.390 72.785 ;
        RECT 51.560 72.035 51.880 72.995 ;
        RECT 52.050 73.035 52.220 73.495 ;
        RECT 52.495 73.415 52.705 73.945 ;
        RECT 52.965 73.205 53.295 73.730 ;
        RECT 53.465 73.335 53.635 73.945 ;
        RECT 53.805 73.290 54.135 73.725 ;
        RECT 53.805 73.205 54.185 73.290 ;
        RECT 53.095 73.035 53.295 73.205 ;
        RECT 53.960 73.165 54.185 73.205 ;
        RECT 52.050 72.705 52.925 73.035 ;
        RECT 53.095 72.705 53.845 73.035 ;
        RECT 50.860 71.565 51.110 71.895 ;
        RECT 52.050 71.865 52.220 72.705 ;
        RECT 53.095 72.500 53.285 72.705 ;
        RECT 54.015 72.585 54.185 73.165 ;
        RECT 53.970 72.535 54.185 72.585 ;
        RECT 52.390 72.125 53.285 72.500 ;
        RECT 53.795 72.455 54.185 72.535 ;
        RECT 54.360 73.205 54.615 73.775 ;
        RECT 54.785 73.545 55.115 73.945 ;
        RECT 55.540 73.410 56.070 73.775 ;
        RECT 55.540 73.375 55.715 73.410 ;
        RECT 54.785 73.205 55.715 73.375 ;
        RECT 54.360 72.535 54.530 73.205 ;
        RECT 54.785 73.035 54.955 73.205 ;
        RECT 54.700 72.705 54.955 73.035 ;
        RECT 55.180 72.705 55.375 73.035 ;
        RECT 51.335 71.695 52.220 71.865 ;
        RECT 52.400 71.395 52.715 71.895 ;
        RECT 52.945 71.565 53.285 72.125 ;
        RECT 53.455 71.395 53.625 72.405 ;
        RECT 53.795 71.610 54.125 72.455 ;
        RECT 54.360 71.565 54.695 72.535 ;
        RECT 54.865 71.395 55.035 72.535 ;
        RECT 55.205 71.735 55.375 72.705 ;
        RECT 55.545 72.075 55.715 73.205 ;
        RECT 55.885 72.415 56.055 73.215 ;
        RECT 56.260 72.925 56.535 73.775 ;
        RECT 56.255 72.755 56.535 72.925 ;
        RECT 56.260 72.615 56.535 72.755 ;
        RECT 56.705 72.415 56.895 73.775 ;
        RECT 57.075 73.410 57.585 73.945 ;
        RECT 57.805 73.135 58.050 73.740 ;
        RECT 58.495 73.205 58.880 73.775 ;
        RECT 59.050 73.485 59.375 73.945 ;
        RECT 59.895 73.315 60.175 73.775 ;
        RECT 57.095 72.965 58.325 73.135 ;
        RECT 55.885 72.245 56.895 72.415 ;
        RECT 57.065 72.400 57.815 72.590 ;
        RECT 55.545 71.905 56.670 72.075 ;
        RECT 57.065 71.735 57.235 72.400 ;
        RECT 57.985 72.155 58.325 72.965 ;
        RECT 55.205 71.565 57.235 71.735 ;
        RECT 57.405 71.395 57.575 72.155 ;
        RECT 57.810 71.745 58.325 72.155 ;
        RECT 58.495 72.535 58.775 73.205 ;
        RECT 59.050 73.145 60.175 73.315 ;
        RECT 59.050 73.035 59.500 73.145 ;
        RECT 58.945 72.705 59.500 73.035 ;
        RECT 60.365 72.975 60.765 73.775 ;
        RECT 61.165 73.485 61.435 73.945 ;
        RECT 61.605 73.315 61.890 73.775 ;
        RECT 58.495 71.565 58.880 72.535 ;
        RECT 59.050 72.245 59.500 72.705 ;
        RECT 59.670 72.415 60.765 72.975 ;
        RECT 59.050 72.025 60.175 72.245 ;
        RECT 59.050 71.395 59.375 71.855 ;
        RECT 59.895 71.565 60.175 72.025 ;
        RECT 60.365 71.565 60.765 72.415 ;
        RECT 60.935 73.145 61.890 73.315 ;
        RECT 62.175 73.195 63.385 73.945 ;
        RECT 63.555 73.220 63.845 73.945 ;
        RECT 64.495 73.475 64.790 73.945 ;
        RECT 64.960 73.305 65.220 73.750 ;
        RECT 65.390 73.475 65.650 73.945 ;
        RECT 65.820 73.305 66.075 73.750 ;
        RECT 66.245 73.475 66.545 73.945 ;
        RECT 60.935 72.245 61.145 73.145 ;
        RECT 61.315 72.415 62.005 72.975 ;
        RECT 62.175 72.655 62.695 73.195 ;
        RECT 64.035 73.135 67.065 73.305 ;
        RECT 67.235 73.145 67.930 73.775 ;
        RECT 68.135 73.145 68.445 73.945 ;
        RECT 68.615 73.145 69.310 73.775 ;
        RECT 69.515 73.145 69.825 73.945 ;
        RECT 62.865 72.485 63.385 73.025 ;
        RECT 64.035 72.570 64.205 73.135 ;
        RECT 64.375 72.740 66.590 72.965 ;
        RECT 66.765 72.570 67.065 73.135 ;
        RECT 67.255 72.705 67.590 72.955 ;
        RECT 60.935 72.025 61.890 72.245 ;
        RECT 61.165 71.395 61.435 71.855 ;
        RECT 61.605 71.565 61.890 72.025 ;
        RECT 62.175 71.395 63.385 72.485 ;
        RECT 63.555 71.395 63.845 72.560 ;
        RECT 64.035 72.400 67.065 72.570 ;
        RECT 67.760 72.545 67.930 73.145 ;
        RECT 68.100 72.705 68.435 72.975 ;
        RECT 68.635 72.705 68.970 72.955 ;
        RECT 69.140 72.545 69.310 73.145 ;
        RECT 70.005 73.135 70.275 73.945 ;
        RECT 70.445 73.135 70.775 73.775 ;
        RECT 70.945 73.135 71.185 73.945 ;
        RECT 72.300 73.180 72.755 73.945 ;
        RECT 73.030 73.565 74.330 73.775 ;
        RECT 74.585 73.585 74.915 73.945 ;
        RECT 74.160 73.415 74.330 73.565 ;
        RECT 75.085 73.445 75.345 73.775 ;
        RECT 75.115 73.435 75.345 73.445 ;
        RECT 69.480 72.705 69.815 72.975 ;
        RECT 69.995 72.705 70.345 72.955 ;
        RECT 64.015 71.395 64.360 72.230 ;
        RECT 64.535 71.595 64.790 72.400 ;
        RECT 64.960 71.395 65.220 72.230 ;
        RECT 65.395 71.595 65.650 72.400 ;
        RECT 65.820 71.395 66.080 72.230 ;
        RECT 66.250 71.595 66.510 72.400 ;
        RECT 66.680 71.395 67.065 72.230 ;
        RECT 67.235 71.395 67.495 72.535 ;
        RECT 67.665 71.565 67.995 72.545 ;
        RECT 68.165 71.395 68.445 72.535 ;
        RECT 68.615 71.395 68.875 72.535 ;
        RECT 69.045 71.565 69.375 72.545 ;
        RECT 70.515 72.535 70.685 73.135 ;
        RECT 73.230 72.955 73.450 73.355 ;
        RECT 70.855 72.705 71.205 72.955 ;
        RECT 72.295 72.755 72.785 72.955 ;
        RECT 72.975 72.745 73.450 72.955 ;
        RECT 73.695 72.955 73.905 73.355 ;
        RECT 74.160 73.290 74.915 73.415 ;
        RECT 74.160 73.245 75.005 73.290 ;
        RECT 74.735 73.125 75.005 73.245 ;
        RECT 73.695 72.745 74.025 72.955 ;
        RECT 74.195 72.685 74.605 72.990 ;
        RECT 69.545 71.395 69.825 72.535 ;
        RECT 70.005 71.395 70.335 72.535 ;
        RECT 70.515 72.365 71.195 72.535 ;
        RECT 70.865 71.580 71.195 72.365 ;
        RECT 72.300 72.515 73.475 72.575 ;
        RECT 74.835 72.550 75.005 73.125 ;
        RECT 74.805 72.515 75.005 72.550 ;
        RECT 72.300 72.405 75.005 72.515 ;
        RECT 72.300 71.785 72.555 72.405 ;
        RECT 73.145 72.345 74.945 72.405 ;
        RECT 73.145 72.315 73.475 72.345 ;
        RECT 75.175 72.245 75.345 73.435 ;
        RECT 75.720 73.165 76.220 73.775 ;
        RECT 75.515 72.705 75.865 72.955 ;
        RECT 76.050 72.535 76.220 73.165 ;
        RECT 76.850 73.295 77.180 73.775 ;
        RECT 77.350 73.485 77.575 73.945 ;
        RECT 77.745 73.295 78.075 73.775 ;
        RECT 76.850 73.125 78.075 73.295 ;
        RECT 78.265 73.145 78.515 73.945 ;
        RECT 78.685 73.145 79.025 73.775 ;
        RECT 76.390 72.755 76.720 72.955 ;
        RECT 76.890 72.755 77.220 72.955 ;
        RECT 77.390 72.755 77.810 72.955 ;
        RECT 77.985 72.785 78.680 72.955 ;
        RECT 77.985 72.535 78.155 72.785 ;
        RECT 78.850 72.535 79.025 73.145 ;
        RECT 79.195 73.175 80.865 73.945 ;
        RECT 81.500 73.205 81.755 73.775 ;
        RECT 81.925 73.545 82.255 73.945 ;
        RECT 82.680 73.410 83.210 73.775 ;
        RECT 82.680 73.375 82.855 73.410 ;
        RECT 81.925 73.205 82.855 73.375 ;
        RECT 79.195 72.655 79.945 73.175 ;
        RECT 72.805 72.145 72.990 72.235 ;
        RECT 73.580 72.145 74.415 72.155 ;
        RECT 72.805 71.945 74.415 72.145 ;
        RECT 72.805 71.905 73.035 71.945 ;
        RECT 72.300 71.565 72.635 71.785 ;
        RECT 73.640 71.395 73.995 71.775 ;
        RECT 74.165 71.565 74.415 71.945 ;
        RECT 74.665 71.395 74.915 72.175 ;
        RECT 75.085 71.565 75.345 72.245 ;
        RECT 75.720 72.365 78.155 72.535 ;
        RECT 75.720 71.565 76.050 72.365 ;
        RECT 76.220 71.395 76.550 72.195 ;
        RECT 76.850 71.565 77.180 72.365 ;
        RECT 77.825 71.395 78.075 72.195 ;
        RECT 78.345 71.395 78.515 72.535 ;
        RECT 78.685 71.565 79.025 72.535 ;
        RECT 80.115 72.485 80.865 73.005 ;
        RECT 79.195 71.395 80.865 72.485 ;
        RECT 81.500 72.535 81.670 73.205 ;
        RECT 81.925 73.035 82.095 73.205 ;
        RECT 81.840 72.705 82.095 73.035 ;
        RECT 82.320 72.705 82.515 73.035 ;
        RECT 81.500 71.565 81.835 72.535 ;
        RECT 82.005 71.395 82.175 72.535 ;
        RECT 82.345 71.735 82.515 72.705 ;
        RECT 82.685 72.075 82.855 73.205 ;
        RECT 83.025 72.415 83.195 73.215 ;
        RECT 83.400 72.925 83.675 73.775 ;
        RECT 83.395 72.755 83.675 72.925 ;
        RECT 83.400 72.615 83.675 72.755 ;
        RECT 83.845 72.415 84.035 73.775 ;
        RECT 84.215 73.410 84.725 73.945 ;
        RECT 84.945 73.135 85.190 73.740 ;
        RECT 85.635 73.205 86.020 73.775 ;
        RECT 86.190 73.485 86.515 73.945 ;
        RECT 87.035 73.315 87.315 73.775 ;
        RECT 84.235 72.965 85.465 73.135 ;
        RECT 83.025 72.245 84.035 72.415 ;
        RECT 84.205 72.400 84.955 72.590 ;
        RECT 82.685 71.905 83.810 72.075 ;
        RECT 84.205 71.735 84.375 72.400 ;
        RECT 85.125 72.155 85.465 72.965 ;
        RECT 82.345 71.565 84.375 71.735 ;
        RECT 84.545 71.395 84.715 72.155 ;
        RECT 84.950 71.745 85.465 72.155 ;
        RECT 85.635 72.535 85.915 73.205 ;
        RECT 86.190 73.145 87.315 73.315 ;
        RECT 86.190 73.035 86.640 73.145 ;
        RECT 86.085 72.705 86.640 73.035 ;
        RECT 87.505 72.975 87.905 73.775 ;
        RECT 88.305 73.485 88.575 73.945 ;
        RECT 88.745 73.315 89.030 73.775 ;
        RECT 85.635 71.565 86.020 72.535 ;
        RECT 86.190 72.245 86.640 72.705 ;
        RECT 86.810 72.415 87.905 72.975 ;
        RECT 86.190 72.025 87.315 72.245 ;
        RECT 86.190 71.395 86.515 71.855 ;
        RECT 87.035 71.565 87.315 72.025 ;
        RECT 87.505 71.565 87.905 72.415 ;
        RECT 88.075 73.145 89.030 73.315 ;
        RECT 89.315 73.195 90.525 73.945 ;
        RECT 88.075 72.245 88.285 73.145 ;
        RECT 88.455 72.415 89.145 72.975 ;
        RECT 89.315 72.485 89.835 73.025 ;
        RECT 90.005 72.655 90.525 73.195 ;
        RECT 88.075 72.025 89.030 72.245 ;
        RECT 88.305 71.395 88.575 71.855 ;
        RECT 88.745 71.565 89.030 72.025 ;
        RECT 89.315 71.395 90.525 72.485 ;
        RECT 11.950 71.225 90.610 71.395 ;
        RECT 12.035 70.135 13.245 71.225 ;
        RECT 13.505 70.555 13.675 71.055 ;
        RECT 13.845 70.725 14.175 71.225 ;
        RECT 13.505 70.385 14.170 70.555 ;
        RECT 12.035 69.425 12.555 69.965 ;
        RECT 12.725 69.595 13.245 70.135 ;
        RECT 13.420 69.565 13.770 70.215 ;
        RECT 12.035 68.675 13.245 69.425 ;
        RECT 13.940 69.395 14.170 70.385 ;
        RECT 13.505 69.225 14.170 69.395 ;
        RECT 13.505 68.935 13.675 69.225 ;
        RECT 13.845 68.675 14.175 69.055 ;
        RECT 14.345 68.935 14.530 71.055 ;
        RECT 14.770 70.765 15.035 71.225 ;
        RECT 15.205 70.630 15.455 71.055 ;
        RECT 15.665 70.780 16.770 70.950 ;
        RECT 15.150 70.500 15.455 70.630 ;
        RECT 14.700 69.305 14.980 70.255 ;
        RECT 15.150 69.395 15.320 70.500 ;
        RECT 15.490 69.715 15.730 70.310 ;
        RECT 15.900 70.245 16.430 70.610 ;
        RECT 15.900 69.545 16.070 70.245 ;
        RECT 16.600 70.165 16.770 70.780 ;
        RECT 16.940 70.425 17.110 71.225 ;
        RECT 17.280 70.725 17.530 71.055 ;
        RECT 17.755 70.755 18.640 70.925 ;
        RECT 16.600 70.075 17.110 70.165 ;
        RECT 15.150 69.265 15.375 69.395 ;
        RECT 15.545 69.325 16.070 69.545 ;
        RECT 16.240 69.905 17.110 70.075 ;
        RECT 14.785 68.675 15.035 69.135 ;
        RECT 15.205 69.125 15.375 69.265 ;
        RECT 16.240 69.125 16.410 69.905 ;
        RECT 16.940 69.835 17.110 69.905 ;
        RECT 16.620 69.655 16.820 69.685 ;
        RECT 17.280 69.655 17.450 70.725 ;
        RECT 17.620 69.835 17.810 70.555 ;
        RECT 16.620 69.355 17.450 69.655 ;
        RECT 17.980 69.625 18.300 70.585 ;
        RECT 15.205 68.955 15.540 69.125 ;
        RECT 15.735 68.955 16.410 69.125 ;
        RECT 16.730 68.675 17.100 69.175 ;
        RECT 17.280 69.125 17.450 69.355 ;
        RECT 17.835 69.295 18.300 69.625 ;
        RECT 18.470 69.915 18.640 70.755 ;
        RECT 18.820 70.725 19.135 71.225 ;
        RECT 19.365 70.495 19.705 71.055 ;
        RECT 18.810 70.120 19.705 70.495 ;
        RECT 19.875 70.215 20.045 71.225 ;
        RECT 19.515 69.915 19.705 70.120 ;
        RECT 20.215 70.165 20.545 71.010 ;
        RECT 20.715 70.310 20.885 71.225 ;
        RECT 20.215 70.085 20.605 70.165 ;
        RECT 21.235 70.135 24.745 71.225 ;
        RECT 20.390 70.035 20.605 70.085 ;
        RECT 18.470 69.585 19.345 69.915 ;
        RECT 19.515 69.585 20.265 69.915 ;
        RECT 18.470 69.125 18.640 69.585 ;
        RECT 19.515 69.415 19.715 69.585 ;
        RECT 20.435 69.455 20.605 70.035 ;
        RECT 20.380 69.415 20.605 69.455 ;
        RECT 17.280 68.955 17.685 69.125 ;
        RECT 17.855 68.955 18.640 69.125 ;
        RECT 18.915 68.675 19.125 69.205 ;
        RECT 19.385 68.890 19.715 69.415 ;
        RECT 20.225 69.330 20.605 69.415 ;
        RECT 21.235 69.445 22.885 69.965 ;
        RECT 23.055 69.615 24.745 70.135 ;
        RECT 24.915 70.060 25.205 71.225 ;
        RECT 25.465 70.555 25.635 71.055 ;
        RECT 25.805 70.725 26.135 71.225 ;
        RECT 25.465 70.385 26.130 70.555 ;
        RECT 25.380 69.565 25.730 70.215 ;
        RECT 19.885 68.675 20.055 69.285 ;
        RECT 20.225 68.895 20.555 69.330 ;
        RECT 20.725 68.675 20.895 69.190 ;
        RECT 21.235 68.675 24.745 69.445 ;
        RECT 24.915 68.675 25.205 69.400 ;
        RECT 25.900 69.395 26.130 70.385 ;
        RECT 25.465 69.225 26.130 69.395 ;
        RECT 25.465 68.935 25.635 69.225 ;
        RECT 25.805 68.675 26.135 69.055 ;
        RECT 26.305 68.935 26.490 71.055 ;
        RECT 26.730 70.765 26.995 71.225 ;
        RECT 27.165 70.630 27.415 71.055 ;
        RECT 27.625 70.780 28.730 70.950 ;
        RECT 27.110 70.500 27.415 70.630 ;
        RECT 26.660 69.305 26.940 70.255 ;
        RECT 27.110 69.395 27.280 70.500 ;
        RECT 27.450 69.715 27.690 70.310 ;
        RECT 27.860 70.245 28.390 70.610 ;
        RECT 27.860 69.545 28.030 70.245 ;
        RECT 28.560 70.165 28.730 70.780 ;
        RECT 28.900 70.425 29.070 71.225 ;
        RECT 29.240 70.725 29.490 71.055 ;
        RECT 29.715 70.755 30.600 70.925 ;
        RECT 28.560 70.075 29.070 70.165 ;
        RECT 27.110 69.265 27.335 69.395 ;
        RECT 27.505 69.325 28.030 69.545 ;
        RECT 28.200 69.905 29.070 70.075 ;
        RECT 26.745 68.675 26.995 69.135 ;
        RECT 27.165 69.125 27.335 69.265 ;
        RECT 28.200 69.125 28.370 69.905 ;
        RECT 28.900 69.835 29.070 69.905 ;
        RECT 28.580 69.655 28.780 69.685 ;
        RECT 29.240 69.655 29.410 70.725 ;
        RECT 29.580 69.835 29.770 70.555 ;
        RECT 28.580 69.355 29.410 69.655 ;
        RECT 29.940 69.625 30.260 70.585 ;
        RECT 27.165 68.955 27.500 69.125 ;
        RECT 27.695 68.955 28.370 69.125 ;
        RECT 28.690 68.675 29.060 69.175 ;
        RECT 29.240 69.125 29.410 69.355 ;
        RECT 29.795 69.295 30.260 69.625 ;
        RECT 30.430 69.915 30.600 70.755 ;
        RECT 30.780 70.725 31.095 71.225 ;
        RECT 31.325 70.495 31.665 71.055 ;
        RECT 30.770 70.120 31.665 70.495 ;
        RECT 31.835 70.215 32.005 71.225 ;
        RECT 31.475 69.915 31.665 70.120 ;
        RECT 32.175 70.165 32.505 71.010 ;
        RECT 32.675 70.310 32.845 71.225 ;
        RECT 32.175 70.085 32.565 70.165 ;
        RECT 33.195 70.135 34.865 71.225 ;
        RECT 32.350 70.035 32.565 70.085 ;
        RECT 30.430 69.585 31.305 69.915 ;
        RECT 31.475 69.585 32.225 69.915 ;
        RECT 30.430 69.125 30.600 69.585 ;
        RECT 31.475 69.415 31.675 69.585 ;
        RECT 32.395 69.455 32.565 70.035 ;
        RECT 32.340 69.415 32.565 69.455 ;
        RECT 29.240 68.955 29.645 69.125 ;
        RECT 29.815 68.955 30.600 69.125 ;
        RECT 30.875 68.675 31.085 69.205 ;
        RECT 31.345 68.890 31.675 69.415 ;
        RECT 32.185 69.330 32.565 69.415 ;
        RECT 33.195 69.445 33.945 69.965 ;
        RECT 34.115 69.615 34.865 70.135 ;
        RECT 35.040 70.085 35.375 71.055 ;
        RECT 35.545 70.085 35.715 71.225 ;
        RECT 35.885 70.885 37.915 71.055 ;
        RECT 31.845 68.675 32.015 69.285 ;
        RECT 32.185 68.895 32.515 69.330 ;
        RECT 32.685 68.675 32.855 69.190 ;
        RECT 33.195 68.675 34.865 69.445 ;
        RECT 35.040 69.415 35.210 70.085 ;
        RECT 35.885 69.915 36.055 70.885 ;
        RECT 35.380 69.585 35.635 69.915 ;
        RECT 35.860 69.585 36.055 69.915 ;
        RECT 36.225 70.545 37.350 70.715 ;
        RECT 35.465 69.415 35.635 69.585 ;
        RECT 36.225 69.415 36.395 70.545 ;
        RECT 35.040 68.845 35.295 69.415 ;
        RECT 35.465 69.245 36.395 69.415 ;
        RECT 36.565 70.205 37.575 70.375 ;
        RECT 36.565 69.405 36.735 70.205 ;
        RECT 36.220 69.210 36.395 69.245 ;
        RECT 35.465 68.675 35.795 69.075 ;
        RECT 36.220 68.845 36.750 69.210 ;
        RECT 36.940 69.185 37.215 70.005 ;
        RECT 36.935 69.015 37.215 69.185 ;
        RECT 36.940 68.845 37.215 69.015 ;
        RECT 37.385 68.845 37.575 70.205 ;
        RECT 37.745 70.220 37.915 70.885 ;
        RECT 38.085 70.465 38.255 71.225 ;
        RECT 38.490 70.465 39.005 70.875 ;
        RECT 37.745 70.030 38.495 70.220 ;
        RECT 38.665 69.655 39.005 70.465 ;
        RECT 39.265 70.555 39.435 71.055 ;
        RECT 39.605 70.725 39.935 71.225 ;
        RECT 39.265 70.385 39.930 70.555 ;
        RECT 37.775 69.485 39.005 69.655 ;
        RECT 39.180 69.565 39.530 70.215 ;
        RECT 37.755 68.675 38.265 69.210 ;
        RECT 38.485 68.880 38.730 69.485 ;
        RECT 39.700 69.395 39.930 70.385 ;
        RECT 39.265 69.225 39.930 69.395 ;
        RECT 39.265 68.935 39.435 69.225 ;
        RECT 39.605 68.675 39.935 69.055 ;
        RECT 40.105 68.935 40.290 71.055 ;
        RECT 40.530 70.765 40.795 71.225 ;
        RECT 40.965 70.630 41.215 71.055 ;
        RECT 41.425 70.780 42.530 70.950 ;
        RECT 40.910 70.500 41.215 70.630 ;
        RECT 40.460 69.305 40.740 70.255 ;
        RECT 40.910 69.395 41.080 70.500 ;
        RECT 41.250 69.715 41.490 70.310 ;
        RECT 41.660 70.245 42.190 70.610 ;
        RECT 41.660 69.545 41.830 70.245 ;
        RECT 42.360 70.165 42.530 70.780 ;
        RECT 42.700 70.425 42.870 71.225 ;
        RECT 43.040 70.725 43.290 71.055 ;
        RECT 43.515 70.755 44.400 70.925 ;
        RECT 42.360 70.075 42.870 70.165 ;
        RECT 40.910 69.265 41.135 69.395 ;
        RECT 41.305 69.325 41.830 69.545 ;
        RECT 42.000 69.905 42.870 70.075 ;
        RECT 40.545 68.675 40.795 69.135 ;
        RECT 40.965 69.125 41.135 69.265 ;
        RECT 42.000 69.125 42.170 69.905 ;
        RECT 42.700 69.835 42.870 69.905 ;
        RECT 42.380 69.655 42.580 69.685 ;
        RECT 43.040 69.655 43.210 70.725 ;
        RECT 43.380 69.835 43.570 70.555 ;
        RECT 42.380 69.355 43.210 69.655 ;
        RECT 43.740 69.625 44.060 70.585 ;
        RECT 40.965 68.955 41.300 69.125 ;
        RECT 41.495 68.955 42.170 69.125 ;
        RECT 42.490 68.675 42.860 69.175 ;
        RECT 43.040 69.125 43.210 69.355 ;
        RECT 43.595 69.295 44.060 69.625 ;
        RECT 44.230 69.915 44.400 70.755 ;
        RECT 44.580 70.725 44.895 71.225 ;
        RECT 45.125 70.495 45.465 71.055 ;
        RECT 44.570 70.120 45.465 70.495 ;
        RECT 45.635 70.215 45.805 71.225 ;
        RECT 45.275 69.915 45.465 70.120 ;
        RECT 45.975 70.165 46.305 71.010 ;
        RECT 45.975 70.085 46.365 70.165 ;
        RECT 46.150 70.035 46.365 70.085 ;
        RECT 44.230 69.585 45.105 69.915 ;
        RECT 45.275 69.585 46.025 69.915 ;
        RECT 44.230 69.125 44.400 69.585 ;
        RECT 45.275 69.415 45.475 69.585 ;
        RECT 46.195 69.455 46.365 70.035 ;
        RECT 46.140 69.415 46.365 69.455 ;
        RECT 43.040 68.955 43.445 69.125 ;
        RECT 43.615 68.955 44.400 69.125 ;
        RECT 44.675 68.675 44.885 69.205 ;
        RECT 45.145 68.890 45.475 69.415 ;
        RECT 45.985 69.330 46.365 69.415 ;
        RECT 46.540 70.085 46.875 71.055 ;
        RECT 47.045 70.085 47.215 71.225 ;
        RECT 47.385 70.885 49.415 71.055 ;
        RECT 46.540 69.415 46.710 70.085 ;
        RECT 47.385 69.915 47.555 70.885 ;
        RECT 46.880 69.585 47.135 69.915 ;
        RECT 47.360 69.585 47.555 69.915 ;
        RECT 47.725 70.545 48.850 70.715 ;
        RECT 46.965 69.415 47.135 69.585 ;
        RECT 47.725 69.415 47.895 70.545 ;
        RECT 45.645 68.675 45.815 69.285 ;
        RECT 45.985 68.895 46.315 69.330 ;
        RECT 46.540 68.845 46.795 69.415 ;
        RECT 46.965 69.245 47.895 69.415 ;
        RECT 48.065 70.205 49.075 70.375 ;
        RECT 48.065 69.405 48.235 70.205 ;
        RECT 47.720 69.210 47.895 69.245 ;
        RECT 46.965 68.675 47.295 69.075 ;
        RECT 47.720 68.845 48.250 69.210 ;
        RECT 48.440 69.185 48.715 70.005 ;
        RECT 48.435 69.015 48.715 69.185 ;
        RECT 48.440 68.845 48.715 69.015 ;
        RECT 48.885 68.845 49.075 70.205 ;
        RECT 49.245 70.220 49.415 70.885 ;
        RECT 49.585 70.465 49.755 71.225 ;
        RECT 49.990 70.465 50.505 70.875 ;
        RECT 49.245 70.030 49.995 70.220 ;
        RECT 50.165 69.655 50.505 70.465 ;
        RECT 50.675 70.060 50.965 71.225 ;
        RECT 51.135 70.085 51.520 71.055 ;
        RECT 51.690 70.765 52.015 71.225 ;
        RECT 52.535 70.595 52.815 71.055 ;
        RECT 51.690 70.375 52.815 70.595 ;
        RECT 49.275 69.485 50.505 69.655 ;
        RECT 49.255 68.675 49.765 69.210 ;
        RECT 49.985 68.880 50.230 69.485 ;
        RECT 51.135 69.415 51.415 70.085 ;
        RECT 51.690 69.915 52.140 70.375 ;
        RECT 53.005 70.205 53.405 71.055 ;
        RECT 53.805 70.765 54.075 71.225 ;
        RECT 54.245 70.595 54.530 71.055 ;
        RECT 51.585 69.585 52.140 69.915 ;
        RECT 52.310 69.645 53.405 70.205 ;
        RECT 51.690 69.475 52.140 69.585 ;
        RECT 50.675 68.675 50.965 69.400 ;
        RECT 51.135 68.845 51.520 69.415 ;
        RECT 51.690 69.305 52.815 69.475 ;
        RECT 51.690 68.675 52.015 69.135 ;
        RECT 52.535 68.845 52.815 69.305 ;
        RECT 53.005 68.845 53.405 69.645 ;
        RECT 53.575 70.375 54.530 70.595 ;
        RECT 53.575 69.475 53.785 70.375 ;
        RECT 53.955 69.645 54.645 70.205 ;
        RECT 54.815 70.135 58.325 71.225 ;
        RECT 53.575 69.305 54.530 69.475 ;
        RECT 53.805 68.675 54.075 69.135 ;
        RECT 54.245 68.845 54.530 69.305 ;
        RECT 54.815 69.445 56.465 69.965 ;
        RECT 56.635 69.615 58.325 70.135 ;
        RECT 59.425 70.115 59.720 71.225 ;
        RECT 59.900 69.915 60.150 71.050 ;
        RECT 60.320 70.115 60.580 71.225 ;
        RECT 60.750 70.325 61.010 71.050 ;
        RECT 61.180 70.495 61.440 71.225 ;
        RECT 61.610 70.325 61.870 71.050 ;
        RECT 62.040 70.495 62.300 71.225 ;
        RECT 62.470 70.325 62.730 71.050 ;
        RECT 62.900 70.495 63.160 71.225 ;
        RECT 63.330 70.325 63.590 71.050 ;
        RECT 63.760 70.495 64.055 71.225 ;
        RECT 64.590 70.595 64.875 71.055 ;
        RECT 65.045 70.765 65.315 71.225 ;
        RECT 64.590 70.375 65.545 70.595 ;
        RECT 60.750 70.085 64.060 70.325 ;
        RECT 54.815 68.675 58.325 69.445 ;
        RECT 59.415 69.305 59.730 69.915 ;
        RECT 59.900 69.665 62.920 69.915 ;
        RECT 59.475 68.675 59.720 69.135 ;
        RECT 59.900 68.855 60.150 69.665 ;
        RECT 63.090 69.495 64.060 70.085 ;
        RECT 64.475 69.645 65.165 70.205 ;
        RECT 60.750 69.325 64.060 69.495 ;
        RECT 65.335 69.475 65.545 70.375 ;
        RECT 60.320 68.675 60.580 69.200 ;
        RECT 60.750 68.870 61.010 69.325 ;
        RECT 61.180 68.675 61.440 69.155 ;
        RECT 61.610 68.870 61.870 69.325 ;
        RECT 62.040 68.675 62.300 69.155 ;
        RECT 62.470 68.870 62.730 69.325 ;
        RECT 62.900 68.675 63.160 69.155 ;
        RECT 63.330 68.870 63.590 69.325 ;
        RECT 64.590 69.305 65.545 69.475 ;
        RECT 65.715 70.205 66.115 71.055 ;
        RECT 66.305 70.595 66.585 71.055 ;
        RECT 67.105 70.765 67.430 71.225 ;
        RECT 66.305 70.375 67.430 70.595 ;
        RECT 65.715 69.645 66.810 70.205 ;
        RECT 66.980 69.915 67.430 70.375 ;
        RECT 67.600 70.085 67.985 71.055 ;
        RECT 63.760 68.675 64.060 69.155 ;
        RECT 64.590 68.845 64.875 69.305 ;
        RECT 65.045 68.675 65.315 69.135 ;
        RECT 65.715 68.845 66.115 69.645 ;
        RECT 66.980 69.585 67.535 69.915 ;
        RECT 66.980 69.475 67.430 69.585 ;
        RECT 66.305 69.305 67.430 69.475 ;
        RECT 67.705 69.415 67.985 70.085 ;
        RECT 66.305 68.845 66.585 69.305 ;
        RECT 67.105 68.675 67.430 69.135 ;
        RECT 67.600 68.845 67.985 69.415 ;
        RECT 68.155 70.505 68.615 71.055 ;
        RECT 68.805 70.505 69.135 71.225 ;
        RECT 68.155 69.135 68.405 70.505 ;
        RECT 69.335 70.335 69.635 70.885 ;
        RECT 69.805 70.555 70.085 71.225 ;
        RECT 68.695 70.165 69.635 70.335 ;
        RECT 68.695 69.915 68.865 70.165 ;
        RECT 70.005 69.915 70.270 70.275 ;
        RECT 70.515 70.085 70.725 71.225 ;
        RECT 68.575 69.585 68.865 69.915 ;
        RECT 69.035 69.665 69.375 69.915 ;
        RECT 69.595 69.665 70.270 69.915 ;
        RECT 70.895 70.075 71.225 71.055 ;
        RECT 71.395 70.085 71.625 71.225 ;
        RECT 71.835 70.085 72.115 71.225 ;
        RECT 72.285 70.075 72.615 71.055 ;
        RECT 72.785 70.085 73.045 71.225 ;
        RECT 73.215 70.715 74.405 71.005 ;
        RECT 73.235 70.375 74.405 70.545 ;
        RECT 74.575 70.425 74.855 71.225 ;
        RECT 73.235 70.085 73.560 70.375 ;
        RECT 74.235 70.255 74.405 70.375 ;
        RECT 68.695 69.495 68.865 69.585 ;
        RECT 68.695 69.305 70.085 69.495 ;
        RECT 68.155 68.845 68.715 69.135 ;
        RECT 68.885 68.675 69.135 69.135 ;
        RECT 69.755 68.945 70.085 69.305 ;
        RECT 70.515 68.675 70.725 69.495 ;
        RECT 70.895 69.475 71.145 70.075 ;
        RECT 71.315 69.665 71.645 69.915 ;
        RECT 71.845 69.645 72.180 69.915 ;
        RECT 70.895 68.845 71.225 69.475 ;
        RECT 71.395 68.675 71.625 69.495 ;
        RECT 72.350 69.475 72.520 70.075 ;
        RECT 73.730 69.915 73.925 70.205 ;
        RECT 74.235 70.085 74.895 70.255 ;
        RECT 75.065 70.085 75.340 71.055 ;
        RECT 74.725 69.915 74.895 70.085 ;
        RECT 72.690 69.665 73.025 69.915 ;
        RECT 73.215 69.585 73.560 69.915 ;
        RECT 73.730 69.585 74.555 69.915 ;
        RECT 74.725 69.585 75.000 69.915 ;
        RECT 71.835 68.675 72.145 69.475 ;
        RECT 72.350 68.845 73.045 69.475 ;
        RECT 74.725 69.415 74.895 69.585 ;
        RECT 73.230 69.245 74.895 69.415 ;
        RECT 75.170 69.350 75.340 70.085 ;
        RECT 76.435 70.060 76.725 71.225 ;
        RECT 77.820 70.835 78.155 71.055 ;
        RECT 79.160 70.845 79.515 71.225 ;
        RECT 77.820 70.215 78.075 70.835 ;
        RECT 78.325 70.675 78.555 70.715 ;
        RECT 79.685 70.675 79.935 71.055 ;
        RECT 78.325 70.475 79.935 70.675 ;
        RECT 78.325 70.385 78.510 70.475 ;
        RECT 79.100 70.465 79.935 70.475 ;
        RECT 80.185 70.445 80.435 71.225 ;
        RECT 80.605 70.375 80.865 71.055 ;
        RECT 78.665 70.275 78.995 70.305 ;
        RECT 78.665 70.215 80.465 70.275 ;
        RECT 77.820 70.105 80.525 70.215 ;
        RECT 77.820 70.045 78.995 70.105 ;
        RECT 80.325 70.070 80.525 70.105 ;
        RECT 77.815 69.665 78.305 69.865 ;
        RECT 78.495 69.665 78.970 69.875 ;
        RECT 73.230 68.895 73.485 69.245 ;
        RECT 73.655 68.675 73.985 69.075 ;
        RECT 74.155 68.895 74.325 69.245 ;
        RECT 74.495 68.675 74.875 69.075 ;
        RECT 75.065 69.005 75.340 69.350 ;
        RECT 76.435 68.675 76.725 69.400 ;
        RECT 77.820 68.675 78.275 69.440 ;
        RECT 78.750 69.265 78.970 69.665 ;
        RECT 79.215 69.665 79.545 69.875 ;
        RECT 79.215 69.265 79.425 69.665 ;
        RECT 79.715 69.630 80.125 69.935 ;
        RECT 80.355 69.495 80.525 70.070 ;
        RECT 80.255 69.375 80.525 69.495 ;
        RECT 79.680 69.330 80.525 69.375 ;
        RECT 79.680 69.205 80.435 69.330 ;
        RECT 79.680 69.055 79.850 69.205 ;
        RECT 80.695 69.185 80.865 70.375 ;
        RECT 81.035 70.135 83.625 71.225 ;
        RECT 80.635 69.175 80.865 69.185 ;
        RECT 78.550 68.845 79.850 69.055 ;
        RECT 80.105 68.675 80.435 69.035 ;
        RECT 80.605 68.845 80.865 69.175 ;
        RECT 81.035 69.445 82.245 69.965 ;
        RECT 82.415 69.615 83.625 70.135 ;
        RECT 83.800 70.075 84.060 71.225 ;
        RECT 84.235 70.150 84.490 71.055 ;
        RECT 84.660 70.465 84.990 71.225 ;
        RECT 85.205 70.295 85.375 71.055 ;
        RECT 81.035 68.675 83.625 69.445 ;
        RECT 83.800 68.675 84.060 69.515 ;
        RECT 84.235 69.420 84.405 70.150 ;
        RECT 84.660 70.125 85.375 70.295 ;
        RECT 84.660 69.915 84.830 70.125 ;
        RECT 85.635 70.085 86.020 71.055 ;
        RECT 86.190 70.765 86.515 71.225 ;
        RECT 87.035 70.595 87.315 71.055 ;
        RECT 86.190 70.375 87.315 70.595 ;
        RECT 84.575 69.585 84.830 69.915 ;
        RECT 84.235 68.845 84.490 69.420 ;
        RECT 84.660 69.395 84.830 69.585 ;
        RECT 85.110 69.575 85.465 69.945 ;
        RECT 85.635 69.415 85.915 70.085 ;
        RECT 86.190 69.915 86.640 70.375 ;
        RECT 87.505 70.205 87.905 71.055 ;
        RECT 88.305 70.765 88.575 71.225 ;
        RECT 88.745 70.595 89.030 71.055 ;
        RECT 86.085 69.585 86.640 69.915 ;
        RECT 86.810 69.645 87.905 70.205 ;
        RECT 86.190 69.475 86.640 69.585 ;
        RECT 84.660 69.225 85.375 69.395 ;
        RECT 84.660 68.675 84.990 69.055 ;
        RECT 85.205 68.845 85.375 69.225 ;
        RECT 85.635 68.845 86.020 69.415 ;
        RECT 86.190 69.305 87.315 69.475 ;
        RECT 86.190 68.675 86.515 69.135 ;
        RECT 87.035 68.845 87.315 69.305 ;
        RECT 87.505 68.845 87.905 69.645 ;
        RECT 88.075 70.375 89.030 70.595 ;
        RECT 88.075 69.475 88.285 70.375 ;
        RECT 88.455 69.645 89.145 70.205 ;
        RECT 89.315 70.135 90.525 71.225 ;
        RECT 89.315 69.595 89.835 70.135 ;
        RECT 88.075 69.305 89.030 69.475 ;
        RECT 90.005 69.425 90.525 69.965 ;
        RECT 88.305 68.675 88.575 69.135 ;
        RECT 88.745 68.845 89.030 69.305 ;
        RECT 89.315 68.675 90.525 69.425 ;
        RECT 11.950 68.505 90.610 68.675 ;
        RECT 12.035 67.755 13.245 68.505 ;
        RECT 12.035 67.215 12.555 67.755 ;
        RECT 13.420 67.665 13.680 68.505 ;
        RECT 13.855 67.760 14.110 68.335 ;
        RECT 14.280 68.125 14.610 68.505 ;
        RECT 14.825 67.955 14.995 68.335 ;
        RECT 14.280 67.785 14.995 67.955 ;
        RECT 16.265 67.955 16.435 68.245 ;
        RECT 16.605 68.125 16.935 68.505 ;
        RECT 16.265 67.785 16.930 67.955 ;
        RECT 12.725 67.045 13.245 67.585 ;
        RECT 12.035 65.955 13.245 67.045 ;
        RECT 13.420 65.955 13.680 67.105 ;
        RECT 13.855 67.030 14.025 67.760 ;
        RECT 14.280 67.595 14.450 67.785 ;
        RECT 14.195 67.265 14.450 67.595 ;
        RECT 14.280 67.055 14.450 67.265 ;
        RECT 14.730 67.235 15.085 67.605 ;
        RECT 13.855 66.125 14.110 67.030 ;
        RECT 14.280 66.885 14.995 67.055 ;
        RECT 16.180 66.965 16.530 67.615 ;
        RECT 14.280 65.955 14.610 66.715 ;
        RECT 14.825 66.125 14.995 66.885 ;
        RECT 16.700 66.795 16.930 67.785 ;
        RECT 16.265 66.625 16.930 66.795 ;
        RECT 16.265 66.125 16.435 66.625 ;
        RECT 16.605 65.955 16.935 66.455 ;
        RECT 17.105 66.125 17.290 68.245 ;
        RECT 17.545 68.045 17.795 68.505 ;
        RECT 17.965 68.055 18.300 68.225 ;
        RECT 18.495 68.055 19.170 68.225 ;
        RECT 17.965 67.915 18.135 68.055 ;
        RECT 17.460 66.925 17.740 67.875 ;
        RECT 17.910 67.785 18.135 67.915 ;
        RECT 17.910 66.680 18.080 67.785 ;
        RECT 18.305 67.635 18.830 67.855 ;
        RECT 18.250 66.870 18.490 67.465 ;
        RECT 18.660 66.935 18.830 67.635 ;
        RECT 19.000 67.275 19.170 68.055 ;
        RECT 19.490 68.005 19.860 68.505 ;
        RECT 20.040 68.055 20.445 68.225 ;
        RECT 20.615 68.055 21.400 68.225 ;
        RECT 20.040 67.825 20.210 68.055 ;
        RECT 19.380 67.525 20.210 67.825 ;
        RECT 20.595 67.555 21.060 67.885 ;
        RECT 19.380 67.495 19.580 67.525 ;
        RECT 19.700 67.275 19.870 67.345 ;
        RECT 19.000 67.105 19.870 67.275 ;
        RECT 19.360 67.015 19.870 67.105 ;
        RECT 17.910 66.550 18.215 66.680 ;
        RECT 18.660 66.570 19.190 66.935 ;
        RECT 17.530 65.955 17.795 66.415 ;
        RECT 17.965 66.125 18.215 66.550 ;
        RECT 19.360 66.400 19.530 67.015 ;
        RECT 18.425 66.230 19.530 66.400 ;
        RECT 19.700 65.955 19.870 66.755 ;
        RECT 20.040 66.455 20.210 67.525 ;
        RECT 20.380 66.625 20.570 67.345 ;
        RECT 20.740 66.595 21.060 67.555 ;
        RECT 21.230 67.595 21.400 68.055 ;
        RECT 21.675 67.975 21.885 68.505 ;
        RECT 22.145 67.765 22.475 68.290 ;
        RECT 22.645 67.895 22.815 68.505 ;
        RECT 22.985 67.850 23.315 68.285 ;
        RECT 23.485 67.990 23.655 68.505 ;
        RECT 22.985 67.765 23.365 67.850 ;
        RECT 22.275 67.595 22.475 67.765 ;
        RECT 23.140 67.725 23.365 67.765 ;
        RECT 21.230 67.265 22.105 67.595 ;
        RECT 22.275 67.265 23.025 67.595 ;
        RECT 20.040 66.125 20.290 66.455 ;
        RECT 21.230 66.425 21.400 67.265 ;
        RECT 22.275 67.060 22.465 67.265 ;
        RECT 23.195 67.145 23.365 67.725 ;
        RECT 24.270 67.695 24.515 68.300 ;
        RECT 24.735 67.970 25.245 68.505 ;
        RECT 23.150 67.095 23.365 67.145 ;
        RECT 21.570 66.685 22.465 67.060 ;
        RECT 22.975 67.015 23.365 67.095 ;
        RECT 23.995 67.525 25.225 67.695 ;
        RECT 20.515 66.255 21.400 66.425 ;
        RECT 21.580 65.955 21.895 66.455 ;
        RECT 22.125 66.125 22.465 66.685 ;
        RECT 22.635 65.955 22.805 66.965 ;
        RECT 22.975 66.170 23.305 67.015 ;
        RECT 23.475 65.955 23.645 66.870 ;
        RECT 23.995 66.715 24.335 67.525 ;
        RECT 24.505 66.960 25.255 67.150 ;
        RECT 23.995 66.305 24.510 66.715 ;
        RECT 24.745 65.955 24.915 66.715 ;
        RECT 25.085 66.295 25.255 66.960 ;
        RECT 25.425 66.975 25.615 68.335 ;
        RECT 25.785 68.165 26.060 68.335 ;
        RECT 25.785 67.995 26.065 68.165 ;
        RECT 25.785 67.175 26.060 67.995 ;
        RECT 26.250 67.970 26.780 68.335 ;
        RECT 27.205 68.105 27.535 68.505 ;
        RECT 26.605 67.935 26.780 67.970 ;
        RECT 26.265 66.975 26.435 67.775 ;
        RECT 25.425 66.805 26.435 66.975 ;
        RECT 26.605 67.765 27.535 67.935 ;
        RECT 27.705 67.765 27.960 68.335 ;
        RECT 28.135 67.960 33.480 68.505 ;
        RECT 26.605 66.635 26.775 67.765 ;
        RECT 27.365 67.595 27.535 67.765 ;
        RECT 25.650 66.465 26.775 66.635 ;
        RECT 26.945 67.265 27.140 67.595 ;
        RECT 27.365 67.265 27.620 67.595 ;
        RECT 26.945 66.295 27.115 67.265 ;
        RECT 27.790 67.095 27.960 67.765 ;
        RECT 29.720 67.130 30.060 67.960 ;
        RECT 33.655 67.735 37.165 68.505 ;
        RECT 37.795 67.780 38.085 68.505 ;
        RECT 38.715 67.765 39.100 68.335 ;
        RECT 39.270 68.045 39.595 68.505 ;
        RECT 40.115 67.875 40.395 68.335 ;
        RECT 25.085 66.125 27.115 66.295 ;
        RECT 27.285 65.955 27.455 67.095 ;
        RECT 27.625 66.125 27.960 67.095 ;
        RECT 31.540 66.390 31.890 67.640 ;
        RECT 33.655 67.215 35.305 67.735 ;
        RECT 35.475 67.045 37.165 67.565 ;
        RECT 28.135 65.955 33.480 66.390 ;
        RECT 33.655 65.955 37.165 67.045 ;
        RECT 37.795 65.955 38.085 67.120 ;
        RECT 38.715 67.095 38.995 67.765 ;
        RECT 39.270 67.705 40.395 67.875 ;
        RECT 39.270 67.595 39.720 67.705 ;
        RECT 39.165 67.265 39.720 67.595 ;
        RECT 40.585 67.535 40.985 68.335 ;
        RECT 41.385 68.045 41.655 68.505 ;
        RECT 41.825 67.875 42.110 68.335 ;
        RECT 38.715 66.125 39.100 67.095 ;
        RECT 39.270 66.805 39.720 67.265 ;
        RECT 39.890 66.975 40.985 67.535 ;
        RECT 39.270 66.585 40.395 66.805 ;
        RECT 39.270 65.955 39.595 66.415 ;
        RECT 40.115 66.125 40.395 66.585 ;
        RECT 40.585 66.125 40.985 66.975 ;
        RECT 41.155 67.705 42.110 67.875 ;
        RECT 42.445 67.965 42.670 68.325 ;
        RECT 42.850 68.135 43.180 68.505 ;
        RECT 43.360 67.965 43.615 68.325 ;
        RECT 44.180 68.135 44.925 68.505 ;
        RECT 42.445 67.775 44.930 67.965 ;
        RECT 41.155 66.805 41.365 67.705 ;
        RECT 41.535 66.975 42.225 67.535 ;
        RECT 42.405 67.265 42.675 67.595 ;
        RECT 42.855 67.265 43.290 67.595 ;
        RECT 43.470 67.265 44.045 67.595 ;
        RECT 44.225 67.265 44.505 67.595 ;
        RECT 44.705 67.085 44.930 67.775 ;
        RECT 42.435 66.905 44.930 67.085 ;
        RECT 45.105 66.905 45.440 68.325 ;
        RECT 45.615 67.755 46.825 68.505 ;
        RECT 46.995 67.765 47.380 68.335 ;
        RECT 47.550 68.045 47.875 68.505 ;
        RECT 48.395 67.875 48.675 68.335 ;
        RECT 45.615 67.215 46.135 67.755 ;
        RECT 46.305 67.045 46.825 67.585 ;
        RECT 41.155 66.585 42.110 66.805 ;
        RECT 41.385 65.955 41.655 66.415 ;
        RECT 41.825 66.125 42.110 66.585 ;
        RECT 42.435 66.135 42.725 66.905 ;
        RECT 43.295 66.495 44.485 66.725 ;
        RECT 43.295 66.135 43.555 66.495 ;
        RECT 43.725 65.955 44.055 66.325 ;
        RECT 44.225 66.135 44.485 66.495 ;
        RECT 44.675 65.955 45.005 66.675 ;
        RECT 45.175 66.135 45.440 66.905 ;
        RECT 45.615 65.955 46.825 67.045 ;
        RECT 46.995 67.095 47.275 67.765 ;
        RECT 47.550 67.705 48.675 67.875 ;
        RECT 47.550 67.595 48.000 67.705 ;
        RECT 47.445 67.265 48.000 67.595 ;
        RECT 48.865 67.535 49.265 68.335 ;
        RECT 49.665 68.045 49.935 68.505 ;
        RECT 50.105 67.875 50.390 68.335 ;
        RECT 46.995 66.125 47.380 67.095 ;
        RECT 47.550 66.805 48.000 67.265 ;
        RECT 48.170 66.975 49.265 67.535 ;
        RECT 47.550 66.585 48.675 66.805 ;
        RECT 47.550 65.955 47.875 66.415 ;
        RECT 48.395 66.125 48.675 66.585 ;
        RECT 48.865 66.125 49.265 66.975 ;
        RECT 49.435 67.705 50.390 67.875 ;
        RECT 51.600 67.765 51.855 68.335 ;
        RECT 52.025 68.105 52.355 68.505 ;
        RECT 52.780 67.970 53.310 68.335 ;
        RECT 52.780 67.935 52.955 67.970 ;
        RECT 52.025 67.765 52.955 67.935 ;
        RECT 49.435 66.805 49.645 67.705 ;
        RECT 49.815 66.975 50.505 67.535 ;
        RECT 51.600 67.095 51.770 67.765 ;
        RECT 52.025 67.595 52.195 67.765 ;
        RECT 51.940 67.265 52.195 67.595 ;
        RECT 52.420 67.265 52.615 67.595 ;
        RECT 49.435 66.585 50.390 66.805 ;
        RECT 49.665 65.955 49.935 66.415 ;
        RECT 50.105 66.125 50.390 66.585 ;
        RECT 51.600 66.125 51.935 67.095 ;
        RECT 52.105 65.955 52.275 67.095 ;
        RECT 52.445 66.295 52.615 67.265 ;
        RECT 52.785 66.635 52.955 67.765 ;
        RECT 53.125 66.975 53.295 67.775 ;
        RECT 53.500 67.485 53.775 68.335 ;
        RECT 53.495 67.315 53.775 67.485 ;
        RECT 53.500 67.175 53.775 67.315 ;
        RECT 53.945 66.975 54.135 68.335 ;
        RECT 54.315 67.970 54.825 68.505 ;
        RECT 55.045 67.695 55.290 68.300 ;
        RECT 55.785 67.850 56.115 68.285 ;
        RECT 56.285 67.895 56.455 68.505 ;
        RECT 55.735 67.765 56.115 67.850 ;
        RECT 56.625 67.765 56.955 68.290 ;
        RECT 57.215 67.975 57.425 68.505 ;
        RECT 57.700 68.055 58.485 68.225 ;
        RECT 58.655 68.055 59.060 68.225 ;
        RECT 55.735 67.725 55.960 67.765 ;
        RECT 54.335 67.525 55.565 67.695 ;
        RECT 53.125 66.805 54.135 66.975 ;
        RECT 54.305 66.960 55.055 67.150 ;
        RECT 52.785 66.465 53.910 66.635 ;
        RECT 54.305 66.295 54.475 66.960 ;
        RECT 55.225 66.715 55.565 67.525 ;
        RECT 55.735 67.145 55.905 67.725 ;
        RECT 56.625 67.595 56.825 67.765 ;
        RECT 57.700 67.595 57.870 68.055 ;
        RECT 56.075 67.265 56.825 67.595 ;
        RECT 56.995 67.265 57.870 67.595 ;
        RECT 55.735 67.095 55.950 67.145 ;
        RECT 55.735 67.015 56.125 67.095 ;
        RECT 52.445 66.125 54.475 66.295 ;
        RECT 54.645 65.955 54.815 66.715 ;
        RECT 55.050 66.305 55.565 66.715 ;
        RECT 55.795 66.170 56.125 67.015 ;
        RECT 56.635 67.060 56.825 67.265 ;
        RECT 56.295 65.955 56.465 66.965 ;
        RECT 56.635 66.685 57.530 67.060 ;
        RECT 56.635 66.125 56.975 66.685 ;
        RECT 57.205 65.955 57.520 66.455 ;
        RECT 57.700 66.425 57.870 67.265 ;
        RECT 58.040 67.555 58.505 67.885 ;
        RECT 58.890 67.825 59.060 68.055 ;
        RECT 59.240 68.005 59.610 68.505 ;
        RECT 59.930 68.055 60.605 68.225 ;
        RECT 60.800 68.055 61.135 68.225 ;
        RECT 58.040 66.595 58.360 67.555 ;
        RECT 58.890 67.525 59.720 67.825 ;
        RECT 58.530 66.625 58.720 67.345 ;
        RECT 58.890 66.455 59.060 67.525 ;
        RECT 59.520 67.495 59.720 67.525 ;
        RECT 59.230 67.275 59.400 67.345 ;
        RECT 59.930 67.275 60.100 68.055 ;
        RECT 60.965 67.915 61.135 68.055 ;
        RECT 61.305 68.045 61.555 68.505 ;
        RECT 59.230 67.105 60.100 67.275 ;
        RECT 60.270 67.635 60.795 67.855 ;
        RECT 60.965 67.785 61.190 67.915 ;
        RECT 59.230 67.015 59.740 67.105 ;
        RECT 57.700 66.255 58.585 66.425 ;
        RECT 58.810 66.125 59.060 66.455 ;
        RECT 59.230 65.955 59.400 66.755 ;
        RECT 59.570 66.400 59.740 67.015 ;
        RECT 60.270 66.935 60.440 67.635 ;
        RECT 59.910 66.570 60.440 66.935 ;
        RECT 60.610 66.870 60.850 67.465 ;
        RECT 61.020 66.680 61.190 67.785 ;
        RECT 61.360 66.925 61.640 67.875 ;
        RECT 60.885 66.550 61.190 66.680 ;
        RECT 59.570 66.230 60.675 66.400 ;
        RECT 60.885 66.125 61.135 66.550 ;
        RECT 61.305 65.955 61.570 66.415 ;
        RECT 61.810 66.125 61.995 68.245 ;
        RECT 62.165 68.125 62.495 68.505 ;
        RECT 62.665 67.955 62.835 68.245 ;
        RECT 62.170 67.785 62.835 67.955 ;
        RECT 62.170 66.795 62.400 67.785 ;
        RECT 63.555 67.780 63.845 68.505 ;
        RECT 64.020 67.765 64.275 68.335 ;
        RECT 64.445 68.105 64.775 68.505 ;
        RECT 65.200 67.970 65.730 68.335 ;
        RECT 65.920 68.165 66.195 68.335 ;
        RECT 65.915 67.995 66.195 68.165 ;
        RECT 65.200 67.935 65.375 67.970 ;
        RECT 64.445 67.765 65.375 67.935 ;
        RECT 62.570 66.965 62.920 67.615 ;
        RECT 62.170 66.625 62.835 66.795 ;
        RECT 62.165 65.955 62.495 66.455 ;
        RECT 62.665 66.125 62.835 66.625 ;
        RECT 63.555 65.955 63.845 67.120 ;
        RECT 64.020 67.095 64.190 67.765 ;
        RECT 64.445 67.595 64.615 67.765 ;
        RECT 64.360 67.265 64.615 67.595 ;
        RECT 64.840 67.265 65.035 67.595 ;
        RECT 64.020 66.125 64.355 67.095 ;
        RECT 64.525 65.955 64.695 67.095 ;
        RECT 64.865 66.295 65.035 67.265 ;
        RECT 65.205 66.635 65.375 67.765 ;
        RECT 65.545 66.975 65.715 67.775 ;
        RECT 65.920 67.175 66.195 67.995 ;
        RECT 66.365 66.975 66.555 68.335 ;
        RECT 66.735 67.970 67.245 68.505 ;
        RECT 67.465 67.695 67.710 68.300 ;
        RECT 68.155 67.735 70.745 68.505 ;
        RECT 71.390 67.935 71.645 68.285 ;
        RECT 71.815 68.105 72.145 68.505 ;
        RECT 72.315 67.935 72.485 68.285 ;
        RECT 72.655 68.105 73.035 68.505 ;
        RECT 71.390 67.765 73.055 67.935 ;
        RECT 73.225 67.830 73.500 68.175 ;
        RECT 66.755 67.525 67.985 67.695 ;
        RECT 65.545 66.805 66.555 66.975 ;
        RECT 66.725 66.960 67.475 67.150 ;
        RECT 65.205 66.465 66.330 66.635 ;
        RECT 66.725 66.295 66.895 66.960 ;
        RECT 67.645 66.715 67.985 67.525 ;
        RECT 68.155 67.215 69.365 67.735 ;
        RECT 72.885 67.595 73.055 67.765 ;
        RECT 69.535 67.045 70.745 67.565 ;
        RECT 71.375 67.265 71.720 67.595 ;
        RECT 71.890 67.265 72.715 67.595 ;
        RECT 72.885 67.265 73.160 67.595 ;
        RECT 64.865 66.125 66.895 66.295 ;
        RECT 67.065 65.955 67.235 66.715 ;
        RECT 67.470 66.305 67.985 66.715 ;
        RECT 68.155 65.955 70.745 67.045 ;
        RECT 71.395 66.805 71.720 67.095 ;
        RECT 71.890 66.975 72.085 67.265 ;
        RECT 72.885 67.095 73.055 67.265 ;
        RECT 73.330 67.095 73.500 67.830 ;
        RECT 73.880 67.725 74.380 68.335 ;
        RECT 73.675 67.265 74.025 67.515 ;
        RECT 74.210 67.095 74.380 67.725 ;
        RECT 75.010 67.855 75.340 68.335 ;
        RECT 75.510 68.045 75.735 68.505 ;
        RECT 75.905 67.855 76.235 68.335 ;
        RECT 75.010 67.685 76.235 67.855 ;
        RECT 76.425 67.705 76.675 68.505 ;
        RECT 76.845 67.705 77.185 68.335 ;
        RECT 77.360 67.740 77.815 68.505 ;
        RECT 78.090 68.125 79.390 68.335 ;
        RECT 79.645 68.145 79.975 68.505 ;
        RECT 79.220 67.975 79.390 68.125 ;
        RECT 80.145 68.005 80.405 68.335 ;
        RECT 74.550 67.315 74.880 67.515 ;
        RECT 75.050 67.315 75.380 67.515 ;
        RECT 75.550 67.315 75.970 67.515 ;
        RECT 76.145 67.345 76.840 67.515 ;
        RECT 76.145 67.095 76.315 67.345 ;
        RECT 77.010 67.095 77.185 67.705 ;
        RECT 78.290 67.515 78.510 67.915 ;
        RECT 77.355 67.315 77.845 67.515 ;
        RECT 78.035 67.305 78.510 67.515 ;
        RECT 78.755 67.515 78.965 67.915 ;
        RECT 79.220 67.850 79.975 67.975 ;
        RECT 79.220 67.805 80.065 67.850 ;
        RECT 79.795 67.685 80.065 67.805 ;
        RECT 78.755 67.305 79.085 67.515 ;
        RECT 79.255 67.245 79.665 67.550 ;
        RECT 72.395 66.925 73.055 67.095 ;
        RECT 72.395 66.805 72.565 66.925 ;
        RECT 71.395 66.635 72.565 66.805 ;
        RECT 71.375 66.175 72.565 66.465 ;
        RECT 72.735 65.955 73.015 66.755 ;
        RECT 73.225 66.125 73.500 67.095 ;
        RECT 73.880 66.925 76.315 67.095 ;
        RECT 73.880 66.125 74.210 66.925 ;
        RECT 74.380 65.955 74.710 66.755 ;
        RECT 75.010 66.125 75.340 66.925 ;
        RECT 75.985 65.955 76.235 66.755 ;
        RECT 76.505 65.955 76.675 67.095 ;
        RECT 76.845 66.125 77.185 67.095 ;
        RECT 77.360 67.075 78.535 67.135 ;
        RECT 79.895 67.110 80.065 67.685 ;
        RECT 79.865 67.075 80.065 67.110 ;
        RECT 77.360 66.965 80.065 67.075 ;
        RECT 77.360 66.345 77.615 66.965 ;
        RECT 78.205 66.905 80.005 66.965 ;
        RECT 78.205 66.875 78.535 66.905 ;
        RECT 80.235 66.805 80.405 68.005 ;
        RECT 80.665 67.955 80.835 68.245 ;
        RECT 81.005 68.125 81.335 68.505 ;
        RECT 80.665 67.785 81.330 67.955 ;
        RECT 80.580 66.965 80.930 67.615 ;
        RECT 77.865 66.705 78.050 66.795 ;
        RECT 78.640 66.705 79.475 66.715 ;
        RECT 77.865 66.505 79.475 66.705 ;
        RECT 77.865 66.465 78.095 66.505 ;
        RECT 77.360 66.125 77.695 66.345 ;
        RECT 78.700 65.955 79.055 66.335 ;
        RECT 79.225 66.125 79.475 66.505 ;
        RECT 79.725 65.955 79.975 66.735 ;
        RECT 80.145 66.125 80.405 66.805 ;
        RECT 81.100 66.795 81.330 67.785 ;
        RECT 80.665 66.625 81.330 66.795 ;
        RECT 80.665 66.125 80.835 66.625 ;
        RECT 81.005 65.955 81.335 66.455 ;
        RECT 81.505 66.125 81.690 68.245 ;
        RECT 81.945 68.045 82.195 68.505 ;
        RECT 82.365 68.055 82.700 68.225 ;
        RECT 82.895 68.055 83.570 68.225 ;
        RECT 82.365 67.915 82.535 68.055 ;
        RECT 81.860 66.925 82.140 67.875 ;
        RECT 82.310 67.785 82.535 67.915 ;
        RECT 82.310 66.680 82.480 67.785 ;
        RECT 82.705 67.635 83.230 67.855 ;
        RECT 82.650 66.870 82.890 67.465 ;
        RECT 83.060 66.935 83.230 67.635 ;
        RECT 83.400 67.275 83.570 68.055 ;
        RECT 83.890 68.005 84.260 68.505 ;
        RECT 84.440 68.055 84.845 68.225 ;
        RECT 85.015 68.055 85.800 68.225 ;
        RECT 84.440 67.825 84.610 68.055 ;
        RECT 83.780 67.525 84.610 67.825 ;
        RECT 84.995 67.555 85.460 67.885 ;
        RECT 83.780 67.495 83.980 67.525 ;
        RECT 84.100 67.275 84.270 67.345 ;
        RECT 83.400 67.105 84.270 67.275 ;
        RECT 83.760 67.015 84.270 67.105 ;
        RECT 82.310 66.550 82.615 66.680 ;
        RECT 83.060 66.570 83.590 66.935 ;
        RECT 81.930 65.955 82.195 66.415 ;
        RECT 82.365 66.125 82.615 66.550 ;
        RECT 83.760 66.400 83.930 67.015 ;
        RECT 82.825 66.230 83.930 66.400 ;
        RECT 84.100 65.955 84.270 66.755 ;
        RECT 84.440 66.455 84.610 67.525 ;
        RECT 84.780 66.625 84.970 67.345 ;
        RECT 85.140 66.595 85.460 67.555 ;
        RECT 85.630 67.595 85.800 68.055 ;
        RECT 86.075 67.975 86.285 68.505 ;
        RECT 86.545 67.765 86.875 68.290 ;
        RECT 87.045 67.895 87.215 68.505 ;
        RECT 87.385 67.850 87.715 68.285 ;
        RECT 87.385 67.765 87.765 67.850 ;
        RECT 86.675 67.595 86.875 67.765 ;
        RECT 87.540 67.725 87.765 67.765 ;
        RECT 85.630 67.265 86.505 67.595 ;
        RECT 86.675 67.265 87.425 67.595 ;
        RECT 84.440 66.125 84.690 66.455 ;
        RECT 85.630 66.425 85.800 67.265 ;
        RECT 86.675 67.060 86.865 67.265 ;
        RECT 87.595 67.145 87.765 67.725 ;
        RECT 87.550 67.095 87.765 67.145 ;
        RECT 85.970 66.685 86.865 67.060 ;
        RECT 87.375 67.015 87.765 67.095 ;
        RECT 87.935 67.830 88.195 68.335 ;
        RECT 88.375 68.125 88.705 68.505 ;
        RECT 88.885 67.955 89.055 68.335 ;
        RECT 87.935 67.030 88.105 67.830 ;
        RECT 88.390 67.785 89.055 67.955 ;
        RECT 88.390 67.530 88.560 67.785 ;
        RECT 89.315 67.755 90.525 68.505 ;
        RECT 88.275 67.200 88.560 67.530 ;
        RECT 88.795 67.235 89.125 67.605 ;
        RECT 88.390 67.055 88.560 67.200 ;
        RECT 84.915 66.255 85.800 66.425 ;
        RECT 85.980 65.955 86.295 66.455 ;
        RECT 86.525 66.125 86.865 66.685 ;
        RECT 87.035 65.955 87.205 66.965 ;
        RECT 87.375 66.170 87.705 67.015 ;
        RECT 87.935 66.125 88.205 67.030 ;
        RECT 88.390 66.885 89.055 67.055 ;
        RECT 88.375 65.955 88.705 66.715 ;
        RECT 88.885 66.125 89.055 66.885 ;
        RECT 89.315 67.045 89.835 67.585 ;
        RECT 90.005 67.215 90.525 67.755 ;
        RECT 89.315 65.955 90.525 67.045 ;
        RECT 11.950 65.785 90.610 65.955 ;
        RECT 12.035 64.695 13.245 65.785 ;
        RECT 12.035 63.985 12.555 64.525 ;
        RECT 12.725 64.155 13.245 64.695 ;
        RECT 13.420 64.635 13.680 65.785 ;
        RECT 13.855 64.710 14.110 65.615 ;
        RECT 14.280 65.025 14.610 65.785 ;
        RECT 14.825 64.855 14.995 65.615 ;
        RECT 12.035 63.235 13.245 63.985 ;
        RECT 13.420 63.235 13.680 64.075 ;
        RECT 13.855 63.980 14.025 64.710 ;
        RECT 14.280 64.685 14.995 64.855 ;
        RECT 14.280 64.475 14.450 64.685 ;
        RECT 15.260 64.635 15.520 65.785 ;
        RECT 15.695 64.710 15.950 65.615 ;
        RECT 16.120 65.025 16.450 65.785 ;
        RECT 16.665 64.855 16.835 65.615 ;
        RECT 14.195 64.145 14.450 64.475 ;
        RECT 13.855 63.405 14.110 63.980 ;
        RECT 14.280 63.955 14.450 64.145 ;
        RECT 14.730 64.135 15.085 64.505 ;
        RECT 14.280 63.785 14.995 63.955 ;
        RECT 14.280 63.235 14.610 63.615 ;
        RECT 14.825 63.405 14.995 63.785 ;
        RECT 15.260 63.235 15.520 64.075 ;
        RECT 15.695 63.980 15.865 64.710 ;
        RECT 16.120 64.685 16.835 64.855 ;
        RECT 17.095 64.695 18.305 65.785 ;
        RECT 16.120 64.475 16.290 64.685 ;
        RECT 16.035 64.145 16.290 64.475 ;
        RECT 15.695 63.405 15.950 63.980 ;
        RECT 16.120 63.955 16.290 64.145 ;
        RECT 16.570 64.135 16.925 64.505 ;
        RECT 17.095 63.985 17.615 64.525 ;
        RECT 17.785 64.155 18.305 64.695 ;
        RECT 18.480 64.635 18.740 65.785 ;
        RECT 18.915 64.710 19.170 65.615 ;
        RECT 19.340 65.025 19.670 65.785 ;
        RECT 19.885 64.855 20.055 65.615 ;
        RECT 16.120 63.785 16.835 63.955 ;
        RECT 16.120 63.235 16.450 63.615 ;
        RECT 16.665 63.405 16.835 63.785 ;
        RECT 17.095 63.235 18.305 63.985 ;
        RECT 18.480 63.235 18.740 64.075 ;
        RECT 18.915 63.980 19.085 64.710 ;
        RECT 19.340 64.685 20.055 64.855 ;
        RECT 20.315 64.695 23.825 65.785 ;
        RECT 19.340 64.475 19.510 64.685 ;
        RECT 19.255 64.145 19.510 64.475 ;
        RECT 18.915 63.405 19.170 63.980 ;
        RECT 19.340 63.955 19.510 64.145 ;
        RECT 19.790 64.135 20.145 64.505 ;
        RECT 20.315 64.005 21.965 64.525 ;
        RECT 22.135 64.175 23.825 64.695 ;
        RECT 24.915 64.620 25.205 65.785 ;
        RECT 25.375 64.645 25.715 65.615 ;
        RECT 25.885 64.645 26.055 65.785 ;
        RECT 26.325 64.985 26.575 65.785 ;
        RECT 27.220 64.815 27.550 65.615 ;
        RECT 27.850 64.985 28.180 65.785 ;
        RECT 28.350 64.815 28.680 65.615 ;
        RECT 26.245 64.645 28.680 64.815 ;
        RECT 29.240 64.815 29.630 64.990 ;
        RECT 30.115 64.985 30.445 65.785 ;
        RECT 30.615 64.995 31.150 65.615 ;
        RECT 29.240 64.645 30.665 64.815 ;
        RECT 25.375 64.035 25.550 64.645 ;
        RECT 26.245 64.395 26.415 64.645 ;
        RECT 25.720 64.225 26.415 64.395 ;
        RECT 26.590 64.225 27.010 64.425 ;
        RECT 27.180 64.225 27.510 64.425 ;
        RECT 27.680 64.225 28.010 64.425 ;
        RECT 19.340 63.785 20.055 63.955 ;
        RECT 19.340 63.235 19.670 63.615 ;
        RECT 19.885 63.405 20.055 63.785 ;
        RECT 20.315 63.235 23.825 64.005 ;
        RECT 24.915 63.235 25.205 63.960 ;
        RECT 25.375 63.405 25.715 64.035 ;
        RECT 25.885 63.235 26.135 64.035 ;
        RECT 26.325 63.885 27.550 64.055 ;
        RECT 26.325 63.405 26.655 63.885 ;
        RECT 26.825 63.235 27.050 63.695 ;
        RECT 27.220 63.405 27.550 63.885 ;
        RECT 28.180 64.015 28.350 64.645 ;
        RECT 28.535 64.225 28.885 64.475 ;
        RECT 28.180 63.405 28.680 64.015 ;
        RECT 29.115 63.915 29.470 64.475 ;
        RECT 29.640 63.745 29.810 64.645 ;
        RECT 29.980 63.915 30.245 64.475 ;
        RECT 30.495 64.145 30.665 64.645 ;
        RECT 30.835 63.975 31.150 64.995 ;
        RECT 31.355 64.695 33.025 65.785 ;
        RECT 33.285 65.115 33.455 65.615 ;
        RECT 33.625 65.285 33.955 65.785 ;
        RECT 33.285 64.945 33.950 65.115 ;
        RECT 29.220 63.235 29.460 63.745 ;
        RECT 29.640 63.415 29.920 63.745 ;
        RECT 30.150 63.235 30.365 63.745 ;
        RECT 30.535 63.405 31.150 63.975 ;
        RECT 31.355 64.005 32.105 64.525 ;
        RECT 32.275 64.175 33.025 64.695 ;
        RECT 33.200 64.125 33.550 64.775 ;
        RECT 31.355 63.235 33.025 64.005 ;
        RECT 33.720 63.955 33.950 64.945 ;
        RECT 33.285 63.785 33.950 63.955 ;
        RECT 33.285 63.495 33.455 63.785 ;
        RECT 33.625 63.235 33.955 63.615 ;
        RECT 34.125 63.495 34.310 65.615 ;
        RECT 34.550 65.325 34.815 65.785 ;
        RECT 34.985 65.190 35.235 65.615 ;
        RECT 35.445 65.340 36.550 65.510 ;
        RECT 34.930 65.060 35.235 65.190 ;
        RECT 34.480 63.865 34.760 64.815 ;
        RECT 34.930 63.955 35.100 65.060 ;
        RECT 35.270 64.275 35.510 64.870 ;
        RECT 35.680 64.805 36.210 65.170 ;
        RECT 35.680 64.105 35.850 64.805 ;
        RECT 36.380 64.725 36.550 65.340 ;
        RECT 36.720 64.985 36.890 65.785 ;
        RECT 37.060 65.285 37.310 65.615 ;
        RECT 37.535 65.315 38.420 65.485 ;
        RECT 36.380 64.635 36.890 64.725 ;
        RECT 34.930 63.825 35.155 63.955 ;
        RECT 35.325 63.885 35.850 64.105 ;
        RECT 36.020 64.465 36.890 64.635 ;
        RECT 34.565 63.235 34.815 63.695 ;
        RECT 34.985 63.685 35.155 63.825 ;
        RECT 36.020 63.685 36.190 64.465 ;
        RECT 36.720 64.395 36.890 64.465 ;
        RECT 36.400 64.215 36.600 64.245 ;
        RECT 37.060 64.215 37.230 65.285 ;
        RECT 37.400 64.395 37.590 65.115 ;
        RECT 36.400 63.915 37.230 64.215 ;
        RECT 37.760 64.185 38.080 65.145 ;
        RECT 34.985 63.515 35.320 63.685 ;
        RECT 35.515 63.515 36.190 63.685 ;
        RECT 36.510 63.235 36.880 63.735 ;
        RECT 37.060 63.685 37.230 63.915 ;
        RECT 37.615 63.855 38.080 64.185 ;
        RECT 38.250 64.475 38.420 65.315 ;
        RECT 38.600 65.285 38.915 65.785 ;
        RECT 39.145 65.055 39.485 65.615 ;
        RECT 38.590 64.680 39.485 65.055 ;
        RECT 39.655 64.775 39.825 65.785 ;
        RECT 39.295 64.475 39.485 64.680 ;
        RECT 39.995 64.725 40.325 65.570 ;
        RECT 39.995 64.645 40.385 64.725 ;
        RECT 40.555 64.695 43.145 65.785 ;
        RECT 40.170 64.595 40.385 64.645 ;
        RECT 38.250 64.145 39.125 64.475 ;
        RECT 39.295 64.145 40.045 64.475 ;
        RECT 38.250 63.685 38.420 64.145 ;
        RECT 39.295 63.975 39.495 64.145 ;
        RECT 40.215 64.015 40.385 64.595 ;
        RECT 40.160 63.975 40.385 64.015 ;
        RECT 37.060 63.515 37.465 63.685 ;
        RECT 37.635 63.515 38.420 63.685 ;
        RECT 38.695 63.235 38.905 63.765 ;
        RECT 39.165 63.450 39.495 63.975 ;
        RECT 40.005 63.890 40.385 63.975 ;
        RECT 40.555 64.005 41.765 64.525 ;
        RECT 41.935 64.175 43.145 64.695 ;
        RECT 43.320 64.645 43.655 65.615 ;
        RECT 43.825 64.645 43.995 65.785 ;
        RECT 44.165 65.445 46.195 65.615 ;
        RECT 39.665 63.235 39.835 63.845 ;
        RECT 40.005 63.455 40.335 63.890 ;
        RECT 40.555 63.235 43.145 64.005 ;
        RECT 43.320 63.975 43.490 64.645 ;
        RECT 44.165 64.475 44.335 65.445 ;
        RECT 43.660 64.145 43.915 64.475 ;
        RECT 44.140 64.145 44.335 64.475 ;
        RECT 44.505 65.105 45.630 65.275 ;
        RECT 43.745 63.975 43.915 64.145 ;
        RECT 44.505 63.975 44.675 65.105 ;
        RECT 43.320 63.405 43.575 63.975 ;
        RECT 43.745 63.805 44.675 63.975 ;
        RECT 44.845 64.765 45.855 64.935 ;
        RECT 44.845 63.965 45.015 64.765 ;
        RECT 45.220 64.425 45.495 64.565 ;
        RECT 45.215 64.255 45.495 64.425 ;
        RECT 44.500 63.770 44.675 63.805 ;
        RECT 43.745 63.235 44.075 63.635 ;
        RECT 44.500 63.405 45.030 63.770 ;
        RECT 45.220 63.405 45.495 64.255 ;
        RECT 45.665 63.405 45.855 64.765 ;
        RECT 46.025 64.780 46.195 65.445 ;
        RECT 46.365 65.025 46.535 65.785 ;
        RECT 46.770 65.025 47.285 65.435 ;
        RECT 46.025 64.590 46.775 64.780 ;
        RECT 46.945 64.215 47.285 65.025 ;
        RECT 47.970 64.915 48.255 65.785 ;
        RECT 48.425 65.155 48.685 65.615 ;
        RECT 48.860 65.325 49.115 65.785 ;
        RECT 49.285 65.155 49.545 65.615 ;
        RECT 48.425 64.985 49.545 65.155 ;
        RECT 49.715 64.985 50.025 65.785 ;
        RECT 48.425 64.735 48.685 64.985 ;
        RECT 50.195 64.815 50.505 65.615 ;
        RECT 46.055 64.045 47.285 64.215 ;
        RECT 47.930 64.565 48.685 64.735 ;
        RECT 49.475 64.645 50.505 64.815 ;
        RECT 47.930 64.055 48.335 64.565 ;
        RECT 49.475 64.395 49.645 64.645 ;
        RECT 48.505 64.225 49.645 64.395 ;
        RECT 46.035 63.235 46.545 63.770 ;
        RECT 46.765 63.440 47.010 64.045 ;
        RECT 47.930 63.885 49.580 64.055 ;
        RECT 49.815 63.905 50.165 64.475 ;
        RECT 47.975 63.235 48.255 63.715 ;
        RECT 48.425 63.495 48.685 63.885 ;
        RECT 48.860 63.235 49.115 63.715 ;
        RECT 49.285 63.495 49.580 63.885 ;
        RECT 50.335 63.735 50.505 64.645 ;
        RECT 50.675 64.620 50.965 65.785 ;
        RECT 51.225 65.115 51.395 65.615 ;
        RECT 51.565 65.285 51.895 65.785 ;
        RECT 51.225 64.945 51.890 65.115 ;
        RECT 51.140 64.125 51.490 64.775 ;
        RECT 49.760 63.235 50.035 63.715 ;
        RECT 50.205 63.405 50.505 63.735 ;
        RECT 50.675 63.235 50.965 63.960 ;
        RECT 51.660 63.955 51.890 64.945 ;
        RECT 51.225 63.785 51.890 63.955 ;
        RECT 51.225 63.495 51.395 63.785 ;
        RECT 51.565 63.235 51.895 63.615 ;
        RECT 52.065 63.495 52.250 65.615 ;
        RECT 52.490 65.325 52.755 65.785 ;
        RECT 52.925 65.190 53.175 65.615 ;
        RECT 53.385 65.340 54.490 65.510 ;
        RECT 52.870 65.060 53.175 65.190 ;
        RECT 52.420 63.865 52.700 64.815 ;
        RECT 52.870 63.955 53.040 65.060 ;
        RECT 53.210 64.275 53.450 64.870 ;
        RECT 53.620 64.805 54.150 65.170 ;
        RECT 53.620 64.105 53.790 64.805 ;
        RECT 54.320 64.725 54.490 65.340 ;
        RECT 54.660 64.985 54.830 65.785 ;
        RECT 55.000 65.285 55.250 65.615 ;
        RECT 55.475 65.315 56.360 65.485 ;
        RECT 54.320 64.635 54.830 64.725 ;
        RECT 52.870 63.825 53.095 63.955 ;
        RECT 53.265 63.885 53.790 64.105 ;
        RECT 53.960 64.465 54.830 64.635 ;
        RECT 52.505 63.235 52.755 63.695 ;
        RECT 52.925 63.685 53.095 63.825 ;
        RECT 53.960 63.685 54.130 64.465 ;
        RECT 54.660 64.395 54.830 64.465 ;
        RECT 54.340 64.215 54.540 64.245 ;
        RECT 55.000 64.215 55.170 65.285 ;
        RECT 55.340 64.395 55.530 65.115 ;
        RECT 54.340 63.915 55.170 64.215 ;
        RECT 55.700 64.185 56.020 65.145 ;
        RECT 52.925 63.515 53.260 63.685 ;
        RECT 53.455 63.515 54.130 63.685 ;
        RECT 54.450 63.235 54.820 63.735 ;
        RECT 55.000 63.685 55.170 63.915 ;
        RECT 55.555 63.855 56.020 64.185 ;
        RECT 56.190 64.475 56.360 65.315 ;
        RECT 56.540 65.285 56.855 65.785 ;
        RECT 57.085 65.055 57.425 65.615 ;
        RECT 56.530 64.680 57.425 65.055 ;
        RECT 57.595 64.775 57.765 65.785 ;
        RECT 57.235 64.475 57.425 64.680 ;
        RECT 57.935 64.725 58.265 65.570 ;
        RECT 57.935 64.645 58.325 64.725 ;
        RECT 58.110 64.595 58.325 64.645 ;
        RECT 56.190 64.145 57.065 64.475 ;
        RECT 57.235 64.145 57.985 64.475 ;
        RECT 56.190 63.685 56.360 64.145 ;
        RECT 57.235 63.975 57.435 64.145 ;
        RECT 58.155 64.015 58.325 64.595 ;
        RECT 58.100 63.975 58.325 64.015 ;
        RECT 55.000 63.515 55.405 63.685 ;
        RECT 55.575 63.515 56.360 63.685 ;
        RECT 56.635 63.235 56.845 63.765 ;
        RECT 57.105 63.450 57.435 63.975 ;
        RECT 57.945 63.890 58.325 63.975 ;
        RECT 58.495 64.645 58.880 65.615 ;
        RECT 59.050 65.325 59.375 65.785 ;
        RECT 59.895 65.155 60.175 65.615 ;
        RECT 59.050 64.935 60.175 65.155 ;
        RECT 58.495 63.975 58.775 64.645 ;
        RECT 59.050 64.475 59.500 64.935 ;
        RECT 60.365 64.765 60.765 65.615 ;
        RECT 61.165 65.325 61.435 65.785 ;
        RECT 61.605 65.155 61.890 65.615 ;
        RECT 58.945 64.145 59.500 64.475 ;
        RECT 59.670 64.205 60.765 64.765 ;
        RECT 59.050 64.035 59.500 64.145 ;
        RECT 57.605 63.235 57.775 63.845 ;
        RECT 57.945 63.455 58.275 63.890 ;
        RECT 58.495 63.405 58.880 63.975 ;
        RECT 59.050 63.865 60.175 64.035 ;
        RECT 59.050 63.235 59.375 63.695 ;
        RECT 59.895 63.405 60.175 63.865 ;
        RECT 60.365 63.405 60.765 64.205 ;
        RECT 60.935 64.935 61.890 65.155 ;
        RECT 62.290 65.155 62.575 65.615 ;
        RECT 62.745 65.325 63.015 65.785 ;
        RECT 62.290 64.935 63.245 65.155 ;
        RECT 60.935 64.035 61.145 64.935 ;
        RECT 61.315 64.205 62.005 64.765 ;
        RECT 62.175 64.205 62.865 64.765 ;
        RECT 63.035 64.035 63.245 64.935 ;
        RECT 60.935 63.865 61.890 64.035 ;
        RECT 61.165 63.235 61.435 63.695 ;
        RECT 61.605 63.405 61.890 63.865 ;
        RECT 62.290 63.865 63.245 64.035 ;
        RECT 63.415 64.765 63.815 65.615 ;
        RECT 64.005 65.155 64.285 65.615 ;
        RECT 64.805 65.325 65.130 65.785 ;
        RECT 64.005 64.935 65.130 65.155 ;
        RECT 63.415 64.205 64.510 64.765 ;
        RECT 64.680 64.475 65.130 64.935 ;
        RECT 65.300 64.645 65.685 65.615 ;
        RECT 65.860 64.985 66.115 65.785 ;
        RECT 66.315 64.935 66.645 65.615 ;
        RECT 62.290 63.405 62.575 63.865 ;
        RECT 62.745 63.235 63.015 63.695 ;
        RECT 63.415 63.405 63.815 64.205 ;
        RECT 64.680 64.145 65.235 64.475 ;
        RECT 64.680 64.035 65.130 64.145 ;
        RECT 64.005 63.865 65.130 64.035 ;
        RECT 65.405 63.975 65.685 64.645 ;
        RECT 65.860 64.445 66.105 64.805 ;
        RECT 66.295 64.655 66.645 64.935 ;
        RECT 66.295 64.275 66.465 64.655 ;
        RECT 66.825 64.475 67.020 65.525 ;
        RECT 67.200 64.645 67.520 65.785 ;
        RECT 68.625 64.675 68.920 65.785 ;
        RECT 69.100 64.475 69.350 65.610 ;
        RECT 69.520 64.675 69.780 65.785 ;
        RECT 69.950 64.885 70.210 65.610 ;
        RECT 70.380 65.055 70.640 65.785 ;
        RECT 70.810 64.885 71.070 65.610 ;
        RECT 71.240 65.055 71.500 65.785 ;
        RECT 71.670 64.885 71.930 65.610 ;
        RECT 72.100 65.055 72.360 65.785 ;
        RECT 72.530 64.885 72.790 65.610 ;
        RECT 72.960 65.055 73.255 65.785 ;
        RECT 69.950 64.645 73.260 64.885 ;
        RECT 74.320 64.815 74.710 64.990 ;
        RECT 75.195 64.985 75.525 65.785 ;
        RECT 75.695 64.995 76.230 65.615 ;
        RECT 74.320 64.645 75.745 64.815 ;
        RECT 64.005 63.405 64.285 63.865 ;
        RECT 64.805 63.235 65.130 63.695 ;
        RECT 65.300 63.405 65.685 63.975 ;
        RECT 65.945 64.105 66.465 64.275 ;
        RECT 66.635 64.145 67.020 64.475 ;
        RECT 67.200 64.425 67.460 64.475 ;
        RECT 67.200 64.255 67.465 64.425 ;
        RECT 67.200 64.145 67.460 64.255 ;
        RECT 65.945 63.745 66.115 64.105 ;
        RECT 65.915 63.575 66.115 63.745 ;
        RECT 65.945 63.540 66.115 63.575 ;
        RECT 66.305 63.765 67.520 63.935 ;
        RECT 68.615 63.865 68.930 64.475 ;
        RECT 69.100 64.225 72.120 64.475 ;
        RECT 66.305 63.460 66.535 63.765 ;
        RECT 66.705 63.235 67.035 63.595 ;
        RECT 67.230 63.415 67.520 63.765 ;
        RECT 68.675 63.235 68.920 63.695 ;
        RECT 69.100 63.415 69.350 64.225 ;
        RECT 72.290 64.055 73.260 64.645 ;
        RECT 69.950 63.885 73.260 64.055 ;
        RECT 74.195 63.915 74.550 64.475 ;
        RECT 69.520 63.235 69.780 63.760 ;
        RECT 69.950 63.430 70.210 63.885 ;
        RECT 70.380 63.235 70.640 63.715 ;
        RECT 70.810 63.430 71.070 63.885 ;
        RECT 71.240 63.235 71.500 63.715 ;
        RECT 71.670 63.430 71.930 63.885 ;
        RECT 72.100 63.235 72.360 63.715 ;
        RECT 72.530 63.430 72.790 63.885 ;
        RECT 74.720 63.745 74.890 64.645 ;
        RECT 75.060 63.915 75.325 64.475 ;
        RECT 75.575 64.145 75.745 64.645 ;
        RECT 75.915 63.975 76.230 64.995 ;
        RECT 76.435 64.620 76.725 65.785 ;
        RECT 76.895 64.695 78.565 65.785 ;
        RECT 78.850 65.155 79.135 65.615 ;
        RECT 79.305 65.325 79.575 65.785 ;
        RECT 78.850 64.935 79.805 65.155 ;
        RECT 72.960 63.235 73.260 63.715 ;
        RECT 74.300 63.235 74.540 63.745 ;
        RECT 74.720 63.415 75.000 63.745 ;
        RECT 75.230 63.235 75.445 63.745 ;
        RECT 75.615 63.405 76.230 63.975 ;
        RECT 76.895 64.005 77.645 64.525 ;
        RECT 77.815 64.175 78.565 64.695 ;
        RECT 78.735 64.205 79.425 64.765 ;
        RECT 79.595 64.035 79.805 64.935 ;
        RECT 76.435 63.235 76.725 63.960 ;
        RECT 76.895 63.235 78.565 64.005 ;
        RECT 78.850 63.865 79.805 64.035 ;
        RECT 79.975 64.765 80.375 65.615 ;
        RECT 80.565 65.155 80.845 65.615 ;
        RECT 81.365 65.325 81.690 65.785 ;
        RECT 80.565 64.935 81.690 65.155 ;
        RECT 79.975 64.205 81.070 64.765 ;
        RECT 81.240 64.475 81.690 64.935 ;
        RECT 81.860 64.645 82.245 65.615 ;
        RECT 78.850 63.405 79.135 63.865 ;
        RECT 79.305 63.235 79.575 63.695 ;
        RECT 79.975 63.405 80.375 64.205 ;
        RECT 81.240 64.145 81.795 64.475 ;
        RECT 81.240 64.035 81.690 64.145 ;
        RECT 80.565 63.865 81.690 64.035 ;
        RECT 81.965 63.975 82.245 64.645 ;
        RECT 80.565 63.405 80.845 63.865 ;
        RECT 81.365 63.235 81.690 63.695 ;
        RECT 81.860 63.405 82.245 63.975 ;
        RECT 82.420 64.645 82.755 65.615 ;
        RECT 82.925 64.645 83.095 65.785 ;
        RECT 83.265 65.445 85.295 65.615 ;
        RECT 82.420 63.975 82.590 64.645 ;
        RECT 83.265 64.475 83.435 65.445 ;
        RECT 82.760 64.145 83.015 64.475 ;
        RECT 83.240 64.145 83.435 64.475 ;
        RECT 83.605 65.105 84.730 65.275 ;
        RECT 82.845 63.975 83.015 64.145 ;
        RECT 83.605 63.975 83.775 65.105 ;
        RECT 82.420 63.405 82.675 63.975 ;
        RECT 82.845 63.805 83.775 63.975 ;
        RECT 83.945 64.765 84.955 64.935 ;
        RECT 83.945 63.965 84.115 64.765 ;
        RECT 84.320 64.085 84.595 64.565 ;
        RECT 84.315 63.915 84.595 64.085 ;
        RECT 83.600 63.770 83.775 63.805 ;
        RECT 82.845 63.235 83.175 63.635 ;
        RECT 83.600 63.405 84.130 63.770 ;
        RECT 84.320 63.405 84.595 63.915 ;
        RECT 84.765 63.405 84.955 64.765 ;
        RECT 85.125 64.780 85.295 65.445 ;
        RECT 85.465 65.025 85.635 65.785 ;
        RECT 85.870 65.025 86.385 65.435 ;
        RECT 85.125 64.590 85.875 64.780 ;
        RECT 86.045 64.215 86.385 65.025 ;
        RECT 87.565 64.855 87.735 65.615 ;
        RECT 87.950 65.025 88.280 65.785 ;
        RECT 87.565 64.685 88.280 64.855 ;
        RECT 88.450 64.710 88.705 65.615 ;
        RECT 85.155 64.045 86.385 64.215 ;
        RECT 87.475 64.135 87.830 64.505 ;
        RECT 88.110 64.475 88.280 64.685 ;
        RECT 88.110 64.145 88.365 64.475 ;
        RECT 85.135 63.235 85.645 63.770 ;
        RECT 85.865 63.440 86.110 64.045 ;
        RECT 88.110 63.955 88.280 64.145 ;
        RECT 88.535 63.980 88.705 64.710 ;
        RECT 88.880 64.635 89.140 65.785 ;
        RECT 89.315 64.695 90.525 65.785 ;
        RECT 89.315 64.155 89.835 64.695 ;
        RECT 87.565 63.785 88.280 63.955 ;
        RECT 87.565 63.405 87.735 63.785 ;
        RECT 87.950 63.235 88.280 63.615 ;
        RECT 88.450 63.405 88.705 63.980 ;
        RECT 88.880 63.235 89.140 64.075 ;
        RECT 90.005 63.985 90.525 64.525 ;
        RECT 89.315 63.235 90.525 63.985 ;
        RECT 11.950 63.065 90.610 63.235 ;
        RECT 12.035 62.315 13.245 63.065 ;
        RECT 13.415 62.315 14.625 63.065 ;
        RECT 14.960 62.555 15.200 63.065 ;
        RECT 15.380 62.555 15.660 62.885 ;
        RECT 15.890 62.555 16.105 63.065 ;
        RECT 12.035 61.775 12.555 62.315 ;
        RECT 12.725 61.605 13.245 62.145 ;
        RECT 13.415 61.775 13.935 62.315 ;
        RECT 14.105 61.605 14.625 62.145 ;
        RECT 14.855 61.825 15.210 62.385 ;
        RECT 15.380 61.655 15.550 62.555 ;
        RECT 15.720 61.825 15.985 62.385 ;
        RECT 16.275 62.325 16.890 62.895 ;
        RECT 16.235 61.655 16.405 62.155 ;
        RECT 12.035 60.515 13.245 61.605 ;
        RECT 13.415 60.515 14.625 61.605 ;
        RECT 14.980 61.485 16.405 61.655 ;
        RECT 14.980 61.310 15.370 61.485 ;
        RECT 15.855 60.515 16.185 61.315 ;
        RECT 16.575 61.305 16.890 62.325 ;
        RECT 17.095 62.315 18.305 63.065 ;
        RECT 18.475 62.325 18.735 62.895 ;
        RECT 18.905 62.665 19.290 63.065 ;
        RECT 19.460 62.495 19.715 62.895 ;
        RECT 18.905 62.325 19.715 62.495 ;
        RECT 19.905 62.325 20.150 62.895 ;
        RECT 20.320 62.665 20.705 63.065 ;
        RECT 20.875 62.495 21.130 62.895 ;
        RECT 20.320 62.325 21.130 62.495 ;
        RECT 21.320 62.325 21.745 62.895 ;
        RECT 21.915 62.665 22.300 63.065 ;
        RECT 22.470 62.495 22.905 62.895 ;
        RECT 21.915 62.325 22.905 62.495 ;
        RECT 23.165 62.515 23.335 62.805 ;
        RECT 23.505 62.685 23.835 63.065 ;
        RECT 23.165 62.345 23.830 62.515 ;
        RECT 17.095 61.775 17.615 62.315 ;
        RECT 17.785 61.605 18.305 62.145 ;
        RECT 16.355 60.685 16.890 61.305 ;
        RECT 17.095 60.515 18.305 61.605 ;
        RECT 18.475 61.655 18.660 62.325 ;
        RECT 18.905 62.155 19.255 62.325 ;
        RECT 19.905 62.155 20.075 62.325 ;
        RECT 20.320 62.155 20.670 62.325 ;
        RECT 21.320 62.155 21.670 62.325 ;
        RECT 21.915 62.155 22.250 62.325 ;
        RECT 18.830 61.825 19.255 62.155 ;
        RECT 18.475 60.685 18.735 61.655 ;
        RECT 18.905 61.305 19.255 61.825 ;
        RECT 19.425 61.655 20.075 62.155 ;
        RECT 20.245 61.825 20.670 62.155 ;
        RECT 19.425 61.475 20.150 61.655 ;
        RECT 18.905 61.110 19.715 61.305 ;
        RECT 18.905 60.515 19.290 60.940 ;
        RECT 19.460 60.685 19.715 61.110 ;
        RECT 19.905 60.685 20.150 61.475 ;
        RECT 20.320 61.305 20.670 61.825 ;
        RECT 20.840 61.655 21.670 62.155 ;
        RECT 21.840 61.825 22.250 62.155 ;
        RECT 20.840 61.475 21.745 61.655 ;
        RECT 20.320 61.110 21.150 61.305 ;
        RECT 20.320 60.515 20.705 60.940 ;
        RECT 20.875 60.685 21.150 61.110 ;
        RECT 21.320 60.685 21.745 61.475 ;
        RECT 21.915 61.280 22.250 61.825 ;
        RECT 22.420 61.450 22.905 62.155 ;
        RECT 23.080 61.525 23.430 62.175 ;
        RECT 23.600 61.355 23.830 62.345 ;
        RECT 21.915 61.110 22.905 61.280 ;
        RECT 21.915 60.515 22.300 60.940 ;
        RECT 22.470 60.685 22.905 61.110 ;
        RECT 23.165 61.185 23.830 61.355 ;
        RECT 23.165 60.685 23.335 61.185 ;
        RECT 23.505 60.515 23.835 61.015 ;
        RECT 24.005 60.685 24.190 62.805 ;
        RECT 24.445 62.605 24.695 63.065 ;
        RECT 24.865 62.615 25.200 62.785 ;
        RECT 25.395 62.615 26.070 62.785 ;
        RECT 24.865 62.475 25.035 62.615 ;
        RECT 24.360 61.485 24.640 62.435 ;
        RECT 24.810 62.345 25.035 62.475 ;
        RECT 24.810 61.240 24.980 62.345 ;
        RECT 25.205 62.195 25.730 62.415 ;
        RECT 25.150 61.430 25.390 62.025 ;
        RECT 25.560 61.495 25.730 62.195 ;
        RECT 25.900 61.835 26.070 62.615 ;
        RECT 26.390 62.565 26.760 63.065 ;
        RECT 26.940 62.615 27.345 62.785 ;
        RECT 27.515 62.615 28.300 62.785 ;
        RECT 26.940 62.385 27.110 62.615 ;
        RECT 26.280 62.085 27.110 62.385 ;
        RECT 27.495 62.115 27.960 62.445 ;
        RECT 26.280 62.055 26.480 62.085 ;
        RECT 26.600 61.835 26.770 61.905 ;
        RECT 25.900 61.665 26.770 61.835 ;
        RECT 26.260 61.575 26.770 61.665 ;
        RECT 24.810 61.110 25.115 61.240 ;
        RECT 25.560 61.130 26.090 61.495 ;
        RECT 24.430 60.515 24.695 60.975 ;
        RECT 24.865 60.685 25.115 61.110 ;
        RECT 26.260 60.960 26.430 61.575 ;
        RECT 25.325 60.790 26.430 60.960 ;
        RECT 26.600 60.515 26.770 61.315 ;
        RECT 26.940 61.015 27.110 62.085 ;
        RECT 27.280 61.185 27.470 61.905 ;
        RECT 27.640 61.155 27.960 62.115 ;
        RECT 28.130 62.155 28.300 62.615 ;
        RECT 28.575 62.535 28.785 63.065 ;
        RECT 29.045 62.325 29.375 62.850 ;
        RECT 29.545 62.455 29.715 63.065 ;
        RECT 29.885 62.410 30.215 62.845 ;
        RECT 30.525 62.515 30.695 62.805 ;
        RECT 30.865 62.685 31.195 63.065 ;
        RECT 29.885 62.325 30.265 62.410 ;
        RECT 30.525 62.345 31.190 62.515 ;
        RECT 29.175 62.155 29.375 62.325 ;
        RECT 30.040 62.285 30.265 62.325 ;
        RECT 28.130 61.825 29.005 62.155 ;
        RECT 29.175 61.825 29.925 62.155 ;
        RECT 26.940 60.685 27.190 61.015 ;
        RECT 28.130 60.985 28.300 61.825 ;
        RECT 29.175 61.620 29.365 61.825 ;
        RECT 30.095 61.705 30.265 62.285 ;
        RECT 30.050 61.655 30.265 61.705 ;
        RECT 28.470 61.245 29.365 61.620 ;
        RECT 29.875 61.575 30.265 61.655 ;
        RECT 27.415 60.815 28.300 60.985 ;
        RECT 28.480 60.515 28.795 61.015 ;
        RECT 29.025 60.685 29.365 61.245 ;
        RECT 29.535 60.515 29.705 61.525 ;
        RECT 29.875 60.730 30.205 61.575 ;
        RECT 30.440 61.525 30.790 62.175 ;
        RECT 30.960 61.355 31.190 62.345 ;
        RECT 30.525 61.185 31.190 61.355 ;
        RECT 30.525 60.685 30.695 61.185 ;
        RECT 30.865 60.515 31.195 61.015 ;
        RECT 31.365 60.685 31.550 62.805 ;
        RECT 31.805 62.605 32.055 63.065 ;
        RECT 32.225 62.615 32.560 62.785 ;
        RECT 32.755 62.615 33.430 62.785 ;
        RECT 32.225 62.475 32.395 62.615 ;
        RECT 31.720 61.485 32.000 62.435 ;
        RECT 32.170 62.345 32.395 62.475 ;
        RECT 32.170 61.240 32.340 62.345 ;
        RECT 32.565 62.195 33.090 62.415 ;
        RECT 32.510 61.430 32.750 62.025 ;
        RECT 32.920 61.495 33.090 62.195 ;
        RECT 33.260 61.835 33.430 62.615 ;
        RECT 33.750 62.565 34.120 63.065 ;
        RECT 34.300 62.615 34.705 62.785 ;
        RECT 34.875 62.615 35.660 62.785 ;
        RECT 34.300 62.385 34.470 62.615 ;
        RECT 33.640 62.085 34.470 62.385 ;
        RECT 34.855 62.115 35.320 62.445 ;
        RECT 33.640 62.055 33.840 62.085 ;
        RECT 33.960 61.835 34.130 61.905 ;
        RECT 33.260 61.665 34.130 61.835 ;
        RECT 33.620 61.575 34.130 61.665 ;
        RECT 32.170 61.110 32.475 61.240 ;
        RECT 32.920 61.130 33.450 61.495 ;
        RECT 31.790 60.515 32.055 60.975 ;
        RECT 32.225 60.685 32.475 61.110 ;
        RECT 33.620 60.960 33.790 61.575 ;
        RECT 32.685 60.790 33.790 60.960 ;
        RECT 33.960 60.515 34.130 61.315 ;
        RECT 34.300 61.015 34.470 62.085 ;
        RECT 34.640 61.185 34.830 61.905 ;
        RECT 35.000 61.155 35.320 62.115 ;
        RECT 35.490 62.155 35.660 62.615 ;
        RECT 35.935 62.535 36.145 63.065 ;
        RECT 36.405 62.325 36.735 62.850 ;
        RECT 36.905 62.455 37.075 63.065 ;
        RECT 37.245 62.410 37.575 62.845 ;
        RECT 37.245 62.325 37.625 62.410 ;
        RECT 37.795 62.340 38.085 63.065 ;
        RECT 36.535 62.155 36.735 62.325 ;
        RECT 37.400 62.285 37.625 62.325 ;
        RECT 35.490 61.825 36.365 62.155 ;
        RECT 36.535 61.825 37.285 62.155 ;
        RECT 34.300 60.685 34.550 61.015 ;
        RECT 35.490 60.985 35.660 61.825 ;
        RECT 36.535 61.620 36.725 61.825 ;
        RECT 37.455 61.705 37.625 62.285 ;
        RECT 38.255 62.295 40.845 63.065 ;
        RECT 41.105 62.515 41.275 62.805 ;
        RECT 41.445 62.685 41.775 63.065 ;
        RECT 41.105 62.345 41.770 62.515 ;
        RECT 38.255 61.775 39.465 62.295 ;
        RECT 37.410 61.655 37.625 61.705 ;
        RECT 35.830 61.245 36.725 61.620 ;
        RECT 37.235 61.575 37.625 61.655 ;
        RECT 34.775 60.815 35.660 60.985 ;
        RECT 35.840 60.515 36.155 61.015 ;
        RECT 36.385 60.685 36.725 61.245 ;
        RECT 36.895 60.515 37.065 61.525 ;
        RECT 37.235 60.730 37.565 61.575 ;
        RECT 37.795 60.515 38.085 61.680 ;
        RECT 39.635 61.605 40.845 62.125 ;
        RECT 38.255 60.515 40.845 61.605 ;
        RECT 41.020 61.525 41.370 62.175 ;
        RECT 41.540 61.355 41.770 62.345 ;
        RECT 41.105 61.185 41.770 61.355 ;
        RECT 41.105 60.685 41.275 61.185 ;
        RECT 41.445 60.515 41.775 61.015 ;
        RECT 41.945 60.685 42.130 62.805 ;
        RECT 42.385 62.605 42.635 63.065 ;
        RECT 42.805 62.615 43.140 62.785 ;
        RECT 43.335 62.615 44.010 62.785 ;
        RECT 42.805 62.475 42.975 62.615 ;
        RECT 42.300 61.485 42.580 62.435 ;
        RECT 42.750 62.345 42.975 62.475 ;
        RECT 42.750 61.240 42.920 62.345 ;
        RECT 43.145 62.195 43.670 62.415 ;
        RECT 43.090 61.430 43.330 62.025 ;
        RECT 43.500 61.495 43.670 62.195 ;
        RECT 43.840 61.835 44.010 62.615 ;
        RECT 44.330 62.565 44.700 63.065 ;
        RECT 44.880 62.615 45.285 62.785 ;
        RECT 45.455 62.615 46.240 62.785 ;
        RECT 44.880 62.385 45.050 62.615 ;
        RECT 44.220 62.085 45.050 62.385 ;
        RECT 45.435 62.115 45.900 62.445 ;
        RECT 44.220 62.055 44.420 62.085 ;
        RECT 44.540 61.835 44.710 61.905 ;
        RECT 43.840 61.665 44.710 61.835 ;
        RECT 44.200 61.575 44.710 61.665 ;
        RECT 42.750 61.110 43.055 61.240 ;
        RECT 43.500 61.130 44.030 61.495 ;
        RECT 42.370 60.515 42.635 60.975 ;
        RECT 42.805 60.685 43.055 61.110 ;
        RECT 44.200 60.960 44.370 61.575 ;
        RECT 43.265 60.790 44.370 60.960 ;
        RECT 44.540 60.515 44.710 61.315 ;
        RECT 44.880 61.015 45.050 62.085 ;
        RECT 45.220 61.185 45.410 61.905 ;
        RECT 45.580 61.155 45.900 62.115 ;
        RECT 46.070 62.155 46.240 62.615 ;
        RECT 46.515 62.535 46.725 63.065 ;
        RECT 46.985 62.325 47.315 62.850 ;
        RECT 47.485 62.455 47.655 63.065 ;
        RECT 47.825 62.410 48.155 62.845 ;
        RECT 47.825 62.325 48.205 62.410 ;
        RECT 47.115 62.155 47.315 62.325 ;
        RECT 47.980 62.285 48.205 62.325 ;
        RECT 46.070 61.825 46.945 62.155 ;
        RECT 47.115 61.825 47.865 62.155 ;
        RECT 44.880 60.685 45.130 61.015 ;
        RECT 46.070 60.985 46.240 61.825 ;
        RECT 47.115 61.620 47.305 61.825 ;
        RECT 48.035 61.705 48.205 62.285 ;
        RECT 48.375 62.295 50.045 63.065 ;
        RECT 48.375 61.775 49.125 62.295 ;
        RECT 50.490 62.255 50.735 62.860 ;
        RECT 50.955 62.530 51.465 63.065 ;
        RECT 47.990 61.655 48.205 61.705 ;
        RECT 46.410 61.245 47.305 61.620 ;
        RECT 47.815 61.575 48.205 61.655 ;
        RECT 49.295 61.605 50.045 62.125 ;
        RECT 45.355 60.815 46.240 60.985 ;
        RECT 46.420 60.515 46.735 61.015 ;
        RECT 46.965 60.685 47.305 61.245 ;
        RECT 47.475 60.515 47.645 61.525 ;
        RECT 47.815 60.730 48.145 61.575 ;
        RECT 48.375 60.515 50.045 61.605 ;
        RECT 50.215 62.085 51.445 62.255 ;
        RECT 50.215 61.275 50.555 62.085 ;
        RECT 50.725 61.520 51.475 61.710 ;
        RECT 50.215 60.865 50.730 61.275 ;
        RECT 50.965 60.515 51.135 61.275 ;
        RECT 51.305 60.855 51.475 61.520 ;
        RECT 51.645 61.535 51.835 62.895 ;
        RECT 52.005 62.385 52.280 62.895 ;
        RECT 52.470 62.530 53.000 62.895 ;
        RECT 53.425 62.665 53.755 63.065 ;
        RECT 52.825 62.495 53.000 62.530 ;
        RECT 52.005 62.215 52.285 62.385 ;
        RECT 52.005 61.735 52.280 62.215 ;
        RECT 52.485 61.535 52.655 62.335 ;
        RECT 51.645 61.365 52.655 61.535 ;
        RECT 52.825 62.325 53.755 62.495 ;
        RECT 53.925 62.325 54.180 62.895 ;
        RECT 52.825 61.195 52.995 62.325 ;
        RECT 53.585 62.155 53.755 62.325 ;
        RECT 51.870 61.025 52.995 61.195 ;
        RECT 53.165 61.825 53.360 62.155 ;
        RECT 53.585 61.825 53.840 62.155 ;
        RECT 53.165 60.855 53.335 61.825 ;
        RECT 54.010 61.655 54.180 62.325 ;
        RECT 54.355 62.295 56.025 63.065 ;
        RECT 56.245 62.410 56.575 62.845 ;
        RECT 56.745 62.455 56.915 63.065 ;
        RECT 56.195 62.325 56.575 62.410 ;
        RECT 57.085 62.325 57.415 62.850 ;
        RECT 57.675 62.535 57.885 63.065 ;
        RECT 58.160 62.615 58.945 62.785 ;
        RECT 59.115 62.615 59.520 62.785 ;
        RECT 54.355 61.775 55.105 62.295 ;
        RECT 56.195 62.285 56.420 62.325 ;
        RECT 51.305 60.685 53.335 60.855 ;
        RECT 53.505 60.515 53.675 61.655 ;
        RECT 53.845 60.685 54.180 61.655 ;
        RECT 55.275 61.605 56.025 62.125 ;
        RECT 54.355 60.515 56.025 61.605 ;
        RECT 56.195 61.705 56.365 62.285 ;
        RECT 57.085 62.155 57.285 62.325 ;
        RECT 58.160 62.155 58.330 62.615 ;
        RECT 56.535 61.825 57.285 62.155 ;
        RECT 57.455 61.825 58.330 62.155 ;
        RECT 56.195 61.655 56.410 61.705 ;
        RECT 56.195 61.575 56.585 61.655 ;
        RECT 56.255 60.730 56.585 61.575 ;
        RECT 57.095 61.620 57.285 61.825 ;
        RECT 56.755 60.515 56.925 61.525 ;
        RECT 57.095 61.245 57.990 61.620 ;
        RECT 57.095 60.685 57.435 61.245 ;
        RECT 57.665 60.515 57.980 61.015 ;
        RECT 58.160 60.985 58.330 61.825 ;
        RECT 58.500 62.115 58.965 62.445 ;
        RECT 59.350 62.385 59.520 62.615 ;
        RECT 59.700 62.565 60.070 63.065 ;
        RECT 60.390 62.615 61.065 62.785 ;
        RECT 61.260 62.615 61.595 62.785 ;
        RECT 58.500 61.155 58.820 62.115 ;
        RECT 59.350 62.085 60.180 62.385 ;
        RECT 58.990 61.185 59.180 61.905 ;
        RECT 59.350 61.015 59.520 62.085 ;
        RECT 59.980 62.055 60.180 62.085 ;
        RECT 59.690 61.835 59.860 61.905 ;
        RECT 60.390 61.835 60.560 62.615 ;
        RECT 61.425 62.475 61.595 62.615 ;
        RECT 61.765 62.605 62.015 63.065 ;
        RECT 59.690 61.665 60.560 61.835 ;
        RECT 60.730 62.195 61.255 62.415 ;
        RECT 61.425 62.345 61.650 62.475 ;
        RECT 59.690 61.575 60.200 61.665 ;
        RECT 58.160 60.815 59.045 60.985 ;
        RECT 59.270 60.685 59.520 61.015 ;
        RECT 59.690 60.515 59.860 61.315 ;
        RECT 60.030 60.960 60.200 61.575 ;
        RECT 60.730 61.495 60.900 62.195 ;
        RECT 60.370 61.130 60.900 61.495 ;
        RECT 61.070 61.430 61.310 62.025 ;
        RECT 61.480 61.240 61.650 62.345 ;
        RECT 61.820 61.485 62.100 62.435 ;
        RECT 61.345 61.110 61.650 61.240 ;
        RECT 60.030 60.790 61.135 60.960 ;
        RECT 61.345 60.685 61.595 61.110 ;
        RECT 61.765 60.515 62.030 60.975 ;
        RECT 62.270 60.685 62.455 62.805 ;
        RECT 62.625 62.685 62.955 63.065 ;
        RECT 63.125 62.515 63.295 62.805 ;
        RECT 62.630 62.345 63.295 62.515 ;
        RECT 62.630 61.355 62.860 62.345 ;
        RECT 63.555 62.340 63.845 63.065 ;
        RECT 64.015 62.565 64.275 62.895 ;
        RECT 64.445 62.705 64.775 63.065 ;
        RECT 65.030 62.685 66.330 62.895 ;
        RECT 64.015 62.555 64.245 62.565 ;
        RECT 63.030 61.525 63.380 62.175 ;
        RECT 62.630 61.185 63.295 61.355 ;
        RECT 62.625 60.515 62.955 61.015 ;
        RECT 63.125 60.685 63.295 61.185 ;
        RECT 63.555 60.515 63.845 61.680 ;
        RECT 64.015 61.365 64.185 62.555 ;
        RECT 65.030 62.535 65.200 62.685 ;
        RECT 64.445 62.410 65.200 62.535 ;
        RECT 64.355 62.365 65.200 62.410 ;
        RECT 64.355 62.245 64.625 62.365 ;
        RECT 64.355 61.670 64.525 62.245 ;
        RECT 64.755 61.805 65.165 62.110 ;
        RECT 65.455 62.075 65.665 62.475 ;
        RECT 65.335 61.865 65.665 62.075 ;
        RECT 65.910 62.075 66.130 62.475 ;
        RECT 66.605 62.300 67.060 63.065 ;
        RECT 67.235 62.265 67.930 62.895 ;
        RECT 68.135 62.265 68.445 63.065 ;
        RECT 68.625 62.415 68.955 62.890 ;
        RECT 69.125 62.585 69.295 63.065 ;
        RECT 69.465 62.415 69.795 62.890 ;
        RECT 69.965 62.585 70.135 63.065 ;
        RECT 70.305 62.415 70.635 62.890 ;
        RECT 70.805 62.585 70.975 63.065 ;
        RECT 71.145 62.415 71.475 62.890 ;
        RECT 71.645 62.585 71.815 63.065 ;
        RECT 71.985 62.415 72.315 62.890 ;
        RECT 72.485 62.585 72.655 63.065 ;
        RECT 72.825 62.890 73.075 62.895 ;
        RECT 72.825 62.415 73.155 62.890 ;
        RECT 73.325 62.585 73.495 63.065 ;
        RECT 73.745 62.890 73.915 62.895 ;
        RECT 73.665 62.415 73.995 62.890 ;
        RECT 74.165 62.585 74.335 63.065 ;
        RECT 74.585 62.890 74.755 62.895 ;
        RECT 74.505 62.415 74.835 62.890 ;
        RECT 75.005 62.585 75.175 63.065 ;
        RECT 75.345 62.415 75.675 62.890 ;
        RECT 75.845 62.585 76.015 63.065 ;
        RECT 76.185 62.415 76.515 62.890 ;
        RECT 76.685 62.585 76.855 63.065 ;
        RECT 77.025 62.415 77.355 62.890 ;
        RECT 77.525 62.585 77.695 63.065 ;
        RECT 77.865 62.415 78.195 62.890 ;
        RECT 78.365 62.585 78.535 63.065 ;
        RECT 78.705 62.415 79.035 62.890 ;
        RECT 79.205 62.585 79.375 63.065 ;
        RECT 65.910 61.865 66.385 62.075 ;
        RECT 66.575 61.875 67.065 62.075 ;
        RECT 67.255 61.825 67.590 62.075 ;
        RECT 64.355 61.635 64.555 61.670 ;
        RECT 65.885 61.635 67.060 61.695 ;
        RECT 67.760 61.665 67.930 62.265 ;
        RECT 68.625 62.245 70.135 62.415 ;
        RECT 70.305 62.245 72.655 62.415 ;
        RECT 72.825 62.245 79.485 62.415 ;
        RECT 79.655 62.265 79.965 63.065 ;
        RECT 80.170 62.265 80.865 62.895 ;
        RECT 81.960 62.325 82.215 62.895 ;
        RECT 82.385 62.665 82.715 63.065 ;
        RECT 83.140 62.530 83.670 62.895 ;
        RECT 83.860 62.725 84.135 62.895 ;
        RECT 83.855 62.555 84.135 62.725 ;
        RECT 83.140 62.495 83.315 62.530 ;
        RECT 82.385 62.325 83.315 62.495 ;
        RECT 68.100 61.825 68.435 62.095 ;
        RECT 69.965 62.075 70.135 62.245 ;
        RECT 72.480 62.075 72.655 62.245 ;
        RECT 68.620 61.875 69.795 62.075 ;
        RECT 69.965 61.875 72.275 62.075 ;
        RECT 72.480 61.875 79.040 62.075 ;
        RECT 69.965 61.705 70.135 61.875 ;
        RECT 72.480 61.705 72.655 61.875 ;
        RECT 79.210 61.705 79.485 62.245 ;
        RECT 79.665 61.825 80.000 62.095 ;
        RECT 64.355 61.525 67.060 61.635 ;
        RECT 64.415 61.465 66.215 61.525 ;
        RECT 65.885 61.435 66.215 61.465 ;
        RECT 64.015 60.685 64.275 61.365 ;
        RECT 64.445 60.515 64.695 61.295 ;
        RECT 64.945 61.265 65.780 61.275 ;
        RECT 66.370 61.265 66.555 61.355 ;
        RECT 64.945 61.065 66.555 61.265 ;
        RECT 64.945 60.685 65.195 61.065 ;
        RECT 66.325 61.025 66.555 61.065 ;
        RECT 66.805 60.905 67.060 61.525 ;
        RECT 65.365 60.515 65.720 60.895 ;
        RECT 66.725 60.685 67.060 60.905 ;
        RECT 67.235 60.515 67.495 61.655 ;
        RECT 67.665 60.685 67.995 61.665 ;
        RECT 68.165 60.515 68.445 61.655 ;
        RECT 68.625 61.535 70.135 61.705 ;
        RECT 70.305 61.535 72.655 61.705 ;
        RECT 72.825 61.535 79.485 61.705 ;
        RECT 80.170 61.665 80.340 62.265 ;
        RECT 80.510 61.825 80.845 62.075 ;
        RECT 68.625 60.685 68.955 61.535 ;
        RECT 69.125 60.515 69.295 61.365 ;
        RECT 69.465 60.685 69.795 61.535 ;
        RECT 69.965 60.515 70.135 61.365 ;
        RECT 70.305 60.685 70.635 61.535 ;
        RECT 70.805 60.515 70.975 61.315 ;
        RECT 71.145 60.685 71.475 61.535 ;
        RECT 71.645 60.515 71.815 61.315 ;
        RECT 71.985 60.685 72.315 61.535 ;
        RECT 72.485 60.515 72.655 61.315 ;
        RECT 72.825 60.685 73.155 61.535 ;
        RECT 73.325 60.515 73.495 61.315 ;
        RECT 73.665 60.685 73.995 61.535 ;
        RECT 74.165 60.515 74.335 61.315 ;
        RECT 74.505 60.685 74.835 61.535 ;
        RECT 75.005 60.515 75.175 61.315 ;
        RECT 75.345 60.685 75.675 61.535 ;
        RECT 75.845 60.515 76.015 61.315 ;
        RECT 76.185 60.685 76.515 61.535 ;
        RECT 76.685 60.515 76.855 61.315 ;
        RECT 77.025 60.685 77.355 61.535 ;
        RECT 77.525 60.515 77.695 61.315 ;
        RECT 77.865 60.685 78.195 61.535 ;
        RECT 78.365 60.515 78.535 61.315 ;
        RECT 78.705 60.685 79.035 61.535 ;
        RECT 79.205 60.515 79.375 61.315 ;
        RECT 79.655 60.515 79.935 61.655 ;
        RECT 80.105 60.685 80.435 61.665 ;
        RECT 81.960 61.655 82.130 62.325 ;
        RECT 82.385 62.155 82.555 62.325 ;
        RECT 82.300 61.825 82.555 62.155 ;
        RECT 82.780 61.825 82.975 62.155 ;
        RECT 80.605 60.515 80.865 61.655 ;
        RECT 81.960 60.685 82.295 61.655 ;
        RECT 82.465 60.515 82.635 61.655 ;
        RECT 82.805 60.855 82.975 61.825 ;
        RECT 83.145 61.195 83.315 62.325 ;
        RECT 83.485 61.535 83.655 62.335 ;
        RECT 83.860 61.735 84.135 62.555 ;
        RECT 84.305 61.535 84.495 62.895 ;
        RECT 84.675 62.530 85.185 63.065 ;
        RECT 85.405 62.255 85.650 62.860 ;
        RECT 86.095 62.390 86.355 62.895 ;
        RECT 86.535 62.685 86.865 63.065 ;
        RECT 87.045 62.515 87.215 62.895 ;
        RECT 84.695 62.085 85.925 62.255 ;
        RECT 83.485 61.365 84.495 61.535 ;
        RECT 84.665 61.520 85.415 61.710 ;
        RECT 83.145 61.025 84.270 61.195 ;
        RECT 84.665 60.855 84.835 61.520 ;
        RECT 85.585 61.275 85.925 62.085 ;
        RECT 82.805 60.685 84.835 60.855 ;
        RECT 85.005 60.515 85.175 61.275 ;
        RECT 85.410 60.865 85.925 61.275 ;
        RECT 86.095 61.590 86.265 62.390 ;
        RECT 86.550 62.345 87.215 62.515 ;
        RECT 87.565 62.515 87.735 62.895 ;
        RECT 87.950 62.685 88.280 63.065 ;
        RECT 87.565 62.345 88.280 62.515 ;
        RECT 86.550 62.090 86.720 62.345 ;
        RECT 86.435 61.760 86.720 62.090 ;
        RECT 86.955 61.795 87.285 62.165 ;
        RECT 87.475 61.795 87.830 62.165 ;
        RECT 88.110 62.155 88.280 62.345 ;
        RECT 88.450 62.320 88.705 62.895 ;
        RECT 88.110 61.825 88.365 62.155 ;
        RECT 86.550 61.615 86.720 61.760 ;
        RECT 88.110 61.615 88.280 61.825 ;
        RECT 86.095 60.685 86.365 61.590 ;
        RECT 86.550 61.445 87.215 61.615 ;
        RECT 86.535 60.515 86.865 61.275 ;
        RECT 87.045 60.685 87.215 61.445 ;
        RECT 87.565 61.445 88.280 61.615 ;
        RECT 88.535 61.590 88.705 62.320 ;
        RECT 88.880 62.225 89.140 63.065 ;
        RECT 89.315 62.315 90.525 63.065 ;
        RECT 87.565 60.685 87.735 61.445 ;
        RECT 87.950 60.515 88.280 61.275 ;
        RECT 88.450 60.685 88.705 61.590 ;
        RECT 88.880 60.515 89.140 61.665 ;
        RECT 89.315 61.605 89.835 62.145 ;
        RECT 90.005 61.775 90.525 62.315 ;
        RECT 89.315 60.515 90.525 61.605 ;
        RECT 11.950 60.345 90.610 60.515 ;
        RECT 12.035 59.255 13.245 60.345 ;
        RECT 12.035 58.545 12.555 59.085 ;
        RECT 12.725 58.715 13.245 59.255 ;
        RECT 13.420 59.195 13.680 60.345 ;
        RECT 13.855 59.270 14.110 60.175 ;
        RECT 14.280 59.585 14.610 60.345 ;
        RECT 14.825 59.415 14.995 60.175 ;
        RECT 15.345 59.675 15.515 60.175 ;
        RECT 15.685 59.845 16.015 60.345 ;
        RECT 15.345 59.505 16.010 59.675 ;
        RECT 12.035 57.795 13.245 58.545 ;
        RECT 13.420 57.795 13.680 58.635 ;
        RECT 13.855 58.540 14.025 59.270 ;
        RECT 14.280 59.245 14.995 59.415 ;
        RECT 14.280 59.035 14.450 59.245 ;
        RECT 14.195 58.705 14.450 59.035 ;
        RECT 13.855 57.965 14.110 58.540 ;
        RECT 14.280 58.515 14.450 58.705 ;
        RECT 14.730 58.695 15.085 59.065 ;
        RECT 15.260 58.685 15.610 59.335 ;
        RECT 15.780 58.515 16.010 59.505 ;
        RECT 14.280 58.345 14.995 58.515 ;
        RECT 14.280 57.795 14.610 58.175 ;
        RECT 14.825 57.965 14.995 58.345 ;
        RECT 15.345 58.345 16.010 58.515 ;
        RECT 15.345 58.055 15.515 58.345 ;
        RECT 15.685 57.795 16.015 58.175 ;
        RECT 16.185 58.055 16.370 60.175 ;
        RECT 16.610 59.885 16.875 60.345 ;
        RECT 17.045 59.750 17.295 60.175 ;
        RECT 17.505 59.900 18.610 60.070 ;
        RECT 16.990 59.620 17.295 59.750 ;
        RECT 16.540 58.425 16.820 59.375 ;
        RECT 16.990 58.515 17.160 59.620 ;
        RECT 17.330 58.835 17.570 59.430 ;
        RECT 17.740 59.365 18.270 59.730 ;
        RECT 17.740 58.665 17.910 59.365 ;
        RECT 18.440 59.285 18.610 59.900 ;
        RECT 18.780 59.545 18.950 60.345 ;
        RECT 19.120 59.845 19.370 60.175 ;
        RECT 19.595 59.875 20.480 60.045 ;
        RECT 18.440 59.195 18.950 59.285 ;
        RECT 16.990 58.385 17.215 58.515 ;
        RECT 17.385 58.445 17.910 58.665 ;
        RECT 18.080 59.025 18.950 59.195 ;
        RECT 16.625 57.795 16.875 58.255 ;
        RECT 17.045 58.245 17.215 58.385 ;
        RECT 18.080 58.245 18.250 59.025 ;
        RECT 18.780 58.955 18.950 59.025 ;
        RECT 18.460 58.775 18.660 58.805 ;
        RECT 19.120 58.775 19.290 59.845 ;
        RECT 19.460 58.955 19.650 59.675 ;
        RECT 18.460 58.475 19.290 58.775 ;
        RECT 19.820 58.745 20.140 59.705 ;
        RECT 17.045 58.075 17.380 58.245 ;
        RECT 17.575 58.075 18.250 58.245 ;
        RECT 18.570 57.795 18.940 58.295 ;
        RECT 19.120 58.245 19.290 58.475 ;
        RECT 19.675 58.415 20.140 58.745 ;
        RECT 20.310 59.035 20.480 59.875 ;
        RECT 20.660 59.845 20.975 60.345 ;
        RECT 21.205 59.615 21.545 60.175 ;
        RECT 20.650 59.240 21.545 59.615 ;
        RECT 21.715 59.335 21.885 60.345 ;
        RECT 21.355 59.035 21.545 59.240 ;
        RECT 22.055 59.285 22.385 60.130 ;
        RECT 22.055 59.205 22.445 59.285 ;
        RECT 22.615 59.255 24.285 60.345 ;
        RECT 22.230 59.155 22.445 59.205 ;
        RECT 20.310 58.705 21.185 59.035 ;
        RECT 21.355 58.705 22.105 59.035 ;
        RECT 20.310 58.245 20.480 58.705 ;
        RECT 21.355 58.535 21.555 58.705 ;
        RECT 22.275 58.575 22.445 59.155 ;
        RECT 22.220 58.535 22.445 58.575 ;
        RECT 19.120 58.075 19.525 58.245 ;
        RECT 19.695 58.075 20.480 58.245 ;
        RECT 20.755 57.795 20.965 58.325 ;
        RECT 21.225 58.010 21.555 58.535 ;
        RECT 22.065 58.450 22.445 58.535 ;
        RECT 22.615 58.565 23.365 59.085 ;
        RECT 23.535 58.735 24.285 59.255 ;
        RECT 24.915 59.180 25.205 60.345 ;
        RECT 25.560 59.375 25.950 59.550 ;
        RECT 26.435 59.545 26.765 60.345 ;
        RECT 26.935 59.555 27.470 60.175 ;
        RECT 25.560 59.205 26.985 59.375 ;
        RECT 21.725 57.795 21.895 58.405 ;
        RECT 22.065 58.015 22.395 58.450 ;
        RECT 22.615 57.795 24.285 58.565 ;
        RECT 24.915 57.795 25.205 58.520 ;
        RECT 25.435 58.475 25.790 59.035 ;
        RECT 25.960 58.305 26.130 59.205 ;
        RECT 26.300 58.475 26.565 59.035 ;
        RECT 26.815 58.705 26.985 59.205 ;
        RECT 27.155 58.535 27.470 59.555 ;
        RECT 28.340 59.375 28.670 60.175 ;
        RECT 28.840 59.545 29.170 60.345 ;
        RECT 29.470 59.375 29.800 60.175 ;
        RECT 30.445 59.545 30.695 60.345 ;
        RECT 28.340 59.205 30.775 59.375 ;
        RECT 30.965 59.205 31.135 60.345 ;
        RECT 31.305 59.205 31.645 60.175 ;
        RECT 31.815 59.255 33.485 60.345 ;
        RECT 33.745 59.675 33.915 60.175 ;
        RECT 34.085 59.845 34.415 60.345 ;
        RECT 33.745 59.505 34.410 59.675 ;
        RECT 28.135 58.785 28.485 59.035 ;
        RECT 28.670 58.575 28.840 59.205 ;
        RECT 29.010 58.785 29.340 58.985 ;
        RECT 29.510 58.785 29.840 58.985 ;
        RECT 30.010 58.785 30.430 58.985 ;
        RECT 30.605 58.955 30.775 59.205 ;
        RECT 30.605 58.785 31.300 58.955 ;
        RECT 25.540 57.795 25.780 58.305 ;
        RECT 25.960 57.975 26.240 58.305 ;
        RECT 26.470 57.795 26.685 58.305 ;
        RECT 26.855 57.965 27.470 58.535 ;
        RECT 28.340 57.965 28.840 58.575 ;
        RECT 29.470 58.445 30.695 58.615 ;
        RECT 31.470 58.595 31.645 59.205 ;
        RECT 29.470 57.965 29.800 58.445 ;
        RECT 29.970 57.795 30.195 58.255 ;
        RECT 30.365 57.965 30.695 58.445 ;
        RECT 30.885 57.795 31.135 58.595 ;
        RECT 31.305 57.965 31.645 58.595 ;
        RECT 31.815 58.565 32.565 59.085 ;
        RECT 32.735 58.735 33.485 59.255 ;
        RECT 33.660 58.685 34.010 59.335 ;
        RECT 31.815 57.795 33.485 58.565 ;
        RECT 34.180 58.515 34.410 59.505 ;
        RECT 33.745 58.345 34.410 58.515 ;
        RECT 33.745 58.055 33.915 58.345 ;
        RECT 34.085 57.795 34.415 58.175 ;
        RECT 34.585 58.055 34.770 60.175 ;
        RECT 35.010 59.885 35.275 60.345 ;
        RECT 35.445 59.750 35.695 60.175 ;
        RECT 35.905 59.900 37.010 60.070 ;
        RECT 35.390 59.620 35.695 59.750 ;
        RECT 34.940 58.425 35.220 59.375 ;
        RECT 35.390 58.515 35.560 59.620 ;
        RECT 35.730 58.835 35.970 59.430 ;
        RECT 36.140 59.365 36.670 59.730 ;
        RECT 36.140 58.665 36.310 59.365 ;
        RECT 36.840 59.285 37.010 59.900 ;
        RECT 37.180 59.545 37.350 60.345 ;
        RECT 37.520 59.845 37.770 60.175 ;
        RECT 37.995 59.875 38.880 60.045 ;
        RECT 36.840 59.195 37.350 59.285 ;
        RECT 35.390 58.385 35.615 58.515 ;
        RECT 35.785 58.445 36.310 58.665 ;
        RECT 36.480 59.025 37.350 59.195 ;
        RECT 35.025 57.795 35.275 58.255 ;
        RECT 35.445 58.245 35.615 58.385 ;
        RECT 36.480 58.245 36.650 59.025 ;
        RECT 37.180 58.955 37.350 59.025 ;
        RECT 36.860 58.775 37.060 58.805 ;
        RECT 37.520 58.775 37.690 59.845 ;
        RECT 37.860 58.955 38.050 59.675 ;
        RECT 36.860 58.475 37.690 58.775 ;
        RECT 38.220 58.745 38.540 59.705 ;
        RECT 35.445 58.075 35.780 58.245 ;
        RECT 35.975 58.075 36.650 58.245 ;
        RECT 36.970 57.795 37.340 58.295 ;
        RECT 37.520 58.245 37.690 58.475 ;
        RECT 38.075 58.415 38.540 58.745 ;
        RECT 38.710 59.035 38.880 59.875 ;
        RECT 39.060 59.845 39.375 60.345 ;
        RECT 39.605 59.615 39.945 60.175 ;
        RECT 39.050 59.240 39.945 59.615 ;
        RECT 40.115 59.335 40.285 60.345 ;
        RECT 39.755 59.035 39.945 59.240 ;
        RECT 40.455 59.285 40.785 60.130 ;
        RECT 40.455 59.205 40.845 59.285 ;
        RECT 40.630 59.155 40.845 59.205 ;
        RECT 38.710 58.705 39.585 59.035 ;
        RECT 39.755 58.705 40.505 59.035 ;
        RECT 38.710 58.245 38.880 58.705 ;
        RECT 39.755 58.535 39.955 58.705 ;
        RECT 40.675 58.575 40.845 59.155 ;
        RECT 40.620 58.535 40.845 58.575 ;
        RECT 37.520 58.075 37.925 58.245 ;
        RECT 38.095 58.075 38.880 58.245 ;
        RECT 39.155 57.795 39.365 58.325 ;
        RECT 39.625 58.010 39.955 58.535 ;
        RECT 40.465 58.450 40.845 58.535 ;
        RECT 41.020 59.205 41.355 60.175 ;
        RECT 41.525 59.205 41.695 60.345 ;
        RECT 41.865 60.005 43.895 60.175 ;
        RECT 41.020 58.535 41.190 59.205 ;
        RECT 41.865 59.035 42.035 60.005 ;
        RECT 41.360 58.705 41.615 59.035 ;
        RECT 41.840 58.705 42.035 59.035 ;
        RECT 42.205 59.665 43.330 59.835 ;
        RECT 41.445 58.535 41.615 58.705 ;
        RECT 42.205 58.535 42.375 59.665 ;
        RECT 40.125 57.795 40.295 58.405 ;
        RECT 40.465 58.015 40.795 58.450 ;
        RECT 41.020 57.965 41.275 58.535 ;
        RECT 41.445 58.365 42.375 58.535 ;
        RECT 42.545 59.325 43.555 59.495 ;
        RECT 42.545 58.525 42.715 59.325 ;
        RECT 42.200 58.330 42.375 58.365 ;
        RECT 41.445 57.795 41.775 58.195 ;
        RECT 42.200 57.965 42.730 58.330 ;
        RECT 42.920 58.305 43.195 59.125 ;
        RECT 42.915 58.135 43.195 58.305 ;
        RECT 42.920 57.965 43.195 58.135 ;
        RECT 43.365 57.965 43.555 59.325 ;
        RECT 43.725 59.340 43.895 60.005 ;
        RECT 44.065 59.585 44.235 60.345 ;
        RECT 44.470 59.585 44.985 59.995 ;
        RECT 43.725 59.150 44.475 59.340 ;
        RECT 44.645 58.775 44.985 59.585 ;
        RECT 43.755 58.605 44.985 58.775 ;
        RECT 45.615 59.585 46.130 59.995 ;
        RECT 46.365 59.585 46.535 60.345 ;
        RECT 46.705 60.005 48.735 60.175 ;
        RECT 45.615 58.775 45.955 59.585 ;
        RECT 46.705 59.340 46.875 60.005 ;
        RECT 47.270 59.665 48.395 59.835 ;
        RECT 46.125 59.150 46.875 59.340 ;
        RECT 47.045 59.325 48.055 59.495 ;
        RECT 45.615 58.605 46.845 58.775 ;
        RECT 43.735 57.795 44.245 58.330 ;
        RECT 44.465 58.000 44.710 58.605 ;
        RECT 45.890 58.000 46.135 58.605 ;
        RECT 46.355 57.795 46.865 58.330 ;
        RECT 47.045 57.965 47.235 59.325 ;
        RECT 47.405 58.985 47.680 59.125 ;
        RECT 47.405 58.815 47.685 58.985 ;
        RECT 47.405 57.965 47.680 58.815 ;
        RECT 47.885 58.525 48.055 59.325 ;
        RECT 48.225 58.535 48.395 59.665 ;
        RECT 48.565 59.035 48.735 60.005 ;
        RECT 48.905 59.205 49.075 60.345 ;
        RECT 49.245 59.205 49.580 60.175 ;
        RECT 48.565 58.705 48.760 59.035 ;
        RECT 48.985 58.705 49.240 59.035 ;
        RECT 48.985 58.535 49.155 58.705 ;
        RECT 49.410 58.535 49.580 59.205 ;
        RECT 50.675 59.180 50.965 60.345 ;
        RECT 51.135 59.255 54.645 60.345 ;
        RECT 48.225 58.365 49.155 58.535 ;
        RECT 48.225 58.330 48.400 58.365 ;
        RECT 47.870 57.965 48.400 58.330 ;
        RECT 48.825 57.795 49.155 58.195 ;
        RECT 49.325 57.965 49.580 58.535 ;
        RECT 51.135 58.565 52.785 59.085 ;
        RECT 52.955 58.735 54.645 59.255 ;
        RECT 54.820 59.205 55.155 60.175 ;
        RECT 55.325 59.205 55.495 60.345 ;
        RECT 55.665 60.005 57.695 60.175 ;
        RECT 50.675 57.795 50.965 58.520 ;
        RECT 51.135 57.795 54.645 58.565 ;
        RECT 54.820 58.535 54.990 59.205 ;
        RECT 55.665 59.035 55.835 60.005 ;
        RECT 55.160 58.705 55.415 59.035 ;
        RECT 55.640 58.705 55.835 59.035 ;
        RECT 56.005 59.665 57.130 59.835 ;
        RECT 55.245 58.535 55.415 58.705 ;
        RECT 56.005 58.535 56.175 59.665 ;
        RECT 54.820 57.965 55.075 58.535 ;
        RECT 55.245 58.365 56.175 58.535 ;
        RECT 56.345 59.325 57.355 59.495 ;
        RECT 56.345 58.525 56.515 59.325 ;
        RECT 56.000 58.330 56.175 58.365 ;
        RECT 55.245 57.795 55.575 58.195 ;
        RECT 56.000 57.965 56.530 58.330 ;
        RECT 56.720 58.305 56.995 59.125 ;
        RECT 56.715 58.135 56.995 58.305 ;
        RECT 56.720 57.965 56.995 58.135 ;
        RECT 57.165 57.965 57.355 59.325 ;
        RECT 57.525 59.340 57.695 60.005 ;
        RECT 57.865 59.585 58.035 60.345 ;
        RECT 58.270 59.585 58.785 59.995 ;
        RECT 58.955 59.910 64.300 60.345 ;
        RECT 57.525 59.150 58.275 59.340 ;
        RECT 58.445 58.775 58.785 59.585 ;
        RECT 57.555 58.605 58.785 58.775 ;
        RECT 57.535 57.795 58.045 58.330 ;
        RECT 58.265 58.000 58.510 58.605 ;
        RECT 60.540 58.340 60.880 59.170 ;
        RECT 62.360 58.660 62.710 59.910 ;
        RECT 64.475 59.495 64.735 60.175 ;
        RECT 64.905 59.565 65.155 60.345 ;
        RECT 65.405 59.795 65.655 60.175 ;
        RECT 65.825 59.965 66.180 60.345 ;
        RECT 67.185 59.955 67.520 60.175 ;
        RECT 66.785 59.795 67.015 59.835 ;
        RECT 65.405 59.595 67.015 59.795 ;
        RECT 65.405 59.585 66.240 59.595 ;
        RECT 66.830 59.505 67.015 59.595 ;
        RECT 58.955 57.795 64.300 58.340 ;
        RECT 64.475 58.305 64.645 59.495 ;
        RECT 66.345 59.395 66.675 59.425 ;
        RECT 64.875 59.335 66.675 59.395 ;
        RECT 67.265 59.335 67.520 59.955 ;
        RECT 64.815 59.225 67.520 59.335 ;
        RECT 64.815 59.190 65.015 59.225 ;
        RECT 64.815 58.615 64.985 59.190 ;
        RECT 66.345 59.165 67.520 59.225 ;
        RECT 67.695 59.205 67.975 60.345 ;
        RECT 68.145 59.195 68.475 60.175 ;
        RECT 68.645 59.205 68.905 60.345 ;
        RECT 69.085 59.285 69.415 60.135 ;
        RECT 68.210 59.155 68.385 59.195 ;
        RECT 65.215 58.750 65.625 59.055 ;
        RECT 65.795 58.785 66.125 58.995 ;
        RECT 64.815 58.495 65.085 58.615 ;
        RECT 64.815 58.450 65.660 58.495 ;
        RECT 64.905 58.325 65.660 58.450 ;
        RECT 65.915 58.385 66.125 58.785 ;
        RECT 66.370 58.785 66.845 58.995 ;
        RECT 67.035 58.785 67.525 58.985 ;
        RECT 66.370 58.385 66.590 58.785 ;
        RECT 67.705 58.765 68.040 59.035 ;
        RECT 68.210 58.595 68.380 59.155 ;
        RECT 68.550 58.785 68.885 59.035 ;
        RECT 64.475 58.295 64.705 58.305 ;
        RECT 64.475 57.965 64.735 58.295 ;
        RECT 65.490 58.175 65.660 58.325 ;
        RECT 64.905 57.795 65.235 58.155 ;
        RECT 65.490 57.965 66.790 58.175 ;
        RECT 67.065 57.795 67.520 58.560 ;
        RECT 67.695 57.795 68.005 58.595 ;
        RECT 68.210 57.965 68.905 58.595 ;
        RECT 69.085 58.520 69.275 59.285 ;
        RECT 69.585 59.205 69.835 60.345 ;
        RECT 70.025 59.705 70.275 60.125 ;
        RECT 70.505 59.875 70.835 60.345 ;
        RECT 71.065 59.705 71.315 60.125 ;
        RECT 70.025 59.535 71.315 59.705 ;
        RECT 71.495 59.705 71.825 60.135 ;
        RECT 71.495 59.535 71.950 59.705 ;
        RECT 70.015 59.035 70.230 59.365 ;
        RECT 69.445 58.705 69.755 59.035 ;
        RECT 69.925 58.705 70.230 59.035 ;
        RECT 70.405 58.705 70.690 59.365 ;
        RECT 70.885 58.705 71.150 59.365 ;
        RECT 71.365 58.705 71.610 59.365 ;
        RECT 69.585 58.535 69.755 58.705 ;
        RECT 71.780 58.535 71.950 59.535 ;
        RECT 72.450 59.335 72.750 60.175 ;
        RECT 72.945 59.505 73.195 60.345 ;
        RECT 73.785 59.755 74.590 60.175 ;
        RECT 73.365 59.585 74.930 59.755 ;
        RECT 73.365 59.335 73.535 59.585 ;
        RECT 72.450 59.165 73.535 59.335 ;
        RECT 72.295 58.705 72.625 58.995 ;
        RECT 72.795 58.535 72.965 59.165 ;
        RECT 73.705 59.035 74.025 59.415 ;
        RECT 74.215 59.325 74.590 59.415 ;
        RECT 74.195 59.155 74.590 59.325 ;
        RECT 74.760 59.335 74.930 59.585 ;
        RECT 75.100 59.505 75.430 60.345 ;
        RECT 75.600 59.585 76.265 60.175 ;
        RECT 74.760 59.165 75.680 59.335 ;
        RECT 73.135 58.785 73.465 58.995 ;
        RECT 73.645 58.785 74.025 59.035 ;
        RECT 74.215 58.995 74.590 59.155 ;
        RECT 75.510 58.995 75.680 59.165 ;
        RECT 74.215 58.785 74.700 58.995 ;
        RECT 74.890 58.785 75.340 58.995 ;
        RECT 75.510 58.785 75.845 58.995 ;
        RECT 76.015 58.615 76.265 59.585 ;
        RECT 76.435 59.180 76.725 60.345 ;
        RECT 76.900 59.955 77.235 60.175 ;
        RECT 78.240 59.965 78.595 60.345 ;
        RECT 76.900 59.335 77.155 59.955 ;
        RECT 77.405 59.795 77.635 59.835 ;
        RECT 78.765 59.795 79.015 60.175 ;
        RECT 77.405 59.595 79.015 59.795 ;
        RECT 77.405 59.505 77.590 59.595 ;
        RECT 78.180 59.585 79.015 59.595 ;
        RECT 79.265 59.565 79.515 60.345 ;
        RECT 79.685 59.495 79.945 60.175 ;
        RECT 80.665 59.675 80.835 60.175 ;
        RECT 81.005 59.845 81.335 60.345 ;
        RECT 80.665 59.505 81.330 59.675 ;
        RECT 77.745 59.395 78.075 59.425 ;
        RECT 77.745 59.335 79.545 59.395 ;
        RECT 76.900 59.225 79.605 59.335 ;
        RECT 76.900 59.165 78.075 59.225 ;
        RECT 79.405 59.190 79.605 59.225 ;
        RECT 76.895 58.785 77.385 58.985 ;
        RECT 77.575 58.785 78.050 58.995 ;
        RECT 69.085 58.010 69.415 58.520 ;
        RECT 69.585 58.365 71.950 58.535 ;
        RECT 69.585 57.795 69.915 58.195 ;
        RECT 70.965 58.025 71.295 58.365 ;
        RECT 72.455 58.355 72.965 58.535 ;
        RECT 73.370 58.445 75.070 58.615 ;
        RECT 73.370 58.355 73.755 58.445 ;
        RECT 71.465 57.795 71.795 58.195 ;
        RECT 72.455 57.965 72.785 58.355 ;
        RECT 72.955 58.015 74.140 58.185 ;
        RECT 74.400 57.795 74.570 58.265 ;
        RECT 74.740 57.980 75.070 58.445 ;
        RECT 75.240 57.795 75.410 58.615 ;
        RECT 75.580 57.975 76.265 58.615 ;
        RECT 76.435 57.795 76.725 58.520 ;
        RECT 76.900 57.795 77.355 58.560 ;
        RECT 77.830 58.385 78.050 58.785 ;
        RECT 78.295 58.785 78.625 58.995 ;
        RECT 78.295 58.385 78.505 58.785 ;
        RECT 78.795 58.750 79.205 59.055 ;
        RECT 79.435 58.615 79.605 59.190 ;
        RECT 79.335 58.495 79.605 58.615 ;
        RECT 78.760 58.450 79.605 58.495 ;
        RECT 78.760 58.325 79.515 58.450 ;
        RECT 78.760 58.175 78.930 58.325 ;
        RECT 79.775 58.295 79.945 59.495 ;
        RECT 80.580 58.685 80.930 59.335 ;
        RECT 81.100 58.515 81.330 59.505 ;
        RECT 77.630 57.965 78.930 58.175 ;
        RECT 79.185 57.795 79.515 58.155 ;
        RECT 79.685 57.965 79.945 58.295 ;
        RECT 80.665 58.345 81.330 58.515 ;
        RECT 80.665 58.055 80.835 58.345 ;
        RECT 81.005 57.795 81.335 58.175 ;
        RECT 81.505 58.055 81.690 60.175 ;
        RECT 81.930 59.885 82.195 60.345 ;
        RECT 82.365 59.750 82.615 60.175 ;
        RECT 82.825 59.900 83.930 60.070 ;
        RECT 82.310 59.620 82.615 59.750 ;
        RECT 81.860 58.425 82.140 59.375 ;
        RECT 82.310 58.515 82.480 59.620 ;
        RECT 82.650 58.835 82.890 59.430 ;
        RECT 83.060 59.365 83.590 59.730 ;
        RECT 83.060 58.665 83.230 59.365 ;
        RECT 83.760 59.285 83.930 59.900 ;
        RECT 84.100 59.545 84.270 60.345 ;
        RECT 84.440 59.845 84.690 60.175 ;
        RECT 84.915 59.875 85.800 60.045 ;
        RECT 83.760 59.195 84.270 59.285 ;
        RECT 82.310 58.385 82.535 58.515 ;
        RECT 82.705 58.445 83.230 58.665 ;
        RECT 83.400 59.025 84.270 59.195 ;
        RECT 81.945 57.795 82.195 58.255 ;
        RECT 82.365 58.245 82.535 58.385 ;
        RECT 83.400 58.245 83.570 59.025 ;
        RECT 84.100 58.955 84.270 59.025 ;
        RECT 83.780 58.775 83.980 58.805 ;
        RECT 84.440 58.775 84.610 59.845 ;
        RECT 84.780 58.955 84.970 59.675 ;
        RECT 83.780 58.475 84.610 58.775 ;
        RECT 85.140 58.745 85.460 59.705 ;
        RECT 82.365 58.075 82.700 58.245 ;
        RECT 82.895 58.075 83.570 58.245 ;
        RECT 83.890 57.795 84.260 58.295 ;
        RECT 84.440 58.245 84.610 58.475 ;
        RECT 84.995 58.415 85.460 58.745 ;
        RECT 85.630 59.035 85.800 59.875 ;
        RECT 85.980 59.845 86.295 60.345 ;
        RECT 86.525 59.615 86.865 60.175 ;
        RECT 85.970 59.240 86.865 59.615 ;
        RECT 87.035 59.335 87.205 60.345 ;
        RECT 86.675 59.035 86.865 59.240 ;
        RECT 87.375 59.285 87.705 60.130 ;
        RECT 87.375 59.205 87.765 59.285 ;
        RECT 87.550 59.155 87.765 59.205 ;
        RECT 85.630 58.705 86.505 59.035 ;
        RECT 86.675 58.705 87.425 59.035 ;
        RECT 85.630 58.245 85.800 58.705 ;
        RECT 86.675 58.535 86.875 58.705 ;
        RECT 87.595 58.575 87.765 59.155 ;
        RECT 87.540 58.535 87.765 58.575 ;
        RECT 84.440 58.075 84.845 58.245 ;
        RECT 85.015 58.075 85.800 58.245 ;
        RECT 86.075 57.795 86.285 58.325 ;
        RECT 86.545 58.010 86.875 58.535 ;
        RECT 87.385 58.450 87.765 58.535 ;
        RECT 87.935 59.270 88.205 60.175 ;
        RECT 88.375 59.585 88.705 60.345 ;
        RECT 88.885 59.415 89.055 60.175 ;
        RECT 87.935 58.470 88.105 59.270 ;
        RECT 88.390 59.245 89.055 59.415 ;
        RECT 89.315 59.255 90.525 60.345 ;
        RECT 88.390 59.100 88.560 59.245 ;
        RECT 88.275 58.770 88.560 59.100 ;
        RECT 88.390 58.515 88.560 58.770 ;
        RECT 88.795 58.695 89.125 59.065 ;
        RECT 89.315 58.715 89.835 59.255 ;
        RECT 90.005 58.545 90.525 59.085 ;
        RECT 87.045 57.795 87.215 58.405 ;
        RECT 87.385 58.015 87.715 58.450 ;
        RECT 87.935 57.965 88.195 58.470 ;
        RECT 88.390 58.345 89.055 58.515 ;
        RECT 88.375 57.795 88.705 58.175 ;
        RECT 88.885 57.965 89.055 58.345 ;
        RECT 89.315 57.795 90.525 58.545 ;
        RECT 11.950 57.625 90.610 57.795 ;
        RECT 12.035 56.875 13.245 57.625 ;
        RECT 13.415 56.875 14.625 57.625 ;
        RECT 12.035 56.335 12.555 56.875 ;
        RECT 12.725 56.165 13.245 56.705 ;
        RECT 13.415 56.335 13.935 56.875 ;
        RECT 14.795 56.825 15.135 57.455 ;
        RECT 15.305 56.825 15.555 57.625 ;
        RECT 15.745 56.975 16.075 57.455 ;
        RECT 16.245 57.165 16.470 57.625 ;
        RECT 16.640 56.975 16.970 57.455 ;
        RECT 14.105 56.165 14.625 56.705 ;
        RECT 12.035 55.075 13.245 56.165 ;
        RECT 13.415 55.075 14.625 56.165 ;
        RECT 14.795 56.215 14.970 56.825 ;
        RECT 15.745 56.805 16.970 56.975 ;
        RECT 17.600 56.845 18.100 57.455 ;
        RECT 15.140 56.465 15.835 56.635 ;
        RECT 15.665 56.215 15.835 56.465 ;
        RECT 16.010 56.435 16.430 56.635 ;
        RECT 16.600 56.435 16.930 56.635 ;
        RECT 17.100 56.435 17.430 56.635 ;
        RECT 17.600 56.215 17.770 56.845 ;
        RECT 18.475 56.825 18.815 57.455 ;
        RECT 18.985 56.825 19.235 57.625 ;
        RECT 19.425 56.975 19.755 57.455 ;
        RECT 19.925 57.165 20.150 57.625 ;
        RECT 20.320 56.975 20.650 57.455 ;
        RECT 17.955 56.385 18.305 56.635 ;
        RECT 18.475 56.215 18.650 56.825 ;
        RECT 19.425 56.805 20.650 56.975 ;
        RECT 21.280 56.845 21.780 57.455 ;
        RECT 22.205 57.085 22.430 57.445 ;
        RECT 22.610 57.255 22.940 57.625 ;
        RECT 23.120 57.085 23.375 57.445 ;
        RECT 23.940 57.255 24.685 57.625 ;
        RECT 22.205 56.895 24.690 57.085 ;
        RECT 18.820 56.465 19.515 56.635 ;
        RECT 19.345 56.215 19.515 56.465 ;
        RECT 19.690 56.435 20.110 56.635 ;
        RECT 20.280 56.435 20.610 56.635 ;
        RECT 20.780 56.435 21.110 56.635 ;
        RECT 21.280 56.215 21.450 56.845 ;
        RECT 21.635 56.385 21.985 56.635 ;
        RECT 22.165 56.385 22.435 56.715 ;
        RECT 22.615 56.385 23.050 56.715 ;
        RECT 23.230 56.385 23.805 56.715 ;
        RECT 23.985 56.385 24.265 56.715 ;
        RECT 14.795 55.245 15.135 56.215 ;
        RECT 15.305 55.075 15.475 56.215 ;
        RECT 15.665 56.045 18.100 56.215 ;
        RECT 15.745 55.075 15.995 55.875 ;
        RECT 16.640 55.245 16.970 56.045 ;
        RECT 17.270 55.075 17.600 55.875 ;
        RECT 17.770 55.245 18.100 56.045 ;
        RECT 18.475 55.245 18.815 56.215 ;
        RECT 18.985 55.075 19.155 56.215 ;
        RECT 19.345 56.045 21.780 56.215 ;
        RECT 24.465 56.205 24.690 56.895 ;
        RECT 19.425 55.075 19.675 55.875 ;
        RECT 20.320 55.245 20.650 56.045 ;
        RECT 20.950 55.075 21.280 55.875 ;
        RECT 21.450 55.245 21.780 56.045 ;
        RECT 22.195 56.025 24.690 56.205 ;
        RECT 24.865 56.025 25.200 57.445 ;
        RECT 25.580 56.845 26.080 57.455 ;
        RECT 25.375 56.385 25.725 56.635 ;
        RECT 25.910 56.215 26.080 56.845 ;
        RECT 26.710 56.975 27.040 57.455 ;
        RECT 27.210 57.165 27.435 57.625 ;
        RECT 27.605 56.975 27.935 57.455 ;
        RECT 26.710 56.805 27.935 56.975 ;
        RECT 28.125 56.825 28.375 57.625 ;
        RECT 28.545 56.825 28.885 57.455 ;
        RECT 29.145 57.075 29.315 57.365 ;
        RECT 29.485 57.245 29.815 57.625 ;
        RECT 29.145 56.905 29.810 57.075 ;
        RECT 28.655 56.775 28.885 56.825 ;
        RECT 26.250 56.435 26.580 56.635 ;
        RECT 26.750 56.435 27.080 56.635 ;
        RECT 27.250 56.435 27.670 56.635 ;
        RECT 27.845 56.465 28.540 56.635 ;
        RECT 27.845 56.215 28.015 56.465 ;
        RECT 28.710 56.215 28.885 56.775 ;
        RECT 22.195 55.255 22.485 56.025 ;
        RECT 23.055 55.615 24.245 55.845 ;
        RECT 23.055 55.255 23.315 55.615 ;
        RECT 23.485 55.075 23.815 55.445 ;
        RECT 23.985 55.255 24.245 55.615 ;
        RECT 24.435 55.075 24.765 55.795 ;
        RECT 24.935 55.255 25.200 56.025 ;
        RECT 25.580 56.045 28.015 56.215 ;
        RECT 25.580 55.245 25.910 56.045 ;
        RECT 26.080 55.075 26.410 55.875 ;
        RECT 26.710 55.245 27.040 56.045 ;
        RECT 27.685 55.075 27.935 55.875 ;
        RECT 28.205 55.075 28.375 56.215 ;
        RECT 28.545 55.245 28.885 56.215 ;
        RECT 29.060 56.085 29.410 56.735 ;
        RECT 29.580 55.915 29.810 56.905 ;
        RECT 29.145 55.745 29.810 55.915 ;
        RECT 29.145 55.245 29.315 55.745 ;
        RECT 29.485 55.075 29.815 55.575 ;
        RECT 29.985 55.245 30.170 57.365 ;
        RECT 30.425 57.165 30.675 57.625 ;
        RECT 30.845 57.175 31.180 57.345 ;
        RECT 31.375 57.175 32.050 57.345 ;
        RECT 30.845 57.035 31.015 57.175 ;
        RECT 30.340 56.045 30.620 56.995 ;
        RECT 30.790 56.905 31.015 57.035 ;
        RECT 30.790 55.800 30.960 56.905 ;
        RECT 31.185 56.755 31.710 56.975 ;
        RECT 31.130 55.990 31.370 56.585 ;
        RECT 31.540 56.055 31.710 56.755 ;
        RECT 31.880 56.395 32.050 57.175 ;
        RECT 32.370 57.125 32.740 57.625 ;
        RECT 32.920 57.175 33.325 57.345 ;
        RECT 33.495 57.175 34.280 57.345 ;
        RECT 32.920 56.945 33.090 57.175 ;
        RECT 32.260 56.645 33.090 56.945 ;
        RECT 33.475 56.675 33.940 57.005 ;
        RECT 32.260 56.615 32.460 56.645 ;
        RECT 32.580 56.395 32.750 56.465 ;
        RECT 31.880 56.225 32.750 56.395 ;
        RECT 32.240 56.135 32.750 56.225 ;
        RECT 30.790 55.670 31.095 55.800 ;
        RECT 31.540 55.690 32.070 56.055 ;
        RECT 30.410 55.075 30.675 55.535 ;
        RECT 30.845 55.245 31.095 55.670 ;
        RECT 32.240 55.520 32.410 56.135 ;
        RECT 31.305 55.350 32.410 55.520 ;
        RECT 32.580 55.075 32.750 55.875 ;
        RECT 32.920 55.575 33.090 56.645 ;
        RECT 33.260 55.745 33.450 56.465 ;
        RECT 33.620 55.715 33.940 56.675 ;
        RECT 34.110 56.715 34.280 57.175 ;
        RECT 34.555 57.095 34.765 57.625 ;
        RECT 35.025 56.885 35.355 57.410 ;
        RECT 35.525 57.015 35.695 57.625 ;
        RECT 35.865 56.970 36.195 57.405 ;
        RECT 35.865 56.885 36.245 56.970 ;
        RECT 35.155 56.715 35.355 56.885 ;
        RECT 36.020 56.845 36.245 56.885 ;
        RECT 34.110 56.385 34.985 56.715 ;
        RECT 35.155 56.385 35.905 56.715 ;
        RECT 32.920 55.245 33.170 55.575 ;
        RECT 34.110 55.545 34.280 56.385 ;
        RECT 35.155 56.180 35.345 56.385 ;
        RECT 36.075 56.265 36.245 56.845 ;
        RECT 36.415 56.875 37.625 57.625 ;
        RECT 37.795 56.900 38.085 57.625 ;
        RECT 38.260 56.885 38.515 57.455 ;
        RECT 38.685 57.225 39.015 57.625 ;
        RECT 39.440 57.090 39.970 57.455 ;
        RECT 39.440 57.055 39.615 57.090 ;
        RECT 38.685 56.885 39.615 57.055 ;
        RECT 36.415 56.335 36.935 56.875 ;
        RECT 36.030 56.215 36.245 56.265 ;
        RECT 34.450 55.805 35.345 56.180 ;
        RECT 35.855 56.135 36.245 56.215 ;
        RECT 37.105 56.165 37.625 56.705 ;
        RECT 33.395 55.375 34.280 55.545 ;
        RECT 34.460 55.075 34.775 55.575 ;
        RECT 35.005 55.245 35.345 55.805 ;
        RECT 35.515 55.075 35.685 56.085 ;
        RECT 35.855 55.290 36.185 56.135 ;
        RECT 36.415 55.075 37.625 56.165 ;
        RECT 37.795 55.075 38.085 56.240 ;
        RECT 38.260 56.215 38.430 56.885 ;
        RECT 38.685 56.715 38.855 56.885 ;
        RECT 38.600 56.385 38.855 56.715 ;
        RECT 39.080 56.385 39.275 56.715 ;
        RECT 38.260 55.245 38.595 56.215 ;
        RECT 38.765 55.075 38.935 56.215 ;
        RECT 39.105 55.415 39.275 56.385 ;
        RECT 39.445 55.755 39.615 56.885 ;
        RECT 39.785 56.095 39.955 56.895 ;
        RECT 40.160 56.605 40.435 57.455 ;
        RECT 40.155 56.435 40.435 56.605 ;
        RECT 40.160 56.295 40.435 56.435 ;
        RECT 40.605 56.095 40.795 57.455 ;
        RECT 40.975 57.090 41.485 57.625 ;
        RECT 41.705 56.815 41.950 57.420 ;
        RECT 42.395 56.885 42.780 57.455 ;
        RECT 42.950 57.165 43.275 57.625 ;
        RECT 43.795 56.995 44.075 57.455 ;
        RECT 40.995 56.645 42.225 56.815 ;
        RECT 39.785 55.925 40.795 56.095 ;
        RECT 40.965 56.080 41.715 56.270 ;
        RECT 39.445 55.585 40.570 55.755 ;
        RECT 40.965 55.415 41.135 56.080 ;
        RECT 41.885 55.835 42.225 56.645 ;
        RECT 39.105 55.245 41.135 55.415 ;
        RECT 41.305 55.075 41.475 55.835 ;
        RECT 41.710 55.425 42.225 55.835 ;
        RECT 42.395 56.215 42.675 56.885 ;
        RECT 42.950 56.825 44.075 56.995 ;
        RECT 42.950 56.715 43.400 56.825 ;
        RECT 42.845 56.385 43.400 56.715 ;
        RECT 44.265 56.655 44.665 57.455 ;
        RECT 45.065 57.165 45.335 57.625 ;
        RECT 45.505 56.995 45.790 57.455 ;
        RECT 42.395 55.245 42.780 56.215 ;
        RECT 42.950 55.925 43.400 56.385 ;
        RECT 43.570 56.095 44.665 56.655 ;
        RECT 42.950 55.705 44.075 55.925 ;
        RECT 42.950 55.075 43.275 55.535 ;
        RECT 43.795 55.245 44.075 55.705 ;
        RECT 44.265 55.245 44.665 56.095 ;
        RECT 44.835 56.825 45.790 56.995 ;
        RECT 44.835 55.925 45.045 56.825 ;
        RECT 45.215 56.095 45.905 56.655 ;
        RECT 46.080 56.025 46.415 57.445 ;
        RECT 46.595 57.255 47.340 57.625 ;
        RECT 47.905 57.085 48.160 57.445 ;
        RECT 48.340 57.255 48.670 57.625 ;
        RECT 48.850 57.085 49.075 57.445 ;
        RECT 46.590 56.895 49.075 57.085 ;
        RECT 46.590 56.205 46.815 56.895 ;
        RECT 49.295 56.855 50.965 57.625 ;
        RECT 51.140 56.885 51.395 57.455 ;
        RECT 51.565 57.225 51.895 57.625 ;
        RECT 52.320 57.090 52.850 57.455 ;
        RECT 52.320 57.055 52.495 57.090 ;
        RECT 51.565 56.885 52.495 57.055 ;
        RECT 47.015 56.385 47.295 56.715 ;
        RECT 47.475 56.385 48.050 56.715 ;
        RECT 48.230 56.385 48.665 56.715 ;
        RECT 48.845 56.385 49.115 56.715 ;
        RECT 49.295 56.335 50.045 56.855 ;
        RECT 46.590 56.025 49.085 56.205 ;
        RECT 50.215 56.165 50.965 56.685 ;
        RECT 44.835 55.705 45.790 55.925 ;
        RECT 45.065 55.075 45.335 55.535 ;
        RECT 45.505 55.245 45.790 55.705 ;
        RECT 46.080 55.255 46.345 56.025 ;
        RECT 46.515 55.075 46.845 55.795 ;
        RECT 47.035 55.615 48.225 55.845 ;
        RECT 47.035 55.255 47.295 55.615 ;
        RECT 47.465 55.075 47.795 55.445 ;
        RECT 47.965 55.255 48.225 55.615 ;
        RECT 48.795 55.255 49.085 56.025 ;
        RECT 49.295 55.075 50.965 56.165 ;
        RECT 51.140 56.215 51.310 56.885 ;
        RECT 51.565 56.715 51.735 56.885 ;
        RECT 51.480 56.385 51.735 56.715 ;
        RECT 51.960 56.385 52.155 56.715 ;
        RECT 51.140 55.245 51.475 56.215 ;
        RECT 51.645 55.075 51.815 56.215 ;
        RECT 51.985 55.415 52.155 56.385 ;
        RECT 52.325 55.755 52.495 56.885 ;
        RECT 52.665 56.095 52.835 56.895 ;
        RECT 53.040 56.605 53.315 57.455 ;
        RECT 53.035 56.435 53.315 56.605 ;
        RECT 53.040 56.295 53.315 56.435 ;
        RECT 53.485 56.095 53.675 57.455 ;
        RECT 53.855 57.090 54.365 57.625 ;
        RECT 54.585 56.815 54.830 57.420 ;
        RECT 55.275 56.885 55.660 57.455 ;
        RECT 55.830 57.165 56.155 57.625 ;
        RECT 56.675 56.995 56.955 57.455 ;
        RECT 53.875 56.645 55.105 56.815 ;
        RECT 52.665 55.925 53.675 56.095 ;
        RECT 53.845 56.080 54.595 56.270 ;
        RECT 52.325 55.585 53.450 55.755 ;
        RECT 53.845 55.415 54.015 56.080 ;
        RECT 54.765 55.835 55.105 56.645 ;
        RECT 51.985 55.245 54.015 55.415 ;
        RECT 54.185 55.075 54.355 55.835 ;
        RECT 54.590 55.425 55.105 55.835 ;
        RECT 55.275 56.215 55.555 56.885 ;
        RECT 55.830 56.825 56.955 56.995 ;
        RECT 55.830 56.715 56.280 56.825 ;
        RECT 55.725 56.385 56.280 56.715 ;
        RECT 57.145 56.655 57.545 57.455 ;
        RECT 57.945 57.165 58.215 57.625 ;
        RECT 58.385 56.995 58.670 57.455 ;
        RECT 55.275 55.245 55.660 56.215 ;
        RECT 55.830 55.925 56.280 56.385 ;
        RECT 56.450 56.095 57.545 56.655 ;
        RECT 55.830 55.705 56.955 55.925 ;
        RECT 55.830 55.075 56.155 55.535 ;
        RECT 56.675 55.245 56.955 55.705 ;
        RECT 57.145 55.245 57.545 56.095 ;
        RECT 57.715 56.825 58.670 56.995 ;
        RECT 59.415 56.885 59.800 57.455 ;
        RECT 59.970 57.165 60.295 57.625 ;
        RECT 60.815 56.995 61.095 57.455 ;
        RECT 57.715 55.925 57.925 56.825 ;
        RECT 58.095 56.095 58.785 56.655 ;
        RECT 59.415 56.215 59.695 56.885 ;
        RECT 59.970 56.825 61.095 56.995 ;
        RECT 59.970 56.715 60.420 56.825 ;
        RECT 59.865 56.385 60.420 56.715 ;
        RECT 61.285 56.655 61.685 57.455 ;
        RECT 62.085 57.165 62.355 57.625 ;
        RECT 62.525 56.995 62.810 57.455 ;
        RECT 57.715 55.705 58.670 55.925 ;
        RECT 57.945 55.075 58.215 55.535 ;
        RECT 58.385 55.245 58.670 55.705 ;
        RECT 59.415 55.245 59.800 56.215 ;
        RECT 59.970 55.925 60.420 56.385 ;
        RECT 60.590 56.095 61.685 56.655 ;
        RECT 59.970 55.705 61.095 55.925 ;
        RECT 59.970 55.075 60.295 55.535 ;
        RECT 60.815 55.245 61.095 55.705 ;
        RECT 61.285 55.245 61.685 56.095 ;
        RECT 61.855 56.825 62.810 56.995 ;
        RECT 63.555 56.900 63.845 57.625 ;
        RECT 64.130 56.995 64.415 57.455 ;
        RECT 64.585 57.165 64.855 57.625 ;
        RECT 64.130 56.825 65.085 56.995 ;
        RECT 61.855 55.925 62.065 56.825 ;
        RECT 62.235 56.095 62.925 56.655 ;
        RECT 61.855 55.705 62.810 55.925 ;
        RECT 62.085 55.075 62.355 55.535 ;
        RECT 62.525 55.245 62.810 55.705 ;
        RECT 63.555 55.075 63.845 56.240 ;
        RECT 64.015 56.095 64.705 56.655 ;
        RECT 64.875 55.925 65.085 56.825 ;
        RECT 64.130 55.705 65.085 55.925 ;
        RECT 65.255 56.655 65.655 57.455 ;
        RECT 65.845 56.995 66.125 57.455 ;
        RECT 66.645 57.165 66.970 57.625 ;
        RECT 65.845 56.825 66.970 56.995 ;
        RECT 67.140 56.885 67.525 57.455 ;
        RECT 67.705 57.115 68.935 57.455 ;
        RECT 69.105 57.135 69.360 57.625 ;
        RECT 67.705 56.885 68.035 57.115 ;
        RECT 66.520 56.715 66.970 56.825 ;
        RECT 65.255 56.095 66.350 56.655 ;
        RECT 66.520 56.385 67.075 56.715 ;
        RECT 64.130 55.245 64.415 55.705 ;
        RECT 64.585 55.075 64.855 55.535 ;
        RECT 65.255 55.245 65.655 56.095 ;
        RECT 66.520 55.925 66.970 56.385 ;
        RECT 67.245 56.215 67.525 56.885 ;
        RECT 67.695 56.385 68.005 56.715 ;
        RECT 68.210 56.385 68.585 56.945 ;
        RECT 68.755 56.215 68.935 57.115 ;
        RECT 69.120 56.385 69.340 56.965 ;
        RECT 69.625 56.945 69.795 57.320 ;
        RECT 69.595 56.775 69.795 56.945 ;
        RECT 69.985 57.095 70.215 57.400 ;
        RECT 70.385 57.265 70.715 57.625 ;
        RECT 70.910 57.095 71.200 57.445 ;
        RECT 72.335 57.115 72.735 57.625 ;
        RECT 69.985 56.925 71.200 57.095 ;
        RECT 73.310 57.010 73.480 57.455 ;
        RECT 73.650 57.225 74.370 57.625 ;
        RECT 74.540 57.055 74.710 57.455 ;
        RECT 74.945 57.180 75.375 57.625 ;
        RECT 69.625 56.755 69.795 56.775 ;
        RECT 69.625 56.585 70.145 56.755 ;
        RECT 65.845 55.705 66.970 55.925 ;
        RECT 65.845 55.245 66.125 55.705 ;
        RECT 66.645 55.075 66.970 55.535 ;
        RECT 67.140 55.245 67.525 56.215 ;
        RECT 67.705 56.045 68.935 56.215 ;
        RECT 67.705 55.245 68.035 56.045 ;
        RECT 68.205 55.075 68.435 55.875 ;
        RECT 68.605 55.245 68.935 56.045 ;
        RECT 69.105 55.075 69.360 56.215 ;
        RECT 69.540 56.055 69.785 56.415 ;
        RECT 69.975 56.205 70.145 56.585 ;
        RECT 70.315 56.385 70.700 56.715 ;
        RECT 70.880 56.605 71.140 56.715 ;
        RECT 70.880 56.435 71.145 56.605 ;
        RECT 70.880 56.385 71.140 56.435 ;
        RECT 69.975 55.925 70.325 56.205 ;
        RECT 69.540 55.075 69.795 55.875 ;
        RECT 69.995 55.245 70.325 55.925 ;
        RECT 70.505 55.335 70.700 56.385 ;
        RECT 70.880 55.075 71.200 56.215 ;
        RECT 72.350 56.055 72.610 56.945 ;
        RECT 72.810 56.355 73.070 56.945 ;
        RECT 73.310 56.840 73.660 57.010 ;
        RECT 72.810 56.055 73.290 56.355 ;
        RECT 72.375 55.705 73.315 55.875 ;
        RECT 72.375 55.245 72.555 55.705 ;
        RECT 72.725 55.075 72.975 55.535 ;
        RECT 73.145 55.455 73.315 55.705 ;
        RECT 73.490 55.815 73.660 56.840 ;
        RECT 73.830 56.885 74.710 57.055 ;
        RECT 75.545 56.900 75.805 57.455 ;
        RECT 73.830 56.165 74.000 56.885 ;
        RECT 74.190 56.335 74.480 56.715 ;
        RECT 73.830 55.995 74.350 56.165 ;
        RECT 74.650 56.095 74.980 56.715 ;
        RECT 75.205 56.385 75.460 56.715 ;
        RECT 73.490 55.645 73.900 55.815 ;
        RECT 74.180 55.805 74.350 55.995 ;
        RECT 75.205 55.905 75.375 56.385 ;
        RECT 75.630 56.185 75.805 56.900 ;
        RECT 75.995 56.895 76.325 57.625 ;
        RECT 76.495 56.715 76.705 57.335 ;
        RECT 76.885 56.915 77.315 57.445 ;
        RECT 76.010 56.365 76.300 56.715 ;
        RECT 76.495 56.365 76.890 56.715 ;
        RECT 77.070 56.665 77.315 56.915 ;
        RECT 77.495 56.845 77.725 57.625 ;
        RECT 77.905 56.995 78.285 57.445 ;
        RECT 79.285 57.075 79.455 57.365 ;
        RECT 79.625 57.245 79.955 57.625 ;
        RECT 77.070 56.365 77.605 56.665 ;
        RECT 77.905 56.545 78.135 56.995 ;
        RECT 79.285 56.905 79.950 57.075 ;
        RECT 73.645 55.510 73.900 55.645 ;
        RECT 74.615 55.735 75.375 55.905 ;
        RECT 74.615 55.510 74.785 55.735 ;
        RECT 73.145 55.285 73.475 55.455 ;
        RECT 73.645 55.340 74.785 55.510 ;
        RECT 73.645 55.245 73.900 55.340 ;
        RECT 75.045 55.075 75.375 55.475 ;
        RECT 75.545 55.245 75.805 56.185 ;
        RECT 76.065 55.985 77.105 56.185 ;
        RECT 76.065 55.255 76.235 55.985 ;
        RECT 76.415 55.075 76.745 55.805 ;
        RECT 76.915 55.255 77.105 55.985 ;
        RECT 77.275 55.255 77.605 56.365 ;
        RECT 77.795 55.865 78.135 56.545 ;
        RECT 78.315 56.045 78.545 56.735 ;
        RECT 79.200 56.085 79.550 56.735 ;
        RECT 79.720 55.915 79.950 56.905 ;
        RECT 77.795 55.665 78.555 55.865 ;
        RECT 77.795 55.075 78.125 55.485 ;
        RECT 78.295 55.275 78.555 55.665 ;
        RECT 79.285 55.745 79.950 55.915 ;
        RECT 79.285 55.245 79.455 55.745 ;
        RECT 79.625 55.075 79.955 55.575 ;
        RECT 80.125 55.245 80.310 57.365 ;
        RECT 80.565 57.165 80.815 57.625 ;
        RECT 80.985 57.175 81.320 57.345 ;
        RECT 81.515 57.175 82.190 57.345 ;
        RECT 80.985 57.035 81.155 57.175 ;
        RECT 80.480 56.045 80.760 56.995 ;
        RECT 80.930 56.905 81.155 57.035 ;
        RECT 80.930 55.800 81.100 56.905 ;
        RECT 81.325 56.755 81.850 56.975 ;
        RECT 81.270 55.990 81.510 56.585 ;
        RECT 81.680 56.055 81.850 56.755 ;
        RECT 82.020 56.395 82.190 57.175 ;
        RECT 82.510 57.125 82.880 57.625 ;
        RECT 83.060 57.175 83.465 57.345 ;
        RECT 83.635 57.175 84.420 57.345 ;
        RECT 83.060 56.945 83.230 57.175 ;
        RECT 82.400 56.645 83.230 56.945 ;
        RECT 83.615 56.675 84.080 57.005 ;
        RECT 82.400 56.615 82.600 56.645 ;
        RECT 82.720 56.395 82.890 56.465 ;
        RECT 82.020 56.225 82.890 56.395 ;
        RECT 82.380 56.135 82.890 56.225 ;
        RECT 80.930 55.670 81.235 55.800 ;
        RECT 81.680 55.690 82.210 56.055 ;
        RECT 80.550 55.075 80.815 55.535 ;
        RECT 80.985 55.245 81.235 55.670 ;
        RECT 82.380 55.520 82.550 56.135 ;
        RECT 81.445 55.350 82.550 55.520 ;
        RECT 82.720 55.075 82.890 55.875 ;
        RECT 83.060 55.575 83.230 56.645 ;
        RECT 83.400 55.745 83.590 56.465 ;
        RECT 83.760 55.715 84.080 56.675 ;
        RECT 84.250 56.715 84.420 57.175 ;
        RECT 84.695 57.095 84.905 57.625 ;
        RECT 85.165 56.885 85.495 57.410 ;
        RECT 85.665 57.015 85.835 57.625 ;
        RECT 86.005 56.970 86.335 57.405 ;
        RECT 87.565 57.075 87.735 57.455 ;
        RECT 87.950 57.245 88.280 57.625 ;
        RECT 86.005 56.885 86.385 56.970 ;
        RECT 87.565 56.905 88.280 57.075 ;
        RECT 85.295 56.715 85.495 56.885 ;
        RECT 86.160 56.845 86.385 56.885 ;
        RECT 84.250 56.385 85.125 56.715 ;
        RECT 85.295 56.385 86.045 56.715 ;
        RECT 83.060 55.245 83.310 55.575 ;
        RECT 84.250 55.545 84.420 56.385 ;
        RECT 85.295 56.180 85.485 56.385 ;
        RECT 86.215 56.265 86.385 56.845 ;
        RECT 87.475 56.355 87.830 56.725 ;
        RECT 88.110 56.715 88.280 56.905 ;
        RECT 88.450 56.880 88.705 57.455 ;
        RECT 88.110 56.385 88.365 56.715 ;
        RECT 86.170 56.215 86.385 56.265 ;
        RECT 84.590 55.805 85.485 56.180 ;
        RECT 85.995 56.135 86.385 56.215 ;
        RECT 88.110 56.175 88.280 56.385 ;
        RECT 83.535 55.375 84.420 55.545 ;
        RECT 84.600 55.075 84.915 55.575 ;
        RECT 85.145 55.245 85.485 55.805 ;
        RECT 85.655 55.075 85.825 56.085 ;
        RECT 85.995 55.290 86.325 56.135 ;
        RECT 87.565 56.005 88.280 56.175 ;
        RECT 88.535 56.150 88.705 56.880 ;
        RECT 88.880 56.785 89.140 57.625 ;
        RECT 89.315 56.875 90.525 57.625 ;
        RECT 87.565 55.245 87.735 56.005 ;
        RECT 87.950 55.075 88.280 55.835 ;
        RECT 88.450 55.245 88.705 56.150 ;
        RECT 88.880 55.075 89.140 56.225 ;
        RECT 89.315 56.165 89.835 56.705 ;
        RECT 90.005 56.335 90.525 56.875 ;
        RECT 89.315 55.075 90.525 56.165 ;
        RECT 11.950 54.905 90.610 55.075 ;
        RECT 12.035 53.815 13.245 54.905 ;
        RECT 12.035 53.105 12.555 53.645 ;
        RECT 12.725 53.275 13.245 53.815 ;
        RECT 13.600 53.935 13.990 54.110 ;
        RECT 14.475 54.105 14.805 54.905 ;
        RECT 14.975 54.115 15.510 54.735 ;
        RECT 13.600 53.765 15.025 53.935 ;
        RECT 12.035 52.355 13.245 53.105 ;
        RECT 13.475 53.035 13.830 53.595 ;
        RECT 14.000 52.865 14.170 53.765 ;
        RECT 14.340 53.035 14.605 53.595 ;
        RECT 14.855 53.265 15.025 53.765 ;
        RECT 15.195 53.095 15.510 54.115 ;
        RECT 15.805 54.235 15.975 54.735 ;
        RECT 16.145 54.405 16.475 54.905 ;
        RECT 15.805 54.065 16.470 54.235 ;
        RECT 15.720 53.245 16.070 53.895 ;
        RECT 13.580 52.355 13.820 52.865 ;
        RECT 14.000 52.535 14.280 52.865 ;
        RECT 14.510 52.355 14.725 52.865 ;
        RECT 14.895 52.525 15.510 53.095 ;
        RECT 16.240 53.075 16.470 54.065 ;
        RECT 15.805 52.905 16.470 53.075 ;
        RECT 15.805 52.615 15.975 52.905 ;
        RECT 16.145 52.355 16.475 52.735 ;
        RECT 16.645 52.615 16.830 54.735 ;
        RECT 17.070 54.445 17.335 54.905 ;
        RECT 17.505 54.310 17.755 54.735 ;
        RECT 17.965 54.460 19.070 54.630 ;
        RECT 17.450 54.180 17.755 54.310 ;
        RECT 17.000 52.985 17.280 53.935 ;
        RECT 17.450 53.075 17.620 54.180 ;
        RECT 17.790 53.395 18.030 53.990 ;
        RECT 18.200 53.925 18.730 54.290 ;
        RECT 18.200 53.225 18.370 53.925 ;
        RECT 18.900 53.845 19.070 54.460 ;
        RECT 19.240 54.105 19.410 54.905 ;
        RECT 19.580 54.405 19.830 54.735 ;
        RECT 20.055 54.435 20.940 54.605 ;
        RECT 18.900 53.755 19.410 53.845 ;
        RECT 17.450 52.945 17.675 53.075 ;
        RECT 17.845 53.005 18.370 53.225 ;
        RECT 18.540 53.585 19.410 53.755 ;
        RECT 17.085 52.355 17.335 52.815 ;
        RECT 17.505 52.805 17.675 52.945 ;
        RECT 18.540 52.805 18.710 53.585 ;
        RECT 19.240 53.515 19.410 53.585 ;
        RECT 18.920 53.335 19.120 53.365 ;
        RECT 19.580 53.335 19.750 54.405 ;
        RECT 19.920 53.515 20.110 54.235 ;
        RECT 18.920 53.035 19.750 53.335 ;
        RECT 20.280 53.305 20.600 54.265 ;
        RECT 17.505 52.635 17.840 52.805 ;
        RECT 18.035 52.635 18.710 52.805 ;
        RECT 19.030 52.355 19.400 52.855 ;
        RECT 19.580 52.805 19.750 53.035 ;
        RECT 20.135 52.975 20.600 53.305 ;
        RECT 20.770 53.595 20.940 54.435 ;
        RECT 21.120 54.405 21.435 54.905 ;
        RECT 21.665 54.175 22.005 54.735 ;
        RECT 21.110 53.800 22.005 54.175 ;
        RECT 22.175 53.895 22.345 54.905 ;
        RECT 21.815 53.595 22.005 53.800 ;
        RECT 22.515 53.845 22.845 54.690 ;
        RECT 22.515 53.765 22.905 53.845 ;
        RECT 23.075 53.815 24.745 54.905 ;
        RECT 22.690 53.715 22.905 53.765 ;
        RECT 20.770 53.265 21.645 53.595 ;
        RECT 21.815 53.265 22.565 53.595 ;
        RECT 20.770 52.805 20.940 53.265 ;
        RECT 21.815 53.095 22.015 53.265 ;
        RECT 22.735 53.135 22.905 53.715 ;
        RECT 22.680 53.095 22.905 53.135 ;
        RECT 19.580 52.635 19.985 52.805 ;
        RECT 20.155 52.635 20.940 52.805 ;
        RECT 21.215 52.355 21.425 52.885 ;
        RECT 21.685 52.570 22.015 53.095 ;
        RECT 22.525 53.010 22.905 53.095 ;
        RECT 23.075 53.125 23.825 53.645 ;
        RECT 23.995 53.295 24.745 53.815 ;
        RECT 24.915 53.740 25.205 54.905 ;
        RECT 25.385 53.795 25.680 54.905 ;
        RECT 25.860 53.595 26.110 54.730 ;
        RECT 26.280 53.795 26.540 54.905 ;
        RECT 26.710 54.005 26.970 54.730 ;
        RECT 27.140 54.175 27.400 54.905 ;
        RECT 27.570 54.005 27.830 54.730 ;
        RECT 28.000 54.175 28.260 54.905 ;
        RECT 28.430 54.005 28.690 54.730 ;
        RECT 28.860 54.175 29.120 54.905 ;
        RECT 29.290 54.005 29.550 54.730 ;
        RECT 29.720 54.175 30.015 54.905 ;
        RECT 26.710 53.765 30.020 54.005 ;
        RECT 30.475 53.955 30.765 54.725 ;
        RECT 31.335 54.365 31.595 54.725 ;
        RECT 31.765 54.535 32.095 54.905 ;
        RECT 32.265 54.365 32.525 54.725 ;
        RECT 31.335 54.135 32.525 54.365 ;
        RECT 32.715 54.185 33.045 54.905 ;
        RECT 33.215 53.955 33.480 54.725 ;
        RECT 33.655 54.470 39.000 54.905 ;
        RECT 39.175 54.470 44.520 54.905 ;
        RECT 30.475 53.775 32.970 53.955 ;
        RECT 22.185 52.355 22.355 52.965 ;
        RECT 22.525 52.575 22.855 53.010 ;
        RECT 23.075 52.355 24.745 53.125 ;
        RECT 24.915 52.355 25.205 53.080 ;
        RECT 25.375 52.985 25.690 53.595 ;
        RECT 25.860 53.345 28.880 53.595 ;
        RECT 25.435 52.355 25.680 52.815 ;
        RECT 25.860 52.535 26.110 53.345 ;
        RECT 29.050 53.175 30.020 53.765 ;
        RECT 30.445 53.265 30.715 53.595 ;
        RECT 30.895 53.265 31.330 53.595 ;
        RECT 31.510 53.265 32.085 53.595 ;
        RECT 32.265 53.265 32.545 53.595 ;
        RECT 26.710 53.005 30.020 53.175 ;
        RECT 32.745 53.085 32.970 53.775 ;
        RECT 26.280 52.355 26.540 52.880 ;
        RECT 26.710 52.550 26.970 53.005 ;
        RECT 27.140 52.355 27.400 52.835 ;
        RECT 27.570 52.550 27.830 53.005 ;
        RECT 28.000 52.355 28.260 52.835 ;
        RECT 28.430 52.550 28.690 53.005 ;
        RECT 28.860 52.355 29.120 52.835 ;
        RECT 29.290 52.550 29.550 53.005 ;
        RECT 30.485 52.895 32.970 53.085 ;
        RECT 29.720 52.355 30.020 52.835 ;
        RECT 30.485 52.535 30.710 52.895 ;
        RECT 30.890 52.355 31.220 52.725 ;
        RECT 31.400 52.535 31.655 52.895 ;
        RECT 32.220 52.355 32.965 52.725 ;
        RECT 33.145 52.535 33.480 53.955 ;
        RECT 35.240 52.900 35.580 53.730 ;
        RECT 37.060 53.220 37.410 54.470 ;
        RECT 40.760 52.900 41.100 53.730 ;
        RECT 42.580 53.220 42.930 54.470 ;
        RECT 44.695 53.815 47.285 54.905 ;
        RECT 44.695 53.125 45.905 53.645 ;
        RECT 46.075 53.295 47.285 53.815 ;
        RECT 47.460 53.955 47.725 54.725 ;
        RECT 47.895 54.185 48.225 54.905 ;
        RECT 48.415 54.365 48.675 54.725 ;
        RECT 48.845 54.535 49.175 54.905 ;
        RECT 49.345 54.365 49.605 54.725 ;
        RECT 48.415 54.135 49.605 54.365 ;
        RECT 50.175 53.955 50.465 54.725 ;
        RECT 33.655 52.355 39.000 52.900 ;
        RECT 39.175 52.355 44.520 52.900 ;
        RECT 44.695 52.355 47.285 53.125 ;
        RECT 47.460 52.535 47.795 53.955 ;
        RECT 47.970 53.775 50.465 53.955 ;
        RECT 47.970 53.085 48.195 53.775 ;
        RECT 50.675 53.740 50.965 54.905 ;
        RECT 52.145 54.235 52.315 54.735 ;
        RECT 52.485 54.405 52.815 54.905 ;
        RECT 52.145 54.065 52.810 54.235 ;
        RECT 48.395 53.265 48.675 53.595 ;
        RECT 48.855 53.265 49.430 53.595 ;
        RECT 49.610 53.265 50.045 53.595 ;
        RECT 50.225 53.265 50.495 53.595 ;
        RECT 52.060 53.245 52.410 53.895 ;
        RECT 47.970 52.895 50.455 53.085 ;
        RECT 47.975 52.355 48.720 52.725 ;
        RECT 49.285 52.535 49.540 52.895 ;
        RECT 49.720 52.355 50.050 52.725 ;
        RECT 50.230 52.535 50.455 52.895 ;
        RECT 50.675 52.355 50.965 53.080 ;
        RECT 52.580 53.075 52.810 54.065 ;
        RECT 52.145 52.905 52.810 53.075 ;
        RECT 52.145 52.615 52.315 52.905 ;
        RECT 52.485 52.355 52.815 52.735 ;
        RECT 52.985 52.615 53.170 54.735 ;
        RECT 53.410 54.445 53.675 54.905 ;
        RECT 53.845 54.310 54.095 54.735 ;
        RECT 54.305 54.460 55.410 54.630 ;
        RECT 53.790 54.180 54.095 54.310 ;
        RECT 53.340 52.985 53.620 53.935 ;
        RECT 53.790 53.075 53.960 54.180 ;
        RECT 54.130 53.395 54.370 53.990 ;
        RECT 54.540 53.925 55.070 54.290 ;
        RECT 54.540 53.225 54.710 53.925 ;
        RECT 55.240 53.845 55.410 54.460 ;
        RECT 55.580 54.105 55.750 54.905 ;
        RECT 55.920 54.405 56.170 54.735 ;
        RECT 56.395 54.435 57.280 54.605 ;
        RECT 55.240 53.755 55.750 53.845 ;
        RECT 53.790 52.945 54.015 53.075 ;
        RECT 54.185 53.005 54.710 53.225 ;
        RECT 54.880 53.585 55.750 53.755 ;
        RECT 53.425 52.355 53.675 52.815 ;
        RECT 53.845 52.805 54.015 52.945 ;
        RECT 54.880 52.805 55.050 53.585 ;
        RECT 55.580 53.515 55.750 53.585 ;
        RECT 55.260 53.335 55.460 53.365 ;
        RECT 55.920 53.335 56.090 54.405 ;
        RECT 56.260 53.515 56.450 54.235 ;
        RECT 55.260 53.035 56.090 53.335 ;
        RECT 56.620 53.305 56.940 54.265 ;
        RECT 53.845 52.635 54.180 52.805 ;
        RECT 54.375 52.635 55.050 52.805 ;
        RECT 55.370 52.355 55.740 52.855 ;
        RECT 55.920 52.805 56.090 53.035 ;
        RECT 56.475 52.975 56.940 53.305 ;
        RECT 57.110 53.595 57.280 54.435 ;
        RECT 57.460 54.405 57.775 54.905 ;
        RECT 58.005 54.175 58.345 54.735 ;
        RECT 57.450 53.800 58.345 54.175 ;
        RECT 58.515 53.895 58.685 54.905 ;
        RECT 58.155 53.595 58.345 53.800 ;
        RECT 58.855 53.845 59.185 54.690 ;
        RECT 59.475 53.845 59.805 54.690 ;
        RECT 59.975 53.895 60.145 54.905 ;
        RECT 60.315 54.175 60.655 54.735 ;
        RECT 60.885 54.405 61.200 54.905 ;
        RECT 61.380 54.435 62.265 54.605 ;
        RECT 58.855 53.765 59.245 53.845 ;
        RECT 59.030 53.715 59.245 53.765 ;
        RECT 57.110 53.265 57.985 53.595 ;
        RECT 58.155 53.265 58.905 53.595 ;
        RECT 57.110 52.805 57.280 53.265 ;
        RECT 58.155 53.095 58.355 53.265 ;
        RECT 59.075 53.135 59.245 53.715 ;
        RECT 59.020 53.095 59.245 53.135 ;
        RECT 55.920 52.635 56.325 52.805 ;
        RECT 56.495 52.635 57.280 52.805 ;
        RECT 57.555 52.355 57.765 52.885 ;
        RECT 58.025 52.570 58.355 53.095 ;
        RECT 58.865 53.010 59.245 53.095 ;
        RECT 59.415 53.765 59.805 53.845 ;
        RECT 60.315 53.800 61.210 54.175 ;
        RECT 59.415 53.715 59.630 53.765 ;
        RECT 59.415 53.135 59.585 53.715 ;
        RECT 60.315 53.595 60.505 53.800 ;
        RECT 61.380 53.595 61.550 54.435 ;
        RECT 62.490 54.405 62.740 54.735 ;
        RECT 59.755 53.265 60.505 53.595 ;
        RECT 60.675 53.265 61.550 53.595 ;
        RECT 59.415 53.095 59.640 53.135 ;
        RECT 60.305 53.095 60.505 53.265 ;
        RECT 59.415 53.010 59.795 53.095 ;
        RECT 58.525 52.355 58.695 52.965 ;
        RECT 58.865 52.575 59.195 53.010 ;
        RECT 59.465 52.575 59.795 53.010 ;
        RECT 59.965 52.355 60.135 52.965 ;
        RECT 60.305 52.570 60.635 53.095 ;
        RECT 60.895 52.355 61.105 52.885 ;
        RECT 61.380 52.805 61.550 53.265 ;
        RECT 61.720 53.305 62.040 54.265 ;
        RECT 62.210 53.515 62.400 54.235 ;
        RECT 62.570 53.335 62.740 54.405 ;
        RECT 62.910 54.105 63.080 54.905 ;
        RECT 63.250 54.460 64.355 54.630 ;
        RECT 63.250 53.845 63.420 54.460 ;
        RECT 64.565 54.310 64.815 54.735 ;
        RECT 64.985 54.445 65.250 54.905 ;
        RECT 63.590 53.925 64.120 54.290 ;
        RECT 64.565 54.180 64.870 54.310 ;
        RECT 62.910 53.755 63.420 53.845 ;
        RECT 62.910 53.585 63.780 53.755 ;
        RECT 62.910 53.515 63.080 53.585 ;
        RECT 63.200 53.335 63.400 53.365 ;
        RECT 61.720 52.975 62.185 53.305 ;
        RECT 62.570 53.035 63.400 53.335 ;
        RECT 62.570 52.805 62.740 53.035 ;
        RECT 61.380 52.635 62.165 52.805 ;
        RECT 62.335 52.635 62.740 52.805 ;
        RECT 62.920 52.355 63.290 52.855 ;
        RECT 63.610 52.805 63.780 53.585 ;
        RECT 63.950 53.225 64.120 53.925 ;
        RECT 64.290 53.395 64.530 53.990 ;
        RECT 63.950 53.005 64.475 53.225 ;
        RECT 64.700 53.075 64.870 54.180 ;
        RECT 64.645 52.945 64.870 53.075 ;
        RECT 65.040 52.985 65.320 53.935 ;
        RECT 64.645 52.805 64.815 52.945 ;
        RECT 63.610 52.635 64.285 52.805 ;
        RECT 64.480 52.635 64.815 52.805 ;
        RECT 64.985 52.355 65.235 52.815 ;
        RECT 65.490 52.615 65.675 54.735 ;
        RECT 65.845 54.405 66.175 54.905 ;
        RECT 66.345 54.235 66.515 54.735 ;
        RECT 65.850 54.065 66.515 54.235 ;
        RECT 65.850 53.075 66.080 54.065 ;
        RECT 66.250 53.245 66.600 53.895 ;
        RECT 66.835 53.845 67.165 54.690 ;
        RECT 67.335 53.895 67.505 54.905 ;
        RECT 67.675 54.175 68.015 54.735 ;
        RECT 68.245 54.405 68.560 54.905 ;
        RECT 68.740 54.435 69.625 54.605 ;
        RECT 66.775 53.765 67.165 53.845 ;
        RECT 67.675 53.800 68.570 54.175 ;
        RECT 66.775 53.715 66.990 53.765 ;
        RECT 66.775 53.135 66.945 53.715 ;
        RECT 67.675 53.595 67.865 53.800 ;
        RECT 68.740 53.595 68.910 54.435 ;
        RECT 69.850 54.405 70.100 54.735 ;
        RECT 67.115 53.265 67.865 53.595 ;
        RECT 68.035 53.265 68.910 53.595 ;
        RECT 66.775 53.095 67.000 53.135 ;
        RECT 67.665 53.095 67.865 53.265 ;
        RECT 65.850 52.905 66.515 53.075 ;
        RECT 66.775 53.010 67.155 53.095 ;
        RECT 65.845 52.355 66.175 52.735 ;
        RECT 66.345 52.615 66.515 52.905 ;
        RECT 66.825 52.575 67.155 53.010 ;
        RECT 67.325 52.355 67.495 52.965 ;
        RECT 67.665 52.570 67.995 53.095 ;
        RECT 68.255 52.355 68.465 52.885 ;
        RECT 68.740 52.805 68.910 53.265 ;
        RECT 69.080 53.305 69.400 54.265 ;
        RECT 69.570 53.515 69.760 54.235 ;
        RECT 69.930 53.335 70.100 54.405 ;
        RECT 70.270 54.105 70.440 54.905 ;
        RECT 70.610 54.460 71.715 54.630 ;
        RECT 70.610 53.845 70.780 54.460 ;
        RECT 71.925 54.310 72.175 54.735 ;
        RECT 72.345 54.445 72.610 54.905 ;
        RECT 70.950 53.925 71.480 54.290 ;
        RECT 71.925 54.180 72.230 54.310 ;
        RECT 70.270 53.755 70.780 53.845 ;
        RECT 70.270 53.585 71.140 53.755 ;
        RECT 70.270 53.515 70.440 53.585 ;
        RECT 70.560 53.335 70.760 53.365 ;
        RECT 69.080 52.975 69.545 53.305 ;
        RECT 69.930 53.035 70.760 53.335 ;
        RECT 69.930 52.805 70.100 53.035 ;
        RECT 68.740 52.635 69.525 52.805 ;
        RECT 69.695 52.635 70.100 52.805 ;
        RECT 70.280 52.355 70.650 52.855 ;
        RECT 70.970 52.805 71.140 53.585 ;
        RECT 71.310 53.225 71.480 53.925 ;
        RECT 71.650 53.395 71.890 53.990 ;
        RECT 71.310 53.005 71.835 53.225 ;
        RECT 72.060 53.075 72.230 54.180 ;
        RECT 72.005 52.945 72.230 53.075 ;
        RECT 72.400 52.985 72.680 53.935 ;
        RECT 72.005 52.805 72.175 52.945 ;
        RECT 70.970 52.635 71.645 52.805 ;
        RECT 71.840 52.635 72.175 52.805 ;
        RECT 72.345 52.355 72.595 52.815 ;
        RECT 72.850 52.615 73.035 54.735 ;
        RECT 73.205 54.405 73.535 54.905 ;
        RECT 73.705 54.235 73.875 54.735 ;
        RECT 73.210 54.065 73.875 54.235 ;
        RECT 73.210 53.075 73.440 54.065 ;
        RECT 73.610 53.245 73.960 53.895 ;
        RECT 74.135 53.765 74.415 54.905 ;
        RECT 74.585 53.755 74.915 54.735 ;
        RECT 75.085 53.765 75.345 54.905 ;
        RECT 74.145 53.325 74.480 53.595 ;
        RECT 74.650 53.155 74.820 53.755 ;
        RECT 76.435 53.740 76.725 54.905 ;
        RECT 76.895 53.765 77.280 54.735 ;
        RECT 77.450 54.445 77.775 54.905 ;
        RECT 78.295 54.275 78.575 54.735 ;
        RECT 77.450 54.055 78.575 54.275 ;
        RECT 74.990 53.345 75.325 53.595 ;
        RECT 73.210 52.905 73.875 53.075 ;
        RECT 73.205 52.355 73.535 52.735 ;
        RECT 73.705 52.615 73.875 52.905 ;
        RECT 74.135 52.355 74.445 53.155 ;
        RECT 74.650 52.525 75.345 53.155 ;
        RECT 76.895 53.095 77.175 53.765 ;
        RECT 77.450 53.595 77.900 54.055 ;
        RECT 78.765 53.885 79.165 54.735 ;
        RECT 79.565 54.445 79.835 54.905 ;
        RECT 80.005 54.275 80.290 54.735 ;
        RECT 77.345 53.265 77.900 53.595 ;
        RECT 78.070 53.325 79.165 53.885 ;
        RECT 77.450 53.155 77.900 53.265 ;
        RECT 76.435 52.355 76.725 53.080 ;
        RECT 76.895 52.525 77.280 53.095 ;
        RECT 77.450 52.985 78.575 53.155 ;
        RECT 77.450 52.355 77.775 52.815 ;
        RECT 78.295 52.525 78.575 52.985 ;
        RECT 78.765 52.525 79.165 53.325 ;
        RECT 79.335 54.055 80.290 54.275 ;
        RECT 79.335 53.155 79.545 54.055 ;
        RECT 79.715 53.325 80.405 53.885 ;
        RECT 81.040 53.765 81.375 54.735 ;
        RECT 81.545 53.765 81.715 54.905 ;
        RECT 81.885 54.565 83.915 54.735 ;
        RECT 79.335 52.985 80.290 53.155 ;
        RECT 79.565 52.355 79.835 52.815 ;
        RECT 80.005 52.525 80.290 52.985 ;
        RECT 81.040 53.095 81.210 53.765 ;
        RECT 81.885 53.595 82.055 54.565 ;
        RECT 81.380 53.265 81.635 53.595 ;
        RECT 81.860 53.265 82.055 53.595 ;
        RECT 82.225 54.225 83.350 54.395 ;
        RECT 81.465 53.095 81.635 53.265 ;
        RECT 82.225 53.095 82.395 54.225 ;
        RECT 81.040 52.525 81.295 53.095 ;
        RECT 81.465 52.925 82.395 53.095 ;
        RECT 82.565 53.885 83.575 54.055 ;
        RECT 82.565 53.085 82.735 53.885 ;
        RECT 82.220 52.890 82.395 52.925 ;
        RECT 81.465 52.355 81.795 52.755 ;
        RECT 82.220 52.525 82.750 52.890 ;
        RECT 82.940 52.865 83.215 53.685 ;
        RECT 82.935 52.695 83.215 52.865 ;
        RECT 82.940 52.525 83.215 52.695 ;
        RECT 83.385 52.525 83.575 53.885 ;
        RECT 83.745 53.900 83.915 54.565 ;
        RECT 84.085 54.145 84.255 54.905 ;
        RECT 84.490 54.145 85.005 54.555 ;
        RECT 83.745 53.710 84.495 53.900 ;
        RECT 84.665 53.335 85.005 54.145 ;
        RECT 83.775 53.165 85.005 53.335 ;
        RECT 85.175 53.765 85.560 54.735 ;
        RECT 85.730 54.445 86.055 54.905 ;
        RECT 86.575 54.275 86.855 54.735 ;
        RECT 85.730 54.055 86.855 54.275 ;
        RECT 83.755 52.355 84.265 52.890 ;
        RECT 84.485 52.560 84.730 53.165 ;
        RECT 85.175 53.095 85.455 53.765 ;
        RECT 85.730 53.595 86.180 54.055 ;
        RECT 87.045 53.885 87.445 54.735 ;
        RECT 87.845 54.445 88.115 54.905 ;
        RECT 88.285 54.275 88.570 54.735 ;
        RECT 85.625 53.265 86.180 53.595 ;
        RECT 86.350 53.325 87.445 53.885 ;
        RECT 85.730 53.155 86.180 53.265 ;
        RECT 85.175 52.525 85.560 53.095 ;
        RECT 85.730 52.985 86.855 53.155 ;
        RECT 85.730 52.355 86.055 52.815 ;
        RECT 86.575 52.525 86.855 52.985 ;
        RECT 87.045 52.525 87.445 53.325 ;
        RECT 87.615 54.055 88.570 54.275 ;
        RECT 87.615 53.155 87.825 54.055 ;
        RECT 87.995 53.325 88.685 53.885 ;
        RECT 89.315 53.815 90.525 54.905 ;
        RECT 89.315 53.275 89.835 53.815 ;
        RECT 87.615 52.985 88.570 53.155 ;
        RECT 90.005 53.105 90.525 53.645 ;
        RECT 87.845 52.355 88.115 52.815 ;
        RECT 88.285 52.525 88.570 52.985 ;
        RECT 89.315 52.355 90.525 53.105 ;
        RECT 11.950 52.185 90.610 52.355 ;
        RECT 12.035 51.435 13.245 52.185 ;
        RECT 12.035 50.895 12.555 51.435 ;
        RECT 13.420 51.345 13.680 52.185 ;
        RECT 13.855 51.440 14.110 52.015 ;
        RECT 14.280 51.805 14.610 52.185 ;
        RECT 14.825 51.635 14.995 52.015 ;
        RECT 14.280 51.465 14.995 51.635 ;
        RECT 12.725 50.725 13.245 51.265 ;
        RECT 12.035 49.635 13.245 50.725 ;
        RECT 13.420 49.635 13.680 50.785 ;
        RECT 13.855 50.710 14.025 51.440 ;
        RECT 14.280 51.275 14.450 51.465 ;
        RECT 15.260 51.345 15.520 52.185 ;
        RECT 15.695 51.440 15.950 52.015 ;
        RECT 16.120 51.805 16.450 52.185 ;
        RECT 16.665 51.635 16.835 52.015 ;
        RECT 17.095 51.640 22.440 52.185 ;
        RECT 23.240 51.675 23.480 52.185 ;
        RECT 23.660 51.675 23.940 52.005 ;
        RECT 24.170 51.675 24.385 52.185 ;
        RECT 16.120 51.465 16.835 51.635 ;
        RECT 14.195 50.945 14.450 51.275 ;
        RECT 14.280 50.735 14.450 50.945 ;
        RECT 14.730 50.915 15.085 51.285 ;
        RECT 13.855 49.805 14.110 50.710 ;
        RECT 14.280 50.565 14.995 50.735 ;
        RECT 14.280 49.635 14.610 50.395 ;
        RECT 14.825 49.805 14.995 50.565 ;
        RECT 15.260 49.635 15.520 50.785 ;
        RECT 15.695 50.710 15.865 51.440 ;
        RECT 16.120 51.275 16.290 51.465 ;
        RECT 16.035 50.945 16.290 51.275 ;
        RECT 16.120 50.735 16.290 50.945 ;
        RECT 16.570 50.915 16.925 51.285 ;
        RECT 18.680 50.810 19.020 51.640 ;
        RECT 15.695 49.805 15.950 50.710 ;
        RECT 16.120 50.565 16.835 50.735 ;
        RECT 16.120 49.635 16.450 50.395 ;
        RECT 16.665 49.805 16.835 50.565 ;
        RECT 20.500 50.070 20.850 51.320 ;
        RECT 23.135 50.945 23.490 51.505 ;
        RECT 23.660 50.775 23.830 51.675 ;
        RECT 24.000 50.945 24.265 51.505 ;
        RECT 24.555 51.445 25.170 52.015 ;
        RECT 25.620 51.705 25.920 52.185 ;
        RECT 26.090 51.535 26.350 51.990 ;
        RECT 26.520 51.705 26.780 52.185 ;
        RECT 26.950 51.535 27.210 51.990 ;
        RECT 27.380 51.705 27.640 52.185 ;
        RECT 27.810 51.535 28.070 51.990 ;
        RECT 28.240 51.705 28.500 52.185 ;
        RECT 28.670 51.535 28.930 51.990 ;
        RECT 29.100 51.660 29.360 52.185 ;
        RECT 24.515 50.775 24.685 51.275 ;
        RECT 23.260 50.605 24.685 50.775 ;
        RECT 23.260 50.430 23.650 50.605 ;
        RECT 17.095 49.635 22.440 50.070 ;
        RECT 24.135 49.635 24.465 50.435 ;
        RECT 24.855 50.425 25.170 51.445 ;
        RECT 25.620 51.365 28.930 51.535 ;
        RECT 25.620 50.775 26.590 51.365 ;
        RECT 29.530 51.195 29.780 52.005 ;
        RECT 29.960 51.725 30.205 52.185 ;
        RECT 30.600 51.675 30.840 52.185 ;
        RECT 31.020 51.675 31.300 52.005 ;
        RECT 31.530 51.675 31.745 52.185 ;
        RECT 26.760 50.945 29.780 51.195 ;
        RECT 29.950 50.945 30.265 51.555 ;
        RECT 30.495 50.945 30.850 51.505 ;
        RECT 25.620 50.535 28.930 50.775 ;
        RECT 24.635 49.805 25.170 50.425 ;
        RECT 25.625 49.635 25.920 50.365 ;
        RECT 26.090 49.810 26.350 50.535 ;
        RECT 26.520 49.635 26.780 50.365 ;
        RECT 26.950 49.810 27.210 50.535 ;
        RECT 27.380 49.635 27.640 50.365 ;
        RECT 27.810 49.810 28.070 50.535 ;
        RECT 28.240 49.635 28.500 50.365 ;
        RECT 28.670 49.810 28.930 50.535 ;
        RECT 29.100 49.635 29.360 50.745 ;
        RECT 29.530 49.810 29.780 50.945 ;
        RECT 31.020 50.775 31.190 51.675 ;
        RECT 31.360 50.945 31.625 51.505 ;
        RECT 31.915 51.445 32.530 52.015 ;
        RECT 31.875 50.775 32.045 51.275 ;
        RECT 29.960 49.635 30.255 50.745 ;
        RECT 30.620 50.605 32.045 50.775 ;
        RECT 30.620 50.430 31.010 50.605 ;
        RECT 31.495 49.635 31.825 50.435 ;
        RECT 32.215 50.425 32.530 51.445 ;
        RECT 32.735 51.415 34.405 52.185 ;
        RECT 35.095 51.715 35.395 52.185 ;
        RECT 35.565 51.545 35.820 51.990 ;
        RECT 35.990 51.715 36.250 52.185 ;
        RECT 36.420 51.545 36.680 51.990 ;
        RECT 36.850 51.715 37.145 52.185 ;
        RECT 32.735 50.895 33.485 51.415 ;
        RECT 34.575 51.375 37.605 51.545 ;
        RECT 37.795 51.460 38.085 52.185 ;
        RECT 33.655 50.725 34.405 51.245 ;
        RECT 31.995 49.805 32.530 50.425 ;
        RECT 32.735 49.635 34.405 50.725 ;
        RECT 34.575 50.810 34.875 51.375 ;
        RECT 35.050 50.980 37.265 51.205 ;
        RECT 37.435 50.810 37.605 51.375 ;
        RECT 34.575 50.640 37.605 50.810 ;
        RECT 34.575 49.635 34.960 50.470 ;
        RECT 35.130 49.835 35.390 50.640 ;
        RECT 35.560 49.635 35.820 50.470 ;
        RECT 35.990 49.835 36.245 50.640 ;
        RECT 36.420 49.635 36.680 50.470 ;
        RECT 36.850 49.835 37.105 50.640 ;
        RECT 37.280 49.635 37.625 50.470 ;
        RECT 37.795 49.635 38.085 50.800 ;
        RECT 38.720 50.585 39.055 52.005 ;
        RECT 39.235 51.815 39.980 52.185 ;
        RECT 40.545 51.645 40.800 52.005 ;
        RECT 40.980 51.815 41.310 52.185 ;
        RECT 41.490 51.645 41.715 52.005 ;
        RECT 39.230 51.455 41.715 51.645 ;
        RECT 42.485 51.635 42.655 51.925 ;
        RECT 42.825 51.805 43.155 52.185 ;
        RECT 42.485 51.465 43.150 51.635 ;
        RECT 39.230 50.765 39.455 51.455 ;
        RECT 39.655 50.945 39.935 51.275 ;
        RECT 40.115 50.945 40.690 51.275 ;
        RECT 40.870 50.945 41.305 51.275 ;
        RECT 41.485 50.945 41.755 51.275 ;
        RECT 39.230 50.585 41.725 50.765 ;
        RECT 42.400 50.645 42.750 51.295 ;
        RECT 38.720 49.815 38.985 50.585 ;
        RECT 39.155 49.635 39.485 50.355 ;
        RECT 39.675 50.175 40.865 50.405 ;
        RECT 39.675 49.815 39.935 50.175 ;
        RECT 40.105 49.635 40.435 50.005 ;
        RECT 40.605 49.815 40.865 50.175 ;
        RECT 41.435 49.815 41.725 50.585 ;
        RECT 42.920 50.475 43.150 51.465 ;
        RECT 42.485 50.305 43.150 50.475 ;
        RECT 42.485 49.805 42.655 50.305 ;
        RECT 42.825 49.635 43.155 50.135 ;
        RECT 43.325 49.805 43.510 51.925 ;
        RECT 43.765 51.725 44.015 52.185 ;
        RECT 44.185 51.735 44.520 51.905 ;
        RECT 44.715 51.735 45.390 51.905 ;
        RECT 44.185 51.595 44.355 51.735 ;
        RECT 43.680 50.605 43.960 51.555 ;
        RECT 44.130 51.465 44.355 51.595 ;
        RECT 44.130 50.360 44.300 51.465 ;
        RECT 44.525 51.315 45.050 51.535 ;
        RECT 44.470 50.550 44.710 51.145 ;
        RECT 44.880 50.615 45.050 51.315 ;
        RECT 45.220 50.955 45.390 51.735 ;
        RECT 45.710 51.685 46.080 52.185 ;
        RECT 46.260 51.735 46.665 51.905 ;
        RECT 46.835 51.735 47.620 51.905 ;
        RECT 46.260 51.505 46.430 51.735 ;
        RECT 45.600 51.205 46.430 51.505 ;
        RECT 46.815 51.235 47.280 51.565 ;
        RECT 45.600 51.175 45.800 51.205 ;
        RECT 45.920 50.955 46.090 51.025 ;
        RECT 45.220 50.785 46.090 50.955 ;
        RECT 45.580 50.695 46.090 50.785 ;
        RECT 44.130 50.230 44.435 50.360 ;
        RECT 44.880 50.250 45.410 50.615 ;
        RECT 43.750 49.635 44.015 50.095 ;
        RECT 44.185 49.805 44.435 50.230 ;
        RECT 45.580 50.080 45.750 50.695 ;
        RECT 44.645 49.910 45.750 50.080 ;
        RECT 45.920 49.635 46.090 50.435 ;
        RECT 46.260 50.135 46.430 51.205 ;
        RECT 46.600 50.305 46.790 51.025 ;
        RECT 46.960 50.275 47.280 51.235 ;
        RECT 47.450 51.275 47.620 51.735 ;
        RECT 47.895 51.655 48.105 52.185 ;
        RECT 48.365 51.445 48.695 51.970 ;
        RECT 48.865 51.575 49.035 52.185 ;
        RECT 49.205 51.530 49.535 51.965 ;
        RECT 49.845 51.635 50.015 51.925 ;
        RECT 50.185 51.805 50.515 52.185 ;
        RECT 49.205 51.445 49.585 51.530 ;
        RECT 49.845 51.465 50.510 51.635 ;
        RECT 48.495 51.275 48.695 51.445 ;
        RECT 49.360 51.405 49.585 51.445 ;
        RECT 47.450 50.945 48.325 51.275 ;
        RECT 48.495 50.945 49.245 51.275 ;
        RECT 46.260 49.805 46.510 50.135 ;
        RECT 47.450 50.105 47.620 50.945 ;
        RECT 48.495 50.740 48.685 50.945 ;
        RECT 49.415 50.825 49.585 51.405 ;
        RECT 49.370 50.775 49.585 50.825 ;
        RECT 47.790 50.365 48.685 50.740 ;
        RECT 49.195 50.695 49.585 50.775 ;
        RECT 46.735 49.935 47.620 50.105 ;
        RECT 47.800 49.635 48.115 50.135 ;
        RECT 48.345 49.805 48.685 50.365 ;
        RECT 48.855 49.635 49.025 50.645 ;
        RECT 49.195 49.850 49.525 50.695 ;
        RECT 49.760 50.645 50.110 51.295 ;
        RECT 50.280 50.475 50.510 51.465 ;
        RECT 49.845 50.305 50.510 50.475 ;
        RECT 49.845 49.805 50.015 50.305 ;
        RECT 50.185 49.635 50.515 50.135 ;
        RECT 50.685 49.805 50.870 51.925 ;
        RECT 51.125 51.725 51.375 52.185 ;
        RECT 51.545 51.735 51.880 51.905 ;
        RECT 52.075 51.735 52.750 51.905 ;
        RECT 51.545 51.595 51.715 51.735 ;
        RECT 51.040 50.605 51.320 51.555 ;
        RECT 51.490 51.465 51.715 51.595 ;
        RECT 51.490 50.360 51.660 51.465 ;
        RECT 51.885 51.315 52.410 51.535 ;
        RECT 51.830 50.550 52.070 51.145 ;
        RECT 52.240 50.615 52.410 51.315 ;
        RECT 52.580 50.955 52.750 51.735 ;
        RECT 53.070 51.685 53.440 52.185 ;
        RECT 53.620 51.735 54.025 51.905 ;
        RECT 54.195 51.735 54.980 51.905 ;
        RECT 53.620 51.505 53.790 51.735 ;
        RECT 52.960 51.205 53.790 51.505 ;
        RECT 54.175 51.235 54.640 51.565 ;
        RECT 52.960 51.175 53.160 51.205 ;
        RECT 53.280 50.955 53.450 51.025 ;
        RECT 52.580 50.785 53.450 50.955 ;
        RECT 52.940 50.695 53.450 50.785 ;
        RECT 51.490 50.230 51.795 50.360 ;
        RECT 52.240 50.250 52.770 50.615 ;
        RECT 51.110 49.635 51.375 50.095 ;
        RECT 51.545 49.805 51.795 50.230 ;
        RECT 52.940 50.080 53.110 50.695 ;
        RECT 52.005 49.910 53.110 50.080 ;
        RECT 53.280 49.635 53.450 50.435 ;
        RECT 53.620 50.135 53.790 51.205 ;
        RECT 53.960 50.305 54.150 51.025 ;
        RECT 54.320 50.275 54.640 51.235 ;
        RECT 54.810 51.275 54.980 51.735 ;
        RECT 55.255 51.655 55.465 52.185 ;
        RECT 55.725 51.445 56.055 51.970 ;
        RECT 56.225 51.575 56.395 52.185 ;
        RECT 56.565 51.530 56.895 51.965 ;
        RECT 56.565 51.445 56.945 51.530 ;
        RECT 55.855 51.275 56.055 51.445 ;
        RECT 56.720 51.405 56.945 51.445 ;
        RECT 54.810 50.945 55.685 51.275 ;
        RECT 55.855 50.945 56.605 51.275 ;
        RECT 53.620 49.805 53.870 50.135 ;
        RECT 54.810 50.105 54.980 50.945 ;
        RECT 55.855 50.740 56.045 50.945 ;
        RECT 56.775 50.825 56.945 51.405 ;
        RECT 56.730 50.775 56.945 50.825 ;
        RECT 55.150 50.365 56.045 50.740 ;
        RECT 56.555 50.695 56.945 50.775 ;
        RECT 57.120 51.445 57.375 52.015 ;
        RECT 57.545 51.785 57.875 52.185 ;
        RECT 58.300 51.650 58.830 52.015 ;
        RECT 59.020 51.845 59.295 52.015 ;
        RECT 59.015 51.675 59.295 51.845 ;
        RECT 58.300 51.615 58.475 51.650 ;
        RECT 57.545 51.445 58.475 51.615 ;
        RECT 57.120 50.775 57.290 51.445 ;
        RECT 57.545 51.275 57.715 51.445 ;
        RECT 57.460 50.945 57.715 51.275 ;
        RECT 57.940 50.945 58.135 51.275 ;
        RECT 54.095 49.935 54.980 50.105 ;
        RECT 55.160 49.635 55.475 50.135 ;
        RECT 55.705 49.805 56.045 50.365 ;
        RECT 56.215 49.635 56.385 50.645 ;
        RECT 56.555 49.850 56.885 50.695 ;
        RECT 57.120 49.805 57.455 50.775 ;
        RECT 57.625 49.635 57.795 50.775 ;
        RECT 57.965 49.975 58.135 50.945 ;
        RECT 58.305 50.315 58.475 51.445 ;
        RECT 58.645 50.655 58.815 51.455 ;
        RECT 59.020 50.855 59.295 51.675 ;
        RECT 59.465 50.655 59.655 52.015 ;
        RECT 59.835 51.650 60.345 52.185 ;
        RECT 60.565 51.375 60.810 51.980 ;
        RECT 61.255 51.415 62.925 52.185 ;
        RECT 63.555 51.460 63.845 52.185 ;
        RECT 64.015 51.640 69.360 52.185 ;
        RECT 69.535 51.640 74.880 52.185 ;
        RECT 59.855 51.205 61.085 51.375 ;
        RECT 58.645 50.485 59.655 50.655 ;
        RECT 59.825 50.640 60.575 50.830 ;
        RECT 58.305 50.145 59.430 50.315 ;
        RECT 59.825 49.975 59.995 50.640 ;
        RECT 60.745 50.395 61.085 51.205 ;
        RECT 61.255 50.895 62.005 51.415 ;
        RECT 62.175 50.725 62.925 51.245 ;
        RECT 65.600 50.810 65.940 51.640 ;
        RECT 57.965 49.805 59.995 49.975 ;
        RECT 60.165 49.635 60.335 50.395 ;
        RECT 60.570 49.985 61.085 50.395 ;
        RECT 61.255 49.635 62.925 50.725 ;
        RECT 63.555 49.635 63.845 50.800 ;
        RECT 67.420 50.070 67.770 51.320 ;
        RECT 71.120 50.810 71.460 51.640 ;
        RECT 75.055 51.415 76.725 52.185 ;
        RECT 72.940 50.070 73.290 51.320 ;
        RECT 75.055 50.895 75.805 51.415 ;
        RECT 76.935 51.365 77.165 52.185 ;
        RECT 77.335 51.385 77.665 52.015 ;
        RECT 75.975 50.725 76.725 51.245 ;
        RECT 76.915 50.945 77.245 51.195 ;
        RECT 77.415 50.785 77.665 51.385 ;
        RECT 77.835 51.365 78.045 52.185 ;
        RECT 78.275 51.640 83.620 52.185 ;
        RECT 79.860 50.810 80.200 51.640 ;
        RECT 83.795 51.415 87.305 52.185 ;
        RECT 87.935 51.510 88.195 52.015 ;
        RECT 88.375 51.805 88.705 52.185 ;
        RECT 88.885 51.635 89.055 52.015 ;
        RECT 64.015 49.635 69.360 50.070 ;
        RECT 69.535 49.635 74.880 50.070 ;
        RECT 75.055 49.635 76.725 50.725 ;
        RECT 76.935 49.635 77.165 50.775 ;
        RECT 77.335 49.805 77.665 50.785 ;
        RECT 77.835 49.635 78.045 50.775 ;
        RECT 81.680 50.070 82.030 51.320 ;
        RECT 83.795 50.895 85.445 51.415 ;
        RECT 85.615 50.725 87.305 51.245 ;
        RECT 78.275 49.635 83.620 50.070 ;
        RECT 83.795 49.635 87.305 50.725 ;
        RECT 87.935 50.710 88.105 51.510 ;
        RECT 88.390 51.465 89.055 51.635 ;
        RECT 88.390 51.210 88.560 51.465 ;
        RECT 89.315 51.435 90.525 52.185 ;
        RECT 88.275 50.880 88.560 51.210 ;
        RECT 88.795 50.915 89.125 51.285 ;
        RECT 88.390 50.735 88.560 50.880 ;
        RECT 87.935 49.805 88.205 50.710 ;
        RECT 88.390 50.565 89.055 50.735 ;
        RECT 88.375 49.635 88.705 50.395 ;
        RECT 88.885 49.805 89.055 50.565 ;
        RECT 89.315 50.725 89.835 51.265 ;
        RECT 90.005 50.895 90.525 51.435 ;
        RECT 89.315 49.635 90.525 50.725 ;
        RECT 11.950 49.465 90.610 49.635 ;
        RECT 12.035 48.375 13.245 49.465 ;
        RECT 12.035 47.665 12.555 48.205 ;
        RECT 12.725 47.835 13.245 48.375 ;
        RECT 13.420 48.315 13.680 49.465 ;
        RECT 13.855 48.390 14.110 49.295 ;
        RECT 14.280 48.705 14.610 49.465 ;
        RECT 14.825 48.535 14.995 49.295 ;
        RECT 12.035 46.915 13.245 47.665 ;
        RECT 13.420 46.915 13.680 47.755 ;
        RECT 13.855 47.660 14.025 48.390 ;
        RECT 14.280 48.365 14.995 48.535 ;
        RECT 16.380 48.495 16.710 49.295 ;
        RECT 16.880 48.665 17.210 49.465 ;
        RECT 17.510 48.495 17.840 49.295 ;
        RECT 18.485 48.665 18.735 49.465 ;
        RECT 14.280 48.155 14.450 48.365 ;
        RECT 16.380 48.325 18.815 48.495 ;
        RECT 19.005 48.325 19.175 49.465 ;
        RECT 19.345 48.325 19.685 49.295 ;
        RECT 14.195 47.825 14.450 48.155 ;
        RECT 13.855 47.085 14.110 47.660 ;
        RECT 14.280 47.635 14.450 47.825 ;
        RECT 14.730 47.815 15.085 48.185 ;
        RECT 16.175 47.905 16.525 48.155 ;
        RECT 16.710 47.695 16.880 48.325 ;
        RECT 17.050 47.905 17.380 48.105 ;
        RECT 17.550 47.905 17.880 48.105 ;
        RECT 18.050 47.905 18.470 48.105 ;
        RECT 18.645 48.075 18.815 48.325 ;
        RECT 18.645 47.905 19.340 48.075 ;
        RECT 14.280 47.465 14.995 47.635 ;
        RECT 14.280 46.915 14.610 47.295 ;
        RECT 14.825 47.085 14.995 47.465 ;
        RECT 16.380 47.085 16.880 47.695 ;
        RECT 17.510 47.565 18.735 47.735 ;
        RECT 19.510 47.715 19.685 48.325 ;
        RECT 19.860 48.315 20.120 49.465 ;
        RECT 20.295 48.390 20.550 49.295 ;
        RECT 20.720 48.705 21.050 49.465 ;
        RECT 21.265 48.535 21.435 49.295 ;
        RECT 17.510 47.085 17.840 47.565 ;
        RECT 18.010 46.915 18.235 47.375 ;
        RECT 18.405 47.085 18.735 47.565 ;
        RECT 18.925 46.915 19.175 47.715 ;
        RECT 19.345 47.085 19.685 47.715 ;
        RECT 19.860 46.915 20.120 47.755 ;
        RECT 20.295 47.660 20.465 48.390 ;
        RECT 20.720 48.365 21.435 48.535 ;
        RECT 21.695 48.375 24.285 49.465 ;
        RECT 20.720 48.155 20.890 48.365 ;
        RECT 20.635 47.825 20.890 48.155 ;
        RECT 20.295 47.085 20.550 47.660 ;
        RECT 20.720 47.635 20.890 47.825 ;
        RECT 21.170 47.815 21.525 48.185 ;
        RECT 21.695 47.685 22.905 48.205 ;
        RECT 23.075 47.855 24.285 48.375 ;
        RECT 24.915 48.300 25.205 49.465 ;
        RECT 26.040 48.495 26.370 49.295 ;
        RECT 26.540 48.665 26.870 49.465 ;
        RECT 27.170 48.495 27.500 49.295 ;
        RECT 28.145 48.665 28.395 49.465 ;
        RECT 26.040 48.325 28.475 48.495 ;
        RECT 28.665 48.325 28.835 49.465 ;
        RECT 29.005 48.325 29.345 49.295 ;
        RECT 29.605 48.795 29.775 49.295 ;
        RECT 29.945 48.965 30.275 49.465 ;
        RECT 29.605 48.625 30.270 48.795 ;
        RECT 25.835 47.905 26.185 48.155 ;
        RECT 26.370 47.695 26.540 48.325 ;
        RECT 26.710 47.905 27.040 48.105 ;
        RECT 27.210 47.905 27.540 48.105 ;
        RECT 27.710 47.905 28.130 48.105 ;
        RECT 28.305 48.075 28.475 48.325 ;
        RECT 28.305 47.905 29.000 48.075 ;
        RECT 29.170 47.765 29.345 48.325 ;
        RECT 29.520 47.805 29.870 48.455 ;
        RECT 20.720 47.465 21.435 47.635 ;
        RECT 20.720 46.915 21.050 47.295 ;
        RECT 21.265 47.085 21.435 47.465 ;
        RECT 21.695 46.915 24.285 47.685 ;
        RECT 24.915 46.915 25.205 47.640 ;
        RECT 26.040 47.085 26.540 47.695 ;
        RECT 27.170 47.565 28.395 47.735 ;
        RECT 29.115 47.715 29.345 47.765 ;
        RECT 27.170 47.085 27.500 47.565 ;
        RECT 27.670 46.915 27.895 47.375 ;
        RECT 28.065 47.085 28.395 47.565 ;
        RECT 28.585 46.915 28.835 47.715 ;
        RECT 29.005 47.085 29.345 47.715 ;
        RECT 30.040 47.635 30.270 48.625 ;
        RECT 29.605 47.465 30.270 47.635 ;
        RECT 29.605 47.175 29.775 47.465 ;
        RECT 29.945 46.915 30.275 47.295 ;
        RECT 30.445 47.175 30.630 49.295 ;
        RECT 30.870 49.005 31.135 49.465 ;
        RECT 31.305 48.870 31.555 49.295 ;
        RECT 31.765 49.020 32.870 49.190 ;
        RECT 31.250 48.740 31.555 48.870 ;
        RECT 30.800 47.545 31.080 48.495 ;
        RECT 31.250 47.635 31.420 48.740 ;
        RECT 31.590 47.955 31.830 48.550 ;
        RECT 32.000 48.485 32.530 48.850 ;
        RECT 32.000 47.785 32.170 48.485 ;
        RECT 32.700 48.405 32.870 49.020 ;
        RECT 33.040 48.665 33.210 49.465 ;
        RECT 33.380 48.965 33.630 49.295 ;
        RECT 33.855 48.995 34.740 49.165 ;
        RECT 32.700 48.315 33.210 48.405 ;
        RECT 31.250 47.505 31.475 47.635 ;
        RECT 31.645 47.565 32.170 47.785 ;
        RECT 32.340 48.145 33.210 48.315 ;
        RECT 30.885 46.915 31.135 47.375 ;
        RECT 31.305 47.365 31.475 47.505 ;
        RECT 32.340 47.365 32.510 48.145 ;
        RECT 33.040 48.075 33.210 48.145 ;
        RECT 32.720 47.895 32.920 47.925 ;
        RECT 33.380 47.895 33.550 48.965 ;
        RECT 33.720 48.075 33.910 48.795 ;
        RECT 32.720 47.595 33.550 47.895 ;
        RECT 34.080 47.865 34.400 48.825 ;
        RECT 31.305 47.195 31.640 47.365 ;
        RECT 31.835 47.195 32.510 47.365 ;
        RECT 32.830 46.915 33.200 47.415 ;
        RECT 33.380 47.365 33.550 47.595 ;
        RECT 33.935 47.535 34.400 47.865 ;
        RECT 34.570 48.155 34.740 48.995 ;
        RECT 34.920 48.965 35.235 49.465 ;
        RECT 35.465 48.735 35.805 49.295 ;
        RECT 34.910 48.360 35.805 48.735 ;
        RECT 35.975 48.455 36.145 49.465 ;
        RECT 35.615 48.155 35.805 48.360 ;
        RECT 36.315 48.405 36.645 49.250 ;
        RECT 36.965 48.795 37.135 49.295 ;
        RECT 37.305 48.965 37.635 49.465 ;
        RECT 36.965 48.625 37.630 48.795 ;
        RECT 36.315 48.325 36.705 48.405 ;
        RECT 36.490 48.275 36.705 48.325 ;
        RECT 34.570 47.825 35.445 48.155 ;
        RECT 35.615 47.825 36.365 48.155 ;
        RECT 34.570 47.365 34.740 47.825 ;
        RECT 35.615 47.655 35.815 47.825 ;
        RECT 36.535 47.695 36.705 48.275 ;
        RECT 36.880 47.805 37.230 48.455 ;
        RECT 36.480 47.655 36.705 47.695 ;
        RECT 33.380 47.195 33.785 47.365 ;
        RECT 33.955 47.195 34.740 47.365 ;
        RECT 35.015 46.915 35.225 47.445 ;
        RECT 35.485 47.130 35.815 47.655 ;
        RECT 36.325 47.570 36.705 47.655 ;
        RECT 37.400 47.635 37.630 48.625 ;
        RECT 35.985 46.915 36.155 47.525 ;
        RECT 36.325 47.135 36.655 47.570 ;
        RECT 36.965 47.465 37.630 47.635 ;
        RECT 36.965 47.175 37.135 47.465 ;
        RECT 37.305 46.915 37.635 47.295 ;
        RECT 37.805 47.175 37.990 49.295 ;
        RECT 38.230 49.005 38.495 49.465 ;
        RECT 38.665 48.870 38.915 49.295 ;
        RECT 39.125 49.020 40.230 49.190 ;
        RECT 38.610 48.740 38.915 48.870 ;
        RECT 38.160 47.545 38.440 48.495 ;
        RECT 38.610 47.635 38.780 48.740 ;
        RECT 38.950 47.955 39.190 48.550 ;
        RECT 39.360 48.485 39.890 48.850 ;
        RECT 39.360 47.785 39.530 48.485 ;
        RECT 40.060 48.405 40.230 49.020 ;
        RECT 40.400 48.665 40.570 49.465 ;
        RECT 40.740 48.965 40.990 49.295 ;
        RECT 41.215 48.995 42.100 49.165 ;
        RECT 40.060 48.315 40.570 48.405 ;
        RECT 38.610 47.505 38.835 47.635 ;
        RECT 39.005 47.565 39.530 47.785 ;
        RECT 39.700 48.145 40.570 48.315 ;
        RECT 38.245 46.915 38.495 47.375 ;
        RECT 38.665 47.365 38.835 47.505 ;
        RECT 39.700 47.365 39.870 48.145 ;
        RECT 40.400 48.075 40.570 48.145 ;
        RECT 40.080 47.895 40.280 47.925 ;
        RECT 40.740 47.895 40.910 48.965 ;
        RECT 41.080 48.075 41.270 48.795 ;
        RECT 40.080 47.595 40.910 47.895 ;
        RECT 41.440 47.865 41.760 48.825 ;
        RECT 38.665 47.195 39.000 47.365 ;
        RECT 39.195 47.195 39.870 47.365 ;
        RECT 40.190 46.915 40.560 47.415 ;
        RECT 40.740 47.365 40.910 47.595 ;
        RECT 41.295 47.535 41.760 47.865 ;
        RECT 41.930 48.155 42.100 48.995 ;
        RECT 42.280 48.965 42.595 49.465 ;
        RECT 42.825 48.735 43.165 49.295 ;
        RECT 42.270 48.360 43.165 48.735 ;
        RECT 43.335 48.455 43.505 49.465 ;
        RECT 42.975 48.155 43.165 48.360 ;
        RECT 43.675 48.405 44.005 49.250 ;
        RECT 43.675 48.325 44.065 48.405 ;
        RECT 43.850 48.275 44.065 48.325 ;
        RECT 41.930 47.825 42.805 48.155 ;
        RECT 42.975 47.825 43.725 48.155 ;
        RECT 41.930 47.365 42.100 47.825 ;
        RECT 42.975 47.655 43.175 47.825 ;
        RECT 43.895 47.695 44.065 48.275 ;
        RECT 43.840 47.655 44.065 47.695 ;
        RECT 40.740 47.195 41.145 47.365 ;
        RECT 41.315 47.195 42.100 47.365 ;
        RECT 42.375 46.915 42.585 47.445 ;
        RECT 42.845 47.130 43.175 47.655 ;
        RECT 43.685 47.570 44.065 47.655 ;
        RECT 44.240 48.325 44.575 49.295 ;
        RECT 44.745 48.325 44.915 49.465 ;
        RECT 45.085 49.125 47.115 49.295 ;
        RECT 44.240 47.655 44.410 48.325 ;
        RECT 45.085 48.155 45.255 49.125 ;
        RECT 44.580 47.825 44.835 48.155 ;
        RECT 45.060 47.825 45.255 48.155 ;
        RECT 45.425 48.785 46.550 48.955 ;
        RECT 44.665 47.655 44.835 47.825 ;
        RECT 45.425 47.655 45.595 48.785 ;
        RECT 43.345 46.915 43.515 47.525 ;
        RECT 43.685 47.135 44.015 47.570 ;
        RECT 44.240 47.085 44.495 47.655 ;
        RECT 44.665 47.485 45.595 47.655 ;
        RECT 45.765 48.445 46.775 48.615 ;
        RECT 45.765 47.645 45.935 48.445 ;
        RECT 46.140 47.765 46.415 48.245 ;
        RECT 46.135 47.595 46.415 47.765 ;
        RECT 45.420 47.450 45.595 47.485 ;
        RECT 44.665 46.915 44.995 47.315 ;
        RECT 45.420 47.085 45.950 47.450 ;
        RECT 46.140 47.085 46.415 47.595 ;
        RECT 46.585 47.085 46.775 48.445 ;
        RECT 46.945 48.460 47.115 49.125 ;
        RECT 47.285 48.705 47.455 49.465 ;
        RECT 47.690 48.705 48.205 49.115 ;
        RECT 46.945 48.270 47.695 48.460 ;
        RECT 47.865 47.895 48.205 48.705 ;
        RECT 48.375 48.375 50.045 49.465 ;
        RECT 46.975 47.725 48.205 47.895 ;
        RECT 46.955 46.915 47.465 47.450 ;
        RECT 47.685 47.120 47.930 47.725 ;
        RECT 48.375 47.685 49.125 48.205 ;
        RECT 49.295 47.855 50.045 48.375 ;
        RECT 50.675 48.300 50.965 49.465 ;
        RECT 51.135 48.325 51.520 49.295 ;
        RECT 51.690 49.005 52.015 49.465 ;
        RECT 52.535 48.835 52.815 49.295 ;
        RECT 51.690 48.615 52.815 48.835 ;
        RECT 48.375 46.915 50.045 47.685 ;
        RECT 51.135 47.655 51.415 48.325 ;
        RECT 51.690 48.155 52.140 48.615 ;
        RECT 53.005 48.445 53.405 49.295 ;
        RECT 53.805 49.005 54.075 49.465 ;
        RECT 54.245 48.835 54.530 49.295 ;
        RECT 54.815 48.960 55.445 49.465 ;
        RECT 51.585 47.825 52.140 48.155 ;
        RECT 52.310 47.885 53.405 48.445 ;
        RECT 51.690 47.715 52.140 47.825 ;
        RECT 50.675 46.915 50.965 47.640 ;
        RECT 51.135 47.085 51.520 47.655 ;
        RECT 51.690 47.545 52.815 47.715 ;
        RECT 51.690 46.915 52.015 47.375 ;
        RECT 52.535 47.085 52.815 47.545 ;
        RECT 53.005 47.085 53.405 47.885 ;
        RECT 53.575 48.615 54.530 48.835 ;
        RECT 53.575 47.715 53.785 48.615 ;
        RECT 53.955 47.885 54.645 48.445 ;
        RECT 54.830 48.425 55.085 48.790 ;
        RECT 55.255 48.785 55.445 48.960 ;
        RECT 55.625 48.955 56.100 49.295 ;
        RECT 55.255 48.595 55.585 48.785 ;
        RECT 55.810 48.425 56.060 48.720 ;
        RECT 56.285 48.620 56.500 49.465 ;
        RECT 56.700 48.625 56.975 49.295 ;
        RECT 54.830 48.255 56.620 48.425 ;
        RECT 56.805 48.275 56.975 48.625 ;
        RECT 57.145 48.455 57.405 49.465 ;
        RECT 57.575 48.495 57.845 49.265 ;
        RECT 58.015 48.685 58.345 49.465 ;
        RECT 58.550 48.860 58.735 49.265 ;
        RECT 58.905 49.040 59.240 49.465 ;
        RECT 58.550 48.685 59.215 48.860 ;
        RECT 57.575 48.325 58.705 48.495 ;
        RECT 53.575 47.545 54.530 47.715 ;
        RECT 54.815 47.595 55.200 48.075 ;
        RECT 53.805 46.915 54.075 47.375 ;
        RECT 54.245 47.085 54.530 47.545 ;
        RECT 55.370 47.400 55.625 48.255 ;
        RECT 54.835 47.135 55.625 47.400 ;
        RECT 55.795 47.580 56.205 48.075 ;
        RECT 56.390 47.825 56.620 48.255 ;
        RECT 56.790 47.755 57.405 48.275 ;
        RECT 55.795 47.135 56.025 47.580 ;
        RECT 56.790 47.545 56.960 47.755 ;
        RECT 56.205 46.915 56.535 47.410 ;
        RECT 56.710 47.085 56.960 47.545 ;
        RECT 57.130 46.915 57.405 47.575 ;
        RECT 57.575 47.415 57.745 48.325 ;
        RECT 57.915 47.575 58.275 48.155 ;
        RECT 58.455 47.825 58.705 48.325 ;
        RECT 58.875 47.655 59.215 48.685 ;
        RECT 59.415 48.375 60.625 49.465 ;
        RECT 58.530 47.485 59.215 47.655 ;
        RECT 59.415 47.665 59.935 48.205 ;
        RECT 60.105 47.835 60.625 48.375 ;
        RECT 60.795 48.615 61.055 49.295 ;
        RECT 61.225 48.685 61.475 49.465 ;
        RECT 61.725 48.915 61.975 49.295 ;
        RECT 62.145 49.085 62.500 49.465 ;
        RECT 63.505 49.075 63.840 49.295 ;
        RECT 63.105 48.915 63.335 48.955 ;
        RECT 61.725 48.715 63.335 48.915 ;
        RECT 61.725 48.705 62.560 48.715 ;
        RECT 63.150 48.625 63.335 48.715 ;
        RECT 57.575 47.085 57.835 47.415 ;
        RECT 58.045 46.915 58.320 47.395 ;
        RECT 58.530 47.085 58.735 47.485 ;
        RECT 58.905 46.915 59.240 47.315 ;
        RECT 59.415 46.915 60.625 47.665 ;
        RECT 60.795 47.415 60.965 48.615 ;
        RECT 62.665 48.515 62.995 48.545 ;
        RECT 61.195 48.455 62.995 48.515 ;
        RECT 63.585 48.455 63.840 49.075 ;
        RECT 64.015 48.870 64.450 49.295 ;
        RECT 64.620 49.040 65.005 49.465 ;
        RECT 64.015 48.700 65.005 48.870 ;
        RECT 61.135 48.345 63.840 48.455 ;
        RECT 61.135 48.310 61.335 48.345 ;
        RECT 61.135 47.735 61.305 48.310 ;
        RECT 62.665 48.285 63.840 48.345 ;
        RECT 61.535 47.870 61.945 48.175 ;
        RECT 62.115 47.905 62.445 48.115 ;
        RECT 61.135 47.615 61.405 47.735 ;
        RECT 61.135 47.570 61.980 47.615 ;
        RECT 61.225 47.445 61.980 47.570 ;
        RECT 62.235 47.505 62.445 47.905 ;
        RECT 62.690 47.905 63.165 48.115 ;
        RECT 63.355 47.905 63.845 48.105 ;
        RECT 62.690 47.505 62.910 47.905 ;
        RECT 64.015 47.825 64.500 48.530 ;
        RECT 64.670 48.155 65.005 48.700 ;
        RECT 65.175 48.505 65.600 49.295 ;
        RECT 65.770 48.870 66.045 49.295 ;
        RECT 66.215 49.040 66.600 49.465 ;
        RECT 65.770 48.675 66.600 48.870 ;
        RECT 65.175 48.325 66.080 48.505 ;
        RECT 64.670 47.825 65.080 48.155 ;
        RECT 65.250 47.825 66.080 48.325 ;
        RECT 66.250 48.155 66.600 48.675 ;
        RECT 66.770 48.505 67.015 49.295 ;
        RECT 67.205 48.870 67.460 49.295 ;
        RECT 67.630 49.040 68.015 49.465 ;
        RECT 67.205 48.675 68.015 48.870 ;
        RECT 66.770 48.325 67.495 48.505 ;
        RECT 66.250 47.825 66.675 48.155 ;
        RECT 66.845 47.825 67.495 48.325 ;
        RECT 67.665 48.155 68.015 48.675 ;
        RECT 68.185 48.325 68.445 49.295 ;
        RECT 67.665 47.825 68.090 48.155 ;
        RECT 60.795 47.085 61.055 47.415 ;
        RECT 61.810 47.295 61.980 47.445 ;
        RECT 61.225 46.915 61.555 47.275 ;
        RECT 61.810 47.085 63.110 47.295 ;
        RECT 63.385 46.915 63.840 47.680 ;
        RECT 64.670 47.655 65.005 47.825 ;
        RECT 65.250 47.655 65.600 47.825 ;
        RECT 66.250 47.655 66.600 47.825 ;
        RECT 66.845 47.655 67.015 47.825 ;
        RECT 67.665 47.655 68.015 47.825 ;
        RECT 68.260 47.655 68.445 48.325 ;
        RECT 68.620 49.075 68.955 49.295 ;
        RECT 69.960 49.085 70.315 49.465 ;
        RECT 68.620 48.455 68.875 49.075 ;
        RECT 69.125 48.915 69.355 48.955 ;
        RECT 70.485 48.915 70.735 49.295 ;
        RECT 69.125 48.715 70.735 48.915 ;
        RECT 69.125 48.625 69.310 48.715 ;
        RECT 69.900 48.705 70.735 48.715 ;
        RECT 70.985 48.685 71.235 49.465 ;
        RECT 71.405 48.615 71.665 49.295 ;
        RECT 69.465 48.515 69.795 48.545 ;
        RECT 69.465 48.455 71.265 48.515 ;
        RECT 68.620 48.345 71.325 48.455 ;
        RECT 68.620 48.285 69.795 48.345 ;
        RECT 71.125 48.310 71.325 48.345 ;
        RECT 68.615 47.905 69.105 48.105 ;
        RECT 69.295 47.905 69.770 48.115 ;
        RECT 64.015 47.485 65.005 47.655 ;
        RECT 64.015 47.085 64.450 47.485 ;
        RECT 64.620 46.915 65.005 47.315 ;
        RECT 65.175 47.085 65.600 47.655 ;
        RECT 65.790 47.485 66.600 47.655 ;
        RECT 65.790 47.085 66.045 47.485 ;
        RECT 66.215 46.915 66.600 47.315 ;
        RECT 66.770 47.085 67.015 47.655 ;
        RECT 67.205 47.485 68.015 47.655 ;
        RECT 67.205 47.085 67.460 47.485 ;
        RECT 67.630 46.915 68.015 47.315 ;
        RECT 68.185 47.085 68.445 47.655 ;
        RECT 68.620 46.915 69.075 47.680 ;
        RECT 69.550 47.505 69.770 47.905 ;
        RECT 70.015 47.905 70.345 48.115 ;
        RECT 70.015 47.505 70.225 47.905 ;
        RECT 70.515 47.870 70.925 48.175 ;
        RECT 71.155 47.735 71.325 48.310 ;
        RECT 71.055 47.615 71.325 47.735 ;
        RECT 70.480 47.570 71.325 47.615 ;
        RECT 70.480 47.445 71.235 47.570 ;
        RECT 70.480 47.295 70.650 47.445 ;
        RECT 71.495 47.415 71.665 48.615 ;
        RECT 69.350 47.085 70.650 47.295 ;
        RECT 70.905 46.915 71.235 47.275 ;
        RECT 71.405 47.085 71.665 47.415 ;
        RECT 71.870 48.675 72.405 49.295 ;
        RECT 71.870 47.655 72.185 48.675 ;
        RECT 72.575 48.665 72.905 49.465 ;
        RECT 73.390 48.495 73.780 48.670 ;
        RECT 72.355 48.325 73.780 48.495 ;
        RECT 74.135 48.375 75.805 49.465 ;
        RECT 72.355 47.825 72.525 48.325 ;
        RECT 71.870 47.085 72.485 47.655 ;
        RECT 72.775 47.595 73.040 48.155 ;
        RECT 73.210 47.425 73.380 48.325 ;
        RECT 73.550 47.595 73.905 48.155 ;
        RECT 74.135 47.685 74.885 48.205 ;
        RECT 75.055 47.855 75.805 48.375 ;
        RECT 76.435 48.300 76.725 49.465 ;
        RECT 77.100 48.495 77.430 49.295 ;
        RECT 77.600 48.665 77.930 49.465 ;
        RECT 78.230 48.495 78.560 49.295 ;
        RECT 79.205 48.665 79.455 49.465 ;
        RECT 77.100 48.325 79.535 48.495 ;
        RECT 79.725 48.325 79.895 49.465 ;
        RECT 80.065 48.325 80.405 49.295 ;
        RECT 80.575 49.030 85.920 49.465 ;
        RECT 76.895 47.905 77.245 48.155 ;
        RECT 77.430 47.695 77.600 48.325 ;
        RECT 77.770 47.905 78.100 48.105 ;
        RECT 78.270 47.905 78.600 48.105 ;
        RECT 78.770 47.905 79.190 48.105 ;
        RECT 79.365 48.075 79.535 48.325 ;
        RECT 79.365 47.905 80.060 48.075 ;
        RECT 72.655 46.915 72.870 47.425 ;
        RECT 73.100 47.095 73.380 47.425 ;
        RECT 73.560 46.915 73.800 47.425 ;
        RECT 74.135 46.915 75.805 47.685 ;
        RECT 76.435 46.915 76.725 47.640 ;
        RECT 77.100 47.085 77.600 47.695 ;
        RECT 78.230 47.565 79.455 47.735 ;
        RECT 80.230 47.715 80.405 48.325 ;
        RECT 78.230 47.085 78.560 47.565 ;
        RECT 78.730 46.915 78.955 47.375 ;
        RECT 79.125 47.085 79.455 47.565 ;
        RECT 79.645 46.915 79.895 47.715 ;
        RECT 80.065 47.085 80.405 47.715 ;
        RECT 82.160 47.460 82.500 48.290 ;
        RECT 83.980 47.780 84.330 49.030 ;
        RECT 86.095 48.375 88.685 49.465 ;
        RECT 86.095 47.685 87.305 48.205 ;
        RECT 87.475 47.855 88.685 48.375 ;
        RECT 89.315 48.375 90.525 49.465 ;
        RECT 89.315 47.835 89.835 48.375 ;
        RECT 80.575 46.915 85.920 47.460 ;
        RECT 86.095 46.915 88.685 47.685 ;
        RECT 90.005 47.665 90.525 48.205 ;
        RECT 89.315 46.915 90.525 47.665 ;
        RECT 11.950 46.745 90.610 46.915 ;
        RECT 12.035 45.995 13.245 46.745 ;
        RECT 13.415 45.995 14.625 46.745 ;
        RECT 14.960 46.235 15.200 46.745 ;
        RECT 15.380 46.235 15.660 46.565 ;
        RECT 15.890 46.235 16.105 46.745 ;
        RECT 12.035 45.455 12.555 45.995 ;
        RECT 12.725 45.285 13.245 45.825 ;
        RECT 13.415 45.455 13.935 45.995 ;
        RECT 14.105 45.285 14.625 45.825 ;
        RECT 14.855 45.505 15.210 46.065 ;
        RECT 15.380 45.335 15.550 46.235 ;
        RECT 15.720 45.505 15.985 46.065 ;
        RECT 16.275 46.005 16.890 46.575 ;
        RECT 17.185 46.195 17.355 46.485 ;
        RECT 17.525 46.365 17.855 46.745 ;
        RECT 17.185 46.025 17.850 46.195 ;
        RECT 16.235 45.335 16.405 45.835 ;
        RECT 12.035 44.195 13.245 45.285 ;
        RECT 13.415 44.195 14.625 45.285 ;
        RECT 14.980 45.165 16.405 45.335 ;
        RECT 14.980 44.990 15.370 45.165 ;
        RECT 15.855 44.195 16.185 44.995 ;
        RECT 16.575 44.985 16.890 46.005 ;
        RECT 17.100 45.205 17.450 45.855 ;
        RECT 17.620 45.035 17.850 46.025 ;
        RECT 16.355 44.365 16.890 44.985 ;
        RECT 17.185 44.865 17.850 45.035 ;
        RECT 17.185 44.365 17.355 44.865 ;
        RECT 17.525 44.195 17.855 44.695 ;
        RECT 18.025 44.365 18.210 46.485 ;
        RECT 18.465 46.285 18.715 46.745 ;
        RECT 18.885 46.295 19.220 46.465 ;
        RECT 19.415 46.295 20.090 46.465 ;
        RECT 18.885 46.155 19.055 46.295 ;
        RECT 18.380 45.165 18.660 46.115 ;
        RECT 18.830 46.025 19.055 46.155 ;
        RECT 18.830 44.920 19.000 46.025 ;
        RECT 19.225 45.875 19.750 46.095 ;
        RECT 19.170 45.110 19.410 45.705 ;
        RECT 19.580 45.175 19.750 45.875 ;
        RECT 19.920 45.515 20.090 46.295 ;
        RECT 20.410 46.245 20.780 46.745 ;
        RECT 20.960 46.295 21.365 46.465 ;
        RECT 21.535 46.295 22.320 46.465 ;
        RECT 20.960 46.065 21.130 46.295 ;
        RECT 20.300 45.765 21.130 46.065 ;
        RECT 21.515 45.795 21.980 46.125 ;
        RECT 20.300 45.735 20.500 45.765 ;
        RECT 20.620 45.515 20.790 45.585 ;
        RECT 19.920 45.345 20.790 45.515 ;
        RECT 20.280 45.255 20.790 45.345 ;
        RECT 18.830 44.790 19.135 44.920 ;
        RECT 19.580 44.810 20.110 45.175 ;
        RECT 18.450 44.195 18.715 44.655 ;
        RECT 18.885 44.365 19.135 44.790 ;
        RECT 20.280 44.640 20.450 45.255 ;
        RECT 19.345 44.470 20.450 44.640 ;
        RECT 20.620 44.195 20.790 44.995 ;
        RECT 20.960 44.695 21.130 45.765 ;
        RECT 21.300 44.865 21.490 45.585 ;
        RECT 21.660 44.835 21.980 45.795 ;
        RECT 22.150 45.835 22.320 46.295 ;
        RECT 22.595 46.215 22.805 46.745 ;
        RECT 23.065 46.005 23.395 46.530 ;
        RECT 23.565 46.135 23.735 46.745 ;
        RECT 23.905 46.090 24.235 46.525 ;
        RECT 24.620 46.235 24.860 46.745 ;
        RECT 25.040 46.235 25.320 46.565 ;
        RECT 25.550 46.235 25.765 46.745 ;
        RECT 23.905 46.005 24.285 46.090 ;
        RECT 23.195 45.835 23.395 46.005 ;
        RECT 24.060 45.965 24.285 46.005 ;
        RECT 22.150 45.505 23.025 45.835 ;
        RECT 23.195 45.505 23.945 45.835 ;
        RECT 20.960 44.365 21.210 44.695 ;
        RECT 22.150 44.665 22.320 45.505 ;
        RECT 23.195 45.300 23.385 45.505 ;
        RECT 24.115 45.385 24.285 45.965 ;
        RECT 24.515 45.505 24.870 46.065 ;
        RECT 24.070 45.335 24.285 45.385 ;
        RECT 25.040 45.335 25.210 46.235 ;
        RECT 25.380 45.505 25.645 46.065 ;
        RECT 25.935 46.005 26.550 46.575 ;
        RECT 25.895 45.335 26.065 45.835 ;
        RECT 22.490 44.925 23.385 45.300 ;
        RECT 23.895 45.255 24.285 45.335 ;
        RECT 21.435 44.495 22.320 44.665 ;
        RECT 22.500 44.195 22.815 44.695 ;
        RECT 23.045 44.365 23.385 44.925 ;
        RECT 23.555 44.195 23.725 45.205 ;
        RECT 23.895 44.410 24.225 45.255 ;
        RECT 24.640 45.165 26.065 45.335 ;
        RECT 24.640 44.990 25.030 45.165 ;
        RECT 25.515 44.195 25.845 44.995 ;
        RECT 26.235 44.985 26.550 46.005 ;
        RECT 26.960 45.965 27.460 46.575 ;
        RECT 26.755 45.505 27.105 45.755 ;
        RECT 27.290 45.335 27.460 45.965 ;
        RECT 28.090 46.095 28.420 46.575 ;
        RECT 28.590 46.285 28.815 46.745 ;
        RECT 28.985 46.095 29.315 46.575 ;
        RECT 28.090 45.925 29.315 46.095 ;
        RECT 29.505 45.945 29.755 46.745 ;
        RECT 29.925 45.945 30.265 46.575 ;
        RECT 30.525 46.195 30.695 46.485 ;
        RECT 30.865 46.365 31.195 46.745 ;
        RECT 30.525 46.025 31.190 46.195 ;
        RECT 27.630 45.555 27.960 45.755 ;
        RECT 28.130 45.555 28.460 45.755 ;
        RECT 28.630 45.555 29.050 45.755 ;
        RECT 29.225 45.585 29.920 45.755 ;
        RECT 29.225 45.335 29.395 45.585 ;
        RECT 30.090 45.385 30.265 45.945 ;
        RECT 30.035 45.335 30.265 45.385 ;
        RECT 26.015 44.365 26.550 44.985 ;
        RECT 26.960 45.165 29.395 45.335 ;
        RECT 26.960 44.365 27.290 45.165 ;
        RECT 27.460 44.195 27.790 44.995 ;
        RECT 28.090 44.365 28.420 45.165 ;
        RECT 29.065 44.195 29.315 44.995 ;
        RECT 29.585 44.195 29.755 45.335 ;
        RECT 29.925 44.365 30.265 45.335 ;
        RECT 30.440 45.205 30.790 45.855 ;
        RECT 30.960 45.035 31.190 46.025 ;
        RECT 30.525 44.865 31.190 45.035 ;
        RECT 30.525 44.365 30.695 44.865 ;
        RECT 30.865 44.195 31.195 44.695 ;
        RECT 31.365 44.365 31.550 46.485 ;
        RECT 31.805 46.285 32.055 46.745 ;
        RECT 32.225 46.295 32.560 46.465 ;
        RECT 32.755 46.295 33.430 46.465 ;
        RECT 32.225 46.155 32.395 46.295 ;
        RECT 31.720 45.165 32.000 46.115 ;
        RECT 32.170 46.025 32.395 46.155 ;
        RECT 32.170 44.920 32.340 46.025 ;
        RECT 32.565 45.875 33.090 46.095 ;
        RECT 32.510 45.110 32.750 45.705 ;
        RECT 32.920 45.175 33.090 45.875 ;
        RECT 33.260 45.515 33.430 46.295 ;
        RECT 33.750 46.245 34.120 46.745 ;
        RECT 34.300 46.295 34.705 46.465 ;
        RECT 34.875 46.295 35.660 46.465 ;
        RECT 34.300 46.065 34.470 46.295 ;
        RECT 33.640 45.765 34.470 46.065 ;
        RECT 34.855 45.795 35.320 46.125 ;
        RECT 33.640 45.735 33.840 45.765 ;
        RECT 33.960 45.515 34.130 45.585 ;
        RECT 33.260 45.345 34.130 45.515 ;
        RECT 33.620 45.255 34.130 45.345 ;
        RECT 32.170 44.790 32.475 44.920 ;
        RECT 32.920 44.810 33.450 45.175 ;
        RECT 31.790 44.195 32.055 44.655 ;
        RECT 32.225 44.365 32.475 44.790 ;
        RECT 33.620 44.640 33.790 45.255 ;
        RECT 32.685 44.470 33.790 44.640 ;
        RECT 33.960 44.195 34.130 44.995 ;
        RECT 34.300 44.695 34.470 45.765 ;
        RECT 34.640 44.865 34.830 45.585 ;
        RECT 35.000 44.835 35.320 45.795 ;
        RECT 35.490 45.835 35.660 46.295 ;
        RECT 35.935 46.215 36.145 46.745 ;
        RECT 36.405 46.005 36.735 46.530 ;
        RECT 36.905 46.135 37.075 46.745 ;
        RECT 37.245 46.090 37.575 46.525 ;
        RECT 37.245 46.005 37.625 46.090 ;
        RECT 37.795 46.020 38.085 46.745 ;
        RECT 38.315 46.285 38.560 46.745 ;
        RECT 36.535 45.835 36.735 46.005 ;
        RECT 37.400 45.965 37.625 46.005 ;
        RECT 35.490 45.505 36.365 45.835 ;
        RECT 36.535 45.505 37.285 45.835 ;
        RECT 34.300 44.365 34.550 44.695 ;
        RECT 35.490 44.665 35.660 45.505 ;
        RECT 36.535 45.300 36.725 45.505 ;
        RECT 37.455 45.385 37.625 45.965 ;
        RECT 38.255 45.505 38.570 46.115 ;
        RECT 38.740 45.755 38.990 46.565 ;
        RECT 39.160 46.220 39.420 46.745 ;
        RECT 39.590 46.095 39.850 46.550 ;
        RECT 40.020 46.265 40.280 46.745 ;
        RECT 40.450 46.095 40.710 46.550 ;
        RECT 40.880 46.265 41.140 46.745 ;
        RECT 41.310 46.095 41.570 46.550 ;
        RECT 41.740 46.265 42.000 46.745 ;
        RECT 42.170 46.095 42.430 46.550 ;
        RECT 42.600 46.265 42.900 46.745 ;
        RECT 39.590 45.925 42.900 46.095 ;
        RECT 38.740 45.505 41.760 45.755 ;
        RECT 37.410 45.335 37.625 45.385 ;
        RECT 35.830 44.925 36.725 45.300 ;
        RECT 37.235 45.255 37.625 45.335 ;
        RECT 34.775 44.495 35.660 44.665 ;
        RECT 35.840 44.195 36.155 44.695 ;
        RECT 36.385 44.365 36.725 44.925 ;
        RECT 36.895 44.195 37.065 45.205 ;
        RECT 37.235 44.410 37.565 45.255 ;
        RECT 37.795 44.195 38.085 45.360 ;
        RECT 38.265 44.195 38.560 45.305 ;
        RECT 38.740 44.370 38.990 45.505 ;
        RECT 41.930 45.335 42.900 45.925 ;
        RECT 39.160 44.195 39.420 45.305 ;
        RECT 39.590 45.095 42.900 45.335 ;
        RECT 43.315 46.005 43.700 46.575 ;
        RECT 43.870 46.285 44.195 46.745 ;
        RECT 44.715 46.115 44.995 46.575 ;
        RECT 43.315 45.335 43.595 46.005 ;
        RECT 43.870 45.945 44.995 46.115 ;
        RECT 43.870 45.835 44.320 45.945 ;
        RECT 43.765 45.505 44.320 45.835 ;
        RECT 45.185 45.775 45.585 46.575 ;
        RECT 45.985 46.285 46.255 46.745 ;
        RECT 46.425 46.115 46.710 46.575 ;
        RECT 39.590 44.370 39.850 45.095 ;
        RECT 40.020 44.195 40.280 44.925 ;
        RECT 40.450 44.370 40.710 45.095 ;
        RECT 40.880 44.195 41.140 44.925 ;
        RECT 41.310 44.370 41.570 45.095 ;
        RECT 41.740 44.195 42.000 44.925 ;
        RECT 42.170 44.370 42.430 45.095 ;
        RECT 42.600 44.195 42.895 44.925 ;
        RECT 43.315 44.365 43.700 45.335 ;
        RECT 43.870 45.045 44.320 45.505 ;
        RECT 44.490 45.215 45.585 45.775 ;
        RECT 43.870 44.825 44.995 45.045 ;
        RECT 43.870 44.195 44.195 44.655 ;
        RECT 44.715 44.365 44.995 44.825 ;
        RECT 45.185 44.365 45.585 45.215 ;
        RECT 45.755 45.945 46.710 46.115 ;
        RECT 46.995 46.245 47.295 46.575 ;
        RECT 47.465 46.265 47.740 46.745 ;
        RECT 45.755 45.045 45.965 45.945 ;
        RECT 46.135 45.215 46.825 45.775 ;
        RECT 46.995 45.335 47.165 46.245 ;
        RECT 47.920 46.095 48.215 46.485 ;
        RECT 48.385 46.265 48.640 46.745 ;
        RECT 48.815 46.095 49.075 46.485 ;
        RECT 49.245 46.265 49.525 46.745 ;
        RECT 47.335 45.505 47.685 46.075 ;
        RECT 47.920 45.925 49.570 46.095 ;
        RECT 49.760 45.925 50.035 46.745 ;
        RECT 50.205 46.105 50.535 46.575 ;
        RECT 50.705 46.275 50.875 46.745 ;
        RECT 51.045 46.105 51.375 46.575 ;
        RECT 51.545 46.275 52.255 46.745 ;
        RECT 52.425 46.105 52.755 46.575 ;
        RECT 52.925 46.275 53.215 46.745 ;
        RECT 50.205 45.925 53.265 46.105 ;
        RECT 47.855 45.585 48.995 45.755 ;
        RECT 47.855 45.335 48.025 45.585 ;
        RECT 49.165 45.415 49.570 45.925 ;
        RECT 49.805 45.545 50.635 45.755 ;
        RECT 50.805 45.545 51.855 45.755 ;
        RECT 52.045 45.545 52.635 45.755 ;
        RECT 46.995 45.165 48.025 45.335 ;
        RECT 48.815 45.245 49.570 45.415 ;
        RECT 45.755 44.825 46.710 45.045 ;
        RECT 45.985 44.195 46.255 44.655 ;
        RECT 46.425 44.365 46.710 44.825 ;
        RECT 46.995 44.365 47.305 45.165 ;
        RECT 48.815 44.995 49.075 45.245 ;
        RECT 49.820 45.205 51.755 45.375 ;
        RECT 52.045 45.205 52.310 45.545 ;
        RECT 52.805 45.375 53.265 45.925 ;
        RECT 53.435 45.975 55.105 46.745 ;
        RECT 55.285 46.255 55.615 46.745 ;
        RECT 55.785 46.150 56.405 46.575 ;
        RECT 53.435 45.455 54.185 45.975 ;
        RECT 52.505 45.205 53.265 45.375 ;
        RECT 54.355 45.285 55.105 45.805 ;
        RECT 55.275 45.505 55.615 46.085 ;
        RECT 55.785 45.815 56.145 46.150 ;
        RECT 56.865 46.055 57.195 46.745 ;
        RECT 59.065 46.365 60.235 46.575 ;
        RECT 59.065 46.345 59.395 46.365 ;
        RECT 58.955 45.925 59.815 46.175 ;
        RECT 59.985 46.115 60.235 46.365 ;
        RECT 60.405 46.285 60.575 46.745 ;
        RECT 60.745 46.115 61.085 46.575 ;
        RECT 59.985 45.945 61.085 46.115 ;
        RECT 61.255 45.975 62.925 46.745 ;
        RECT 63.555 46.020 63.845 46.745 ;
        RECT 64.015 45.975 65.685 46.745 ;
        RECT 65.860 46.275 66.190 46.745 ;
        RECT 66.360 46.105 66.585 46.550 ;
        RECT 66.755 46.220 67.050 46.745 ;
        RECT 67.755 46.285 68.000 46.745 ;
        RECT 55.785 45.535 57.205 45.815 ;
        RECT 47.475 44.195 47.785 44.995 ;
        RECT 47.955 44.825 49.075 44.995 ;
        RECT 47.955 44.365 48.215 44.825 ;
        RECT 48.385 44.195 48.640 44.655 ;
        RECT 48.815 44.365 49.075 44.825 ;
        RECT 49.245 44.195 49.530 45.065 ;
        RECT 49.820 44.365 50.075 45.205 ;
        RECT 50.245 44.195 50.495 45.035 ;
        RECT 50.665 44.365 50.915 45.205 ;
        RECT 51.085 44.535 51.335 45.035 ;
        RECT 51.505 44.705 51.755 45.205 ;
        RECT 52.085 44.535 52.295 45.035 ;
        RECT 52.505 44.705 52.715 45.205 ;
        RECT 52.885 44.535 53.135 45.035 ;
        RECT 51.085 44.365 53.135 44.535 ;
        RECT 53.435 44.195 55.105 45.285 ;
        RECT 55.285 44.195 55.615 45.335 ;
        RECT 55.785 44.365 56.145 45.535 ;
        RECT 56.345 44.195 56.675 45.365 ;
        RECT 56.875 44.365 57.205 45.535 ;
        RECT 57.405 44.195 57.735 45.365 ;
        RECT 58.955 45.335 59.235 45.925 ;
        RECT 59.405 45.505 60.155 45.755 ;
        RECT 60.325 45.505 61.085 45.755 ;
        RECT 61.255 45.455 62.005 45.975 ;
        RECT 58.955 45.165 60.655 45.335 ;
        RECT 59.060 44.195 59.315 44.995 ;
        RECT 59.485 44.365 59.815 45.165 ;
        RECT 59.985 44.195 60.155 44.995 ;
        RECT 60.325 44.365 60.655 45.165 ;
        RECT 60.825 44.195 61.085 45.335 ;
        RECT 62.175 45.285 62.925 45.805 ;
        RECT 64.015 45.455 64.765 45.975 ;
        RECT 65.855 45.935 66.585 46.105 ;
        RECT 61.255 44.195 62.925 45.285 ;
        RECT 63.555 44.195 63.845 45.360 ;
        RECT 64.935 45.285 65.685 45.805 ;
        RECT 64.015 44.195 65.685 45.285 ;
        RECT 65.855 45.370 66.135 45.935 ;
        RECT 66.305 45.540 67.525 45.765 ;
        RECT 67.695 45.505 68.010 46.115 ;
        RECT 68.180 45.755 68.430 46.565 ;
        RECT 68.600 46.220 68.860 46.745 ;
        RECT 69.030 46.095 69.290 46.550 ;
        RECT 69.460 46.265 69.720 46.745 ;
        RECT 69.890 46.095 70.150 46.550 ;
        RECT 70.320 46.265 70.580 46.745 ;
        RECT 70.750 46.095 71.010 46.550 ;
        RECT 71.180 46.265 71.440 46.745 ;
        RECT 71.610 46.095 71.870 46.550 ;
        RECT 72.040 46.265 72.340 46.745 ;
        RECT 72.845 46.195 73.015 46.485 ;
        RECT 73.185 46.365 73.515 46.745 ;
        RECT 69.030 45.925 72.340 46.095 ;
        RECT 72.845 46.025 73.510 46.195 ;
        RECT 68.180 45.505 71.200 45.755 ;
        RECT 65.855 45.200 67.455 45.370 ;
        RECT 65.915 44.195 66.170 45.030 ;
        RECT 66.340 44.395 66.600 45.200 ;
        RECT 66.770 44.195 67.030 45.030 ;
        RECT 67.200 44.395 67.455 45.200 ;
        RECT 67.705 44.195 68.000 45.305 ;
        RECT 68.180 44.370 68.430 45.505 ;
        RECT 71.370 45.335 72.340 45.925 ;
        RECT 68.600 44.195 68.860 45.305 ;
        RECT 69.030 45.095 72.340 45.335 ;
        RECT 72.760 45.205 73.110 45.855 ;
        RECT 69.030 44.370 69.290 45.095 ;
        RECT 69.460 44.195 69.720 44.925 ;
        RECT 69.890 44.370 70.150 45.095 ;
        RECT 70.320 44.195 70.580 44.925 ;
        RECT 70.750 44.370 71.010 45.095 ;
        RECT 71.180 44.195 71.440 44.925 ;
        RECT 71.610 44.370 71.870 45.095 ;
        RECT 73.280 45.035 73.510 46.025 ;
        RECT 72.040 44.195 72.335 44.925 ;
        RECT 72.845 44.865 73.510 45.035 ;
        RECT 72.845 44.365 73.015 44.865 ;
        RECT 73.185 44.195 73.515 44.695 ;
        RECT 73.685 44.365 73.870 46.485 ;
        RECT 74.125 46.285 74.375 46.745 ;
        RECT 74.545 46.295 74.880 46.465 ;
        RECT 75.075 46.295 75.750 46.465 ;
        RECT 74.545 46.155 74.715 46.295 ;
        RECT 74.040 45.165 74.320 46.115 ;
        RECT 74.490 46.025 74.715 46.155 ;
        RECT 74.490 44.920 74.660 46.025 ;
        RECT 74.885 45.875 75.410 46.095 ;
        RECT 74.830 45.110 75.070 45.705 ;
        RECT 75.240 45.175 75.410 45.875 ;
        RECT 75.580 45.515 75.750 46.295 ;
        RECT 76.070 46.245 76.440 46.745 ;
        RECT 76.620 46.295 77.025 46.465 ;
        RECT 77.195 46.295 77.980 46.465 ;
        RECT 76.620 46.065 76.790 46.295 ;
        RECT 75.960 45.765 76.790 46.065 ;
        RECT 77.175 45.795 77.640 46.125 ;
        RECT 75.960 45.735 76.160 45.765 ;
        RECT 76.280 45.515 76.450 45.585 ;
        RECT 75.580 45.345 76.450 45.515 ;
        RECT 75.940 45.255 76.450 45.345 ;
        RECT 74.490 44.790 74.795 44.920 ;
        RECT 75.240 44.810 75.770 45.175 ;
        RECT 74.110 44.195 74.375 44.655 ;
        RECT 74.545 44.365 74.795 44.790 ;
        RECT 75.940 44.640 76.110 45.255 ;
        RECT 75.005 44.470 76.110 44.640 ;
        RECT 76.280 44.195 76.450 44.995 ;
        RECT 76.620 44.695 76.790 45.765 ;
        RECT 76.960 44.865 77.150 45.585 ;
        RECT 77.320 44.835 77.640 45.795 ;
        RECT 77.810 45.835 77.980 46.295 ;
        RECT 78.255 46.215 78.465 46.745 ;
        RECT 78.725 46.005 79.055 46.530 ;
        RECT 79.225 46.135 79.395 46.745 ;
        RECT 79.565 46.090 79.895 46.525 ;
        RECT 80.115 46.200 85.460 46.745 ;
        RECT 79.565 46.005 79.945 46.090 ;
        RECT 78.855 45.835 79.055 46.005 ;
        RECT 79.720 45.965 79.945 46.005 ;
        RECT 77.810 45.505 78.685 45.835 ;
        RECT 78.855 45.505 79.605 45.835 ;
        RECT 76.620 44.365 76.870 44.695 ;
        RECT 77.810 44.665 77.980 45.505 ;
        RECT 78.855 45.300 79.045 45.505 ;
        RECT 79.775 45.385 79.945 45.965 ;
        RECT 79.730 45.335 79.945 45.385 ;
        RECT 81.700 45.370 82.040 46.200 ;
        RECT 85.635 45.975 87.305 46.745 ;
        RECT 87.565 46.195 87.735 46.575 ;
        RECT 87.950 46.365 88.280 46.745 ;
        RECT 87.565 46.025 88.280 46.195 ;
        RECT 78.150 44.925 79.045 45.300 ;
        RECT 79.555 45.255 79.945 45.335 ;
        RECT 77.095 44.495 77.980 44.665 ;
        RECT 78.160 44.195 78.475 44.695 ;
        RECT 78.705 44.365 79.045 44.925 ;
        RECT 79.215 44.195 79.385 45.205 ;
        RECT 79.555 44.410 79.885 45.255 ;
        RECT 83.520 44.630 83.870 45.880 ;
        RECT 85.635 45.455 86.385 45.975 ;
        RECT 86.555 45.285 87.305 45.805 ;
        RECT 87.475 45.475 87.830 45.845 ;
        RECT 88.110 45.835 88.280 46.025 ;
        RECT 88.450 46.000 88.705 46.575 ;
        RECT 88.110 45.505 88.365 45.835 ;
        RECT 88.110 45.295 88.280 45.505 ;
        RECT 80.115 44.195 85.460 44.630 ;
        RECT 85.635 44.195 87.305 45.285 ;
        RECT 87.565 45.125 88.280 45.295 ;
        RECT 88.535 45.270 88.705 46.000 ;
        RECT 88.880 45.905 89.140 46.745 ;
        RECT 89.315 45.995 90.525 46.745 ;
        RECT 87.565 44.365 87.735 45.125 ;
        RECT 87.950 44.195 88.280 44.955 ;
        RECT 88.450 44.365 88.705 45.270 ;
        RECT 88.880 44.195 89.140 45.345 ;
        RECT 89.315 45.285 89.835 45.825 ;
        RECT 90.005 45.455 90.525 45.995 ;
        RECT 89.315 44.195 90.525 45.285 ;
        RECT 11.950 44.025 90.610 44.195 ;
        RECT 12.035 42.935 13.245 44.025 ;
        RECT 13.505 43.355 13.675 43.855 ;
        RECT 13.845 43.525 14.175 44.025 ;
        RECT 13.505 43.185 14.170 43.355 ;
        RECT 12.035 42.225 12.555 42.765 ;
        RECT 12.725 42.395 13.245 42.935 ;
        RECT 13.420 42.365 13.770 43.015 ;
        RECT 12.035 41.475 13.245 42.225 ;
        RECT 13.940 42.195 14.170 43.185 ;
        RECT 13.505 42.025 14.170 42.195 ;
        RECT 13.505 41.735 13.675 42.025 ;
        RECT 13.845 41.475 14.175 41.855 ;
        RECT 14.345 41.735 14.530 43.855 ;
        RECT 14.770 43.565 15.035 44.025 ;
        RECT 15.205 43.430 15.455 43.855 ;
        RECT 15.665 43.580 16.770 43.750 ;
        RECT 15.150 43.300 15.455 43.430 ;
        RECT 14.700 42.105 14.980 43.055 ;
        RECT 15.150 42.195 15.320 43.300 ;
        RECT 15.490 42.515 15.730 43.110 ;
        RECT 15.900 43.045 16.430 43.410 ;
        RECT 15.900 42.345 16.070 43.045 ;
        RECT 16.600 42.965 16.770 43.580 ;
        RECT 16.940 43.225 17.110 44.025 ;
        RECT 17.280 43.525 17.530 43.855 ;
        RECT 17.755 43.555 18.640 43.725 ;
        RECT 16.600 42.875 17.110 42.965 ;
        RECT 15.150 42.065 15.375 42.195 ;
        RECT 15.545 42.125 16.070 42.345 ;
        RECT 16.240 42.705 17.110 42.875 ;
        RECT 14.785 41.475 15.035 41.935 ;
        RECT 15.205 41.925 15.375 42.065 ;
        RECT 16.240 41.925 16.410 42.705 ;
        RECT 16.940 42.635 17.110 42.705 ;
        RECT 16.620 42.455 16.820 42.485 ;
        RECT 17.280 42.455 17.450 43.525 ;
        RECT 17.620 42.635 17.810 43.355 ;
        RECT 16.620 42.155 17.450 42.455 ;
        RECT 17.980 42.425 18.300 43.385 ;
        RECT 15.205 41.755 15.540 41.925 ;
        RECT 15.735 41.755 16.410 41.925 ;
        RECT 16.730 41.475 17.100 41.975 ;
        RECT 17.280 41.925 17.450 42.155 ;
        RECT 17.835 42.095 18.300 42.425 ;
        RECT 18.470 42.715 18.640 43.555 ;
        RECT 18.820 43.525 19.135 44.025 ;
        RECT 19.365 43.295 19.705 43.855 ;
        RECT 18.810 42.920 19.705 43.295 ;
        RECT 19.875 43.015 20.045 44.025 ;
        RECT 19.515 42.715 19.705 42.920 ;
        RECT 20.215 42.965 20.545 43.810 ;
        RECT 20.215 42.885 20.605 42.965 ;
        RECT 20.390 42.835 20.605 42.885 ;
        RECT 20.780 42.875 21.040 44.025 ;
        RECT 21.215 42.950 21.470 43.855 ;
        RECT 21.640 43.265 21.970 44.025 ;
        RECT 22.185 43.095 22.355 43.855 ;
        RECT 18.470 42.385 19.345 42.715 ;
        RECT 19.515 42.385 20.265 42.715 ;
        RECT 18.470 41.925 18.640 42.385 ;
        RECT 19.515 42.215 19.715 42.385 ;
        RECT 20.435 42.255 20.605 42.835 ;
        RECT 20.380 42.215 20.605 42.255 ;
        RECT 17.280 41.755 17.685 41.925 ;
        RECT 17.855 41.755 18.640 41.925 ;
        RECT 18.915 41.475 19.125 42.005 ;
        RECT 19.385 41.690 19.715 42.215 ;
        RECT 20.225 42.130 20.605 42.215 ;
        RECT 19.885 41.475 20.055 42.085 ;
        RECT 20.225 41.695 20.555 42.130 ;
        RECT 20.780 41.475 21.040 42.315 ;
        RECT 21.215 42.220 21.385 42.950 ;
        RECT 21.640 42.925 22.355 43.095 ;
        RECT 22.615 42.935 24.285 44.025 ;
        RECT 21.640 42.715 21.810 42.925 ;
        RECT 21.555 42.385 21.810 42.715 ;
        RECT 21.215 41.645 21.470 42.220 ;
        RECT 21.640 42.195 21.810 42.385 ;
        RECT 22.090 42.375 22.445 42.745 ;
        RECT 22.615 42.245 23.365 42.765 ;
        RECT 23.535 42.415 24.285 42.935 ;
        RECT 24.915 42.860 25.205 44.025 ;
        RECT 25.415 43.075 25.705 43.845 ;
        RECT 26.275 43.485 26.535 43.845 ;
        RECT 26.705 43.655 27.035 44.025 ;
        RECT 27.205 43.485 27.465 43.845 ;
        RECT 26.275 43.255 27.465 43.485 ;
        RECT 27.655 43.305 27.985 44.025 ;
        RECT 28.155 43.075 28.420 43.845 ;
        RECT 28.700 43.565 28.870 44.025 ;
        RECT 29.040 43.395 29.370 43.855 ;
        RECT 25.415 42.895 27.910 43.075 ;
        RECT 25.385 42.385 25.655 42.715 ;
        RECT 25.835 42.385 26.270 42.715 ;
        RECT 26.450 42.385 27.025 42.715 ;
        RECT 27.205 42.385 27.485 42.715 ;
        RECT 21.640 42.025 22.355 42.195 ;
        RECT 21.640 41.475 21.970 41.855 ;
        RECT 22.185 41.645 22.355 42.025 ;
        RECT 22.615 41.475 24.285 42.245 ;
        RECT 27.685 42.205 27.910 42.895 ;
        RECT 24.915 41.475 25.205 42.200 ;
        RECT 25.425 42.015 27.910 42.205 ;
        RECT 25.425 41.655 25.650 42.015 ;
        RECT 25.830 41.475 26.160 41.845 ;
        RECT 26.340 41.655 26.595 42.015 ;
        RECT 27.160 41.475 27.905 41.845 ;
        RECT 28.085 41.655 28.420 43.075 ;
        RECT 28.595 43.225 29.370 43.395 ;
        RECT 29.540 43.225 29.710 44.025 ;
        RECT 28.595 42.215 29.025 43.225 ;
        RECT 30.295 43.055 30.655 43.230 ;
        RECT 29.195 42.885 30.655 43.055 ;
        RECT 30.935 42.885 31.165 44.025 ;
        RECT 29.195 42.385 29.365 42.885 ;
        RECT 28.595 42.045 29.290 42.215 ;
        RECT 29.535 42.155 29.945 42.715 ;
        RECT 28.620 41.475 28.950 41.875 ;
        RECT 29.120 41.775 29.290 42.045 ;
        RECT 30.115 41.985 30.295 42.885 ;
        RECT 31.335 42.875 31.665 43.855 ;
        RECT 31.835 42.885 32.045 44.025 ;
        RECT 32.275 43.590 37.620 44.025 ;
        RECT 30.465 42.665 30.660 42.715 ;
        RECT 30.465 42.495 30.665 42.665 ;
        RECT 30.465 42.155 30.660 42.495 ;
        RECT 30.915 42.465 31.245 42.715 ;
        RECT 29.460 41.475 29.775 41.985 ;
        RECT 30.005 41.645 30.295 41.985 ;
        RECT 30.465 41.475 30.705 41.985 ;
        RECT 30.935 41.475 31.165 42.295 ;
        RECT 31.415 42.275 31.665 42.875 ;
        RECT 31.335 41.645 31.665 42.275 ;
        RECT 31.835 41.475 32.045 42.295 ;
        RECT 33.860 42.020 34.200 42.850 ;
        RECT 35.680 42.340 36.030 43.590 ;
        RECT 38.260 42.885 38.595 43.855 ;
        RECT 38.765 42.885 38.935 44.025 ;
        RECT 39.105 43.685 41.135 43.855 ;
        RECT 38.260 42.215 38.430 42.885 ;
        RECT 39.105 42.715 39.275 43.685 ;
        RECT 38.600 42.385 38.855 42.715 ;
        RECT 39.080 42.385 39.275 42.715 ;
        RECT 39.445 43.345 40.570 43.515 ;
        RECT 38.685 42.215 38.855 42.385 ;
        RECT 39.445 42.215 39.615 43.345 ;
        RECT 32.275 41.475 37.620 42.020 ;
        RECT 38.260 41.645 38.515 42.215 ;
        RECT 38.685 42.045 39.615 42.215 ;
        RECT 39.785 43.005 40.795 43.175 ;
        RECT 39.785 42.205 39.955 43.005 ;
        RECT 40.160 42.665 40.435 42.805 ;
        RECT 40.155 42.495 40.435 42.665 ;
        RECT 39.440 42.010 39.615 42.045 ;
        RECT 38.685 41.475 39.015 41.875 ;
        RECT 39.440 41.645 39.970 42.010 ;
        RECT 40.160 41.645 40.435 42.495 ;
        RECT 40.605 41.645 40.795 43.005 ;
        RECT 40.965 43.020 41.135 43.685 ;
        RECT 41.305 43.265 41.475 44.025 ;
        RECT 41.710 43.265 42.225 43.675 ;
        RECT 40.965 42.830 41.715 43.020 ;
        RECT 41.885 42.455 42.225 43.265 ;
        RECT 43.405 43.355 43.575 43.855 ;
        RECT 43.745 43.525 44.075 44.025 ;
        RECT 43.405 43.185 44.070 43.355 ;
        RECT 40.995 42.285 42.225 42.455 ;
        RECT 43.320 42.365 43.670 43.015 ;
        RECT 40.975 41.475 41.485 42.010 ;
        RECT 41.705 41.680 41.950 42.285 ;
        RECT 43.840 42.195 44.070 43.185 ;
        RECT 43.405 42.025 44.070 42.195 ;
        RECT 43.405 41.735 43.575 42.025 ;
        RECT 43.745 41.475 44.075 41.855 ;
        RECT 44.245 41.735 44.430 43.855 ;
        RECT 44.670 43.565 44.935 44.025 ;
        RECT 45.105 43.430 45.355 43.855 ;
        RECT 45.565 43.580 46.670 43.750 ;
        RECT 45.050 43.300 45.355 43.430 ;
        RECT 44.600 42.105 44.880 43.055 ;
        RECT 45.050 42.195 45.220 43.300 ;
        RECT 45.390 42.515 45.630 43.110 ;
        RECT 45.800 43.045 46.330 43.410 ;
        RECT 45.800 42.345 45.970 43.045 ;
        RECT 46.500 42.965 46.670 43.580 ;
        RECT 46.840 43.225 47.010 44.025 ;
        RECT 47.180 43.525 47.430 43.855 ;
        RECT 47.655 43.555 48.540 43.725 ;
        RECT 46.500 42.875 47.010 42.965 ;
        RECT 45.050 42.065 45.275 42.195 ;
        RECT 45.445 42.125 45.970 42.345 ;
        RECT 46.140 42.705 47.010 42.875 ;
        RECT 44.685 41.475 44.935 41.935 ;
        RECT 45.105 41.925 45.275 42.065 ;
        RECT 46.140 41.925 46.310 42.705 ;
        RECT 46.840 42.635 47.010 42.705 ;
        RECT 46.520 42.455 46.720 42.485 ;
        RECT 47.180 42.455 47.350 43.525 ;
        RECT 47.520 42.635 47.710 43.355 ;
        RECT 46.520 42.155 47.350 42.455 ;
        RECT 47.880 42.425 48.200 43.385 ;
        RECT 45.105 41.755 45.440 41.925 ;
        RECT 45.635 41.755 46.310 41.925 ;
        RECT 46.630 41.475 47.000 41.975 ;
        RECT 47.180 41.925 47.350 42.155 ;
        RECT 47.735 42.095 48.200 42.425 ;
        RECT 48.370 42.715 48.540 43.555 ;
        RECT 48.720 43.525 49.035 44.025 ;
        RECT 49.265 43.295 49.605 43.855 ;
        RECT 48.710 42.920 49.605 43.295 ;
        RECT 49.775 43.015 49.945 44.025 ;
        RECT 49.415 42.715 49.605 42.920 ;
        RECT 50.115 42.965 50.445 43.810 ;
        RECT 50.115 42.885 50.505 42.965 ;
        RECT 50.290 42.835 50.505 42.885 ;
        RECT 50.675 42.860 50.965 44.025 ;
        RECT 51.175 42.885 51.405 44.025 ;
        RECT 51.575 42.875 51.905 43.855 ;
        RECT 52.075 42.885 52.285 44.025 ;
        RECT 52.605 43.355 52.775 43.855 ;
        RECT 52.945 43.525 53.275 44.025 ;
        RECT 52.605 43.185 53.270 43.355 ;
        RECT 48.370 42.385 49.245 42.715 ;
        RECT 49.415 42.385 50.165 42.715 ;
        RECT 48.370 41.925 48.540 42.385 ;
        RECT 49.415 42.215 49.615 42.385 ;
        RECT 50.335 42.255 50.505 42.835 ;
        RECT 51.155 42.465 51.485 42.715 ;
        RECT 50.280 42.215 50.505 42.255 ;
        RECT 47.180 41.755 47.585 41.925 ;
        RECT 47.755 41.755 48.540 41.925 ;
        RECT 48.815 41.475 49.025 42.005 ;
        RECT 49.285 41.690 49.615 42.215 ;
        RECT 50.125 42.130 50.505 42.215 ;
        RECT 49.785 41.475 49.955 42.085 ;
        RECT 50.125 41.695 50.455 42.130 ;
        RECT 50.675 41.475 50.965 42.200 ;
        RECT 51.175 41.475 51.405 42.295 ;
        RECT 51.655 42.275 51.905 42.875 ;
        RECT 52.520 42.365 52.870 43.015 ;
        RECT 51.575 41.645 51.905 42.275 ;
        RECT 52.075 41.475 52.285 42.295 ;
        RECT 53.040 42.195 53.270 43.185 ;
        RECT 52.605 42.025 53.270 42.195 ;
        RECT 52.605 41.735 52.775 42.025 ;
        RECT 52.945 41.475 53.275 41.855 ;
        RECT 53.445 41.735 53.630 43.855 ;
        RECT 53.870 43.565 54.135 44.025 ;
        RECT 54.305 43.430 54.555 43.855 ;
        RECT 54.765 43.580 55.870 43.750 ;
        RECT 54.250 43.300 54.555 43.430 ;
        RECT 53.800 42.105 54.080 43.055 ;
        RECT 54.250 42.195 54.420 43.300 ;
        RECT 54.590 42.515 54.830 43.110 ;
        RECT 55.000 43.045 55.530 43.410 ;
        RECT 55.000 42.345 55.170 43.045 ;
        RECT 55.700 42.965 55.870 43.580 ;
        RECT 56.040 43.225 56.210 44.025 ;
        RECT 56.380 43.525 56.630 43.855 ;
        RECT 56.855 43.555 57.740 43.725 ;
        RECT 55.700 42.875 56.210 42.965 ;
        RECT 54.250 42.065 54.475 42.195 ;
        RECT 54.645 42.125 55.170 42.345 ;
        RECT 55.340 42.705 56.210 42.875 ;
        RECT 53.885 41.475 54.135 41.935 ;
        RECT 54.305 41.925 54.475 42.065 ;
        RECT 55.340 41.925 55.510 42.705 ;
        RECT 56.040 42.635 56.210 42.705 ;
        RECT 55.720 42.455 55.920 42.485 ;
        RECT 56.380 42.455 56.550 43.525 ;
        RECT 56.720 42.635 56.910 43.355 ;
        RECT 55.720 42.155 56.550 42.455 ;
        RECT 57.080 42.425 57.400 43.385 ;
        RECT 54.305 41.755 54.640 41.925 ;
        RECT 54.835 41.755 55.510 41.925 ;
        RECT 55.830 41.475 56.200 41.975 ;
        RECT 56.380 41.925 56.550 42.155 ;
        RECT 56.935 42.095 57.400 42.425 ;
        RECT 57.570 42.715 57.740 43.555 ;
        RECT 57.920 43.525 58.235 44.025 ;
        RECT 58.465 43.295 58.805 43.855 ;
        RECT 57.910 42.920 58.805 43.295 ;
        RECT 58.975 43.015 59.145 44.025 ;
        RECT 58.615 42.715 58.805 42.920 ;
        RECT 59.315 42.965 59.645 43.810 ;
        RECT 60.885 43.355 61.055 43.855 ;
        RECT 61.225 43.525 61.555 44.025 ;
        RECT 60.885 43.185 61.550 43.355 ;
        RECT 59.315 42.885 59.705 42.965 ;
        RECT 59.490 42.835 59.705 42.885 ;
        RECT 57.570 42.385 58.445 42.715 ;
        RECT 58.615 42.385 59.365 42.715 ;
        RECT 57.570 41.925 57.740 42.385 ;
        RECT 58.615 42.215 58.815 42.385 ;
        RECT 59.535 42.255 59.705 42.835 ;
        RECT 60.800 42.365 61.150 43.015 ;
        RECT 59.480 42.215 59.705 42.255 ;
        RECT 56.380 41.755 56.785 41.925 ;
        RECT 56.955 41.755 57.740 41.925 ;
        RECT 58.015 41.475 58.225 42.005 ;
        RECT 58.485 41.690 58.815 42.215 ;
        RECT 59.325 42.130 59.705 42.215 ;
        RECT 61.320 42.195 61.550 43.185 ;
        RECT 58.985 41.475 59.155 42.085 ;
        RECT 59.325 41.695 59.655 42.130 ;
        RECT 60.885 42.025 61.550 42.195 ;
        RECT 60.885 41.735 61.055 42.025 ;
        RECT 61.225 41.475 61.555 41.855 ;
        RECT 61.725 41.735 61.910 43.855 ;
        RECT 62.150 43.565 62.415 44.025 ;
        RECT 62.585 43.430 62.835 43.855 ;
        RECT 63.045 43.580 64.150 43.750 ;
        RECT 62.530 43.300 62.835 43.430 ;
        RECT 62.080 42.105 62.360 43.055 ;
        RECT 62.530 42.195 62.700 43.300 ;
        RECT 62.870 42.515 63.110 43.110 ;
        RECT 63.280 43.045 63.810 43.410 ;
        RECT 63.280 42.345 63.450 43.045 ;
        RECT 63.980 42.965 64.150 43.580 ;
        RECT 64.320 43.225 64.490 44.025 ;
        RECT 64.660 43.525 64.910 43.855 ;
        RECT 65.135 43.555 66.020 43.725 ;
        RECT 63.980 42.875 64.490 42.965 ;
        RECT 62.530 42.065 62.755 42.195 ;
        RECT 62.925 42.125 63.450 42.345 ;
        RECT 63.620 42.705 64.490 42.875 ;
        RECT 62.165 41.475 62.415 41.935 ;
        RECT 62.585 41.925 62.755 42.065 ;
        RECT 63.620 41.925 63.790 42.705 ;
        RECT 64.320 42.635 64.490 42.705 ;
        RECT 64.000 42.455 64.200 42.485 ;
        RECT 64.660 42.455 64.830 43.525 ;
        RECT 65.000 42.635 65.190 43.355 ;
        RECT 64.000 42.155 64.830 42.455 ;
        RECT 65.360 42.425 65.680 43.385 ;
        RECT 62.585 41.755 62.920 41.925 ;
        RECT 63.115 41.755 63.790 41.925 ;
        RECT 64.110 41.475 64.480 41.975 ;
        RECT 64.660 41.925 64.830 42.155 ;
        RECT 65.215 42.095 65.680 42.425 ;
        RECT 65.850 42.715 66.020 43.555 ;
        RECT 66.200 43.525 66.515 44.025 ;
        RECT 66.745 43.295 67.085 43.855 ;
        RECT 66.190 42.920 67.085 43.295 ;
        RECT 67.255 43.015 67.425 44.025 ;
        RECT 66.895 42.715 67.085 42.920 ;
        RECT 67.595 42.965 67.925 43.810 ;
        RECT 69.280 43.055 69.610 43.855 ;
        RECT 69.780 43.225 70.110 44.025 ;
        RECT 70.410 43.055 70.740 43.855 ;
        RECT 71.385 43.225 71.635 44.025 ;
        RECT 67.595 42.885 67.985 42.965 ;
        RECT 69.280 42.885 71.715 43.055 ;
        RECT 71.905 42.885 72.075 44.025 ;
        RECT 72.245 42.885 72.585 43.855 ;
        RECT 72.940 43.055 73.330 43.230 ;
        RECT 73.815 43.225 74.145 44.025 ;
        RECT 74.315 43.235 74.850 43.855 ;
        RECT 72.940 42.885 74.365 43.055 ;
        RECT 67.770 42.835 67.985 42.885 ;
        RECT 65.850 42.385 66.725 42.715 ;
        RECT 66.895 42.385 67.645 42.715 ;
        RECT 65.850 41.925 66.020 42.385 ;
        RECT 66.895 42.215 67.095 42.385 ;
        RECT 67.815 42.255 67.985 42.835 ;
        RECT 69.075 42.465 69.425 42.715 ;
        RECT 69.610 42.255 69.780 42.885 ;
        RECT 69.950 42.465 70.280 42.665 ;
        RECT 70.450 42.465 70.780 42.665 ;
        RECT 70.950 42.465 71.370 42.665 ;
        RECT 71.545 42.635 71.715 42.885 ;
        RECT 71.545 42.465 72.240 42.635 ;
        RECT 67.760 42.215 67.985 42.255 ;
        RECT 64.660 41.755 65.065 41.925 ;
        RECT 65.235 41.755 66.020 41.925 ;
        RECT 66.295 41.475 66.505 42.005 ;
        RECT 66.765 41.690 67.095 42.215 ;
        RECT 67.605 42.130 67.985 42.215 ;
        RECT 67.265 41.475 67.435 42.085 ;
        RECT 67.605 41.695 67.935 42.130 ;
        RECT 69.280 41.645 69.780 42.255 ;
        RECT 70.410 42.125 71.635 42.295 ;
        RECT 72.410 42.275 72.585 42.885 ;
        RECT 70.410 41.645 70.740 42.125 ;
        RECT 70.910 41.475 71.135 41.935 ;
        RECT 71.305 41.645 71.635 42.125 ;
        RECT 71.825 41.475 72.075 42.275 ;
        RECT 72.245 41.645 72.585 42.275 ;
        RECT 72.815 42.155 73.170 42.715 ;
        RECT 73.340 41.985 73.510 42.885 ;
        RECT 73.680 42.155 73.945 42.715 ;
        RECT 74.195 42.385 74.365 42.885 ;
        RECT 74.535 42.215 74.850 43.235 ;
        RECT 75.055 42.935 76.265 44.025 ;
        RECT 72.920 41.475 73.160 41.985 ;
        RECT 73.340 41.655 73.620 41.985 ;
        RECT 73.850 41.475 74.065 41.985 ;
        RECT 74.235 41.645 74.850 42.215 ;
        RECT 75.055 42.225 75.575 42.765 ;
        RECT 75.745 42.395 76.265 42.935 ;
        RECT 76.435 42.860 76.725 44.025 ;
        RECT 76.985 43.355 77.155 43.855 ;
        RECT 77.325 43.525 77.655 44.025 ;
        RECT 76.985 43.185 77.650 43.355 ;
        RECT 76.900 42.365 77.250 43.015 ;
        RECT 75.055 41.475 76.265 42.225 ;
        RECT 76.435 41.475 76.725 42.200 ;
        RECT 77.420 42.195 77.650 43.185 ;
        RECT 76.985 42.025 77.650 42.195 ;
        RECT 76.985 41.735 77.155 42.025 ;
        RECT 77.325 41.475 77.655 41.855 ;
        RECT 77.825 41.735 78.010 43.855 ;
        RECT 78.250 43.565 78.515 44.025 ;
        RECT 78.685 43.430 78.935 43.855 ;
        RECT 79.145 43.580 80.250 43.750 ;
        RECT 78.630 43.300 78.935 43.430 ;
        RECT 78.180 42.105 78.460 43.055 ;
        RECT 78.630 42.195 78.800 43.300 ;
        RECT 78.970 42.515 79.210 43.110 ;
        RECT 79.380 43.045 79.910 43.410 ;
        RECT 79.380 42.345 79.550 43.045 ;
        RECT 80.080 42.965 80.250 43.580 ;
        RECT 80.420 43.225 80.590 44.025 ;
        RECT 80.760 43.525 81.010 43.855 ;
        RECT 81.235 43.555 82.120 43.725 ;
        RECT 80.080 42.875 80.590 42.965 ;
        RECT 78.630 42.065 78.855 42.195 ;
        RECT 79.025 42.125 79.550 42.345 ;
        RECT 79.720 42.705 80.590 42.875 ;
        RECT 78.265 41.475 78.515 41.935 ;
        RECT 78.685 41.925 78.855 42.065 ;
        RECT 79.720 41.925 79.890 42.705 ;
        RECT 80.420 42.635 80.590 42.705 ;
        RECT 80.100 42.455 80.300 42.485 ;
        RECT 80.760 42.455 80.930 43.525 ;
        RECT 81.100 42.635 81.290 43.355 ;
        RECT 80.100 42.155 80.930 42.455 ;
        RECT 81.460 42.425 81.780 43.385 ;
        RECT 78.685 41.755 79.020 41.925 ;
        RECT 79.215 41.755 79.890 41.925 ;
        RECT 80.210 41.475 80.580 41.975 ;
        RECT 80.760 41.925 80.930 42.155 ;
        RECT 81.315 42.095 81.780 42.425 ;
        RECT 81.950 42.715 82.120 43.555 ;
        RECT 82.300 43.525 82.615 44.025 ;
        RECT 82.845 43.295 83.185 43.855 ;
        RECT 82.290 42.920 83.185 43.295 ;
        RECT 83.355 43.015 83.525 44.025 ;
        RECT 82.995 42.715 83.185 42.920 ;
        RECT 83.695 42.965 84.025 43.810 ;
        RECT 83.695 42.885 84.085 42.965 ;
        RECT 84.255 42.935 87.765 44.025 ;
        RECT 87.935 42.935 89.145 44.025 ;
        RECT 83.870 42.835 84.085 42.885 ;
        RECT 81.950 42.385 82.825 42.715 ;
        RECT 82.995 42.385 83.745 42.715 ;
        RECT 81.950 41.925 82.120 42.385 ;
        RECT 82.995 42.215 83.195 42.385 ;
        RECT 83.915 42.255 84.085 42.835 ;
        RECT 83.860 42.215 84.085 42.255 ;
        RECT 80.760 41.755 81.165 41.925 ;
        RECT 81.335 41.755 82.120 41.925 ;
        RECT 82.395 41.475 82.605 42.005 ;
        RECT 82.865 41.690 83.195 42.215 ;
        RECT 83.705 42.130 84.085 42.215 ;
        RECT 84.255 42.245 85.905 42.765 ;
        RECT 86.075 42.415 87.765 42.935 ;
        RECT 83.365 41.475 83.535 42.085 ;
        RECT 83.705 41.695 84.035 42.130 ;
        RECT 84.255 41.475 87.765 42.245 ;
        RECT 87.935 42.225 88.455 42.765 ;
        RECT 88.625 42.395 89.145 42.935 ;
        RECT 89.315 42.935 90.525 44.025 ;
        RECT 89.315 42.395 89.835 42.935 ;
        RECT 90.005 42.225 90.525 42.765 ;
        RECT 87.935 41.475 89.145 42.225 ;
        RECT 89.315 41.475 90.525 42.225 ;
        RECT 11.950 41.305 90.610 41.475 ;
        RECT 12.035 40.555 13.245 41.305 ;
        RECT 12.035 40.015 12.555 40.555 ;
        RECT 14.335 40.505 14.675 41.135 ;
        RECT 14.845 40.505 15.095 41.305 ;
        RECT 15.285 40.655 15.615 41.135 ;
        RECT 15.785 40.845 16.010 41.305 ;
        RECT 16.180 40.655 16.510 41.135 ;
        RECT 12.725 39.845 13.245 40.385 ;
        RECT 12.035 38.755 13.245 39.845 ;
        RECT 14.335 39.895 14.510 40.505 ;
        RECT 15.285 40.485 16.510 40.655 ;
        RECT 17.140 40.525 17.640 41.135 ;
        RECT 18.050 40.565 18.665 41.135 ;
        RECT 18.835 40.795 19.050 41.305 ;
        RECT 19.280 40.795 19.560 41.125 ;
        RECT 19.740 40.795 19.980 41.305 ;
        RECT 14.680 40.145 15.375 40.315 ;
        RECT 15.205 39.895 15.375 40.145 ;
        RECT 15.550 40.115 15.970 40.315 ;
        RECT 16.140 40.115 16.470 40.315 ;
        RECT 16.640 40.115 16.970 40.315 ;
        RECT 17.140 39.895 17.310 40.525 ;
        RECT 17.495 40.065 17.845 40.315 ;
        RECT 14.335 38.925 14.675 39.895 ;
        RECT 14.845 38.755 15.015 39.895 ;
        RECT 15.205 39.725 17.640 39.895 ;
        RECT 15.285 38.755 15.535 39.555 ;
        RECT 16.180 38.925 16.510 39.725 ;
        RECT 16.810 38.755 17.140 39.555 ;
        RECT 17.310 38.925 17.640 39.725 ;
        RECT 18.050 39.545 18.365 40.565 ;
        RECT 18.535 39.895 18.705 40.395 ;
        RECT 18.955 40.065 19.220 40.625 ;
        RECT 19.390 39.895 19.560 40.795 ;
        RECT 19.730 40.065 20.085 40.625 ;
        RECT 20.320 40.540 20.775 41.305 ;
        RECT 21.050 40.925 22.350 41.135 ;
        RECT 22.605 40.945 22.935 41.305 ;
        RECT 22.180 40.775 22.350 40.925 ;
        RECT 23.105 40.805 23.365 41.135 ;
        RECT 23.135 40.795 23.365 40.805 ;
        RECT 21.250 40.315 21.470 40.715 ;
        RECT 20.315 40.115 20.805 40.315 ;
        RECT 20.995 40.105 21.470 40.315 ;
        RECT 21.715 40.315 21.925 40.715 ;
        RECT 22.180 40.650 22.935 40.775 ;
        RECT 22.180 40.605 23.025 40.650 ;
        RECT 22.755 40.485 23.025 40.605 ;
        RECT 21.715 40.105 22.045 40.315 ;
        RECT 22.215 40.045 22.625 40.350 ;
        RECT 18.535 39.725 19.960 39.895 ;
        RECT 18.050 38.925 18.585 39.545 ;
        RECT 18.755 38.755 19.085 39.555 ;
        RECT 19.570 39.550 19.960 39.725 ;
        RECT 20.320 39.875 21.495 39.935 ;
        RECT 22.855 39.910 23.025 40.485 ;
        RECT 22.825 39.875 23.025 39.910 ;
        RECT 20.320 39.765 23.025 39.875 ;
        RECT 20.320 39.145 20.575 39.765 ;
        RECT 21.165 39.705 22.965 39.765 ;
        RECT 21.165 39.675 21.495 39.705 ;
        RECT 23.195 39.605 23.365 40.795 ;
        RECT 23.535 40.535 27.045 41.305 ;
        RECT 23.535 40.015 25.185 40.535 ;
        RECT 27.695 40.495 27.935 41.305 ;
        RECT 28.105 40.495 28.435 41.135 ;
        RECT 28.605 40.495 28.875 41.305 ;
        RECT 29.055 40.555 30.265 41.305 ;
        RECT 30.435 40.845 30.995 41.135 ;
        RECT 31.165 40.845 31.415 41.305 ;
        RECT 25.355 39.845 27.045 40.365 ;
        RECT 27.675 40.065 28.025 40.315 ;
        RECT 28.195 39.895 28.365 40.495 ;
        RECT 28.535 40.065 28.885 40.315 ;
        RECT 29.055 40.015 29.575 40.555 ;
        RECT 20.825 39.505 21.010 39.595 ;
        RECT 21.600 39.505 22.435 39.515 ;
        RECT 20.825 39.305 22.435 39.505 ;
        RECT 20.825 39.265 21.055 39.305 ;
        RECT 20.320 38.925 20.655 39.145 ;
        RECT 21.660 38.755 22.015 39.135 ;
        RECT 22.185 38.925 22.435 39.305 ;
        RECT 22.685 38.755 22.935 39.535 ;
        RECT 23.105 38.925 23.365 39.605 ;
        RECT 23.535 38.755 27.045 39.845 ;
        RECT 27.685 39.725 28.365 39.895 ;
        RECT 27.685 38.940 28.015 39.725 ;
        RECT 28.545 38.755 28.875 39.895 ;
        RECT 29.745 39.845 30.265 40.385 ;
        RECT 29.055 38.755 30.265 39.845 ;
        RECT 30.435 39.475 30.685 40.845 ;
        RECT 32.035 40.675 32.365 41.035 ;
        RECT 30.975 40.485 32.365 40.675 ;
        RECT 32.735 40.535 36.245 41.305 ;
        RECT 36.415 40.555 37.625 41.305 ;
        RECT 37.795 40.580 38.085 41.305 ;
        RECT 30.975 40.395 31.145 40.485 ;
        RECT 30.855 40.065 31.145 40.395 ;
        RECT 31.315 40.065 31.655 40.315 ;
        RECT 31.875 40.065 32.550 40.315 ;
        RECT 30.975 39.815 31.145 40.065 ;
        RECT 30.975 39.645 31.915 39.815 ;
        RECT 32.285 39.705 32.550 40.065 ;
        RECT 32.735 40.015 34.385 40.535 ;
        RECT 34.555 39.845 36.245 40.365 ;
        RECT 36.415 40.015 36.935 40.555 ;
        RECT 38.255 40.535 39.925 41.305 ;
        RECT 37.105 39.845 37.625 40.385 ;
        RECT 38.255 40.015 39.005 40.535 ;
        RECT 30.435 38.925 30.895 39.475 ;
        RECT 31.085 38.755 31.415 39.475 ;
        RECT 31.615 39.095 31.915 39.645 ;
        RECT 32.085 38.755 32.365 39.425 ;
        RECT 32.735 38.755 36.245 39.845 ;
        RECT 36.415 38.755 37.625 39.845 ;
        RECT 37.795 38.755 38.085 39.920 ;
        RECT 39.175 39.845 39.925 40.365 ;
        RECT 38.255 38.755 39.925 39.845 ;
        RECT 40.100 39.705 40.435 41.125 ;
        RECT 40.615 40.935 41.360 41.305 ;
        RECT 41.925 40.765 42.180 41.125 ;
        RECT 42.360 40.935 42.690 41.305 ;
        RECT 42.870 40.765 43.095 41.125 ;
        RECT 40.610 40.575 43.095 40.765 ;
        RECT 40.610 39.885 40.835 40.575 ;
        RECT 43.315 40.535 45.905 41.305 ;
        RECT 46.540 40.565 46.795 41.135 ;
        RECT 46.965 40.905 47.295 41.305 ;
        RECT 47.720 40.770 48.250 41.135 ;
        RECT 48.440 40.965 48.715 41.135 ;
        RECT 48.435 40.795 48.715 40.965 ;
        RECT 47.720 40.735 47.895 40.770 ;
        RECT 46.965 40.565 47.895 40.735 ;
        RECT 41.035 40.065 41.315 40.395 ;
        RECT 41.495 40.065 42.070 40.395 ;
        RECT 42.250 40.065 42.685 40.395 ;
        RECT 42.865 40.065 43.135 40.395 ;
        RECT 43.315 40.015 44.525 40.535 ;
        RECT 40.610 39.705 43.105 39.885 ;
        RECT 44.695 39.845 45.905 40.365 ;
        RECT 40.100 38.935 40.365 39.705 ;
        RECT 40.535 38.755 40.865 39.475 ;
        RECT 41.055 39.295 42.245 39.525 ;
        RECT 41.055 38.935 41.315 39.295 ;
        RECT 41.485 38.755 41.815 39.125 ;
        RECT 41.985 38.935 42.245 39.295 ;
        RECT 42.815 38.935 43.105 39.705 ;
        RECT 43.315 38.755 45.905 39.845 ;
        RECT 46.540 39.895 46.710 40.565 ;
        RECT 46.965 40.395 47.135 40.565 ;
        RECT 46.880 40.065 47.135 40.395 ;
        RECT 47.360 40.065 47.555 40.395 ;
        RECT 46.540 38.925 46.875 39.895 ;
        RECT 47.045 38.755 47.215 39.895 ;
        RECT 47.385 39.095 47.555 40.065 ;
        RECT 47.725 39.435 47.895 40.565 ;
        RECT 48.065 39.775 48.235 40.575 ;
        RECT 48.440 39.975 48.715 40.795 ;
        RECT 48.885 39.775 49.075 41.135 ;
        RECT 49.255 40.770 49.765 41.305 ;
        RECT 49.985 40.495 50.230 41.100 ;
        RECT 50.675 40.645 50.950 41.305 ;
        RECT 51.120 40.675 51.370 41.135 ;
        RECT 51.545 40.810 51.875 41.305 ;
        RECT 49.275 40.325 50.505 40.495 ;
        RECT 51.120 40.465 51.290 40.675 ;
        RECT 52.055 40.640 52.285 41.085 ;
        RECT 48.065 39.605 49.075 39.775 ;
        RECT 49.245 39.760 49.995 39.950 ;
        RECT 47.725 39.265 48.850 39.435 ;
        RECT 49.245 39.095 49.415 39.760 ;
        RECT 50.165 39.515 50.505 40.325 ;
        RECT 50.675 39.945 51.290 40.465 ;
        RECT 51.460 39.965 51.690 40.395 ;
        RECT 51.875 40.145 52.285 40.640 ;
        RECT 52.455 40.820 53.245 41.085 ;
        RECT 52.455 39.965 52.710 40.820 ;
        RECT 52.880 40.145 53.265 40.625 ;
        RECT 53.955 40.485 54.165 41.305 ;
        RECT 54.335 40.505 54.665 41.135 ;
        RECT 47.385 38.925 49.415 39.095 ;
        RECT 49.585 38.755 49.755 39.515 ;
        RECT 49.990 39.105 50.505 39.515 ;
        RECT 50.675 38.755 50.935 39.765 ;
        RECT 51.105 39.595 51.275 39.945 ;
        RECT 51.460 39.795 53.250 39.965 ;
        RECT 54.335 39.905 54.585 40.505 ;
        RECT 54.835 40.485 55.065 41.305 ;
        RECT 55.520 40.825 55.820 41.305 ;
        RECT 55.990 40.655 56.250 41.110 ;
        RECT 56.420 40.825 56.680 41.305 ;
        RECT 56.850 40.655 57.110 41.110 ;
        RECT 57.280 40.825 57.540 41.305 ;
        RECT 57.710 40.655 57.970 41.110 ;
        RECT 58.140 40.825 58.400 41.305 ;
        RECT 58.570 40.655 58.830 41.110 ;
        RECT 59.000 40.780 59.260 41.305 ;
        RECT 55.520 40.485 58.830 40.655 ;
        RECT 54.755 40.065 55.085 40.315 ;
        RECT 51.105 38.925 51.380 39.595 ;
        RECT 51.580 38.755 51.795 39.600 ;
        RECT 52.020 39.500 52.270 39.795 ;
        RECT 52.495 39.435 52.825 39.625 ;
        RECT 51.980 38.925 52.455 39.265 ;
        RECT 52.635 39.260 52.825 39.435 ;
        RECT 52.995 39.430 53.250 39.795 ;
        RECT 52.635 38.755 53.265 39.260 ;
        RECT 53.955 38.755 54.165 39.895 ;
        RECT 54.335 38.925 54.665 39.905 ;
        RECT 55.520 39.895 56.490 40.485 ;
        RECT 59.430 40.315 59.680 41.125 ;
        RECT 59.860 40.845 60.105 41.305 ;
        RECT 60.535 40.675 60.865 41.035 ;
        RECT 61.495 40.845 61.745 41.305 ;
        RECT 61.915 40.845 62.465 41.135 ;
        RECT 56.660 40.065 59.680 40.315 ;
        RECT 59.850 40.065 60.165 40.675 ;
        RECT 60.535 40.485 61.925 40.675 ;
        RECT 61.755 40.395 61.925 40.485 ;
        RECT 60.335 40.065 61.025 40.315 ;
        RECT 61.255 40.065 61.585 40.315 ;
        RECT 61.755 40.065 62.045 40.395 ;
        RECT 54.835 38.755 55.065 39.895 ;
        RECT 55.520 39.655 58.830 39.895 ;
        RECT 55.525 38.755 55.820 39.485 ;
        RECT 55.990 38.930 56.250 39.655 ;
        RECT 56.420 38.755 56.680 39.485 ;
        RECT 56.850 38.930 57.110 39.655 ;
        RECT 57.280 38.755 57.540 39.485 ;
        RECT 57.710 38.930 57.970 39.655 ;
        RECT 58.140 38.755 58.400 39.485 ;
        RECT 58.570 38.930 58.830 39.655 ;
        RECT 59.000 38.755 59.260 39.865 ;
        RECT 59.430 38.930 59.680 40.065 ;
        RECT 59.860 38.755 60.155 39.865 ;
        RECT 60.335 39.625 60.650 40.065 ;
        RECT 61.755 39.815 61.925 40.065 ;
        RECT 60.985 39.645 61.925 39.815 ;
        RECT 60.535 38.755 60.815 39.425 ;
        RECT 60.985 39.095 61.285 39.645 ;
        RECT 62.215 39.475 62.465 40.845 ;
        RECT 62.635 40.505 62.925 41.305 ;
        RECT 63.555 40.580 63.845 41.305 ;
        RECT 64.015 40.505 64.355 41.135 ;
        RECT 64.525 40.505 64.775 41.305 ;
        RECT 64.965 40.655 65.295 41.135 ;
        RECT 65.465 40.845 65.690 41.305 ;
        RECT 65.860 40.655 66.190 41.135 ;
        RECT 61.495 38.755 61.825 39.475 ;
        RECT 62.015 38.925 62.465 39.475 ;
        RECT 62.635 38.755 62.925 39.895 ;
        RECT 63.555 38.755 63.845 39.920 ;
        RECT 64.015 39.895 64.190 40.505 ;
        RECT 64.965 40.485 66.190 40.655 ;
        RECT 66.820 40.525 67.320 41.135 ;
        RECT 68.320 40.795 68.560 41.305 ;
        RECT 68.740 40.795 69.020 41.125 ;
        RECT 69.250 40.795 69.465 41.305 ;
        RECT 64.360 40.145 65.055 40.315 ;
        RECT 64.885 39.895 65.055 40.145 ;
        RECT 65.230 40.115 65.650 40.315 ;
        RECT 65.820 40.115 66.150 40.315 ;
        RECT 66.320 40.115 66.650 40.315 ;
        RECT 66.820 39.895 66.990 40.525 ;
        RECT 67.175 40.065 67.525 40.315 ;
        RECT 68.215 40.065 68.570 40.625 ;
        RECT 68.740 39.895 68.910 40.795 ;
        RECT 69.080 40.065 69.345 40.625 ;
        RECT 69.635 40.565 70.250 41.135 ;
        RECT 69.595 39.895 69.765 40.395 ;
        RECT 64.015 38.925 64.355 39.895 ;
        RECT 64.525 38.755 64.695 39.895 ;
        RECT 64.885 39.725 67.320 39.895 ;
        RECT 64.965 38.755 65.215 39.555 ;
        RECT 65.860 38.925 66.190 39.725 ;
        RECT 66.490 38.755 66.820 39.555 ;
        RECT 66.990 38.925 67.320 39.725 ;
        RECT 68.340 39.725 69.765 39.895 ;
        RECT 68.340 39.550 68.730 39.725 ;
        RECT 69.215 38.755 69.545 39.555 ;
        RECT 69.935 39.545 70.250 40.565 ;
        RECT 70.455 40.675 70.795 41.135 ;
        RECT 70.965 40.845 71.135 41.305 ;
        RECT 71.305 40.925 72.475 41.135 ;
        RECT 71.305 40.675 71.555 40.925 ;
        RECT 72.145 40.905 72.475 40.925 ;
        RECT 70.455 40.505 71.555 40.675 ;
        RECT 71.725 40.485 72.585 40.735 ;
        RECT 72.955 40.675 73.285 41.035 ;
        RECT 73.905 40.845 74.155 41.305 ;
        RECT 74.325 40.845 74.885 41.135 ;
        RECT 72.955 40.485 74.345 40.675 ;
        RECT 70.455 40.065 71.215 40.315 ;
        RECT 71.385 40.065 72.135 40.315 ;
        RECT 72.305 39.895 72.585 40.485 ;
        RECT 74.175 40.395 74.345 40.485 ;
        RECT 69.715 38.925 70.250 39.545 ;
        RECT 70.455 38.755 70.715 39.895 ;
        RECT 70.885 39.725 72.585 39.895 ;
        RECT 72.770 40.065 73.445 40.315 ;
        RECT 73.665 40.065 74.005 40.315 ;
        RECT 74.175 40.065 74.465 40.395 ;
        RECT 70.885 38.925 71.215 39.725 ;
        RECT 71.385 38.755 71.555 39.555 ;
        RECT 71.725 38.925 72.055 39.725 ;
        RECT 72.770 39.705 73.035 40.065 ;
        RECT 74.175 39.815 74.345 40.065 ;
        RECT 73.405 39.645 74.345 39.815 ;
        RECT 72.225 38.755 72.480 39.555 ;
        RECT 72.955 38.755 73.235 39.425 ;
        RECT 73.405 39.095 73.705 39.645 ;
        RECT 74.635 39.475 74.885 40.845 ;
        RECT 75.055 40.535 78.565 41.305 ;
        RECT 75.055 40.015 76.705 40.535 ;
        RECT 78.940 40.525 79.440 41.135 ;
        RECT 76.875 39.845 78.565 40.365 ;
        RECT 78.735 40.065 79.085 40.315 ;
        RECT 79.270 39.895 79.440 40.525 ;
        RECT 80.070 40.655 80.400 41.135 ;
        RECT 80.570 40.845 80.795 41.305 ;
        RECT 80.965 40.655 81.295 41.135 ;
        RECT 80.070 40.485 81.295 40.655 ;
        RECT 81.485 40.505 81.735 41.305 ;
        RECT 81.905 40.505 82.245 41.135 ;
        RECT 79.610 40.115 79.940 40.315 ;
        RECT 80.110 40.115 80.440 40.315 ;
        RECT 80.610 40.115 81.030 40.315 ;
        RECT 81.205 40.145 81.900 40.315 ;
        RECT 81.205 39.895 81.375 40.145 ;
        RECT 82.070 39.895 82.245 40.505 ;
        RECT 73.905 38.755 74.235 39.475 ;
        RECT 74.425 38.925 74.885 39.475 ;
        RECT 75.055 38.755 78.565 39.845 ;
        RECT 78.940 39.725 81.375 39.895 ;
        RECT 78.940 38.925 79.270 39.725 ;
        RECT 79.440 38.755 79.770 39.555 ;
        RECT 80.070 38.925 80.400 39.725 ;
        RECT 81.045 38.755 81.295 39.555 ;
        RECT 81.565 38.755 81.735 39.895 ;
        RECT 81.905 38.925 82.245 39.895 ;
        RECT 82.415 40.630 82.675 41.135 ;
        RECT 82.855 40.925 83.185 41.305 ;
        RECT 83.365 40.755 83.535 41.135 ;
        RECT 83.795 40.760 89.140 41.305 ;
        RECT 82.415 39.830 82.595 40.630 ;
        RECT 82.870 40.585 83.535 40.755 ;
        RECT 82.870 40.330 83.040 40.585 ;
        RECT 82.765 40.000 83.040 40.330 ;
        RECT 83.265 40.035 83.605 40.405 ;
        RECT 82.870 39.855 83.040 40.000 ;
        RECT 85.380 39.930 85.720 40.760 ;
        RECT 89.315 40.555 90.525 41.305 ;
        RECT 82.415 38.925 82.685 39.830 ;
        RECT 82.870 39.685 83.545 39.855 ;
        RECT 82.855 38.755 83.185 39.515 ;
        RECT 83.365 38.925 83.545 39.685 ;
        RECT 87.200 39.190 87.550 40.440 ;
        RECT 89.315 39.845 89.835 40.385 ;
        RECT 90.005 40.015 90.525 40.555 ;
        RECT 83.795 38.755 89.140 39.190 ;
        RECT 89.315 38.755 90.525 39.845 ;
        RECT 11.950 38.585 90.610 38.755 ;
        RECT 12.035 37.495 13.245 38.585 ;
        RECT 13.415 37.495 16.005 38.585 ;
        RECT 16.725 37.915 16.895 38.415 ;
        RECT 17.065 38.085 17.395 38.585 ;
        RECT 16.725 37.745 17.390 37.915 ;
        RECT 12.035 36.785 12.555 37.325 ;
        RECT 12.725 36.955 13.245 37.495 ;
        RECT 13.415 36.805 14.625 37.325 ;
        RECT 14.795 36.975 16.005 37.495 ;
        RECT 16.640 36.925 16.990 37.575 ;
        RECT 12.035 36.035 13.245 36.785 ;
        RECT 13.415 36.035 16.005 36.805 ;
        RECT 17.160 36.755 17.390 37.745 ;
        RECT 16.725 36.585 17.390 36.755 ;
        RECT 16.725 36.295 16.895 36.585 ;
        RECT 17.065 36.035 17.395 36.415 ;
        RECT 17.565 36.295 17.750 38.415 ;
        RECT 17.990 38.125 18.255 38.585 ;
        RECT 18.425 37.990 18.675 38.415 ;
        RECT 18.885 38.140 19.990 38.310 ;
        RECT 18.370 37.860 18.675 37.990 ;
        RECT 17.920 36.665 18.200 37.615 ;
        RECT 18.370 36.755 18.540 37.860 ;
        RECT 18.710 37.075 18.950 37.670 ;
        RECT 19.120 37.605 19.650 37.970 ;
        RECT 19.120 36.905 19.290 37.605 ;
        RECT 19.820 37.525 19.990 38.140 ;
        RECT 20.160 37.785 20.330 38.585 ;
        RECT 20.500 38.085 20.750 38.415 ;
        RECT 20.975 38.115 21.860 38.285 ;
        RECT 19.820 37.435 20.330 37.525 ;
        RECT 18.370 36.625 18.595 36.755 ;
        RECT 18.765 36.685 19.290 36.905 ;
        RECT 19.460 37.265 20.330 37.435 ;
        RECT 18.005 36.035 18.255 36.495 ;
        RECT 18.425 36.485 18.595 36.625 ;
        RECT 19.460 36.485 19.630 37.265 ;
        RECT 20.160 37.195 20.330 37.265 ;
        RECT 19.840 37.015 20.040 37.045 ;
        RECT 20.500 37.015 20.670 38.085 ;
        RECT 20.840 37.195 21.030 37.915 ;
        RECT 19.840 36.715 20.670 37.015 ;
        RECT 21.200 36.985 21.520 37.945 ;
        RECT 18.425 36.315 18.760 36.485 ;
        RECT 18.955 36.315 19.630 36.485 ;
        RECT 19.950 36.035 20.320 36.535 ;
        RECT 20.500 36.485 20.670 36.715 ;
        RECT 21.055 36.655 21.520 36.985 ;
        RECT 21.690 37.275 21.860 38.115 ;
        RECT 22.040 38.085 22.355 38.585 ;
        RECT 22.585 37.855 22.925 38.415 ;
        RECT 22.030 37.480 22.925 37.855 ;
        RECT 23.095 37.575 23.265 38.585 ;
        RECT 22.735 37.275 22.925 37.480 ;
        RECT 23.435 37.525 23.765 38.370 ;
        RECT 23.435 37.445 23.825 37.525 ;
        RECT 23.610 37.395 23.825 37.445 ;
        RECT 24.915 37.420 25.205 38.585 ;
        RECT 25.410 37.795 25.945 38.415 ;
        RECT 21.690 36.945 22.565 37.275 ;
        RECT 22.735 36.945 23.485 37.275 ;
        RECT 21.690 36.485 21.860 36.945 ;
        RECT 22.735 36.775 22.935 36.945 ;
        RECT 23.655 36.815 23.825 37.395 ;
        RECT 23.600 36.775 23.825 36.815 ;
        RECT 20.500 36.315 20.905 36.485 ;
        RECT 21.075 36.315 21.860 36.485 ;
        RECT 22.135 36.035 22.345 36.565 ;
        RECT 22.605 36.250 22.935 36.775 ;
        RECT 23.445 36.690 23.825 36.775 ;
        RECT 25.410 36.775 25.725 37.795 ;
        RECT 26.115 37.785 26.445 38.585 ;
        RECT 26.930 37.615 27.320 37.790 ;
        RECT 25.895 37.445 27.320 37.615 ;
        RECT 28.800 37.615 29.130 38.415 ;
        RECT 29.300 37.785 29.630 38.585 ;
        RECT 29.930 37.615 30.260 38.415 ;
        RECT 30.905 37.785 31.155 38.585 ;
        RECT 28.800 37.445 31.235 37.615 ;
        RECT 31.425 37.445 31.595 38.585 ;
        RECT 31.765 37.445 32.105 38.415 ;
        RECT 32.380 37.785 32.635 38.585 ;
        RECT 32.805 37.615 33.135 38.415 ;
        RECT 33.305 37.785 33.475 38.585 ;
        RECT 33.645 37.615 33.975 38.415 ;
        RECT 25.895 36.945 26.065 37.445 ;
        RECT 23.105 36.035 23.275 36.645 ;
        RECT 23.445 36.255 23.775 36.690 ;
        RECT 24.915 36.035 25.205 36.760 ;
        RECT 25.410 36.205 26.025 36.775 ;
        RECT 26.315 36.715 26.580 37.275 ;
        RECT 26.750 36.545 26.920 37.445 ;
        RECT 27.090 36.715 27.445 37.275 ;
        RECT 28.595 37.025 28.945 37.275 ;
        RECT 29.130 36.815 29.300 37.445 ;
        RECT 29.470 37.025 29.800 37.225 ;
        RECT 29.970 37.025 30.300 37.225 ;
        RECT 30.470 37.025 30.890 37.225 ;
        RECT 31.065 37.195 31.235 37.445 ;
        RECT 31.065 37.025 31.760 37.195 ;
        RECT 26.195 36.035 26.410 36.545 ;
        RECT 26.640 36.215 26.920 36.545 ;
        RECT 27.100 36.035 27.340 36.545 ;
        RECT 28.800 36.205 29.300 36.815 ;
        RECT 29.930 36.685 31.155 36.855 ;
        RECT 31.930 36.835 32.105 37.445 ;
        RECT 29.930 36.205 30.260 36.685 ;
        RECT 30.430 36.035 30.655 36.495 ;
        RECT 30.825 36.205 31.155 36.685 ;
        RECT 31.345 36.035 31.595 36.835 ;
        RECT 31.765 36.205 32.105 36.835 ;
        RECT 32.275 37.445 33.975 37.615 ;
        RECT 34.145 37.445 34.405 38.585 ;
        RECT 34.575 37.495 36.245 38.585 ;
        RECT 36.475 37.525 36.805 38.370 ;
        RECT 36.975 37.575 37.145 38.585 ;
        RECT 37.315 37.855 37.655 38.415 ;
        RECT 37.885 38.085 38.200 38.585 ;
        RECT 38.380 38.115 39.265 38.285 ;
        RECT 32.275 36.855 32.555 37.445 ;
        RECT 32.725 37.025 33.475 37.275 ;
        RECT 33.645 37.025 34.405 37.275 ;
        RECT 32.275 36.605 33.135 36.855 ;
        RECT 33.305 36.665 34.405 36.835 ;
        RECT 32.385 36.415 32.715 36.435 ;
        RECT 33.305 36.415 33.555 36.665 ;
        RECT 32.385 36.205 33.555 36.415 ;
        RECT 33.725 36.035 33.895 36.495 ;
        RECT 34.065 36.205 34.405 36.665 ;
        RECT 34.575 36.805 35.325 37.325 ;
        RECT 35.495 36.975 36.245 37.495 ;
        RECT 36.415 37.445 36.805 37.525 ;
        RECT 37.315 37.480 38.210 37.855 ;
        RECT 36.415 37.395 36.630 37.445 ;
        RECT 36.415 36.815 36.585 37.395 ;
        RECT 37.315 37.275 37.505 37.480 ;
        RECT 38.380 37.275 38.550 38.115 ;
        RECT 39.490 38.085 39.740 38.415 ;
        RECT 36.755 36.945 37.505 37.275 ;
        RECT 37.675 36.945 38.550 37.275 ;
        RECT 34.575 36.035 36.245 36.805 ;
        RECT 36.415 36.775 36.640 36.815 ;
        RECT 37.305 36.775 37.505 36.945 ;
        RECT 36.415 36.690 36.795 36.775 ;
        RECT 36.465 36.255 36.795 36.690 ;
        RECT 36.965 36.035 37.135 36.645 ;
        RECT 37.305 36.250 37.635 36.775 ;
        RECT 37.895 36.035 38.105 36.565 ;
        RECT 38.380 36.485 38.550 36.945 ;
        RECT 38.720 36.985 39.040 37.945 ;
        RECT 39.210 37.195 39.400 37.915 ;
        RECT 39.570 37.015 39.740 38.085 ;
        RECT 39.910 37.785 40.080 38.585 ;
        RECT 40.250 38.140 41.355 38.310 ;
        RECT 40.250 37.525 40.420 38.140 ;
        RECT 41.565 37.990 41.815 38.415 ;
        RECT 41.985 38.125 42.250 38.585 ;
        RECT 40.590 37.605 41.120 37.970 ;
        RECT 41.565 37.860 41.870 37.990 ;
        RECT 39.910 37.435 40.420 37.525 ;
        RECT 39.910 37.265 40.780 37.435 ;
        RECT 39.910 37.195 40.080 37.265 ;
        RECT 40.200 37.015 40.400 37.045 ;
        RECT 38.720 36.655 39.185 36.985 ;
        RECT 39.570 36.715 40.400 37.015 ;
        RECT 39.570 36.485 39.740 36.715 ;
        RECT 38.380 36.315 39.165 36.485 ;
        RECT 39.335 36.315 39.740 36.485 ;
        RECT 39.920 36.035 40.290 36.535 ;
        RECT 40.610 36.485 40.780 37.265 ;
        RECT 40.950 36.905 41.120 37.605 ;
        RECT 41.290 37.075 41.530 37.670 ;
        RECT 40.950 36.685 41.475 36.905 ;
        RECT 41.700 36.755 41.870 37.860 ;
        RECT 41.645 36.625 41.870 36.755 ;
        RECT 42.040 36.665 42.320 37.615 ;
        RECT 41.645 36.485 41.815 36.625 ;
        RECT 40.610 36.315 41.285 36.485 ;
        RECT 41.480 36.315 41.815 36.485 ;
        RECT 41.985 36.035 42.235 36.495 ;
        RECT 42.490 36.295 42.675 38.415 ;
        RECT 42.845 38.085 43.175 38.585 ;
        RECT 43.345 37.915 43.515 38.415 ;
        RECT 42.850 37.745 43.515 37.915 ;
        RECT 42.850 36.755 43.080 37.745 ;
        RECT 43.250 36.925 43.600 37.575 ;
        RECT 43.775 37.445 44.115 38.415 ;
        RECT 44.285 37.445 44.455 38.585 ;
        RECT 44.725 37.785 44.975 38.585 ;
        RECT 45.620 37.615 45.950 38.415 ;
        RECT 46.250 37.785 46.580 38.585 ;
        RECT 46.750 37.615 47.080 38.415 ;
        RECT 44.645 37.445 47.080 37.615 ;
        RECT 47.455 37.495 50.045 38.585 ;
        RECT 43.775 36.885 43.950 37.445 ;
        RECT 44.645 37.195 44.815 37.445 ;
        RECT 44.120 37.025 44.815 37.195 ;
        RECT 44.990 37.025 45.410 37.225 ;
        RECT 45.580 37.025 45.910 37.225 ;
        RECT 46.080 37.025 46.410 37.225 ;
        RECT 43.775 36.835 44.005 36.885 ;
        RECT 42.850 36.585 43.515 36.755 ;
        RECT 42.845 36.035 43.175 36.415 ;
        RECT 43.345 36.295 43.515 36.585 ;
        RECT 43.775 36.205 44.115 36.835 ;
        RECT 44.285 36.035 44.535 36.835 ;
        RECT 44.725 36.685 45.950 36.855 ;
        RECT 44.725 36.205 45.055 36.685 ;
        RECT 45.225 36.035 45.450 36.495 ;
        RECT 45.620 36.205 45.950 36.685 ;
        RECT 46.580 36.815 46.750 37.445 ;
        RECT 46.935 37.025 47.285 37.275 ;
        RECT 46.580 36.205 47.080 36.815 ;
        RECT 47.455 36.805 48.665 37.325 ;
        RECT 48.835 36.975 50.045 37.495 ;
        RECT 50.675 37.420 50.965 38.585 ;
        RECT 51.135 37.495 53.725 38.585 ;
        RECT 51.135 36.805 52.345 37.325 ;
        RECT 52.515 36.975 53.725 37.495 ;
        RECT 53.900 37.445 54.235 38.415 ;
        RECT 54.405 37.445 54.575 38.585 ;
        RECT 54.745 38.245 56.775 38.415 ;
        RECT 47.455 36.035 50.045 36.805 ;
        RECT 50.675 36.035 50.965 36.760 ;
        RECT 51.135 36.035 53.725 36.805 ;
        RECT 53.900 36.775 54.070 37.445 ;
        RECT 54.745 37.275 54.915 38.245 ;
        RECT 54.240 36.945 54.495 37.275 ;
        RECT 54.720 36.945 54.915 37.275 ;
        RECT 55.085 37.905 56.210 38.075 ;
        RECT 54.325 36.775 54.495 36.945 ;
        RECT 55.085 36.775 55.255 37.905 ;
        RECT 53.900 36.205 54.155 36.775 ;
        RECT 54.325 36.605 55.255 36.775 ;
        RECT 55.425 37.565 56.435 37.735 ;
        RECT 55.425 36.765 55.595 37.565 ;
        RECT 55.800 36.885 56.075 37.365 ;
        RECT 55.795 36.715 56.075 36.885 ;
        RECT 55.080 36.570 55.255 36.605 ;
        RECT 54.325 36.035 54.655 36.435 ;
        RECT 55.080 36.205 55.610 36.570 ;
        RECT 55.800 36.205 56.075 36.715 ;
        RECT 56.245 36.205 56.435 37.565 ;
        RECT 56.605 37.580 56.775 38.245 ;
        RECT 56.945 37.825 57.115 38.585 ;
        RECT 57.350 37.825 57.865 38.235 ;
        RECT 56.605 37.390 57.355 37.580 ;
        RECT 57.525 37.015 57.865 37.825 ;
        RECT 56.635 36.845 57.865 37.015 ;
        RECT 58.035 37.445 58.420 38.415 ;
        RECT 58.590 38.125 58.915 38.585 ;
        RECT 59.435 37.955 59.715 38.415 ;
        RECT 58.590 37.735 59.715 37.955 ;
        RECT 56.615 36.035 57.125 36.570 ;
        RECT 57.345 36.240 57.590 36.845 ;
        RECT 58.035 36.775 58.315 37.445 ;
        RECT 58.590 37.275 59.040 37.735 ;
        RECT 59.905 37.565 60.305 38.415 ;
        RECT 60.705 38.125 60.975 38.585 ;
        RECT 61.145 37.955 61.430 38.415 ;
        RECT 58.485 36.945 59.040 37.275 ;
        RECT 59.210 37.005 60.305 37.565 ;
        RECT 58.590 36.835 59.040 36.945 ;
        RECT 58.035 36.205 58.420 36.775 ;
        RECT 58.590 36.665 59.715 36.835 ;
        RECT 58.590 36.035 58.915 36.495 ;
        RECT 59.435 36.205 59.715 36.665 ;
        RECT 59.905 36.205 60.305 37.005 ;
        RECT 60.475 37.735 61.430 37.955 ;
        RECT 60.475 36.835 60.685 37.735 ;
        RECT 61.715 37.615 61.985 38.385 ;
        RECT 62.155 37.805 62.485 38.585 ;
        RECT 62.690 37.980 62.875 38.385 ;
        RECT 63.045 38.160 63.380 38.585 ;
        RECT 63.555 38.150 68.900 38.585 ;
        RECT 62.690 37.805 63.355 37.980 ;
        RECT 60.855 37.005 61.545 37.565 ;
        RECT 61.715 37.445 62.845 37.615 ;
        RECT 60.475 36.665 61.430 36.835 ;
        RECT 60.705 36.035 60.975 36.495 ;
        RECT 61.145 36.205 61.430 36.665 ;
        RECT 61.715 36.535 61.885 37.445 ;
        RECT 62.055 36.695 62.415 37.275 ;
        RECT 62.595 36.945 62.845 37.445 ;
        RECT 63.015 36.775 63.355 37.805 ;
        RECT 62.670 36.605 63.355 36.775 ;
        RECT 61.715 36.205 61.975 36.535 ;
        RECT 62.185 36.035 62.460 36.515 ;
        RECT 62.670 36.205 62.875 36.605 ;
        RECT 65.140 36.580 65.480 37.410 ;
        RECT 66.960 36.900 67.310 38.150 ;
        RECT 69.075 37.495 72.585 38.585 ;
        RECT 72.755 37.495 73.965 38.585 ;
        RECT 69.075 36.805 70.725 37.325 ;
        RECT 70.895 36.975 72.585 37.495 ;
        RECT 63.045 36.035 63.380 36.435 ;
        RECT 63.555 36.035 68.900 36.580 ;
        RECT 69.075 36.035 72.585 36.805 ;
        RECT 72.755 36.785 73.275 37.325 ;
        RECT 73.445 36.955 73.965 37.495 ;
        RECT 74.320 37.615 74.710 37.790 ;
        RECT 75.195 37.785 75.525 38.585 ;
        RECT 75.695 37.795 76.230 38.415 ;
        RECT 74.320 37.445 75.745 37.615 ;
        RECT 72.755 36.035 73.965 36.785 ;
        RECT 74.195 36.715 74.550 37.275 ;
        RECT 74.720 36.545 74.890 37.445 ;
        RECT 75.060 36.715 75.325 37.275 ;
        RECT 75.575 36.945 75.745 37.445 ;
        RECT 75.915 36.775 76.230 37.795 ;
        RECT 76.435 37.420 76.725 38.585 ;
        RECT 78.020 37.615 78.350 38.415 ;
        RECT 78.520 37.785 78.850 38.585 ;
        RECT 79.150 37.615 79.480 38.415 ;
        RECT 80.125 37.785 80.375 38.585 ;
        RECT 78.020 37.445 80.455 37.615 ;
        RECT 80.645 37.445 80.815 38.585 ;
        RECT 80.985 37.445 81.325 38.415 ;
        RECT 81.585 37.915 81.755 38.415 ;
        RECT 81.925 38.085 82.255 38.585 ;
        RECT 81.585 37.745 82.250 37.915 ;
        RECT 77.815 37.025 78.165 37.275 ;
        RECT 78.350 36.815 78.520 37.445 ;
        RECT 78.690 37.025 79.020 37.225 ;
        RECT 79.190 37.025 79.520 37.225 ;
        RECT 79.690 37.025 80.110 37.225 ;
        RECT 80.285 37.195 80.455 37.445 ;
        RECT 80.285 37.025 80.980 37.195 ;
        RECT 81.150 36.885 81.325 37.445 ;
        RECT 81.500 36.925 81.850 37.575 ;
        RECT 74.300 36.035 74.540 36.545 ;
        RECT 74.720 36.215 75.000 36.545 ;
        RECT 75.230 36.035 75.445 36.545 ;
        RECT 75.615 36.205 76.230 36.775 ;
        RECT 76.435 36.035 76.725 36.760 ;
        RECT 78.020 36.205 78.520 36.815 ;
        RECT 79.150 36.685 80.375 36.855 ;
        RECT 81.095 36.835 81.325 36.885 ;
        RECT 79.150 36.205 79.480 36.685 ;
        RECT 79.650 36.035 79.875 36.495 ;
        RECT 80.045 36.205 80.375 36.685 ;
        RECT 80.565 36.035 80.815 36.835 ;
        RECT 80.985 36.205 81.325 36.835 ;
        RECT 82.020 36.755 82.250 37.745 ;
        RECT 81.585 36.585 82.250 36.755 ;
        RECT 81.585 36.295 81.755 36.585 ;
        RECT 81.925 36.035 82.255 36.415 ;
        RECT 82.425 36.295 82.610 38.415 ;
        RECT 82.850 38.125 83.115 38.585 ;
        RECT 83.285 37.990 83.535 38.415 ;
        RECT 83.745 38.140 84.850 38.310 ;
        RECT 83.230 37.860 83.535 37.990 ;
        RECT 82.780 36.665 83.060 37.615 ;
        RECT 83.230 36.755 83.400 37.860 ;
        RECT 83.570 37.075 83.810 37.670 ;
        RECT 83.980 37.605 84.510 37.970 ;
        RECT 83.980 36.905 84.150 37.605 ;
        RECT 84.680 37.525 84.850 38.140 ;
        RECT 85.020 37.785 85.190 38.585 ;
        RECT 85.360 38.085 85.610 38.415 ;
        RECT 85.835 38.115 86.720 38.285 ;
        RECT 84.680 37.435 85.190 37.525 ;
        RECT 83.230 36.625 83.455 36.755 ;
        RECT 83.625 36.685 84.150 36.905 ;
        RECT 84.320 37.265 85.190 37.435 ;
        RECT 82.865 36.035 83.115 36.495 ;
        RECT 83.285 36.485 83.455 36.625 ;
        RECT 84.320 36.485 84.490 37.265 ;
        RECT 85.020 37.195 85.190 37.265 ;
        RECT 84.700 37.015 84.900 37.045 ;
        RECT 85.360 37.015 85.530 38.085 ;
        RECT 85.700 37.195 85.890 37.915 ;
        RECT 84.700 36.715 85.530 37.015 ;
        RECT 86.060 36.985 86.380 37.945 ;
        RECT 83.285 36.315 83.620 36.485 ;
        RECT 83.815 36.315 84.490 36.485 ;
        RECT 84.810 36.035 85.180 36.535 ;
        RECT 85.360 36.485 85.530 36.715 ;
        RECT 85.915 36.655 86.380 36.985 ;
        RECT 86.550 37.275 86.720 38.115 ;
        RECT 86.900 38.085 87.215 38.585 ;
        RECT 87.445 37.855 87.785 38.415 ;
        RECT 86.890 37.480 87.785 37.855 ;
        RECT 87.955 37.575 88.125 38.585 ;
        RECT 87.595 37.275 87.785 37.480 ;
        RECT 88.295 37.525 88.625 38.370 ;
        RECT 88.295 37.445 88.685 37.525 ;
        RECT 88.470 37.395 88.685 37.445 ;
        RECT 86.550 36.945 87.425 37.275 ;
        RECT 87.595 36.945 88.345 37.275 ;
        RECT 86.550 36.485 86.720 36.945 ;
        RECT 87.595 36.775 87.795 36.945 ;
        RECT 88.515 36.815 88.685 37.395 ;
        RECT 89.315 37.495 90.525 38.585 ;
        RECT 89.315 36.955 89.835 37.495 ;
        RECT 88.460 36.775 88.685 36.815 ;
        RECT 90.005 36.785 90.525 37.325 ;
        RECT 85.360 36.315 85.765 36.485 ;
        RECT 85.935 36.315 86.720 36.485 ;
        RECT 86.995 36.035 87.205 36.565 ;
        RECT 87.465 36.250 87.795 36.775 ;
        RECT 88.305 36.690 88.685 36.775 ;
        RECT 87.965 36.035 88.135 36.645 ;
        RECT 88.305 36.255 88.635 36.690 ;
        RECT 89.315 36.035 90.525 36.785 ;
        RECT 11.950 35.865 90.610 36.035 ;
        RECT 12.035 35.115 13.245 35.865 ;
        RECT 13.415 35.320 18.760 35.865 ;
        RECT 12.035 34.575 12.555 35.115 ;
        RECT 12.725 34.405 13.245 34.945 ;
        RECT 15.000 34.490 15.340 35.320 ;
        RECT 19.855 35.065 20.195 35.695 ;
        RECT 20.365 35.065 20.615 35.865 ;
        RECT 20.805 35.215 21.135 35.695 ;
        RECT 21.305 35.405 21.530 35.865 ;
        RECT 21.700 35.215 22.030 35.695 ;
        RECT 12.035 33.315 13.245 34.405 ;
        RECT 16.820 33.750 17.170 35.000 ;
        RECT 19.855 34.455 20.030 35.065 ;
        RECT 20.805 35.045 22.030 35.215 ;
        RECT 22.660 35.085 23.160 35.695 ;
        RECT 23.625 35.315 23.795 35.695 ;
        RECT 24.010 35.485 24.340 35.865 ;
        RECT 23.625 35.145 24.340 35.315 ;
        RECT 20.200 34.705 20.895 34.875 ;
        RECT 20.725 34.455 20.895 34.705 ;
        RECT 21.070 34.675 21.490 34.875 ;
        RECT 21.660 34.675 21.990 34.875 ;
        RECT 22.160 34.675 22.490 34.875 ;
        RECT 22.660 34.455 22.830 35.085 ;
        RECT 23.015 34.625 23.365 34.875 ;
        RECT 23.535 34.595 23.890 34.965 ;
        RECT 24.170 34.955 24.340 35.145 ;
        RECT 24.510 35.120 24.765 35.695 ;
        RECT 24.170 34.625 24.425 34.955 ;
        RECT 13.415 33.315 18.760 33.750 ;
        RECT 19.855 33.485 20.195 34.455 ;
        RECT 20.365 33.315 20.535 34.455 ;
        RECT 20.725 34.285 23.160 34.455 ;
        RECT 24.170 34.415 24.340 34.625 ;
        RECT 20.805 33.315 21.055 34.115 ;
        RECT 21.700 33.485 22.030 34.285 ;
        RECT 22.330 33.315 22.660 34.115 ;
        RECT 22.830 33.485 23.160 34.285 ;
        RECT 23.625 34.245 24.340 34.415 ;
        RECT 24.595 34.390 24.765 35.120 ;
        RECT 24.940 35.025 25.200 35.865 ;
        RECT 25.375 35.095 27.045 35.865 ;
        RECT 27.380 35.355 27.620 35.865 ;
        RECT 27.800 35.355 28.080 35.685 ;
        RECT 28.310 35.355 28.525 35.865 ;
        RECT 25.375 34.575 26.125 35.095 ;
        RECT 23.625 33.485 23.795 34.245 ;
        RECT 24.010 33.315 24.340 34.075 ;
        RECT 24.510 33.485 24.765 34.390 ;
        RECT 24.940 33.315 25.200 34.465 ;
        RECT 26.295 34.405 27.045 34.925 ;
        RECT 27.275 34.625 27.630 35.185 ;
        RECT 27.800 34.455 27.970 35.355 ;
        RECT 28.140 34.625 28.405 35.185 ;
        RECT 28.695 35.125 29.310 35.695 ;
        RECT 29.605 35.315 29.775 35.605 ;
        RECT 29.945 35.485 30.275 35.865 ;
        RECT 29.605 35.145 30.270 35.315 ;
        RECT 28.655 34.455 28.825 34.955 ;
        RECT 25.375 33.315 27.045 34.405 ;
        RECT 27.400 34.285 28.825 34.455 ;
        RECT 27.400 34.110 27.790 34.285 ;
        RECT 28.275 33.315 28.605 34.115 ;
        RECT 28.995 34.105 29.310 35.125 ;
        RECT 29.520 34.325 29.870 34.975 ;
        RECT 30.040 34.155 30.270 35.145 ;
        RECT 28.775 33.485 29.310 34.105 ;
        RECT 29.605 33.985 30.270 34.155 ;
        RECT 29.605 33.485 29.775 33.985 ;
        RECT 29.945 33.315 30.275 33.815 ;
        RECT 30.445 33.485 30.630 35.605 ;
        RECT 30.885 35.405 31.135 35.865 ;
        RECT 31.305 35.415 31.640 35.585 ;
        RECT 31.835 35.415 32.510 35.585 ;
        RECT 31.305 35.275 31.475 35.415 ;
        RECT 30.800 34.285 31.080 35.235 ;
        RECT 31.250 35.145 31.475 35.275 ;
        RECT 31.250 34.040 31.420 35.145 ;
        RECT 31.645 34.995 32.170 35.215 ;
        RECT 31.590 34.230 31.830 34.825 ;
        RECT 32.000 34.295 32.170 34.995 ;
        RECT 32.340 34.635 32.510 35.415 ;
        RECT 32.830 35.365 33.200 35.865 ;
        RECT 33.380 35.415 33.785 35.585 ;
        RECT 33.955 35.415 34.740 35.585 ;
        RECT 33.380 35.185 33.550 35.415 ;
        RECT 32.720 34.885 33.550 35.185 ;
        RECT 33.935 34.915 34.400 35.245 ;
        RECT 32.720 34.855 32.920 34.885 ;
        RECT 33.040 34.635 33.210 34.705 ;
        RECT 32.340 34.465 33.210 34.635 ;
        RECT 32.700 34.375 33.210 34.465 ;
        RECT 31.250 33.910 31.555 34.040 ;
        RECT 32.000 33.930 32.530 34.295 ;
        RECT 30.870 33.315 31.135 33.775 ;
        RECT 31.305 33.485 31.555 33.910 ;
        RECT 32.700 33.760 32.870 34.375 ;
        RECT 31.765 33.590 32.870 33.760 ;
        RECT 33.040 33.315 33.210 34.115 ;
        RECT 33.380 33.815 33.550 34.885 ;
        RECT 33.720 33.985 33.910 34.705 ;
        RECT 34.080 33.955 34.400 34.915 ;
        RECT 34.570 34.955 34.740 35.415 ;
        RECT 35.015 35.335 35.225 35.865 ;
        RECT 35.485 35.125 35.815 35.650 ;
        RECT 35.985 35.255 36.155 35.865 ;
        RECT 36.325 35.210 36.655 35.645 ;
        RECT 36.325 35.125 36.705 35.210 ;
        RECT 37.795 35.140 38.085 35.865 ;
        RECT 35.615 34.955 35.815 35.125 ;
        RECT 36.480 35.085 36.705 35.125 ;
        RECT 38.260 35.100 38.715 35.865 ;
        RECT 38.990 35.485 40.290 35.695 ;
        RECT 40.545 35.505 40.875 35.865 ;
        RECT 40.120 35.335 40.290 35.485 ;
        RECT 41.045 35.365 41.305 35.695 ;
        RECT 41.075 35.355 41.305 35.365 ;
        RECT 41.640 35.355 41.880 35.865 ;
        RECT 42.060 35.355 42.340 35.685 ;
        RECT 42.570 35.355 42.785 35.865 ;
        RECT 34.570 34.625 35.445 34.955 ;
        RECT 35.615 34.625 36.365 34.955 ;
        RECT 33.380 33.485 33.630 33.815 ;
        RECT 34.570 33.785 34.740 34.625 ;
        RECT 35.615 34.420 35.805 34.625 ;
        RECT 36.535 34.505 36.705 35.085 ;
        RECT 39.190 34.875 39.410 35.275 ;
        RECT 38.255 34.675 38.745 34.875 ;
        RECT 38.935 34.665 39.410 34.875 ;
        RECT 39.655 34.875 39.865 35.275 ;
        RECT 40.120 35.210 40.875 35.335 ;
        RECT 40.120 35.165 40.965 35.210 ;
        RECT 40.695 35.045 40.965 35.165 ;
        RECT 39.655 34.665 39.985 34.875 ;
        RECT 40.155 34.605 40.565 34.910 ;
        RECT 36.490 34.455 36.705 34.505 ;
        RECT 34.910 34.045 35.805 34.420 ;
        RECT 36.315 34.375 36.705 34.455 ;
        RECT 33.855 33.615 34.740 33.785 ;
        RECT 34.920 33.315 35.235 33.815 ;
        RECT 35.465 33.485 35.805 34.045 ;
        RECT 35.975 33.315 36.145 34.325 ;
        RECT 36.315 33.530 36.645 34.375 ;
        RECT 37.795 33.315 38.085 34.480 ;
        RECT 38.260 34.435 39.435 34.495 ;
        RECT 40.795 34.470 40.965 35.045 ;
        RECT 40.765 34.435 40.965 34.470 ;
        RECT 38.260 34.325 40.965 34.435 ;
        RECT 38.260 33.705 38.515 34.325 ;
        RECT 39.105 34.265 40.905 34.325 ;
        RECT 39.105 34.235 39.435 34.265 ;
        RECT 41.135 34.165 41.305 35.355 ;
        RECT 41.535 34.625 41.890 35.185 ;
        RECT 42.060 34.455 42.230 35.355 ;
        RECT 42.400 34.625 42.665 35.185 ;
        RECT 42.955 35.125 43.570 35.695 ;
        RECT 43.775 35.320 49.120 35.865 ;
        RECT 42.915 34.455 43.085 34.955 ;
        RECT 38.765 34.065 38.950 34.155 ;
        RECT 39.540 34.065 40.375 34.075 ;
        RECT 38.765 33.865 40.375 34.065 ;
        RECT 38.765 33.825 38.995 33.865 ;
        RECT 38.260 33.485 38.595 33.705 ;
        RECT 39.600 33.315 39.955 33.695 ;
        RECT 40.125 33.485 40.375 33.865 ;
        RECT 40.625 33.315 40.875 34.095 ;
        RECT 41.045 33.485 41.305 34.165 ;
        RECT 41.660 34.285 43.085 34.455 ;
        RECT 41.660 34.110 42.050 34.285 ;
        RECT 42.535 33.315 42.865 34.115 ;
        RECT 43.255 34.105 43.570 35.125 ;
        RECT 45.360 34.490 45.700 35.320 ;
        RECT 49.295 35.095 50.965 35.865 ;
        RECT 43.035 33.485 43.570 34.105 ;
        RECT 47.180 33.750 47.530 35.000 ;
        RECT 49.295 34.575 50.045 35.095 ;
        RECT 51.140 35.045 51.415 35.865 ;
        RECT 51.585 35.225 51.915 35.695 ;
        RECT 52.085 35.395 52.255 35.865 ;
        RECT 52.425 35.225 52.755 35.695 ;
        RECT 52.925 35.395 53.635 35.865 ;
        RECT 53.805 35.225 54.135 35.695 ;
        RECT 54.305 35.395 54.595 35.865 ;
        RECT 51.585 35.045 54.645 35.225 ;
        RECT 50.215 34.405 50.965 34.925 ;
        RECT 51.185 34.665 52.015 34.875 ;
        RECT 52.185 34.665 53.235 34.875 ;
        RECT 53.425 34.665 54.015 34.875 ;
        RECT 43.775 33.315 49.120 33.750 ;
        RECT 49.295 33.315 50.965 34.405 ;
        RECT 51.200 34.325 53.135 34.495 ;
        RECT 53.425 34.325 53.690 34.665 ;
        RECT 54.185 34.495 54.645 35.045 ;
        RECT 54.815 35.115 56.025 35.865 ;
        RECT 56.285 35.315 56.455 35.605 ;
        RECT 56.625 35.485 56.955 35.865 ;
        RECT 56.285 35.145 56.950 35.315 ;
        RECT 54.815 34.575 55.335 35.115 ;
        RECT 53.885 34.325 54.645 34.495 ;
        RECT 55.505 34.405 56.025 34.945 ;
        RECT 51.200 33.485 51.455 34.325 ;
        RECT 51.625 33.315 51.875 34.155 ;
        RECT 52.045 33.485 52.295 34.325 ;
        RECT 52.465 33.655 52.715 34.155 ;
        RECT 52.885 33.825 53.135 34.325 ;
        RECT 53.465 33.655 53.675 34.155 ;
        RECT 53.885 33.825 54.095 34.325 ;
        RECT 54.265 33.655 54.515 34.155 ;
        RECT 52.465 33.485 54.515 33.655 ;
        RECT 54.815 33.315 56.025 34.405 ;
        RECT 56.200 34.325 56.550 34.975 ;
        RECT 56.720 34.155 56.950 35.145 ;
        RECT 56.285 33.985 56.950 34.155 ;
        RECT 56.285 33.485 56.455 33.985 ;
        RECT 56.625 33.315 56.955 33.815 ;
        RECT 57.125 33.485 57.310 35.605 ;
        RECT 57.565 35.405 57.815 35.865 ;
        RECT 57.985 35.415 58.320 35.585 ;
        RECT 58.515 35.415 59.190 35.585 ;
        RECT 57.985 35.275 58.155 35.415 ;
        RECT 57.480 34.285 57.760 35.235 ;
        RECT 57.930 35.145 58.155 35.275 ;
        RECT 57.930 34.040 58.100 35.145 ;
        RECT 58.325 34.995 58.850 35.215 ;
        RECT 58.270 34.230 58.510 34.825 ;
        RECT 58.680 34.295 58.850 34.995 ;
        RECT 59.020 34.635 59.190 35.415 ;
        RECT 59.510 35.365 59.880 35.865 ;
        RECT 60.060 35.415 60.465 35.585 ;
        RECT 60.635 35.415 61.420 35.585 ;
        RECT 60.060 35.185 60.230 35.415 ;
        RECT 59.400 34.885 60.230 35.185 ;
        RECT 60.615 34.915 61.080 35.245 ;
        RECT 59.400 34.855 59.600 34.885 ;
        RECT 59.720 34.635 59.890 34.705 ;
        RECT 59.020 34.465 59.890 34.635 ;
        RECT 59.380 34.375 59.890 34.465 ;
        RECT 57.930 33.910 58.235 34.040 ;
        RECT 58.680 33.930 59.210 34.295 ;
        RECT 57.550 33.315 57.815 33.775 ;
        RECT 57.985 33.485 58.235 33.910 ;
        RECT 59.380 33.760 59.550 34.375 ;
        RECT 58.445 33.590 59.550 33.760 ;
        RECT 59.720 33.315 59.890 34.115 ;
        RECT 60.060 33.815 60.230 34.885 ;
        RECT 60.400 33.985 60.590 34.705 ;
        RECT 60.760 33.955 61.080 34.915 ;
        RECT 61.250 34.955 61.420 35.415 ;
        RECT 61.695 35.335 61.905 35.865 ;
        RECT 62.165 35.125 62.495 35.650 ;
        RECT 62.665 35.255 62.835 35.865 ;
        RECT 63.005 35.210 63.335 35.645 ;
        RECT 63.005 35.125 63.385 35.210 ;
        RECT 63.555 35.140 63.845 35.865 ;
        RECT 62.295 34.955 62.495 35.125 ;
        RECT 63.160 35.085 63.385 35.125 ;
        RECT 61.250 34.625 62.125 34.955 ;
        RECT 62.295 34.625 63.045 34.955 ;
        RECT 60.060 33.485 60.310 33.815 ;
        RECT 61.250 33.785 61.420 34.625 ;
        RECT 62.295 34.420 62.485 34.625 ;
        RECT 63.215 34.505 63.385 35.085 ;
        RECT 64.015 35.095 67.525 35.865 ;
        RECT 64.015 34.575 65.665 35.095 ;
        RECT 68.155 35.065 68.445 35.865 ;
        RECT 68.615 35.405 69.165 35.695 ;
        RECT 69.335 35.405 69.585 35.865 ;
        RECT 63.170 34.455 63.385 34.505 ;
        RECT 61.590 34.045 62.485 34.420 ;
        RECT 62.995 34.375 63.385 34.455 ;
        RECT 60.535 33.615 61.420 33.785 ;
        RECT 61.600 33.315 61.915 33.815 ;
        RECT 62.145 33.485 62.485 34.045 ;
        RECT 62.655 33.315 62.825 34.325 ;
        RECT 62.995 33.530 63.325 34.375 ;
        RECT 63.555 33.315 63.845 34.480 ;
        RECT 65.835 34.405 67.525 34.925 ;
        RECT 64.015 33.315 67.525 34.405 ;
        RECT 68.155 33.315 68.445 34.455 ;
        RECT 68.615 34.035 68.865 35.405 ;
        RECT 70.215 35.235 70.545 35.595 ;
        RECT 69.155 35.045 70.545 35.235 ;
        RECT 70.915 35.235 71.255 35.695 ;
        RECT 71.425 35.405 71.595 35.865 ;
        RECT 71.765 35.485 72.935 35.695 ;
        RECT 71.765 35.235 72.015 35.485 ;
        RECT 72.605 35.465 72.935 35.485 ;
        RECT 70.915 35.065 72.015 35.235 ;
        RECT 72.185 35.045 73.045 35.295 ;
        RECT 69.155 34.955 69.325 35.045 ;
        RECT 69.035 34.625 69.325 34.955 ;
        RECT 69.495 34.625 69.825 34.875 ;
        RECT 70.055 34.625 70.745 34.875 ;
        RECT 70.915 34.625 71.675 34.875 ;
        RECT 71.845 34.625 72.595 34.875 ;
        RECT 69.155 34.375 69.325 34.625 ;
        RECT 69.155 34.205 70.095 34.375 ;
        RECT 68.615 33.485 69.065 34.035 ;
        RECT 69.255 33.315 69.585 34.035 ;
        RECT 69.795 33.655 70.095 34.205 ;
        RECT 70.430 34.185 70.745 34.625 ;
        RECT 72.765 34.455 73.045 35.045 ;
        RECT 73.215 35.095 74.885 35.865 ;
        RECT 75.680 35.355 75.920 35.865 ;
        RECT 76.100 35.355 76.380 35.685 ;
        RECT 76.610 35.355 76.825 35.865 ;
        RECT 73.215 34.575 73.965 35.095 ;
        RECT 70.265 33.315 70.545 33.985 ;
        RECT 70.915 33.315 71.175 34.455 ;
        RECT 71.345 34.285 73.045 34.455 ;
        RECT 74.135 34.405 74.885 34.925 ;
        RECT 75.575 34.625 75.930 35.185 ;
        RECT 76.100 34.455 76.270 35.355 ;
        RECT 76.440 34.625 76.705 35.185 ;
        RECT 76.995 35.125 77.610 35.695 ;
        RECT 76.955 34.455 77.125 34.955 ;
        RECT 71.345 33.485 71.675 34.285 ;
        RECT 71.845 33.315 72.015 34.115 ;
        RECT 72.185 33.485 72.515 34.285 ;
        RECT 72.685 33.315 72.940 34.115 ;
        RECT 73.215 33.315 74.885 34.405 ;
        RECT 75.700 34.285 77.125 34.455 ;
        RECT 75.700 34.110 76.090 34.285 ;
        RECT 76.575 33.315 76.905 34.115 ;
        RECT 77.295 34.105 77.610 35.125 ;
        RECT 77.075 33.485 77.610 34.105 ;
        RECT 77.815 35.365 78.075 35.695 ;
        RECT 78.245 35.505 78.575 35.865 ;
        RECT 78.830 35.485 80.130 35.695 ;
        RECT 77.815 34.165 77.985 35.365 ;
        RECT 78.830 35.335 79.000 35.485 ;
        RECT 78.245 35.210 79.000 35.335 ;
        RECT 78.155 35.165 79.000 35.210 ;
        RECT 78.155 35.045 78.425 35.165 ;
        RECT 78.155 34.470 78.325 35.045 ;
        RECT 78.555 34.605 78.965 34.910 ;
        RECT 79.255 34.875 79.465 35.275 ;
        RECT 79.135 34.665 79.465 34.875 ;
        RECT 79.710 34.875 79.930 35.275 ;
        RECT 80.405 35.100 80.860 35.865 ;
        RECT 82.045 35.315 82.215 35.605 ;
        RECT 82.385 35.485 82.715 35.865 ;
        RECT 82.045 35.145 82.710 35.315 ;
        RECT 79.710 34.665 80.185 34.875 ;
        RECT 80.375 34.675 80.865 34.875 ;
        RECT 78.155 34.435 78.355 34.470 ;
        RECT 79.685 34.435 80.860 34.495 ;
        RECT 78.155 34.325 80.860 34.435 ;
        RECT 81.960 34.325 82.310 34.975 ;
        RECT 78.215 34.265 80.015 34.325 ;
        RECT 79.685 34.235 80.015 34.265 ;
        RECT 77.815 33.485 78.075 34.165 ;
        RECT 78.245 33.315 78.495 34.095 ;
        RECT 78.745 34.065 79.580 34.075 ;
        RECT 80.170 34.065 80.355 34.155 ;
        RECT 78.745 33.865 80.355 34.065 ;
        RECT 78.745 33.485 78.995 33.865 ;
        RECT 80.125 33.825 80.355 33.865 ;
        RECT 80.605 33.705 80.860 34.325 ;
        RECT 82.480 34.155 82.710 35.145 ;
        RECT 79.165 33.315 79.520 33.695 ;
        RECT 80.525 33.485 80.860 33.705 ;
        RECT 82.045 33.985 82.710 34.155 ;
        RECT 82.045 33.485 82.215 33.985 ;
        RECT 82.385 33.315 82.715 33.815 ;
        RECT 82.885 33.485 83.070 35.605 ;
        RECT 83.325 35.405 83.575 35.865 ;
        RECT 83.745 35.415 84.080 35.585 ;
        RECT 84.275 35.415 84.950 35.585 ;
        RECT 83.745 35.275 83.915 35.415 ;
        RECT 83.240 34.285 83.520 35.235 ;
        RECT 83.690 35.145 83.915 35.275 ;
        RECT 83.690 34.040 83.860 35.145 ;
        RECT 84.085 34.995 84.610 35.215 ;
        RECT 84.030 34.230 84.270 34.825 ;
        RECT 84.440 34.295 84.610 34.995 ;
        RECT 84.780 34.635 84.950 35.415 ;
        RECT 85.270 35.365 85.640 35.865 ;
        RECT 85.820 35.415 86.225 35.585 ;
        RECT 86.395 35.415 87.180 35.585 ;
        RECT 85.820 35.185 85.990 35.415 ;
        RECT 85.160 34.885 85.990 35.185 ;
        RECT 86.375 34.915 86.840 35.245 ;
        RECT 85.160 34.855 85.360 34.885 ;
        RECT 85.480 34.635 85.650 34.705 ;
        RECT 84.780 34.465 85.650 34.635 ;
        RECT 85.140 34.375 85.650 34.465 ;
        RECT 83.690 33.910 83.995 34.040 ;
        RECT 84.440 33.930 84.970 34.295 ;
        RECT 83.310 33.315 83.575 33.775 ;
        RECT 83.745 33.485 83.995 33.910 ;
        RECT 85.140 33.760 85.310 34.375 ;
        RECT 84.205 33.590 85.310 33.760 ;
        RECT 85.480 33.315 85.650 34.115 ;
        RECT 85.820 33.815 85.990 34.885 ;
        RECT 86.160 33.985 86.350 34.705 ;
        RECT 86.520 33.955 86.840 34.915 ;
        RECT 87.010 34.955 87.180 35.415 ;
        RECT 87.455 35.335 87.665 35.865 ;
        RECT 87.925 35.125 88.255 35.650 ;
        RECT 88.425 35.255 88.595 35.865 ;
        RECT 88.765 35.210 89.095 35.645 ;
        RECT 88.765 35.125 89.145 35.210 ;
        RECT 88.055 34.955 88.255 35.125 ;
        RECT 88.920 35.085 89.145 35.125 ;
        RECT 89.315 35.115 90.525 35.865 ;
        RECT 87.010 34.625 87.885 34.955 ;
        RECT 88.055 34.625 88.805 34.955 ;
        RECT 85.820 33.485 86.070 33.815 ;
        RECT 87.010 33.785 87.180 34.625 ;
        RECT 88.055 34.420 88.245 34.625 ;
        RECT 88.975 34.505 89.145 35.085 ;
        RECT 88.930 34.455 89.145 34.505 ;
        RECT 87.350 34.045 88.245 34.420 ;
        RECT 88.755 34.375 89.145 34.455 ;
        RECT 89.315 34.405 89.835 34.945 ;
        RECT 90.005 34.575 90.525 35.115 ;
        RECT 86.295 33.615 87.180 33.785 ;
        RECT 87.360 33.315 87.675 33.815 ;
        RECT 87.905 33.485 88.245 34.045 ;
        RECT 88.415 33.315 88.585 34.325 ;
        RECT 88.755 33.530 89.085 34.375 ;
        RECT 89.315 33.315 90.525 34.405 ;
        RECT 11.950 33.145 90.610 33.315 ;
        RECT 12.035 32.055 13.245 33.145 ;
        RECT 12.035 31.345 12.555 31.885 ;
        RECT 12.725 31.515 13.245 32.055 ;
        RECT 13.420 31.995 13.680 33.145 ;
        RECT 13.855 32.070 14.110 32.975 ;
        RECT 14.280 32.385 14.610 33.145 ;
        RECT 14.825 32.215 14.995 32.975 ;
        RECT 12.035 30.595 13.245 31.345 ;
        RECT 13.420 30.595 13.680 31.435 ;
        RECT 13.855 31.340 14.025 32.070 ;
        RECT 14.280 32.045 14.995 32.215 ;
        RECT 15.750 32.355 16.285 32.975 ;
        RECT 14.280 31.835 14.450 32.045 ;
        RECT 14.195 31.505 14.450 31.835 ;
        RECT 13.855 30.765 14.110 31.340 ;
        RECT 14.280 31.315 14.450 31.505 ;
        RECT 14.730 31.495 15.085 31.865 ;
        RECT 15.750 31.335 16.065 32.355 ;
        RECT 16.455 32.345 16.785 33.145 ;
        RECT 17.270 32.175 17.660 32.350 ;
        RECT 16.235 32.005 17.660 32.175 ;
        RECT 18.015 32.055 19.685 33.145 ;
        RECT 16.235 31.505 16.405 32.005 ;
        RECT 14.280 31.145 14.995 31.315 ;
        RECT 14.280 30.595 14.610 30.975 ;
        RECT 14.825 30.765 14.995 31.145 ;
        RECT 15.750 30.765 16.365 31.335 ;
        RECT 16.655 31.275 16.920 31.835 ;
        RECT 17.090 31.105 17.260 32.005 ;
        RECT 17.430 31.275 17.785 31.835 ;
        RECT 18.015 31.365 18.765 31.885 ;
        RECT 18.935 31.535 19.685 32.055 ;
        RECT 20.315 32.005 20.655 32.975 ;
        RECT 20.825 32.005 20.995 33.145 ;
        RECT 21.265 32.345 21.515 33.145 ;
        RECT 22.160 32.175 22.490 32.975 ;
        RECT 22.790 32.345 23.120 33.145 ;
        RECT 23.290 32.175 23.620 32.975 ;
        RECT 21.185 32.005 23.620 32.175 ;
        RECT 20.315 31.395 20.490 32.005 ;
        RECT 21.185 31.755 21.355 32.005 ;
        RECT 20.660 31.585 21.355 31.755 ;
        RECT 21.530 31.585 21.950 31.785 ;
        RECT 22.120 31.585 22.450 31.785 ;
        RECT 22.620 31.585 22.950 31.785 ;
        RECT 16.535 30.595 16.750 31.105 ;
        RECT 16.980 30.775 17.260 31.105 ;
        RECT 17.440 30.595 17.680 31.105 ;
        RECT 18.015 30.595 19.685 31.365 ;
        RECT 20.315 30.765 20.655 31.395 ;
        RECT 20.825 30.595 21.075 31.395 ;
        RECT 21.265 31.245 22.490 31.415 ;
        RECT 21.265 30.765 21.595 31.245 ;
        RECT 21.765 30.595 21.990 31.055 ;
        RECT 22.160 30.765 22.490 31.245 ;
        RECT 23.120 31.375 23.290 32.005 ;
        RECT 24.915 31.980 25.205 33.145 ;
        RECT 25.375 32.710 30.720 33.145 ;
        RECT 30.895 32.710 36.240 33.145 ;
        RECT 36.415 32.710 41.760 33.145 ;
        RECT 23.475 31.585 23.825 31.835 ;
        RECT 23.120 30.765 23.620 31.375 ;
        RECT 24.915 30.595 25.205 31.320 ;
        RECT 26.960 31.140 27.300 31.970 ;
        RECT 28.780 31.460 29.130 32.710 ;
        RECT 32.480 31.140 32.820 31.970 ;
        RECT 34.300 31.460 34.650 32.710 ;
        RECT 38.000 31.140 38.340 31.970 ;
        RECT 39.820 31.460 40.170 32.710 ;
        RECT 43.040 32.175 43.430 32.350 ;
        RECT 43.915 32.345 44.245 33.145 ;
        RECT 44.415 32.355 44.950 32.975 ;
        RECT 43.040 32.005 44.465 32.175 ;
        RECT 42.915 31.275 43.270 31.835 ;
        RECT 25.375 30.595 30.720 31.140 ;
        RECT 30.895 30.595 36.240 31.140 ;
        RECT 36.415 30.595 41.760 31.140 ;
        RECT 43.440 31.105 43.610 32.005 ;
        RECT 43.780 31.275 44.045 31.835 ;
        RECT 44.295 31.505 44.465 32.005 ;
        RECT 44.635 31.335 44.950 32.355 ;
        RECT 45.155 32.055 46.825 33.145 ;
        RECT 43.020 30.595 43.260 31.105 ;
        RECT 43.440 30.775 43.720 31.105 ;
        RECT 43.950 30.595 44.165 31.105 ;
        RECT 44.335 30.765 44.950 31.335 ;
        RECT 45.155 31.365 45.905 31.885 ;
        RECT 46.075 31.535 46.825 32.055 ;
        RECT 47.460 32.755 47.795 32.975 ;
        RECT 48.800 32.765 49.155 33.145 ;
        RECT 47.460 32.135 47.715 32.755 ;
        RECT 47.965 32.595 48.195 32.635 ;
        RECT 49.325 32.595 49.575 32.975 ;
        RECT 47.965 32.395 49.575 32.595 ;
        RECT 47.965 32.305 48.150 32.395 ;
        RECT 48.740 32.385 49.575 32.395 ;
        RECT 49.825 32.365 50.075 33.145 ;
        RECT 50.245 32.295 50.505 32.975 ;
        RECT 48.305 32.195 48.635 32.225 ;
        RECT 48.305 32.135 50.105 32.195 ;
        RECT 47.460 32.025 50.165 32.135 ;
        RECT 47.460 31.965 48.635 32.025 ;
        RECT 49.965 31.990 50.165 32.025 ;
        RECT 47.455 31.585 47.945 31.785 ;
        RECT 48.135 31.585 48.610 31.795 ;
        RECT 45.155 30.595 46.825 31.365 ;
        RECT 47.460 30.595 47.915 31.360 ;
        RECT 48.390 31.185 48.610 31.585 ;
        RECT 48.855 31.585 49.185 31.795 ;
        RECT 48.855 31.185 49.065 31.585 ;
        RECT 49.355 31.550 49.765 31.855 ;
        RECT 49.995 31.415 50.165 31.990 ;
        RECT 49.895 31.295 50.165 31.415 ;
        RECT 49.320 31.250 50.165 31.295 ;
        RECT 49.320 31.125 50.075 31.250 ;
        RECT 49.320 30.975 49.490 31.125 ;
        RECT 50.335 31.095 50.505 32.295 ;
        RECT 50.675 31.980 50.965 33.145 ;
        RECT 51.135 32.055 52.345 33.145 ;
        RECT 51.135 31.345 51.655 31.885 ;
        RECT 51.825 31.515 52.345 32.055 ;
        RECT 52.720 32.175 53.050 32.975 ;
        RECT 53.220 32.345 53.550 33.145 ;
        RECT 53.850 32.175 54.180 32.975 ;
        RECT 54.825 32.345 55.075 33.145 ;
        RECT 52.720 32.005 55.155 32.175 ;
        RECT 55.345 32.005 55.515 33.145 ;
        RECT 55.685 32.005 56.025 32.975 ;
        RECT 52.515 31.585 52.865 31.835 ;
        RECT 53.050 31.375 53.220 32.005 ;
        RECT 53.390 31.585 53.720 31.785 ;
        RECT 53.890 31.585 54.220 31.785 ;
        RECT 54.390 31.585 54.810 31.785 ;
        RECT 54.985 31.755 55.155 32.005 ;
        RECT 54.985 31.585 55.680 31.755 ;
        RECT 48.190 30.765 49.490 30.975 ;
        RECT 49.745 30.595 50.075 30.955 ;
        RECT 50.245 30.765 50.505 31.095 ;
        RECT 50.675 30.595 50.965 31.320 ;
        RECT 51.135 30.595 52.345 31.345 ;
        RECT 52.720 30.765 53.220 31.375 ;
        RECT 53.850 31.245 55.075 31.415 ;
        RECT 55.850 31.395 56.025 32.005 ;
        RECT 53.850 30.765 54.180 31.245 ;
        RECT 54.350 30.595 54.575 31.055 ;
        RECT 54.745 30.765 55.075 31.245 ;
        RECT 55.265 30.595 55.515 31.395 ;
        RECT 55.685 30.765 56.025 31.395 ;
        RECT 56.230 32.355 56.765 32.975 ;
        RECT 56.230 31.335 56.545 32.355 ;
        RECT 56.935 32.345 57.265 33.145 ;
        RECT 58.585 32.475 58.755 32.975 ;
        RECT 58.925 32.645 59.255 33.145 ;
        RECT 57.750 32.175 58.140 32.350 ;
        RECT 58.585 32.305 59.250 32.475 ;
        RECT 56.715 32.005 58.140 32.175 ;
        RECT 56.715 31.505 56.885 32.005 ;
        RECT 56.230 30.765 56.845 31.335 ;
        RECT 57.135 31.275 57.400 31.835 ;
        RECT 57.570 31.105 57.740 32.005 ;
        RECT 57.910 31.275 58.265 31.835 ;
        RECT 58.500 31.485 58.850 32.135 ;
        RECT 59.020 31.315 59.250 32.305 ;
        RECT 58.585 31.145 59.250 31.315 ;
        RECT 57.015 30.595 57.230 31.105 ;
        RECT 57.460 30.775 57.740 31.105 ;
        RECT 57.920 30.595 58.160 31.105 ;
        RECT 58.585 30.855 58.755 31.145 ;
        RECT 58.925 30.595 59.255 30.975 ;
        RECT 59.425 30.855 59.610 32.975 ;
        RECT 59.850 32.685 60.115 33.145 ;
        RECT 60.285 32.550 60.535 32.975 ;
        RECT 60.745 32.700 61.850 32.870 ;
        RECT 60.230 32.420 60.535 32.550 ;
        RECT 59.780 31.225 60.060 32.175 ;
        RECT 60.230 31.315 60.400 32.420 ;
        RECT 60.570 31.635 60.810 32.230 ;
        RECT 60.980 32.165 61.510 32.530 ;
        RECT 60.980 31.465 61.150 32.165 ;
        RECT 61.680 32.085 61.850 32.700 ;
        RECT 62.020 32.345 62.190 33.145 ;
        RECT 62.360 32.645 62.610 32.975 ;
        RECT 62.835 32.675 63.720 32.845 ;
        RECT 61.680 31.995 62.190 32.085 ;
        RECT 60.230 31.185 60.455 31.315 ;
        RECT 60.625 31.245 61.150 31.465 ;
        RECT 61.320 31.825 62.190 31.995 ;
        RECT 59.865 30.595 60.115 31.055 ;
        RECT 60.285 31.045 60.455 31.185 ;
        RECT 61.320 31.045 61.490 31.825 ;
        RECT 62.020 31.755 62.190 31.825 ;
        RECT 61.700 31.575 61.900 31.605 ;
        RECT 62.360 31.575 62.530 32.645 ;
        RECT 62.700 31.755 62.890 32.475 ;
        RECT 61.700 31.275 62.530 31.575 ;
        RECT 63.060 31.545 63.380 32.505 ;
        RECT 60.285 30.875 60.620 31.045 ;
        RECT 60.815 30.875 61.490 31.045 ;
        RECT 61.810 30.595 62.180 31.095 ;
        RECT 62.360 31.045 62.530 31.275 ;
        RECT 62.915 31.215 63.380 31.545 ;
        RECT 63.550 31.835 63.720 32.675 ;
        RECT 63.900 32.645 64.215 33.145 ;
        RECT 64.445 32.415 64.785 32.975 ;
        RECT 63.890 32.040 64.785 32.415 ;
        RECT 64.955 32.135 65.125 33.145 ;
        RECT 64.595 31.835 64.785 32.040 ;
        RECT 65.295 32.085 65.625 32.930 ;
        RECT 65.890 32.355 66.425 32.975 ;
        RECT 65.295 32.005 65.685 32.085 ;
        RECT 65.470 31.955 65.685 32.005 ;
        RECT 63.550 31.505 64.425 31.835 ;
        RECT 64.595 31.505 65.345 31.835 ;
        RECT 63.550 31.045 63.720 31.505 ;
        RECT 64.595 31.335 64.795 31.505 ;
        RECT 65.515 31.375 65.685 31.955 ;
        RECT 65.460 31.335 65.685 31.375 ;
        RECT 62.360 30.875 62.765 31.045 ;
        RECT 62.935 30.875 63.720 31.045 ;
        RECT 63.995 30.595 64.205 31.125 ;
        RECT 64.465 30.810 64.795 31.335 ;
        RECT 65.305 31.250 65.685 31.335 ;
        RECT 65.890 31.335 66.205 32.355 ;
        RECT 66.595 32.345 66.925 33.145 ;
        RECT 68.245 32.475 68.415 32.975 ;
        RECT 68.585 32.645 68.915 33.145 ;
        RECT 67.410 32.175 67.800 32.350 ;
        RECT 68.245 32.305 68.910 32.475 ;
        RECT 66.375 32.005 67.800 32.175 ;
        RECT 66.375 31.505 66.545 32.005 ;
        RECT 64.965 30.595 65.135 31.205 ;
        RECT 65.305 30.815 65.635 31.250 ;
        RECT 65.890 30.765 66.505 31.335 ;
        RECT 66.795 31.275 67.060 31.835 ;
        RECT 67.230 31.105 67.400 32.005 ;
        RECT 67.570 31.275 67.925 31.835 ;
        RECT 68.160 31.485 68.510 32.135 ;
        RECT 68.680 31.315 68.910 32.305 ;
        RECT 68.245 31.145 68.910 31.315 ;
        RECT 66.675 30.595 66.890 31.105 ;
        RECT 67.120 30.775 67.400 31.105 ;
        RECT 67.580 30.595 67.820 31.105 ;
        RECT 68.245 30.855 68.415 31.145 ;
        RECT 68.585 30.595 68.915 30.975 ;
        RECT 69.085 30.855 69.270 32.975 ;
        RECT 69.510 32.685 69.775 33.145 ;
        RECT 69.945 32.550 70.195 32.975 ;
        RECT 70.405 32.700 71.510 32.870 ;
        RECT 69.890 32.420 70.195 32.550 ;
        RECT 69.440 31.225 69.720 32.175 ;
        RECT 69.890 31.315 70.060 32.420 ;
        RECT 70.230 31.635 70.470 32.230 ;
        RECT 70.640 32.165 71.170 32.530 ;
        RECT 70.640 31.465 70.810 32.165 ;
        RECT 71.340 32.085 71.510 32.700 ;
        RECT 71.680 32.345 71.850 33.145 ;
        RECT 72.020 32.645 72.270 32.975 ;
        RECT 72.495 32.675 73.380 32.845 ;
        RECT 71.340 31.995 71.850 32.085 ;
        RECT 69.890 31.185 70.115 31.315 ;
        RECT 70.285 31.245 70.810 31.465 ;
        RECT 70.980 31.825 71.850 31.995 ;
        RECT 69.525 30.595 69.775 31.055 ;
        RECT 69.945 31.045 70.115 31.185 ;
        RECT 70.980 31.045 71.150 31.825 ;
        RECT 71.680 31.755 71.850 31.825 ;
        RECT 71.360 31.575 71.560 31.605 ;
        RECT 72.020 31.575 72.190 32.645 ;
        RECT 72.360 31.755 72.550 32.475 ;
        RECT 71.360 31.275 72.190 31.575 ;
        RECT 72.720 31.545 73.040 32.505 ;
        RECT 69.945 30.875 70.280 31.045 ;
        RECT 70.475 30.875 71.150 31.045 ;
        RECT 71.470 30.595 71.840 31.095 ;
        RECT 72.020 31.045 72.190 31.275 ;
        RECT 72.575 31.215 73.040 31.545 ;
        RECT 73.210 31.835 73.380 32.675 ;
        RECT 73.560 32.645 73.875 33.145 ;
        RECT 74.105 32.415 74.445 32.975 ;
        RECT 73.550 32.040 74.445 32.415 ;
        RECT 74.615 32.135 74.785 33.145 ;
        RECT 74.255 31.835 74.445 32.040 ;
        RECT 74.955 32.085 75.285 32.930 ;
        RECT 74.955 32.005 75.345 32.085 ;
        RECT 75.130 31.955 75.345 32.005 ;
        RECT 76.435 31.980 76.725 33.145 ;
        RECT 77.540 32.175 77.930 32.350 ;
        RECT 78.415 32.345 78.745 33.145 ;
        RECT 78.915 32.355 79.450 32.975 ;
        RECT 79.655 32.710 85.000 33.145 ;
        RECT 77.540 32.005 78.965 32.175 ;
        RECT 73.210 31.505 74.085 31.835 ;
        RECT 74.255 31.505 75.005 31.835 ;
        RECT 73.210 31.045 73.380 31.505 ;
        RECT 74.255 31.335 74.455 31.505 ;
        RECT 75.175 31.375 75.345 31.955 ;
        RECT 75.120 31.335 75.345 31.375 ;
        RECT 72.020 30.875 72.425 31.045 ;
        RECT 72.595 30.875 73.380 31.045 ;
        RECT 73.655 30.595 73.865 31.125 ;
        RECT 74.125 30.810 74.455 31.335 ;
        RECT 74.965 31.250 75.345 31.335 ;
        RECT 74.625 30.595 74.795 31.205 ;
        RECT 74.965 30.815 75.295 31.250 ;
        RECT 76.435 30.595 76.725 31.320 ;
        RECT 77.415 31.275 77.770 31.835 ;
        RECT 77.940 31.105 78.110 32.005 ;
        RECT 78.280 31.275 78.545 31.835 ;
        RECT 78.795 31.505 78.965 32.005 ;
        RECT 79.135 31.335 79.450 32.355 ;
        RECT 77.520 30.595 77.760 31.105 ;
        RECT 77.940 30.775 78.220 31.105 ;
        RECT 78.450 30.595 78.665 31.105 ;
        RECT 78.835 30.765 79.450 31.335 ;
        RECT 81.240 31.140 81.580 31.970 ;
        RECT 83.060 31.460 83.410 32.710 ;
        RECT 85.175 32.055 86.845 33.145 ;
        RECT 85.175 31.365 85.925 31.885 ;
        RECT 86.095 31.535 86.845 32.055 ;
        RECT 87.565 32.215 87.735 32.975 ;
        RECT 87.950 32.385 88.280 33.145 ;
        RECT 87.565 32.045 88.280 32.215 ;
        RECT 88.450 32.070 88.705 32.975 ;
        RECT 87.475 31.495 87.830 31.865 ;
        RECT 88.110 31.835 88.280 32.045 ;
        RECT 88.110 31.505 88.365 31.835 ;
        RECT 79.655 30.595 85.000 31.140 ;
        RECT 85.175 30.595 86.845 31.365 ;
        RECT 88.110 31.315 88.280 31.505 ;
        RECT 88.535 31.340 88.705 32.070 ;
        RECT 88.880 31.995 89.140 33.145 ;
        RECT 89.315 32.055 90.525 33.145 ;
        RECT 89.315 31.515 89.835 32.055 ;
        RECT 87.565 31.145 88.280 31.315 ;
        RECT 87.565 30.765 87.735 31.145 ;
        RECT 87.950 30.595 88.280 30.975 ;
        RECT 88.450 30.765 88.705 31.340 ;
        RECT 88.880 30.595 89.140 31.435 ;
        RECT 90.005 31.345 90.525 31.885 ;
        RECT 89.315 30.595 90.525 31.345 ;
        RECT 11.950 30.425 90.610 30.595 ;
        RECT 12.035 29.675 13.245 30.425 ;
        RECT 12.035 29.135 12.555 29.675 ;
        RECT 13.875 29.625 14.215 30.255 ;
        RECT 14.385 29.625 14.635 30.425 ;
        RECT 14.825 29.775 15.155 30.255 ;
        RECT 15.325 29.965 15.550 30.425 ;
        RECT 15.720 29.775 16.050 30.255 ;
        RECT 12.725 28.965 13.245 29.505 ;
        RECT 12.035 27.875 13.245 28.965 ;
        RECT 13.875 29.015 14.050 29.625 ;
        RECT 14.825 29.605 16.050 29.775 ;
        RECT 16.680 29.645 17.180 30.255 ;
        RECT 17.645 29.875 17.815 30.165 ;
        RECT 17.985 30.045 18.315 30.425 ;
        RECT 17.645 29.705 18.310 29.875 ;
        RECT 14.220 29.265 14.915 29.435 ;
        RECT 14.745 29.015 14.915 29.265 ;
        RECT 15.090 29.235 15.510 29.435 ;
        RECT 15.680 29.235 16.010 29.435 ;
        RECT 16.180 29.235 16.510 29.435 ;
        RECT 16.680 29.015 16.850 29.645 ;
        RECT 17.035 29.185 17.385 29.435 ;
        RECT 13.875 28.045 14.215 29.015 ;
        RECT 14.385 27.875 14.555 29.015 ;
        RECT 14.745 28.845 17.180 29.015 ;
        RECT 17.560 28.885 17.910 29.535 ;
        RECT 14.825 27.875 15.075 28.675 ;
        RECT 15.720 28.045 16.050 28.845 ;
        RECT 16.350 27.875 16.680 28.675 ;
        RECT 16.850 28.045 17.180 28.845 ;
        RECT 18.080 28.715 18.310 29.705 ;
        RECT 17.645 28.545 18.310 28.715 ;
        RECT 17.645 28.045 17.815 28.545 ;
        RECT 17.985 27.875 18.315 28.375 ;
        RECT 18.485 28.045 18.670 30.165 ;
        RECT 18.925 29.965 19.175 30.425 ;
        RECT 19.345 29.975 19.680 30.145 ;
        RECT 19.875 29.975 20.550 30.145 ;
        RECT 19.345 29.835 19.515 29.975 ;
        RECT 18.840 28.845 19.120 29.795 ;
        RECT 19.290 29.705 19.515 29.835 ;
        RECT 19.290 28.600 19.460 29.705 ;
        RECT 19.685 29.555 20.210 29.775 ;
        RECT 19.630 28.790 19.870 29.385 ;
        RECT 20.040 28.855 20.210 29.555 ;
        RECT 20.380 29.195 20.550 29.975 ;
        RECT 20.870 29.925 21.240 30.425 ;
        RECT 21.420 29.975 21.825 30.145 ;
        RECT 21.995 29.975 22.780 30.145 ;
        RECT 21.420 29.745 21.590 29.975 ;
        RECT 20.760 29.445 21.590 29.745 ;
        RECT 21.975 29.475 22.440 29.805 ;
        RECT 20.760 29.415 20.960 29.445 ;
        RECT 21.080 29.195 21.250 29.265 ;
        RECT 20.380 29.025 21.250 29.195 ;
        RECT 20.740 28.935 21.250 29.025 ;
        RECT 19.290 28.470 19.595 28.600 ;
        RECT 20.040 28.490 20.570 28.855 ;
        RECT 18.910 27.875 19.175 28.335 ;
        RECT 19.345 28.045 19.595 28.470 ;
        RECT 20.740 28.320 20.910 28.935 ;
        RECT 19.805 28.150 20.910 28.320 ;
        RECT 21.080 27.875 21.250 28.675 ;
        RECT 21.420 28.375 21.590 29.445 ;
        RECT 21.760 28.545 21.950 29.265 ;
        RECT 22.120 28.515 22.440 29.475 ;
        RECT 22.610 29.515 22.780 29.975 ;
        RECT 23.055 29.895 23.265 30.425 ;
        RECT 23.525 29.685 23.855 30.210 ;
        RECT 24.025 29.815 24.195 30.425 ;
        RECT 24.365 29.770 24.695 30.205 ;
        RECT 24.365 29.685 24.745 29.770 ;
        RECT 23.655 29.515 23.855 29.685 ;
        RECT 24.520 29.645 24.745 29.685 ;
        RECT 22.610 29.185 23.485 29.515 ;
        RECT 23.655 29.185 24.405 29.515 ;
        RECT 21.420 28.045 21.670 28.375 ;
        RECT 22.610 28.345 22.780 29.185 ;
        RECT 23.655 28.980 23.845 29.185 ;
        RECT 24.575 29.065 24.745 29.645 ;
        RECT 24.530 29.015 24.745 29.065 ;
        RECT 22.950 28.605 23.845 28.980 ;
        RECT 24.355 28.935 24.745 29.015 ;
        RECT 24.950 29.685 25.565 30.255 ;
        RECT 25.735 29.915 25.950 30.425 ;
        RECT 26.180 29.915 26.460 30.245 ;
        RECT 26.640 29.915 26.880 30.425 ;
        RECT 21.895 28.175 22.780 28.345 ;
        RECT 22.960 27.875 23.275 28.375 ;
        RECT 23.505 28.045 23.845 28.605 ;
        RECT 24.015 27.875 24.185 28.885 ;
        RECT 24.355 28.090 24.685 28.935 ;
        RECT 24.950 28.665 25.265 29.685 ;
        RECT 25.435 29.015 25.605 29.515 ;
        RECT 25.855 29.185 26.120 29.745 ;
        RECT 26.290 29.015 26.460 29.915 ;
        RECT 26.630 29.185 26.985 29.745 ;
        RECT 27.675 29.625 28.015 30.255 ;
        RECT 28.185 29.625 28.435 30.425 ;
        RECT 28.625 29.775 28.955 30.255 ;
        RECT 29.125 29.965 29.350 30.425 ;
        RECT 29.520 29.775 29.850 30.255 ;
        RECT 27.675 29.015 27.850 29.625 ;
        RECT 28.625 29.605 29.850 29.775 ;
        RECT 30.480 29.645 30.980 30.255 ;
        RECT 32.020 29.645 32.520 30.255 ;
        RECT 28.020 29.265 28.715 29.435 ;
        RECT 28.545 29.015 28.715 29.265 ;
        RECT 28.890 29.235 29.310 29.435 ;
        RECT 29.480 29.235 29.810 29.435 ;
        RECT 29.980 29.235 30.310 29.435 ;
        RECT 30.480 29.015 30.650 29.645 ;
        RECT 30.835 29.185 31.185 29.435 ;
        RECT 31.815 29.185 32.165 29.435 ;
        RECT 32.350 29.015 32.520 29.645 ;
        RECT 33.150 29.775 33.480 30.255 ;
        RECT 33.650 29.965 33.875 30.425 ;
        RECT 34.045 29.775 34.375 30.255 ;
        RECT 33.150 29.605 34.375 29.775 ;
        RECT 34.565 29.625 34.815 30.425 ;
        RECT 34.985 29.625 35.325 30.255 ;
        RECT 35.660 29.915 35.900 30.425 ;
        RECT 36.080 29.915 36.360 30.245 ;
        RECT 36.590 29.915 36.805 30.425 ;
        RECT 32.690 29.235 33.020 29.435 ;
        RECT 33.190 29.235 33.520 29.435 ;
        RECT 33.690 29.235 34.110 29.435 ;
        RECT 34.285 29.265 34.980 29.435 ;
        RECT 34.285 29.015 34.455 29.265 ;
        RECT 35.150 29.015 35.325 29.625 ;
        RECT 35.555 29.185 35.910 29.745 ;
        RECT 36.080 29.015 36.250 29.915 ;
        RECT 36.420 29.185 36.685 29.745 ;
        RECT 36.975 29.685 37.590 30.255 ;
        RECT 37.795 29.700 38.085 30.425 ;
        RECT 36.935 29.015 37.105 29.515 ;
        RECT 25.435 28.845 26.860 29.015 ;
        RECT 24.950 28.045 25.485 28.665 ;
        RECT 25.655 27.875 25.985 28.675 ;
        RECT 26.470 28.670 26.860 28.845 ;
        RECT 27.675 28.045 28.015 29.015 ;
        RECT 28.185 27.875 28.355 29.015 ;
        RECT 28.545 28.845 30.980 29.015 ;
        RECT 28.625 27.875 28.875 28.675 ;
        RECT 29.520 28.045 29.850 28.845 ;
        RECT 30.150 27.875 30.480 28.675 ;
        RECT 30.650 28.045 30.980 28.845 ;
        RECT 32.020 28.845 34.455 29.015 ;
        RECT 32.020 28.045 32.350 28.845 ;
        RECT 32.520 27.875 32.850 28.675 ;
        RECT 33.150 28.045 33.480 28.845 ;
        RECT 34.125 27.875 34.375 28.675 ;
        RECT 34.645 27.875 34.815 29.015 ;
        RECT 34.985 28.045 35.325 29.015 ;
        RECT 35.680 28.845 37.105 29.015 ;
        RECT 35.680 28.670 36.070 28.845 ;
        RECT 36.555 27.875 36.885 28.675 ;
        RECT 37.275 28.665 37.590 29.685 ;
        RECT 38.255 29.655 40.845 30.425 ;
        RECT 41.105 29.875 41.275 30.165 ;
        RECT 41.445 30.045 41.775 30.425 ;
        RECT 41.105 29.705 41.770 29.875 ;
        RECT 38.255 29.135 39.465 29.655 ;
        RECT 37.055 28.045 37.590 28.665 ;
        RECT 37.795 27.875 38.085 29.040 ;
        RECT 39.635 28.965 40.845 29.485 ;
        RECT 38.255 27.875 40.845 28.965 ;
        RECT 41.020 28.885 41.370 29.535 ;
        RECT 41.540 28.715 41.770 29.705 ;
        RECT 41.105 28.545 41.770 28.715 ;
        RECT 41.105 28.045 41.275 28.545 ;
        RECT 41.445 27.875 41.775 28.375 ;
        RECT 41.945 28.045 42.130 30.165 ;
        RECT 42.385 29.965 42.635 30.425 ;
        RECT 42.805 29.975 43.140 30.145 ;
        RECT 43.335 29.975 44.010 30.145 ;
        RECT 42.805 29.835 42.975 29.975 ;
        RECT 42.300 28.845 42.580 29.795 ;
        RECT 42.750 29.705 42.975 29.835 ;
        RECT 42.750 28.600 42.920 29.705 ;
        RECT 43.145 29.555 43.670 29.775 ;
        RECT 43.090 28.790 43.330 29.385 ;
        RECT 43.500 28.855 43.670 29.555 ;
        RECT 43.840 29.195 44.010 29.975 ;
        RECT 44.330 29.925 44.700 30.425 ;
        RECT 44.880 29.975 45.285 30.145 ;
        RECT 45.455 29.975 46.240 30.145 ;
        RECT 44.880 29.745 45.050 29.975 ;
        RECT 44.220 29.445 45.050 29.745 ;
        RECT 45.435 29.475 45.900 29.805 ;
        RECT 44.220 29.415 44.420 29.445 ;
        RECT 44.540 29.195 44.710 29.265 ;
        RECT 43.840 29.025 44.710 29.195 ;
        RECT 44.200 28.935 44.710 29.025 ;
        RECT 42.750 28.470 43.055 28.600 ;
        RECT 43.500 28.490 44.030 28.855 ;
        RECT 42.370 27.875 42.635 28.335 ;
        RECT 42.805 28.045 43.055 28.470 ;
        RECT 44.200 28.320 44.370 28.935 ;
        RECT 43.265 28.150 44.370 28.320 ;
        RECT 44.540 27.875 44.710 28.675 ;
        RECT 44.880 28.375 45.050 29.445 ;
        RECT 45.220 28.545 45.410 29.265 ;
        RECT 45.580 28.515 45.900 29.475 ;
        RECT 46.070 29.515 46.240 29.975 ;
        RECT 46.515 29.895 46.725 30.425 ;
        RECT 46.985 29.685 47.315 30.210 ;
        RECT 47.485 29.815 47.655 30.425 ;
        RECT 47.825 29.770 48.155 30.205 ;
        RECT 47.825 29.685 48.205 29.770 ;
        RECT 47.115 29.515 47.315 29.685 ;
        RECT 47.980 29.645 48.205 29.685 ;
        RECT 46.070 29.185 46.945 29.515 ;
        RECT 47.115 29.185 47.865 29.515 ;
        RECT 44.880 28.045 45.130 28.375 ;
        RECT 46.070 28.345 46.240 29.185 ;
        RECT 47.115 28.980 47.305 29.185 ;
        RECT 48.035 29.065 48.205 29.645 ;
        RECT 48.375 29.675 49.585 30.425 ;
        RECT 49.845 29.875 50.015 30.165 ;
        RECT 50.185 30.045 50.515 30.425 ;
        RECT 49.845 29.705 50.510 29.875 ;
        RECT 48.375 29.135 48.895 29.675 ;
        RECT 47.990 29.015 48.205 29.065 ;
        RECT 46.410 28.605 47.305 28.980 ;
        RECT 47.815 28.935 48.205 29.015 ;
        RECT 49.065 28.965 49.585 29.505 ;
        RECT 45.355 28.175 46.240 28.345 ;
        RECT 46.420 27.875 46.735 28.375 ;
        RECT 46.965 28.045 47.305 28.605 ;
        RECT 47.475 27.875 47.645 28.885 ;
        RECT 47.815 28.090 48.145 28.935 ;
        RECT 48.375 27.875 49.585 28.965 ;
        RECT 49.760 28.885 50.110 29.535 ;
        RECT 50.280 28.715 50.510 29.705 ;
        RECT 49.845 28.545 50.510 28.715 ;
        RECT 49.845 28.045 50.015 28.545 ;
        RECT 50.185 27.875 50.515 28.375 ;
        RECT 50.685 28.045 50.870 30.165 ;
        RECT 51.125 29.965 51.375 30.425 ;
        RECT 51.545 29.975 51.880 30.145 ;
        RECT 52.075 29.975 52.750 30.145 ;
        RECT 51.545 29.835 51.715 29.975 ;
        RECT 51.040 28.845 51.320 29.795 ;
        RECT 51.490 29.705 51.715 29.835 ;
        RECT 51.490 28.600 51.660 29.705 ;
        RECT 51.885 29.555 52.410 29.775 ;
        RECT 51.830 28.790 52.070 29.385 ;
        RECT 52.240 28.855 52.410 29.555 ;
        RECT 52.580 29.195 52.750 29.975 ;
        RECT 53.070 29.925 53.440 30.425 ;
        RECT 53.620 29.975 54.025 30.145 ;
        RECT 54.195 29.975 54.980 30.145 ;
        RECT 53.620 29.745 53.790 29.975 ;
        RECT 52.960 29.445 53.790 29.745 ;
        RECT 54.175 29.475 54.640 29.805 ;
        RECT 52.960 29.415 53.160 29.445 ;
        RECT 53.280 29.195 53.450 29.265 ;
        RECT 52.580 29.025 53.450 29.195 ;
        RECT 52.940 28.935 53.450 29.025 ;
        RECT 51.490 28.470 51.795 28.600 ;
        RECT 52.240 28.490 52.770 28.855 ;
        RECT 51.110 27.875 51.375 28.335 ;
        RECT 51.545 28.045 51.795 28.470 ;
        RECT 52.940 28.320 53.110 28.935 ;
        RECT 52.005 28.150 53.110 28.320 ;
        RECT 53.280 27.875 53.450 28.675 ;
        RECT 53.620 28.375 53.790 29.445 ;
        RECT 53.960 28.545 54.150 29.265 ;
        RECT 54.320 28.515 54.640 29.475 ;
        RECT 54.810 29.515 54.980 29.975 ;
        RECT 55.255 29.895 55.465 30.425 ;
        RECT 55.725 29.685 56.055 30.210 ;
        RECT 56.225 29.815 56.395 30.425 ;
        RECT 56.565 29.770 56.895 30.205 ;
        RECT 56.565 29.685 56.945 29.770 ;
        RECT 55.855 29.515 56.055 29.685 ;
        RECT 56.720 29.645 56.945 29.685 ;
        RECT 54.810 29.185 55.685 29.515 ;
        RECT 55.855 29.185 56.605 29.515 ;
        RECT 53.620 28.045 53.870 28.375 ;
        RECT 54.810 28.345 54.980 29.185 ;
        RECT 55.855 28.980 56.045 29.185 ;
        RECT 56.775 29.065 56.945 29.645 ;
        RECT 56.730 29.015 56.945 29.065 ;
        RECT 55.150 28.605 56.045 28.980 ;
        RECT 56.555 28.935 56.945 29.015 ;
        RECT 57.575 29.625 57.915 30.255 ;
        RECT 58.085 29.625 58.335 30.425 ;
        RECT 58.525 29.775 58.855 30.255 ;
        RECT 59.025 29.965 59.250 30.425 ;
        RECT 59.420 29.775 59.750 30.255 ;
        RECT 57.575 29.015 57.750 29.625 ;
        RECT 58.525 29.605 59.750 29.775 ;
        RECT 60.380 29.645 60.880 30.255 ;
        RECT 61.290 29.685 61.905 30.255 ;
        RECT 62.075 29.915 62.290 30.425 ;
        RECT 62.520 29.915 62.800 30.245 ;
        RECT 62.980 29.915 63.220 30.425 ;
        RECT 57.920 29.265 58.615 29.435 ;
        RECT 58.445 29.015 58.615 29.265 ;
        RECT 58.790 29.235 59.210 29.435 ;
        RECT 59.380 29.235 59.710 29.435 ;
        RECT 59.880 29.235 60.210 29.435 ;
        RECT 60.380 29.015 60.550 29.645 ;
        RECT 60.735 29.185 61.085 29.435 ;
        RECT 54.095 28.175 54.980 28.345 ;
        RECT 55.160 27.875 55.475 28.375 ;
        RECT 55.705 28.045 56.045 28.605 ;
        RECT 56.215 27.875 56.385 28.885 ;
        RECT 56.555 28.090 56.885 28.935 ;
        RECT 57.575 28.045 57.915 29.015 ;
        RECT 58.085 27.875 58.255 29.015 ;
        RECT 58.445 28.845 60.880 29.015 ;
        RECT 58.525 27.875 58.775 28.675 ;
        RECT 59.420 28.045 59.750 28.845 ;
        RECT 60.050 27.875 60.380 28.675 ;
        RECT 60.550 28.045 60.880 28.845 ;
        RECT 61.290 28.665 61.605 29.685 ;
        RECT 61.775 29.015 61.945 29.515 ;
        RECT 62.195 29.185 62.460 29.745 ;
        RECT 62.630 29.015 62.800 29.915 ;
        RECT 62.970 29.185 63.325 29.745 ;
        RECT 63.555 29.700 63.845 30.425 ;
        RECT 64.935 29.925 65.195 30.255 ;
        RECT 65.365 30.065 65.695 30.425 ;
        RECT 65.950 30.045 67.250 30.255 ;
        RECT 64.935 29.915 65.165 29.925 ;
        RECT 61.775 28.845 63.200 29.015 ;
        RECT 61.290 28.045 61.825 28.665 ;
        RECT 61.995 27.875 62.325 28.675 ;
        RECT 62.810 28.670 63.200 28.845 ;
        RECT 63.555 27.875 63.845 29.040 ;
        RECT 64.935 28.725 65.105 29.915 ;
        RECT 65.950 29.895 66.120 30.045 ;
        RECT 65.365 29.770 66.120 29.895 ;
        RECT 65.275 29.725 66.120 29.770 ;
        RECT 65.275 29.605 65.545 29.725 ;
        RECT 65.275 29.030 65.445 29.605 ;
        RECT 65.675 29.165 66.085 29.470 ;
        RECT 66.375 29.435 66.585 29.835 ;
        RECT 66.255 29.225 66.585 29.435 ;
        RECT 66.830 29.435 67.050 29.835 ;
        RECT 67.525 29.660 67.980 30.425 ;
        RECT 68.360 29.645 68.860 30.255 ;
        RECT 66.830 29.225 67.305 29.435 ;
        RECT 67.495 29.235 67.985 29.435 ;
        RECT 68.155 29.185 68.505 29.435 ;
        RECT 65.275 28.995 65.475 29.030 ;
        RECT 66.805 28.995 67.980 29.055 ;
        RECT 68.690 29.015 68.860 29.645 ;
        RECT 69.490 29.775 69.820 30.255 ;
        RECT 69.990 29.965 70.215 30.425 ;
        RECT 70.385 29.775 70.715 30.255 ;
        RECT 69.490 29.605 70.715 29.775 ;
        RECT 70.905 29.625 71.155 30.425 ;
        RECT 71.325 29.625 71.665 30.255 ;
        RECT 69.030 29.235 69.360 29.435 ;
        RECT 69.530 29.235 69.860 29.435 ;
        RECT 70.030 29.235 70.450 29.435 ;
        RECT 70.625 29.265 71.320 29.435 ;
        RECT 70.625 29.015 70.795 29.265 ;
        RECT 71.490 29.015 71.665 29.625 ;
        RECT 71.835 29.655 73.505 30.425 ;
        RECT 74.225 29.875 74.395 30.165 ;
        RECT 74.565 30.045 74.895 30.425 ;
        RECT 74.225 29.705 74.890 29.875 ;
        RECT 71.835 29.135 72.585 29.655 ;
        RECT 65.275 28.885 67.980 28.995 ;
        RECT 65.335 28.825 67.135 28.885 ;
        RECT 66.805 28.795 67.135 28.825 ;
        RECT 64.935 28.045 65.195 28.725 ;
        RECT 65.365 27.875 65.615 28.655 ;
        RECT 65.865 28.625 66.700 28.635 ;
        RECT 67.290 28.625 67.475 28.715 ;
        RECT 65.865 28.425 67.475 28.625 ;
        RECT 65.865 28.045 66.115 28.425 ;
        RECT 67.245 28.385 67.475 28.425 ;
        RECT 67.725 28.265 67.980 28.885 ;
        RECT 66.285 27.875 66.640 28.255 ;
        RECT 67.645 28.045 67.980 28.265 ;
        RECT 68.360 28.845 70.795 29.015 ;
        RECT 68.360 28.045 68.690 28.845 ;
        RECT 68.860 27.875 69.190 28.675 ;
        RECT 69.490 28.045 69.820 28.845 ;
        RECT 70.465 27.875 70.715 28.675 ;
        RECT 70.985 27.875 71.155 29.015 ;
        RECT 71.325 28.045 71.665 29.015 ;
        RECT 72.755 28.965 73.505 29.485 ;
        RECT 71.835 27.875 73.505 28.965 ;
        RECT 74.140 28.885 74.490 29.535 ;
        RECT 74.660 28.715 74.890 29.705 ;
        RECT 74.225 28.545 74.890 28.715 ;
        RECT 74.225 28.045 74.395 28.545 ;
        RECT 74.565 27.875 74.895 28.375 ;
        RECT 75.065 28.045 75.250 30.165 ;
        RECT 75.505 29.965 75.755 30.425 ;
        RECT 75.925 29.975 76.260 30.145 ;
        RECT 76.455 29.975 77.130 30.145 ;
        RECT 75.925 29.835 76.095 29.975 ;
        RECT 75.420 28.845 75.700 29.795 ;
        RECT 75.870 29.705 76.095 29.835 ;
        RECT 75.870 28.600 76.040 29.705 ;
        RECT 76.265 29.555 76.790 29.775 ;
        RECT 76.210 28.790 76.450 29.385 ;
        RECT 76.620 28.855 76.790 29.555 ;
        RECT 76.960 29.195 77.130 29.975 ;
        RECT 77.450 29.925 77.820 30.425 ;
        RECT 78.000 29.975 78.405 30.145 ;
        RECT 78.575 29.975 79.360 30.145 ;
        RECT 78.000 29.745 78.170 29.975 ;
        RECT 77.340 29.445 78.170 29.745 ;
        RECT 78.555 29.475 79.020 29.805 ;
        RECT 77.340 29.415 77.540 29.445 ;
        RECT 77.660 29.195 77.830 29.265 ;
        RECT 76.960 29.025 77.830 29.195 ;
        RECT 77.320 28.935 77.830 29.025 ;
        RECT 75.870 28.470 76.175 28.600 ;
        RECT 76.620 28.490 77.150 28.855 ;
        RECT 75.490 27.875 75.755 28.335 ;
        RECT 75.925 28.045 76.175 28.470 ;
        RECT 77.320 28.320 77.490 28.935 ;
        RECT 76.385 28.150 77.490 28.320 ;
        RECT 77.660 27.875 77.830 28.675 ;
        RECT 78.000 28.375 78.170 29.445 ;
        RECT 78.340 28.545 78.530 29.265 ;
        RECT 78.700 28.515 79.020 29.475 ;
        RECT 79.190 29.515 79.360 29.975 ;
        RECT 79.635 29.895 79.845 30.425 ;
        RECT 80.105 29.685 80.435 30.210 ;
        RECT 80.605 29.815 80.775 30.425 ;
        RECT 80.945 29.770 81.275 30.205 ;
        RECT 81.495 29.925 81.755 30.255 ;
        RECT 81.925 30.065 82.255 30.425 ;
        RECT 82.510 30.045 83.810 30.255 ;
        RECT 80.945 29.685 81.325 29.770 ;
        RECT 80.235 29.515 80.435 29.685 ;
        RECT 81.100 29.645 81.325 29.685 ;
        RECT 79.190 29.185 80.065 29.515 ;
        RECT 80.235 29.185 80.985 29.515 ;
        RECT 78.000 28.045 78.250 28.375 ;
        RECT 79.190 28.345 79.360 29.185 ;
        RECT 80.235 28.980 80.425 29.185 ;
        RECT 81.155 29.065 81.325 29.645 ;
        RECT 81.110 29.015 81.325 29.065 ;
        RECT 79.530 28.605 80.425 28.980 ;
        RECT 80.935 28.935 81.325 29.015 ;
        RECT 78.475 28.175 79.360 28.345 ;
        RECT 79.540 27.875 79.855 28.375 ;
        RECT 80.085 28.045 80.425 28.605 ;
        RECT 80.595 27.875 80.765 28.885 ;
        RECT 80.935 28.090 81.265 28.935 ;
        RECT 81.495 28.725 81.665 29.925 ;
        RECT 82.510 29.895 82.680 30.045 ;
        RECT 81.925 29.770 82.680 29.895 ;
        RECT 81.835 29.725 82.680 29.770 ;
        RECT 81.835 29.605 82.105 29.725 ;
        RECT 81.835 29.030 82.005 29.605 ;
        RECT 82.235 29.165 82.645 29.470 ;
        RECT 82.935 29.435 83.145 29.835 ;
        RECT 82.815 29.225 83.145 29.435 ;
        RECT 83.390 29.435 83.610 29.835 ;
        RECT 84.085 29.660 84.540 30.425 ;
        RECT 84.715 29.655 88.225 30.425 ;
        RECT 89.315 29.675 90.525 30.425 ;
        RECT 83.390 29.225 83.865 29.435 ;
        RECT 84.055 29.235 84.545 29.435 ;
        RECT 84.715 29.135 86.365 29.655 ;
        RECT 81.835 28.995 82.035 29.030 ;
        RECT 83.365 28.995 84.540 29.055 ;
        RECT 81.835 28.885 84.540 28.995 ;
        RECT 86.535 28.965 88.225 29.485 ;
        RECT 81.895 28.825 83.695 28.885 ;
        RECT 83.365 28.795 83.695 28.825 ;
        RECT 81.495 28.045 81.755 28.725 ;
        RECT 81.925 27.875 82.175 28.655 ;
        RECT 82.425 28.625 83.260 28.635 ;
        RECT 83.850 28.625 84.035 28.715 ;
        RECT 82.425 28.425 84.035 28.625 ;
        RECT 82.425 28.045 82.675 28.425 ;
        RECT 83.805 28.385 84.035 28.425 ;
        RECT 84.285 28.265 84.540 28.885 ;
        RECT 82.845 27.875 83.200 28.255 ;
        RECT 84.205 28.045 84.540 28.265 ;
        RECT 84.715 27.875 88.225 28.965 ;
        RECT 89.315 28.965 89.835 29.505 ;
        RECT 90.005 29.135 90.525 29.675 ;
        RECT 89.315 27.875 90.525 28.965 ;
        RECT 11.950 27.705 90.610 27.875 ;
        RECT 12.035 26.615 13.245 27.705 ;
        RECT 13.505 27.035 13.675 27.535 ;
        RECT 13.845 27.205 14.175 27.705 ;
        RECT 13.505 26.865 14.170 27.035 ;
        RECT 12.035 25.905 12.555 26.445 ;
        RECT 12.725 26.075 13.245 26.615 ;
        RECT 13.420 26.045 13.770 26.695 ;
        RECT 12.035 25.155 13.245 25.905 ;
        RECT 13.940 25.875 14.170 26.865 ;
        RECT 13.505 25.705 14.170 25.875 ;
        RECT 13.505 25.415 13.675 25.705 ;
        RECT 13.845 25.155 14.175 25.535 ;
        RECT 14.345 25.415 14.530 27.535 ;
        RECT 14.770 27.245 15.035 27.705 ;
        RECT 15.205 27.110 15.455 27.535 ;
        RECT 15.665 27.260 16.770 27.430 ;
        RECT 15.150 26.980 15.455 27.110 ;
        RECT 14.700 25.785 14.980 26.735 ;
        RECT 15.150 25.875 15.320 26.980 ;
        RECT 15.490 26.195 15.730 26.790 ;
        RECT 15.900 26.725 16.430 27.090 ;
        RECT 15.900 26.025 16.070 26.725 ;
        RECT 16.600 26.645 16.770 27.260 ;
        RECT 16.940 26.905 17.110 27.705 ;
        RECT 17.280 27.205 17.530 27.535 ;
        RECT 17.755 27.235 18.640 27.405 ;
        RECT 16.600 26.555 17.110 26.645 ;
        RECT 15.150 25.745 15.375 25.875 ;
        RECT 15.545 25.805 16.070 26.025 ;
        RECT 16.240 26.385 17.110 26.555 ;
        RECT 14.785 25.155 15.035 25.615 ;
        RECT 15.205 25.605 15.375 25.745 ;
        RECT 16.240 25.605 16.410 26.385 ;
        RECT 16.940 26.315 17.110 26.385 ;
        RECT 16.620 26.135 16.820 26.165 ;
        RECT 17.280 26.135 17.450 27.205 ;
        RECT 17.620 26.315 17.810 27.035 ;
        RECT 16.620 25.835 17.450 26.135 ;
        RECT 17.980 26.105 18.300 27.065 ;
        RECT 15.205 25.435 15.540 25.605 ;
        RECT 15.735 25.435 16.410 25.605 ;
        RECT 16.730 25.155 17.100 25.655 ;
        RECT 17.280 25.605 17.450 25.835 ;
        RECT 17.835 25.775 18.300 26.105 ;
        RECT 18.470 26.395 18.640 27.235 ;
        RECT 18.820 27.205 19.135 27.705 ;
        RECT 19.365 26.975 19.705 27.535 ;
        RECT 18.810 26.600 19.705 26.975 ;
        RECT 19.875 26.695 20.045 27.705 ;
        RECT 19.515 26.395 19.705 26.600 ;
        RECT 20.215 26.645 20.545 27.490 ;
        RECT 20.780 27.315 21.115 27.535 ;
        RECT 22.120 27.325 22.475 27.705 ;
        RECT 20.780 26.695 21.035 27.315 ;
        RECT 21.285 27.155 21.515 27.195 ;
        RECT 22.645 27.155 22.895 27.535 ;
        RECT 21.285 26.955 22.895 27.155 ;
        RECT 21.285 26.865 21.470 26.955 ;
        RECT 22.060 26.945 22.895 26.955 ;
        RECT 23.145 26.925 23.395 27.705 ;
        RECT 23.565 26.855 23.825 27.535 ;
        RECT 21.625 26.755 21.955 26.785 ;
        RECT 21.625 26.695 23.425 26.755 ;
        RECT 20.215 26.565 20.605 26.645 ;
        RECT 20.390 26.515 20.605 26.565 ;
        RECT 20.780 26.585 23.485 26.695 ;
        RECT 20.780 26.525 21.955 26.585 ;
        RECT 23.285 26.550 23.485 26.585 ;
        RECT 18.470 26.065 19.345 26.395 ;
        RECT 19.515 26.065 20.265 26.395 ;
        RECT 18.470 25.605 18.640 26.065 ;
        RECT 19.515 25.895 19.715 26.065 ;
        RECT 20.435 25.935 20.605 26.515 ;
        RECT 20.775 26.145 21.265 26.345 ;
        RECT 21.455 26.145 21.930 26.355 ;
        RECT 20.380 25.895 20.605 25.935 ;
        RECT 17.280 25.435 17.685 25.605 ;
        RECT 17.855 25.435 18.640 25.605 ;
        RECT 18.915 25.155 19.125 25.685 ;
        RECT 19.385 25.370 19.715 25.895 ;
        RECT 20.225 25.810 20.605 25.895 ;
        RECT 19.885 25.155 20.055 25.765 ;
        RECT 20.225 25.375 20.555 25.810 ;
        RECT 20.780 25.155 21.235 25.920 ;
        RECT 21.710 25.745 21.930 26.145 ;
        RECT 22.175 26.145 22.505 26.355 ;
        RECT 22.175 25.745 22.385 26.145 ;
        RECT 22.675 26.110 23.085 26.415 ;
        RECT 23.315 25.975 23.485 26.550 ;
        RECT 23.215 25.855 23.485 25.975 ;
        RECT 22.640 25.810 23.485 25.855 ;
        RECT 22.640 25.685 23.395 25.810 ;
        RECT 22.640 25.535 22.810 25.685 ;
        RECT 23.655 25.655 23.825 26.855 ;
        RECT 24.915 26.540 25.205 27.705 ;
        RECT 25.375 26.615 26.585 27.705 ;
        RECT 26.845 27.035 27.015 27.535 ;
        RECT 27.185 27.205 27.515 27.705 ;
        RECT 26.845 26.865 27.510 27.035 ;
        RECT 25.375 25.905 25.895 26.445 ;
        RECT 26.065 26.075 26.585 26.615 ;
        RECT 26.760 26.045 27.110 26.695 ;
        RECT 21.510 25.325 22.810 25.535 ;
        RECT 23.065 25.155 23.395 25.515 ;
        RECT 23.565 25.325 23.825 25.655 ;
        RECT 24.915 25.155 25.205 25.880 ;
        RECT 25.375 25.155 26.585 25.905 ;
        RECT 27.280 25.875 27.510 26.865 ;
        RECT 26.845 25.705 27.510 25.875 ;
        RECT 26.845 25.415 27.015 25.705 ;
        RECT 27.185 25.155 27.515 25.535 ;
        RECT 27.685 25.415 27.870 27.535 ;
        RECT 28.110 27.245 28.375 27.705 ;
        RECT 28.545 27.110 28.795 27.535 ;
        RECT 29.005 27.260 30.110 27.430 ;
        RECT 28.490 26.980 28.795 27.110 ;
        RECT 28.040 25.785 28.320 26.735 ;
        RECT 28.490 25.875 28.660 26.980 ;
        RECT 28.830 26.195 29.070 26.790 ;
        RECT 29.240 26.725 29.770 27.090 ;
        RECT 29.240 26.025 29.410 26.725 ;
        RECT 29.940 26.645 30.110 27.260 ;
        RECT 30.280 26.905 30.450 27.705 ;
        RECT 30.620 27.205 30.870 27.535 ;
        RECT 31.095 27.235 31.980 27.405 ;
        RECT 29.940 26.555 30.450 26.645 ;
        RECT 28.490 25.745 28.715 25.875 ;
        RECT 28.885 25.805 29.410 26.025 ;
        RECT 29.580 26.385 30.450 26.555 ;
        RECT 28.125 25.155 28.375 25.615 ;
        RECT 28.545 25.605 28.715 25.745 ;
        RECT 29.580 25.605 29.750 26.385 ;
        RECT 30.280 26.315 30.450 26.385 ;
        RECT 29.960 26.135 30.160 26.165 ;
        RECT 30.620 26.135 30.790 27.205 ;
        RECT 30.960 26.315 31.150 27.035 ;
        RECT 29.960 25.835 30.790 26.135 ;
        RECT 31.320 26.105 31.640 27.065 ;
        RECT 28.545 25.435 28.880 25.605 ;
        RECT 29.075 25.435 29.750 25.605 ;
        RECT 30.070 25.155 30.440 25.655 ;
        RECT 30.620 25.605 30.790 25.835 ;
        RECT 31.175 25.775 31.640 26.105 ;
        RECT 31.810 26.395 31.980 27.235 ;
        RECT 32.160 27.205 32.475 27.705 ;
        RECT 32.705 26.975 33.045 27.535 ;
        RECT 32.150 26.600 33.045 26.975 ;
        RECT 33.215 26.695 33.385 27.705 ;
        RECT 32.855 26.395 33.045 26.600 ;
        RECT 33.555 26.645 33.885 27.490 ;
        RECT 34.205 27.035 34.375 27.535 ;
        RECT 34.545 27.205 34.875 27.705 ;
        RECT 34.205 26.865 34.870 27.035 ;
        RECT 33.555 26.565 33.945 26.645 ;
        RECT 33.730 26.515 33.945 26.565 ;
        RECT 31.810 26.065 32.685 26.395 ;
        RECT 32.855 26.065 33.605 26.395 ;
        RECT 31.810 25.605 31.980 26.065 ;
        RECT 32.855 25.895 33.055 26.065 ;
        RECT 33.775 25.935 33.945 26.515 ;
        RECT 34.120 26.045 34.470 26.695 ;
        RECT 33.720 25.895 33.945 25.935 ;
        RECT 30.620 25.435 31.025 25.605 ;
        RECT 31.195 25.435 31.980 25.605 ;
        RECT 32.255 25.155 32.465 25.685 ;
        RECT 32.725 25.370 33.055 25.895 ;
        RECT 33.565 25.810 33.945 25.895 ;
        RECT 34.640 25.875 34.870 26.865 ;
        RECT 33.225 25.155 33.395 25.765 ;
        RECT 33.565 25.375 33.895 25.810 ;
        RECT 34.205 25.705 34.870 25.875 ;
        RECT 34.205 25.415 34.375 25.705 ;
        RECT 34.545 25.155 34.875 25.535 ;
        RECT 35.045 25.415 35.230 27.535 ;
        RECT 35.470 27.245 35.735 27.705 ;
        RECT 35.905 27.110 36.155 27.535 ;
        RECT 36.365 27.260 37.470 27.430 ;
        RECT 35.850 26.980 36.155 27.110 ;
        RECT 35.400 25.785 35.680 26.735 ;
        RECT 35.850 25.875 36.020 26.980 ;
        RECT 36.190 26.195 36.430 26.790 ;
        RECT 36.600 26.725 37.130 27.090 ;
        RECT 36.600 26.025 36.770 26.725 ;
        RECT 37.300 26.645 37.470 27.260 ;
        RECT 37.640 26.905 37.810 27.705 ;
        RECT 37.980 27.205 38.230 27.535 ;
        RECT 38.455 27.235 39.340 27.405 ;
        RECT 37.300 26.555 37.810 26.645 ;
        RECT 35.850 25.745 36.075 25.875 ;
        RECT 36.245 25.805 36.770 26.025 ;
        RECT 36.940 26.385 37.810 26.555 ;
        RECT 35.485 25.155 35.735 25.615 ;
        RECT 35.905 25.605 36.075 25.745 ;
        RECT 36.940 25.605 37.110 26.385 ;
        RECT 37.640 26.315 37.810 26.385 ;
        RECT 37.320 26.135 37.520 26.165 ;
        RECT 37.980 26.135 38.150 27.205 ;
        RECT 38.320 26.315 38.510 27.035 ;
        RECT 37.320 25.835 38.150 26.135 ;
        RECT 38.680 26.105 39.000 27.065 ;
        RECT 35.905 25.435 36.240 25.605 ;
        RECT 36.435 25.435 37.110 25.605 ;
        RECT 37.430 25.155 37.800 25.655 ;
        RECT 37.980 25.605 38.150 25.835 ;
        RECT 38.535 25.775 39.000 26.105 ;
        RECT 39.170 26.395 39.340 27.235 ;
        RECT 39.520 27.205 39.835 27.705 ;
        RECT 40.065 26.975 40.405 27.535 ;
        RECT 39.510 26.600 40.405 26.975 ;
        RECT 40.575 26.695 40.745 27.705 ;
        RECT 40.215 26.395 40.405 26.600 ;
        RECT 40.915 26.645 41.245 27.490 ;
        RECT 40.915 26.565 41.305 26.645 ;
        RECT 41.090 26.515 41.305 26.565 ;
        RECT 39.170 26.065 40.045 26.395 ;
        RECT 40.215 26.065 40.965 26.395 ;
        RECT 39.170 25.605 39.340 26.065 ;
        RECT 40.215 25.895 40.415 26.065 ;
        RECT 41.135 25.935 41.305 26.515 ;
        RECT 41.080 25.895 41.305 25.935 ;
        RECT 37.980 25.435 38.385 25.605 ;
        RECT 38.555 25.435 39.340 25.605 ;
        RECT 39.615 25.155 39.825 25.685 ;
        RECT 40.085 25.370 40.415 25.895 ;
        RECT 40.925 25.810 41.305 25.895 ;
        RECT 42.395 26.565 42.735 27.535 ;
        RECT 42.905 26.565 43.075 27.705 ;
        RECT 43.345 26.905 43.595 27.705 ;
        RECT 44.240 26.735 44.570 27.535 ;
        RECT 44.870 26.905 45.200 27.705 ;
        RECT 45.370 26.735 45.700 27.535 ;
        RECT 43.265 26.565 45.700 26.735 ;
        RECT 46.075 26.615 47.745 27.705 ;
        RECT 42.395 25.955 42.570 26.565 ;
        RECT 43.265 26.315 43.435 26.565 ;
        RECT 42.740 26.145 43.435 26.315 ;
        RECT 43.610 26.145 44.030 26.345 ;
        RECT 44.200 26.145 44.530 26.345 ;
        RECT 44.700 26.145 45.030 26.345 ;
        RECT 40.585 25.155 40.755 25.765 ;
        RECT 40.925 25.375 41.255 25.810 ;
        RECT 42.395 25.325 42.735 25.955 ;
        RECT 42.905 25.155 43.155 25.955 ;
        RECT 43.345 25.805 44.570 25.975 ;
        RECT 43.345 25.325 43.675 25.805 ;
        RECT 43.845 25.155 44.070 25.615 ;
        RECT 44.240 25.325 44.570 25.805 ;
        RECT 45.200 25.935 45.370 26.565 ;
        RECT 45.555 26.145 45.905 26.395 ;
        RECT 45.200 25.325 45.700 25.935 ;
        RECT 46.075 25.925 46.825 26.445 ;
        RECT 46.995 26.095 47.745 26.615 ;
        RECT 48.560 26.735 48.950 26.910 ;
        RECT 49.435 26.905 49.765 27.705 ;
        RECT 49.935 26.915 50.470 27.535 ;
        RECT 48.560 26.565 49.985 26.735 ;
        RECT 46.075 25.155 47.745 25.925 ;
        RECT 48.435 25.835 48.790 26.395 ;
        RECT 48.960 25.665 49.130 26.565 ;
        RECT 49.300 25.835 49.565 26.395 ;
        RECT 49.815 26.065 49.985 26.565 ;
        RECT 50.155 25.895 50.470 26.915 ;
        RECT 50.675 26.540 50.965 27.705 ;
        RECT 51.135 26.565 51.475 27.535 ;
        RECT 51.645 26.565 51.815 27.705 ;
        RECT 52.085 26.905 52.335 27.705 ;
        RECT 52.980 26.735 53.310 27.535 ;
        RECT 53.610 26.905 53.940 27.705 ;
        RECT 54.110 26.735 54.440 27.535 ;
        RECT 52.005 26.565 54.440 26.735 ;
        RECT 54.815 26.615 56.485 27.705 ;
        RECT 48.540 25.155 48.780 25.665 ;
        RECT 48.960 25.335 49.240 25.665 ;
        RECT 49.470 25.155 49.685 25.665 ;
        RECT 49.855 25.325 50.470 25.895 ;
        RECT 51.135 25.955 51.310 26.565 ;
        RECT 52.005 26.315 52.175 26.565 ;
        RECT 51.480 26.145 52.175 26.315 ;
        RECT 52.350 26.145 52.770 26.345 ;
        RECT 52.940 26.145 53.270 26.345 ;
        RECT 53.440 26.145 53.770 26.345 ;
        RECT 50.675 25.155 50.965 25.880 ;
        RECT 51.135 25.325 51.475 25.955 ;
        RECT 51.645 25.155 51.895 25.955 ;
        RECT 52.085 25.805 53.310 25.975 ;
        RECT 52.085 25.325 52.415 25.805 ;
        RECT 52.585 25.155 52.810 25.615 ;
        RECT 52.980 25.325 53.310 25.805 ;
        RECT 53.940 25.935 54.110 26.565 ;
        RECT 54.295 26.145 54.645 26.395 ;
        RECT 53.940 25.325 54.440 25.935 ;
        RECT 54.815 25.925 55.565 26.445 ;
        RECT 55.735 26.095 56.485 26.615 ;
        RECT 56.660 26.555 56.920 27.705 ;
        RECT 57.095 26.630 57.350 27.535 ;
        RECT 57.520 26.945 57.850 27.705 ;
        RECT 58.065 26.775 58.235 27.535 ;
        RECT 58.495 27.270 63.840 27.705 ;
        RECT 64.015 27.270 69.360 27.705 ;
        RECT 54.815 25.155 56.485 25.925 ;
        RECT 56.660 25.155 56.920 25.995 ;
        RECT 57.095 25.900 57.265 26.630 ;
        RECT 57.520 26.605 58.235 26.775 ;
        RECT 57.520 26.395 57.690 26.605 ;
        RECT 57.435 26.065 57.690 26.395 ;
        RECT 57.095 25.325 57.350 25.900 ;
        RECT 57.520 25.875 57.690 26.065 ;
        RECT 57.970 26.055 58.325 26.425 ;
        RECT 57.520 25.705 58.235 25.875 ;
        RECT 57.520 25.155 57.850 25.535 ;
        RECT 58.065 25.325 58.235 25.705 ;
        RECT 60.080 25.700 60.420 26.530 ;
        RECT 61.900 26.020 62.250 27.270 ;
        RECT 65.600 25.700 65.940 26.530 ;
        RECT 67.420 26.020 67.770 27.270 ;
        RECT 69.535 26.615 73.045 27.705 ;
        RECT 69.535 25.925 71.185 26.445 ;
        RECT 71.355 26.095 73.045 26.615 ;
        RECT 74.320 26.735 74.710 26.910 ;
        RECT 75.195 26.905 75.525 27.705 ;
        RECT 75.695 26.915 76.230 27.535 ;
        RECT 74.320 26.565 75.745 26.735 ;
        RECT 58.495 25.155 63.840 25.700 ;
        RECT 64.015 25.155 69.360 25.700 ;
        RECT 69.535 25.155 73.045 25.925 ;
        RECT 74.195 25.835 74.550 26.395 ;
        RECT 74.720 25.665 74.890 26.565 ;
        RECT 75.060 25.835 75.325 26.395 ;
        RECT 75.575 26.065 75.745 26.565 ;
        RECT 75.915 25.895 76.230 26.915 ;
        RECT 76.435 26.540 76.725 27.705 ;
        RECT 76.895 26.565 77.235 27.535 ;
        RECT 77.405 26.565 77.575 27.705 ;
        RECT 77.845 26.905 78.095 27.705 ;
        RECT 78.740 26.735 79.070 27.535 ;
        RECT 79.370 26.905 79.700 27.705 ;
        RECT 79.870 26.735 80.200 27.535 ;
        RECT 77.765 26.565 80.200 26.735 ;
        RECT 80.575 26.615 81.785 27.705 ;
        RECT 82.045 27.035 82.215 27.535 ;
        RECT 82.385 27.205 82.715 27.705 ;
        RECT 82.045 26.865 82.710 27.035 ;
        RECT 74.300 25.155 74.540 25.665 ;
        RECT 74.720 25.335 75.000 25.665 ;
        RECT 75.230 25.155 75.445 25.665 ;
        RECT 75.615 25.325 76.230 25.895 ;
        RECT 76.895 25.955 77.070 26.565 ;
        RECT 77.765 26.315 77.935 26.565 ;
        RECT 77.240 26.145 77.935 26.315 ;
        RECT 78.110 26.145 78.530 26.345 ;
        RECT 78.700 26.145 79.030 26.345 ;
        RECT 79.200 26.145 79.530 26.345 ;
        RECT 76.435 25.155 76.725 25.880 ;
        RECT 76.895 25.325 77.235 25.955 ;
        RECT 77.405 25.155 77.655 25.955 ;
        RECT 77.845 25.805 79.070 25.975 ;
        RECT 77.845 25.325 78.175 25.805 ;
        RECT 78.345 25.155 78.570 25.615 ;
        RECT 78.740 25.325 79.070 25.805 ;
        RECT 79.700 25.935 79.870 26.565 ;
        RECT 80.055 26.145 80.405 26.395 ;
        RECT 79.700 25.325 80.200 25.935 ;
        RECT 80.575 25.905 81.095 26.445 ;
        RECT 81.265 26.075 81.785 26.615 ;
        RECT 81.960 26.045 82.310 26.695 ;
        RECT 80.575 25.155 81.785 25.905 ;
        RECT 82.480 25.875 82.710 26.865 ;
        RECT 82.045 25.705 82.710 25.875 ;
        RECT 82.045 25.415 82.215 25.705 ;
        RECT 82.385 25.155 82.715 25.535 ;
        RECT 82.885 25.415 83.070 27.535 ;
        RECT 83.310 27.245 83.575 27.705 ;
        RECT 83.745 27.110 83.995 27.535 ;
        RECT 84.205 27.260 85.310 27.430 ;
        RECT 83.690 26.980 83.995 27.110 ;
        RECT 83.240 25.785 83.520 26.735 ;
        RECT 83.690 25.875 83.860 26.980 ;
        RECT 84.030 26.195 84.270 26.790 ;
        RECT 84.440 26.725 84.970 27.090 ;
        RECT 84.440 26.025 84.610 26.725 ;
        RECT 85.140 26.645 85.310 27.260 ;
        RECT 85.480 26.905 85.650 27.705 ;
        RECT 85.820 27.205 86.070 27.535 ;
        RECT 86.295 27.235 87.180 27.405 ;
        RECT 85.140 26.555 85.650 26.645 ;
        RECT 83.690 25.745 83.915 25.875 ;
        RECT 84.085 25.805 84.610 26.025 ;
        RECT 84.780 26.385 85.650 26.555 ;
        RECT 83.325 25.155 83.575 25.615 ;
        RECT 83.745 25.605 83.915 25.745 ;
        RECT 84.780 25.605 84.950 26.385 ;
        RECT 85.480 26.315 85.650 26.385 ;
        RECT 85.160 26.135 85.360 26.165 ;
        RECT 85.820 26.135 85.990 27.205 ;
        RECT 86.160 26.315 86.350 27.035 ;
        RECT 85.160 25.835 85.990 26.135 ;
        RECT 86.520 26.105 86.840 27.065 ;
        RECT 83.745 25.435 84.080 25.605 ;
        RECT 84.275 25.435 84.950 25.605 ;
        RECT 85.270 25.155 85.640 25.655 ;
        RECT 85.820 25.605 85.990 25.835 ;
        RECT 86.375 25.775 86.840 26.105 ;
        RECT 87.010 26.395 87.180 27.235 ;
        RECT 87.360 27.205 87.675 27.705 ;
        RECT 87.905 26.975 88.245 27.535 ;
        RECT 87.350 26.600 88.245 26.975 ;
        RECT 88.415 26.695 88.585 27.705 ;
        RECT 88.055 26.395 88.245 26.600 ;
        RECT 88.755 26.645 89.085 27.490 ;
        RECT 88.755 26.565 89.145 26.645 ;
        RECT 88.930 26.515 89.145 26.565 ;
        RECT 87.010 26.065 87.885 26.395 ;
        RECT 88.055 26.065 88.805 26.395 ;
        RECT 87.010 25.605 87.180 26.065 ;
        RECT 88.055 25.895 88.255 26.065 ;
        RECT 88.975 25.935 89.145 26.515 ;
        RECT 89.315 26.615 90.525 27.705 ;
        RECT 89.315 26.075 89.835 26.615 ;
        RECT 88.920 25.895 89.145 25.935 ;
        RECT 90.005 25.905 90.525 26.445 ;
        RECT 85.820 25.435 86.225 25.605 ;
        RECT 86.395 25.435 87.180 25.605 ;
        RECT 87.455 25.155 87.665 25.685 ;
        RECT 87.925 25.370 88.255 25.895 ;
        RECT 88.765 25.810 89.145 25.895 ;
        RECT 88.425 25.155 88.595 25.765 ;
        RECT 88.765 25.375 89.095 25.810 ;
        RECT 89.315 25.155 90.525 25.905 ;
        RECT 11.950 24.985 90.610 25.155 ;
        RECT 12.035 24.235 13.245 24.985 ;
        RECT 12.035 23.695 12.555 24.235 ;
        RECT 13.420 24.145 13.680 24.985 ;
        RECT 13.855 24.240 14.110 24.815 ;
        RECT 14.280 24.605 14.610 24.985 ;
        RECT 14.825 24.435 14.995 24.815 ;
        RECT 14.280 24.265 14.995 24.435 ;
        RECT 12.725 23.525 13.245 24.065 ;
        RECT 12.035 22.435 13.245 23.525 ;
        RECT 13.420 22.435 13.680 23.585 ;
        RECT 13.855 23.510 14.025 24.240 ;
        RECT 14.280 24.075 14.450 24.265 ;
        RECT 15.255 24.235 16.465 24.985 ;
        RECT 14.195 23.745 14.450 24.075 ;
        RECT 14.280 23.535 14.450 23.745 ;
        RECT 14.730 23.715 15.085 24.085 ;
        RECT 15.255 23.695 15.775 24.235 ;
        RECT 16.640 24.145 16.900 24.985 ;
        RECT 17.075 24.240 17.330 24.815 ;
        RECT 17.500 24.605 17.830 24.985 ;
        RECT 18.045 24.435 18.215 24.815 ;
        RECT 17.500 24.265 18.215 24.435 ;
        RECT 13.855 22.605 14.110 23.510 ;
        RECT 14.280 23.365 14.995 23.535 ;
        RECT 15.945 23.525 16.465 24.065 ;
        RECT 14.280 22.435 14.610 23.195 ;
        RECT 14.825 22.605 14.995 23.365 ;
        RECT 15.255 22.435 16.465 23.525 ;
        RECT 16.640 22.435 16.900 23.585 ;
        RECT 17.075 23.510 17.245 24.240 ;
        RECT 17.500 24.075 17.670 24.265 ;
        RECT 18.480 24.145 18.740 24.985 ;
        RECT 18.915 24.240 19.170 24.815 ;
        RECT 19.340 24.605 19.670 24.985 ;
        RECT 19.885 24.435 20.055 24.815 ;
        RECT 19.340 24.265 20.055 24.435 ;
        RECT 17.415 23.745 17.670 24.075 ;
        RECT 17.500 23.535 17.670 23.745 ;
        RECT 17.950 23.715 18.305 24.085 ;
        RECT 17.075 22.605 17.330 23.510 ;
        RECT 17.500 23.365 18.215 23.535 ;
        RECT 17.500 22.435 17.830 23.195 ;
        RECT 18.045 22.605 18.215 23.365 ;
        RECT 18.480 22.435 18.740 23.585 ;
        RECT 18.915 23.510 19.085 24.240 ;
        RECT 19.340 24.075 19.510 24.265 ;
        RECT 21.240 24.220 21.695 24.985 ;
        RECT 21.970 24.605 23.270 24.815 ;
        RECT 23.525 24.625 23.855 24.985 ;
        RECT 23.100 24.455 23.270 24.605 ;
        RECT 24.025 24.485 24.285 24.815 ;
        RECT 19.255 23.745 19.510 24.075 ;
        RECT 19.340 23.535 19.510 23.745 ;
        RECT 19.790 23.715 20.145 24.085 ;
        RECT 22.170 23.995 22.390 24.395 ;
        RECT 21.235 23.795 21.725 23.995 ;
        RECT 21.915 23.785 22.390 23.995 ;
        RECT 22.635 23.995 22.845 24.395 ;
        RECT 23.100 24.330 23.855 24.455 ;
        RECT 23.100 24.285 23.945 24.330 ;
        RECT 23.675 24.165 23.945 24.285 ;
        RECT 22.635 23.785 22.965 23.995 ;
        RECT 23.135 23.725 23.545 24.030 ;
        RECT 21.240 23.555 22.415 23.615 ;
        RECT 23.775 23.590 23.945 24.165 ;
        RECT 23.745 23.555 23.945 23.590 ;
        RECT 18.915 22.605 19.170 23.510 ;
        RECT 19.340 23.365 20.055 23.535 ;
        RECT 19.340 22.435 19.670 23.195 ;
        RECT 19.885 22.605 20.055 23.365 ;
        RECT 21.240 23.445 23.945 23.555 ;
        RECT 21.240 22.825 21.495 23.445 ;
        RECT 22.085 23.385 23.885 23.445 ;
        RECT 22.085 23.355 22.415 23.385 ;
        RECT 24.115 23.285 24.285 24.485 ;
        RECT 24.545 24.435 24.715 24.815 ;
        RECT 24.930 24.605 25.260 24.985 ;
        RECT 24.545 24.265 25.260 24.435 ;
        RECT 24.455 23.715 24.810 24.085 ;
        RECT 25.090 24.075 25.260 24.265 ;
        RECT 25.430 24.240 25.685 24.815 ;
        RECT 25.090 23.745 25.345 24.075 ;
        RECT 25.090 23.535 25.260 23.745 ;
        RECT 21.745 23.185 21.930 23.275 ;
        RECT 22.520 23.185 23.355 23.195 ;
        RECT 21.745 22.985 23.355 23.185 ;
        RECT 21.745 22.945 21.975 22.985 ;
        RECT 21.240 22.605 21.575 22.825 ;
        RECT 22.580 22.435 22.935 22.815 ;
        RECT 23.105 22.605 23.355 22.985 ;
        RECT 23.605 22.435 23.855 23.215 ;
        RECT 24.025 22.605 24.285 23.285 ;
        RECT 24.545 23.365 25.260 23.535 ;
        RECT 25.515 23.510 25.685 24.240 ;
        RECT 25.860 24.145 26.120 24.985 ;
        RECT 27.380 24.475 27.620 24.985 ;
        RECT 27.800 24.475 28.080 24.805 ;
        RECT 28.310 24.475 28.525 24.985 ;
        RECT 27.275 23.745 27.630 24.305 ;
        RECT 24.545 22.605 24.715 23.365 ;
        RECT 24.930 22.435 25.260 23.195 ;
        RECT 25.430 22.605 25.685 23.510 ;
        RECT 25.860 22.435 26.120 23.585 ;
        RECT 27.800 23.575 27.970 24.475 ;
        RECT 28.140 23.745 28.405 24.305 ;
        RECT 28.695 24.245 29.310 24.815 ;
        RECT 29.515 24.440 34.860 24.985 ;
        RECT 28.655 23.575 28.825 24.075 ;
        RECT 27.400 23.405 28.825 23.575 ;
        RECT 27.400 23.230 27.790 23.405 ;
        RECT 28.275 22.435 28.605 23.235 ;
        RECT 28.995 23.225 29.310 24.245 ;
        RECT 31.100 23.610 31.440 24.440 ;
        RECT 35.035 24.215 37.625 24.985 ;
        RECT 37.795 24.260 38.085 24.985 ;
        RECT 38.255 24.215 39.925 24.985 ;
        RECT 40.100 24.220 40.555 24.985 ;
        RECT 40.830 24.605 42.130 24.815 ;
        RECT 42.385 24.625 42.715 24.985 ;
        RECT 41.960 24.455 42.130 24.605 ;
        RECT 42.885 24.485 43.145 24.815 ;
        RECT 28.775 22.605 29.310 23.225 ;
        RECT 32.920 22.870 33.270 24.120 ;
        RECT 35.035 23.695 36.245 24.215 ;
        RECT 36.415 23.525 37.625 24.045 ;
        RECT 38.255 23.695 39.005 24.215 ;
        RECT 29.515 22.435 34.860 22.870 ;
        RECT 35.035 22.435 37.625 23.525 ;
        RECT 37.795 22.435 38.085 23.600 ;
        RECT 39.175 23.525 39.925 24.045 ;
        RECT 41.030 23.995 41.250 24.395 ;
        RECT 40.095 23.795 40.585 23.995 ;
        RECT 40.775 23.785 41.250 23.995 ;
        RECT 41.495 23.995 41.705 24.395 ;
        RECT 41.960 24.330 42.715 24.455 ;
        RECT 41.960 24.285 42.805 24.330 ;
        RECT 42.535 24.165 42.805 24.285 ;
        RECT 41.495 23.785 41.825 23.995 ;
        RECT 41.995 23.725 42.405 24.030 ;
        RECT 38.255 22.435 39.925 23.525 ;
        RECT 40.100 23.555 41.275 23.615 ;
        RECT 42.635 23.590 42.805 24.165 ;
        RECT 42.605 23.555 42.805 23.590 ;
        RECT 40.100 23.445 42.805 23.555 ;
        RECT 40.100 22.825 40.355 23.445 ;
        RECT 40.945 23.385 42.745 23.445 ;
        RECT 40.945 23.355 41.275 23.385 ;
        RECT 42.975 23.285 43.145 24.485 ;
        RECT 43.315 24.235 44.525 24.985 ;
        RECT 43.315 23.695 43.835 24.235 ;
        RECT 44.700 24.220 45.155 24.985 ;
        RECT 45.430 24.605 46.730 24.815 ;
        RECT 46.985 24.625 47.315 24.985 ;
        RECT 46.560 24.455 46.730 24.605 ;
        RECT 47.485 24.485 47.745 24.815 ;
        RECT 44.005 23.525 44.525 24.065 ;
        RECT 45.630 23.995 45.850 24.395 ;
        RECT 44.695 23.795 45.185 23.995 ;
        RECT 45.375 23.785 45.850 23.995 ;
        RECT 46.095 23.995 46.305 24.395 ;
        RECT 46.560 24.330 47.315 24.455 ;
        RECT 46.560 24.285 47.405 24.330 ;
        RECT 47.135 24.165 47.405 24.285 ;
        RECT 46.095 23.785 46.425 23.995 ;
        RECT 46.595 23.725 47.005 24.030 ;
        RECT 40.605 23.185 40.790 23.275 ;
        RECT 41.380 23.185 42.215 23.195 ;
        RECT 40.605 22.985 42.215 23.185 ;
        RECT 40.605 22.945 40.835 22.985 ;
        RECT 40.100 22.605 40.435 22.825 ;
        RECT 41.440 22.435 41.795 22.815 ;
        RECT 41.965 22.605 42.215 22.985 ;
        RECT 42.465 22.435 42.715 23.215 ;
        RECT 42.885 22.605 43.145 23.285 ;
        RECT 43.315 22.435 44.525 23.525 ;
        RECT 44.700 23.555 45.875 23.615 ;
        RECT 47.235 23.590 47.405 24.165 ;
        RECT 47.205 23.555 47.405 23.590 ;
        RECT 44.700 23.445 47.405 23.555 ;
        RECT 44.700 22.825 44.955 23.445 ;
        RECT 45.545 23.385 47.345 23.445 ;
        RECT 45.545 23.355 45.875 23.385 ;
        RECT 47.575 23.285 47.745 24.485 ;
        RECT 47.915 24.440 53.260 24.985 ;
        RECT 49.500 23.610 49.840 24.440 ;
        RECT 53.435 24.215 56.945 24.985 ;
        RECT 45.205 23.185 45.390 23.275 ;
        RECT 45.980 23.185 46.815 23.195 ;
        RECT 45.205 22.985 46.815 23.185 ;
        RECT 45.205 22.945 45.435 22.985 ;
        RECT 44.700 22.605 45.035 22.825 ;
        RECT 46.040 22.435 46.395 22.815 ;
        RECT 46.565 22.605 46.815 22.985 ;
        RECT 47.065 22.435 47.315 23.215 ;
        RECT 47.485 22.605 47.745 23.285 ;
        RECT 51.320 22.870 51.670 24.120 ;
        RECT 53.435 23.695 55.085 24.215 ;
        RECT 57.575 24.185 57.915 24.815 ;
        RECT 58.085 24.185 58.335 24.985 ;
        RECT 58.525 24.335 58.855 24.815 ;
        RECT 59.025 24.525 59.250 24.985 ;
        RECT 59.420 24.335 59.750 24.815 ;
        RECT 55.255 23.525 56.945 24.045 ;
        RECT 47.915 22.435 53.260 22.870 ;
        RECT 53.435 22.435 56.945 23.525 ;
        RECT 57.575 23.575 57.750 24.185 ;
        RECT 58.525 24.165 59.750 24.335 ;
        RECT 60.380 24.205 60.880 24.815 ;
        RECT 61.290 24.245 61.905 24.815 ;
        RECT 62.075 24.475 62.290 24.985 ;
        RECT 62.520 24.475 62.800 24.805 ;
        RECT 62.980 24.475 63.220 24.985 ;
        RECT 57.920 23.825 58.615 23.995 ;
        RECT 58.445 23.575 58.615 23.825 ;
        RECT 58.790 23.795 59.210 23.995 ;
        RECT 59.380 23.795 59.710 23.995 ;
        RECT 59.880 23.795 60.210 23.995 ;
        RECT 60.380 23.575 60.550 24.205 ;
        RECT 60.735 23.745 61.085 23.995 ;
        RECT 57.575 22.605 57.915 23.575 ;
        RECT 58.085 22.435 58.255 23.575 ;
        RECT 58.445 23.405 60.880 23.575 ;
        RECT 58.525 22.435 58.775 23.235 ;
        RECT 59.420 22.605 59.750 23.405 ;
        RECT 60.050 22.435 60.380 23.235 ;
        RECT 60.550 22.605 60.880 23.405 ;
        RECT 61.290 23.225 61.605 24.245 ;
        RECT 61.775 23.575 61.945 24.075 ;
        RECT 62.195 23.745 62.460 24.305 ;
        RECT 62.630 23.575 62.800 24.475 ;
        RECT 62.970 23.745 63.325 24.305 ;
        RECT 63.555 24.260 63.845 24.985 ;
        RECT 64.015 24.485 64.275 24.815 ;
        RECT 64.445 24.625 64.775 24.985 ;
        RECT 65.030 24.605 66.330 24.815 ;
        RECT 61.775 23.405 63.200 23.575 ;
        RECT 61.290 22.605 61.825 23.225 ;
        RECT 61.995 22.435 62.325 23.235 ;
        RECT 62.810 23.230 63.200 23.405 ;
        RECT 63.555 22.435 63.845 23.600 ;
        RECT 64.015 23.285 64.185 24.485 ;
        RECT 65.030 24.455 65.200 24.605 ;
        RECT 64.445 24.330 65.200 24.455 ;
        RECT 64.355 24.285 65.200 24.330 ;
        RECT 64.355 24.165 64.625 24.285 ;
        RECT 64.355 23.590 64.525 24.165 ;
        RECT 64.755 23.725 65.165 24.030 ;
        RECT 65.455 23.995 65.665 24.395 ;
        RECT 65.335 23.785 65.665 23.995 ;
        RECT 65.910 23.995 66.130 24.395 ;
        RECT 66.605 24.220 67.060 24.985 ;
        RECT 67.235 24.185 67.575 24.815 ;
        RECT 67.745 24.185 67.995 24.985 ;
        RECT 68.185 24.335 68.515 24.815 ;
        RECT 68.685 24.525 68.910 24.985 ;
        RECT 69.080 24.335 69.410 24.815 ;
        RECT 65.910 23.785 66.385 23.995 ;
        RECT 66.575 23.795 67.065 23.995 ;
        RECT 64.355 23.555 64.555 23.590 ;
        RECT 65.885 23.555 67.060 23.615 ;
        RECT 64.355 23.445 67.060 23.555 ;
        RECT 64.415 23.385 66.215 23.445 ;
        RECT 65.885 23.355 66.215 23.385 ;
        RECT 64.015 22.605 64.275 23.285 ;
        RECT 64.445 22.435 64.695 23.215 ;
        RECT 64.945 23.185 65.780 23.195 ;
        RECT 66.370 23.185 66.555 23.275 ;
        RECT 64.945 22.985 66.555 23.185 ;
        RECT 64.945 22.605 65.195 22.985 ;
        RECT 66.325 22.945 66.555 22.985 ;
        RECT 66.805 22.825 67.060 23.445 ;
        RECT 65.365 22.435 65.720 22.815 ;
        RECT 66.725 22.605 67.060 22.825 ;
        RECT 67.235 23.575 67.410 24.185 ;
        RECT 68.185 24.165 69.410 24.335 ;
        RECT 70.040 24.205 70.540 24.815 ;
        RECT 70.950 24.245 71.565 24.815 ;
        RECT 71.735 24.475 71.950 24.985 ;
        RECT 72.180 24.475 72.460 24.805 ;
        RECT 72.640 24.475 72.880 24.985 ;
        RECT 67.580 23.825 68.275 23.995 ;
        RECT 68.105 23.575 68.275 23.825 ;
        RECT 68.450 23.795 68.870 23.995 ;
        RECT 69.040 23.795 69.370 23.995 ;
        RECT 69.540 23.795 69.870 23.995 ;
        RECT 70.040 23.575 70.210 24.205 ;
        RECT 70.395 23.745 70.745 23.995 ;
        RECT 67.235 22.605 67.575 23.575 ;
        RECT 67.745 22.435 67.915 23.575 ;
        RECT 68.105 23.405 70.540 23.575 ;
        RECT 68.185 22.435 68.435 23.235 ;
        RECT 69.080 22.605 69.410 23.405 ;
        RECT 69.710 22.435 70.040 23.235 ;
        RECT 70.210 22.605 70.540 23.405 ;
        RECT 70.950 23.225 71.265 24.245 ;
        RECT 71.435 23.575 71.605 24.075 ;
        RECT 71.855 23.745 72.120 24.305 ;
        RECT 72.290 23.575 72.460 24.475 ;
        RECT 72.630 23.745 72.985 24.305 ;
        RECT 73.215 24.215 74.885 24.985 ;
        RECT 75.515 24.485 75.775 24.815 ;
        RECT 75.945 24.625 76.275 24.985 ;
        RECT 76.530 24.605 77.830 24.815 ;
        RECT 73.215 23.695 73.965 24.215 ;
        RECT 71.435 23.405 72.860 23.575 ;
        RECT 74.135 23.525 74.885 24.045 ;
        RECT 70.950 22.605 71.485 23.225 ;
        RECT 71.655 22.435 71.985 23.235 ;
        RECT 72.470 23.230 72.860 23.405 ;
        RECT 73.215 22.435 74.885 23.525 ;
        RECT 75.515 23.285 75.685 24.485 ;
        RECT 76.530 24.455 76.700 24.605 ;
        RECT 75.945 24.330 76.700 24.455 ;
        RECT 75.855 24.285 76.700 24.330 ;
        RECT 75.855 24.165 76.125 24.285 ;
        RECT 75.855 23.590 76.025 24.165 ;
        RECT 76.255 23.725 76.665 24.030 ;
        RECT 76.955 23.995 77.165 24.395 ;
        RECT 76.835 23.785 77.165 23.995 ;
        RECT 77.410 23.995 77.630 24.395 ;
        RECT 78.105 24.220 78.560 24.985 ;
        RECT 78.940 24.205 79.440 24.815 ;
        RECT 77.410 23.785 77.885 23.995 ;
        RECT 78.075 23.795 78.565 23.995 ;
        RECT 78.735 23.745 79.085 23.995 ;
        RECT 75.855 23.555 76.055 23.590 ;
        RECT 77.385 23.555 78.560 23.615 ;
        RECT 79.270 23.575 79.440 24.205 ;
        RECT 80.070 24.335 80.400 24.815 ;
        RECT 80.570 24.525 80.795 24.985 ;
        RECT 80.965 24.335 81.295 24.815 ;
        RECT 80.070 24.165 81.295 24.335 ;
        RECT 81.485 24.185 81.735 24.985 ;
        RECT 81.905 24.185 82.245 24.815 ;
        RECT 79.610 23.795 79.940 23.995 ;
        RECT 80.110 23.795 80.440 23.995 ;
        RECT 80.610 23.795 81.030 23.995 ;
        RECT 81.205 23.825 81.900 23.995 ;
        RECT 81.205 23.575 81.375 23.825 ;
        RECT 82.070 23.625 82.245 24.185 ;
        RECT 82.415 24.235 83.625 24.985 ;
        RECT 83.885 24.435 84.055 24.815 ;
        RECT 84.270 24.605 84.600 24.985 ;
        RECT 83.885 24.265 84.600 24.435 ;
        RECT 82.415 23.695 82.935 24.235 ;
        RECT 82.015 23.575 82.245 23.625 ;
        RECT 75.855 23.445 78.560 23.555 ;
        RECT 75.915 23.385 77.715 23.445 ;
        RECT 77.385 23.355 77.715 23.385 ;
        RECT 75.515 22.605 75.775 23.285 ;
        RECT 75.945 22.435 76.195 23.215 ;
        RECT 76.445 23.185 77.280 23.195 ;
        RECT 77.870 23.185 78.055 23.275 ;
        RECT 76.445 22.985 78.055 23.185 ;
        RECT 76.445 22.605 76.695 22.985 ;
        RECT 77.825 22.945 78.055 22.985 ;
        RECT 78.305 22.825 78.560 23.445 ;
        RECT 76.865 22.435 77.220 22.815 ;
        RECT 78.225 22.605 78.560 22.825 ;
        RECT 78.940 23.405 81.375 23.575 ;
        RECT 78.940 22.605 79.270 23.405 ;
        RECT 79.440 22.435 79.770 23.235 ;
        RECT 80.070 22.605 80.400 23.405 ;
        RECT 81.045 22.435 81.295 23.235 ;
        RECT 81.565 22.435 81.735 23.575 ;
        RECT 81.905 22.605 82.245 23.575 ;
        RECT 83.105 23.525 83.625 24.065 ;
        RECT 83.795 23.715 84.150 24.085 ;
        RECT 84.430 24.075 84.600 24.265 ;
        RECT 84.770 24.240 85.025 24.815 ;
        RECT 84.430 23.745 84.685 24.075 ;
        RECT 84.430 23.535 84.600 23.745 ;
        RECT 82.415 22.435 83.625 23.525 ;
        RECT 83.885 23.365 84.600 23.535 ;
        RECT 84.855 23.510 85.025 24.240 ;
        RECT 85.200 24.145 85.460 24.985 ;
        RECT 85.725 24.435 85.895 24.815 ;
        RECT 86.110 24.605 86.440 24.985 ;
        RECT 85.725 24.265 86.440 24.435 ;
        RECT 85.635 23.715 85.990 24.085 ;
        RECT 86.270 24.075 86.440 24.265 ;
        RECT 86.610 24.240 86.865 24.815 ;
        RECT 86.270 23.745 86.525 24.075 ;
        RECT 83.885 22.605 84.055 23.365 ;
        RECT 84.270 22.435 84.600 23.195 ;
        RECT 84.770 22.605 85.025 23.510 ;
        RECT 85.200 22.435 85.460 23.585 ;
        RECT 86.270 23.535 86.440 23.745 ;
        RECT 85.725 23.365 86.440 23.535 ;
        RECT 86.695 23.510 86.865 24.240 ;
        RECT 87.040 24.145 87.300 24.985 ;
        RECT 87.480 24.145 87.740 24.985 ;
        RECT 87.915 24.240 88.170 24.815 ;
        RECT 88.340 24.605 88.670 24.985 ;
        RECT 88.885 24.435 89.055 24.815 ;
        RECT 88.340 24.265 89.055 24.435 ;
        RECT 85.725 22.605 85.895 23.365 ;
        RECT 86.110 22.435 86.440 23.195 ;
        RECT 86.610 22.605 86.865 23.510 ;
        RECT 87.040 22.435 87.300 23.585 ;
        RECT 87.480 22.435 87.740 23.585 ;
        RECT 87.915 23.510 88.085 24.240 ;
        RECT 88.340 24.075 88.510 24.265 ;
        RECT 89.315 24.235 90.525 24.985 ;
        RECT 88.255 23.745 88.510 24.075 ;
        RECT 88.340 23.535 88.510 23.745 ;
        RECT 88.790 23.715 89.145 24.085 ;
        RECT 87.915 22.605 88.170 23.510 ;
        RECT 88.340 23.365 89.055 23.535 ;
        RECT 88.340 22.435 88.670 23.195 ;
        RECT 88.885 22.605 89.055 23.365 ;
        RECT 89.315 23.525 89.835 24.065 ;
        RECT 90.005 23.695 90.525 24.235 ;
        RECT 89.315 22.435 90.525 23.525 ;
        RECT 11.950 22.265 90.610 22.435 ;
        RECT 12.035 21.175 13.245 22.265 ;
        RECT 12.035 20.465 12.555 21.005 ;
        RECT 12.725 20.635 13.245 21.175 ;
        RECT 13.875 21.125 14.215 22.095 ;
        RECT 14.385 21.125 14.555 22.265 ;
        RECT 14.825 21.465 15.075 22.265 ;
        RECT 15.720 21.295 16.050 22.095 ;
        RECT 16.350 21.465 16.680 22.265 ;
        RECT 16.850 21.295 17.180 22.095 ;
        RECT 14.745 21.125 17.180 21.295 ;
        RECT 13.875 20.515 14.050 21.125 ;
        RECT 14.745 20.875 14.915 21.125 ;
        RECT 14.220 20.705 14.915 20.875 ;
        RECT 15.090 20.705 15.510 20.905 ;
        RECT 15.680 20.705 16.010 20.905 ;
        RECT 16.180 20.705 16.510 20.905 ;
        RECT 12.035 19.715 13.245 20.465 ;
        RECT 13.875 19.885 14.215 20.515 ;
        RECT 14.385 19.715 14.635 20.515 ;
        RECT 14.825 20.365 16.050 20.535 ;
        RECT 14.825 19.885 15.155 20.365 ;
        RECT 15.325 19.715 15.550 20.175 ;
        RECT 15.720 19.885 16.050 20.365 ;
        RECT 16.680 20.495 16.850 21.125 ;
        RECT 18.480 21.115 18.740 22.265 ;
        RECT 18.915 21.190 19.170 22.095 ;
        RECT 19.340 21.505 19.670 22.265 ;
        RECT 19.885 21.335 20.055 22.095 ;
        RECT 17.035 20.705 17.385 20.955 ;
        RECT 16.680 19.885 17.180 20.495 ;
        RECT 18.480 19.715 18.740 20.555 ;
        RECT 18.915 20.460 19.085 21.190 ;
        RECT 19.340 21.165 20.055 21.335 ;
        RECT 19.340 20.955 19.510 21.165 ;
        RECT 20.315 21.125 20.655 22.095 ;
        RECT 20.825 21.125 20.995 22.265 ;
        RECT 21.265 21.465 21.515 22.265 ;
        RECT 22.160 21.295 22.490 22.095 ;
        RECT 22.790 21.465 23.120 22.265 ;
        RECT 23.290 21.295 23.620 22.095 ;
        RECT 21.185 21.125 23.620 21.295 ;
        RECT 19.255 20.625 19.510 20.955 ;
        RECT 18.915 19.885 19.170 20.460 ;
        RECT 19.340 20.435 19.510 20.625 ;
        RECT 19.790 20.615 20.145 20.985 ;
        RECT 20.315 20.515 20.490 21.125 ;
        RECT 21.185 20.875 21.355 21.125 ;
        RECT 20.660 20.705 21.355 20.875 ;
        RECT 21.530 20.705 21.950 20.905 ;
        RECT 22.120 20.705 22.450 20.905 ;
        RECT 22.620 20.705 22.950 20.905 ;
        RECT 19.340 20.265 20.055 20.435 ;
        RECT 19.340 19.715 19.670 20.095 ;
        RECT 19.885 19.885 20.055 20.265 ;
        RECT 20.315 19.885 20.655 20.515 ;
        RECT 20.825 19.715 21.075 20.515 ;
        RECT 21.265 20.365 22.490 20.535 ;
        RECT 21.265 19.885 21.595 20.365 ;
        RECT 21.765 19.715 21.990 20.175 ;
        RECT 22.160 19.885 22.490 20.365 ;
        RECT 23.120 20.495 23.290 21.125 ;
        RECT 24.915 21.100 25.205 22.265 ;
        RECT 26.040 21.295 26.370 22.095 ;
        RECT 26.540 21.465 26.870 22.265 ;
        RECT 27.170 21.295 27.500 22.095 ;
        RECT 28.145 21.465 28.395 22.265 ;
        RECT 26.040 21.125 28.475 21.295 ;
        RECT 28.665 21.125 28.835 22.265 ;
        RECT 29.005 21.125 29.345 22.095 ;
        RECT 29.720 21.295 30.050 22.095 ;
        RECT 30.220 21.465 30.550 22.265 ;
        RECT 30.850 21.295 31.180 22.095 ;
        RECT 31.825 21.465 32.075 22.265 ;
        RECT 29.720 21.125 32.155 21.295 ;
        RECT 32.345 21.125 32.515 22.265 ;
        RECT 32.685 21.125 33.025 22.095 ;
        RECT 33.285 21.595 33.455 22.095 ;
        RECT 33.625 21.765 33.955 22.265 ;
        RECT 33.285 21.425 33.950 21.595 ;
        RECT 23.475 20.705 23.825 20.955 ;
        RECT 25.835 20.705 26.185 20.955 ;
        RECT 26.370 20.495 26.540 21.125 ;
        RECT 26.710 20.705 27.040 20.905 ;
        RECT 27.210 20.705 27.540 20.905 ;
        RECT 27.710 20.705 28.130 20.905 ;
        RECT 28.305 20.875 28.475 21.125 ;
        RECT 28.305 20.705 29.000 20.875 ;
        RECT 23.120 19.885 23.620 20.495 ;
        RECT 24.915 19.715 25.205 20.440 ;
        RECT 26.040 19.885 26.540 20.495 ;
        RECT 27.170 20.365 28.395 20.535 ;
        RECT 29.170 20.515 29.345 21.125 ;
        RECT 29.515 20.705 29.865 20.955 ;
        RECT 27.170 19.885 27.500 20.365 ;
        RECT 27.670 19.715 27.895 20.175 ;
        RECT 28.065 19.885 28.395 20.365 ;
        RECT 28.585 19.715 28.835 20.515 ;
        RECT 29.005 19.885 29.345 20.515 ;
        RECT 30.050 20.495 30.220 21.125 ;
        RECT 30.390 20.705 30.720 20.905 ;
        RECT 30.890 20.705 31.220 20.905 ;
        RECT 31.390 20.705 31.810 20.905 ;
        RECT 31.985 20.875 32.155 21.125 ;
        RECT 31.985 20.705 32.680 20.875 ;
        RECT 32.850 20.565 33.025 21.125 ;
        RECT 33.200 20.605 33.550 21.255 ;
        RECT 29.720 19.885 30.220 20.495 ;
        RECT 30.850 20.365 32.075 20.535 ;
        RECT 32.795 20.515 33.025 20.565 ;
        RECT 30.850 19.885 31.180 20.365 ;
        RECT 31.350 19.715 31.575 20.175 ;
        RECT 31.745 19.885 32.075 20.365 ;
        RECT 32.265 19.715 32.515 20.515 ;
        RECT 32.685 19.885 33.025 20.515 ;
        RECT 33.720 20.435 33.950 21.425 ;
        RECT 33.285 20.265 33.950 20.435 ;
        RECT 33.285 19.975 33.455 20.265 ;
        RECT 33.625 19.715 33.955 20.095 ;
        RECT 34.125 19.975 34.310 22.095 ;
        RECT 34.550 21.805 34.815 22.265 ;
        RECT 34.985 21.670 35.235 22.095 ;
        RECT 35.445 21.820 36.550 21.990 ;
        RECT 34.930 21.540 35.235 21.670 ;
        RECT 34.480 20.345 34.760 21.295 ;
        RECT 34.930 20.435 35.100 21.540 ;
        RECT 35.270 20.755 35.510 21.350 ;
        RECT 35.680 21.285 36.210 21.650 ;
        RECT 35.680 20.585 35.850 21.285 ;
        RECT 36.380 21.205 36.550 21.820 ;
        RECT 36.720 21.465 36.890 22.265 ;
        RECT 37.060 21.765 37.310 22.095 ;
        RECT 37.535 21.795 38.420 21.965 ;
        RECT 36.380 21.115 36.890 21.205 ;
        RECT 34.930 20.305 35.155 20.435 ;
        RECT 35.325 20.365 35.850 20.585 ;
        RECT 36.020 20.945 36.890 21.115 ;
        RECT 34.565 19.715 34.815 20.175 ;
        RECT 34.985 20.165 35.155 20.305 ;
        RECT 36.020 20.165 36.190 20.945 ;
        RECT 36.720 20.875 36.890 20.945 ;
        RECT 36.400 20.695 36.600 20.725 ;
        RECT 37.060 20.695 37.230 21.765 ;
        RECT 37.400 20.875 37.590 21.595 ;
        RECT 36.400 20.395 37.230 20.695 ;
        RECT 37.760 20.665 38.080 21.625 ;
        RECT 34.985 19.995 35.320 20.165 ;
        RECT 35.515 19.995 36.190 20.165 ;
        RECT 36.510 19.715 36.880 20.215 ;
        RECT 37.060 20.165 37.230 20.395 ;
        RECT 37.615 20.335 38.080 20.665 ;
        RECT 38.250 20.955 38.420 21.795 ;
        RECT 38.600 21.765 38.915 22.265 ;
        RECT 39.145 21.535 39.485 22.095 ;
        RECT 38.590 21.160 39.485 21.535 ;
        RECT 39.655 21.255 39.825 22.265 ;
        RECT 39.295 20.955 39.485 21.160 ;
        RECT 39.995 21.205 40.325 22.050 ;
        RECT 39.995 21.125 40.385 21.205 ;
        RECT 40.170 21.075 40.385 21.125 ;
        RECT 38.250 20.625 39.125 20.955 ;
        RECT 39.295 20.625 40.045 20.955 ;
        RECT 38.250 20.165 38.420 20.625 ;
        RECT 39.295 20.455 39.495 20.625 ;
        RECT 40.215 20.495 40.385 21.075 ;
        RECT 40.160 20.455 40.385 20.495 ;
        RECT 37.060 19.995 37.465 20.165 ;
        RECT 37.635 19.995 38.420 20.165 ;
        RECT 38.695 19.715 38.905 20.245 ;
        RECT 39.165 19.930 39.495 20.455 ;
        RECT 40.005 20.370 40.385 20.455 ;
        RECT 41.475 21.125 41.815 22.095 ;
        RECT 41.985 21.125 42.155 22.265 ;
        RECT 42.425 21.465 42.675 22.265 ;
        RECT 43.320 21.295 43.650 22.095 ;
        RECT 43.950 21.465 44.280 22.265 ;
        RECT 44.450 21.295 44.780 22.095 ;
        RECT 42.345 21.125 44.780 21.295 ;
        RECT 45.155 21.175 46.825 22.265 ;
        RECT 41.475 20.515 41.650 21.125 ;
        RECT 42.345 20.875 42.515 21.125 ;
        RECT 41.820 20.705 42.515 20.875 ;
        RECT 42.690 20.705 43.110 20.905 ;
        RECT 43.280 20.705 43.610 20.905 ;
        RECT 43.780 20.705 44.110 20.905 ;
        RECT 39.665 19.715 39.835 20.325 ;
        RECT 40.005 19.935 40.335 20.370 ;
        RECT 41.475 19.885 41.815 20.515 ;
        RECT 41.985 19.715 42.235 20.515 ;
        RECT 42.425 20.365 43.650 20.535 ;
        RECT 42.425 19.885 42.755 20.365 ;
        RECT 42.925 19.715 43.150 20.175 ;
        RECT 43.320 19.885 43.650 20.365 ;
        RECT 44.280 20.495 44.450 21.125 ;
        RECT 44.635 20.705 44.985 20.955 ;
        RECT 44.280 19.885 44.780 20.495 ;
        RECT 45.155 20.485 45.905 21.005 ;
        RECT 46.075 20.655 46.825 21.175 ;
        RECT 46.995 21.125 47.335 22.095 ;
        RECT 47.505 21.125 47.675 22.265 ;
        RECT 47.945 21.465 48.195 22.265 ;
        RECT 48.840 21.295 49.170 22.095 ;
        RECT 49.470 21.465 49.800 22.265 ;
        RECT 49.970 21.295 50.300 22.095 ;
        RECT 47.865 21.125 50.300 21.295 ;
        RECT 46.995 20.515 47.170 21.125 ;
        RECT 47.865 20.875 48.035 21.125 ;
        RECT 47.340 20.705 48.035 20.875 ;
        RECT 48.210 20.705 48.630 20.905 ;
        RECT 48.800 20.705 49.130 20.905 ;
        RECT 49.300 20.705 49.630 20.905 ;
        RECT 45.155 19.715 46.825 20.485 ;
        RECT 46.995 19.885 47.335 20.515 ;
        RECT 47.505 19.715 47.755 20.515 ;
        RECT 47.945 20.365 49.170 20.535 ;
        RECT 47.945 19.885 48.275 20.365 ;
        RECT 48.445 19.715 48.670 20.175 ;
        RECT 48.840 19.885 49.170 20.365 ;
        RECT 49.800 20.495 49.970 21.125 ;
        RECT 50.675 21.100 50.965 22.265 ;
        RECT 51.135 21.175 52.805 22.265 ;
        RECT 50.155 20.705 50.505 20.955 ;
        RECT 49.800 19.885 50.300 20.495 ;
        RECT 51.135 20.485 51.885 21.005 ;
        RECT 52.055 20.655 52.805 21.175 ;
        RECT 53.435 21.125 53.775 22.095 ;
        RECT 53.945 21.125 54.115 22.265 ;
        RECT 54.385 21.465 54.635 22.265 ;
        RECT 55.280 21.295 55.610 22.095 ;
        RECT 55.910 21.465 56.240 22.265 ;
        RECT 56.410 21.295 56.740 22.095 ;
        RECT 57.205 21.595 57.375 22.095 ;
        RECT 57.545 21.765 57.875 22.265 ;
        RECT 57.205 21.425 57.870 21.595 ;
        RECT 54.305 21.125 56.740 21.295 ;
        RECT 53.435 20.515 53.610 21.125 ;
        RECT 54.305 20.875 54.475 21.125 ;
        RECT 53.780 20.705 54.475 20.875 ;
        RECT 54.650 20.705 55.070 20.905 ;
        RECT 55.240 20.705 55.570 20.905 ;
        RECT 55.740 20.705 56.070 20.905 ;
        RECT 50.675 19.715 50.965 20.440 ;
        RECT 51.135 19.715 52.805 20.485 ;
        RECT 53.435 19.885 53.775 20.515 ;
        RECT 53.945 19.715 54.195 20.515 ;
        RECT 54.385 20.365 55.610 20.535 ;
        RECT 54.385 19.885 54.715 20.365 ;
        RECT 54.885 19.715 55.110 20.175 ;
        RECT 55.280 19.885 55.610 20.365 ;
        RECT 56.240 20.495 56.410 21.125 ;
        RECT 56.595 20.705 56.945 20.955 ;
        RECT 57.120 20.605 57.470 21.255 ;
        RECT 56.240 19.885 56.740 20.495 ;
        RECT 57.640 20.435 57.870 21.425 ;
        RECT 57.205 20.265 57.870 20.435 ;
        RECT 57.205 19.975 57.375 20.265 ;
        RECT 57.545 19.715 57.875 20.095 ;
        RECT 58.045 19.975 58.230 22.095 ;
        RECT 58.470 21.805 58.735 22.265 ;
        RECT 58.905 21.670 59.155 22.095 ;
        RECT 59.365 21.820 60.470 21.990 ;
        RECT 58.850 21.540 59.155 21.670 ;
        RECT 58.400 20.345 58.680 21.295 ;
        RECT 58.850 20.435 59.020 21.540 ;
        RECT 59.190 20.755 59.430 21.350 ;
        RECT 59.600 21.285 60.130 21.650 ;
        RECT 59.600 20.585 59.770 21.285 ;
        RECT 60.300 21.205 60.470 21.820 ;
        RECT 60.640 21.465 60.810 22.265 ;
        RECT 60.980 21.765 61.230 22.095 ;
        RECT 61.455 21.795 62.340 21.965 ;
        RECT 60.300 21.115 60.810 21.205 ;
        RECT 58.850 20.305 59.075 20.435 ;
        RECT 59.245 20.365 59.770 20.585 ;
        RECT 59.940 20.945 60.810 21.115 ;
        RECT 58.485 19.715 58.735 20.175 ;
        RECT 58.905 20.165 59.075 20.305 ;
        RECT 59.940 20.165 60.110 20.945 ;
        RECT 60.640 20.875 60.810 20.945 ;
        RECT 60.320 20.695 60.520 20.725 ;
        RECT 60.980 20.695 61.150 21.765 ;
        RECT 61.320 20.875 61.510 21.595 ;
        RECT 60.320 20.395 61.150 20.695 ;
        RECT 61.680 20.665 62.000 21.625 ;
        RECT 58.905 19.995 59.240 20.165 ;
        RECT 59.435 19.995 60.110 20.165 ;
        RECT 60.430 19.715 60.800 20.215 ;
        RECT 60.980 20.165 61.150 20.395 ;
        RECT 61.535 20.335 62.000 20.665 ;
        RECT 62.170 20.955 62.340 21.795 ;
        RECT 62.520 21.765 62.835 22.265 ;
        RECT 63.065 21.535 63.405 22.095 ;
        RECT 62.510 21.160 63.405 21.535 ;
        RECT 63.575 21.255 63.745 22.265 ;
        RECT 63.215 20.955 63.405 21.160 ;
        RECT 63.915 21.205 64.245 22.050 ;
        RECT 64.565 21.595 64.735 22.095 ;
        RECT 64.905 21.765 65.235 22.265 ;
        RECT 64.565 21.425 65.230 21.595 ;
        RECT 63.915 21.125 64.305 21.205 ;
        RECT 64.090 21.075 64.305 21.125 ;
        RECT 62.170 20.625 63.045 20.955 ;
        RECT 63.215 20.625 63.965 20.955 ;
        RECT 62.170 20.165 62.340 20.625 ;
        RECT 63.215 20.455 63.415 20.625 ;
        RECT 64.135 20.495 64.305 21.075 ;
        RECT 64.480 20.605 64.830 21.255 ;
        RECT 64.080 20.455 64.305 20.495 ;
        RECT 60.980 19.995 61.385 20.165 ;
        RECT 61.555 19.995 62.340 20.165 ;
        RECT 62.615 19.715 62.825 20.245 ;
        RECT 63.085 19.930 63.415 20.455 ;
        RECT 63.925 20.370 64.305 20.455 ;
        RECT 65.000 20.435 65.230 21.425 ;
        RECT 63.585 19.715 63.755 20.325 ;
        RECT 63.925 19.935 64.255 20.370 ;
        RECT 64.565 20.265 65.230 20.435 ;
        RECT 64.565 19.975 64.735 20.265 ;
        RECT 64.905 19.715 65.235 20.095 ;
        RECT 65.405 19.975 65.590 22.095 ;
        RECT 65.830 21.805 66.095 22.265 ;
        RECT 66.265 21.670 66.515 22.095 ;
        RECT 66.725 21.820 67.830 21.990 ;
        RECT 66.210 21.540 66.515 21.670 ;
        RECT 65.760 20.345 66.040 21.295 ;
        RECT 66.210 20.435 66.380 21.540 ;
        RECT 66.550 20.755 66.790 21.350 ;
        RECT 66.960 21.285 67.490 21.650 ;
        RECT 66.960 20.585 67.130 21.285 ;
        RECT 67.660 21.205 67.830 21.820 ;
        RECT 68.000 21.465 68.170 22.265 ;
        RECT 68.340 21.765 68.590 22.095 ;
        RECT 68.815 21.795 69.700 21.965 ;
        RECT 67.660 21.115 68.170 21.205 ;
        RECT 66.210 20.305 66.435 20.435 ;
        RECT 66.605 20.365 67.130 20.585 ;
        RECT 67.300 20.945 68.170 21.115 ;
        RECT 65.845 19.715 66.095 20.175 ;
        RECT 66.265 20.165 66.435 20.305 ;
        RECT 67.300 20.165 67.470 20.945 ;
        RECT 68.000 20.875 68.170 20.945 ;
        RECT 67.680 20.695 67.880 20.725 ;
        RECT 68.340 20.695 68.510 21.765 ;
        RECT 68.680 20.875 68.870 21.595 ;
        RECT 67.680 20.395 68.510 20.695 ;
        RECT 69.040 20.665 69.360 21.625 ;
        RECT 66.265 19.995 66.600 20.165 ;
        RECT 66.795 19.995 67.470 20.165 ;
        RECT 67.790 19.715 68.160 20.215 ;
        RECT 68.340 20.165 68.510 20.395 ;
        RECT 68.895 20.335 69.360 20.665 ;
        RECT 69.530 20.955 69.700 21.795 ;
        RECT 69.880 21.765 70.195 22.265 ;
        RECT 70.425 21.535 70.765 22.095 ;
        RECT 69.870 21.160 70.765 21.535 ;
        RECT 70.935 21.255 71.105 22.265 ;
        RECT 70.575 20.955 70.765 21.160 ;
        RECT 71.275 21.205 71.605 22.050 ;
        RECT 71.275 21.125 71.665 21.205 ;
        RECT 71.450 21.075 71.665 21.125 ;
        RECT 69.530 20.625 70.405 20.955 ;
        RECT 70.575 20.625 71.325 20.955 ;
        RECT 69.530 20.165 69.700 20.625 ;
        RECT 70.575 20.455 70.775 20.625 ;
        RECT 71.495 20.495 71.665 21.075 ;
        RECT 71.440 20.455 71.665 20.495 ;
        RECT 68.340 19.995 68.745 20.165 ;
        RECT 68.915 19.995 69.700 20.165 ;
        RECT 69.975 19.715 70.185 20.245 ;
        RECT 70.445 19.930 70.775 20.455 ;
        RECT 71.285 20.370 71.665 20.455 ;
        RECT 71.835 21.125 72.175 22.095 ;
        RECT 72.345 21.125 72.515 22.265 ;
        RECT 72.785 21.465 73.035 22.265 ;
        RECT 73.680 21.295 74.010 22.095 ;
        RECT 74.310 21.465 74.640 22.265 ;
        RECT 74.810 21.295 75.140 22.095 ;
        RECT 72.705 21.125 75.140 21.295 ;
        RECT 71.835 20.515 72.010 21.125 ;
        RECT 72.705 20.875 72.875 21.125 ;
        RECT 72.180 20.705 72.875 20.875 ;
        RECT 73.050 20.705 73.470 20.905 ;
        RECT 73.640 20.705 73.970 20.905 ;
        RECT 74.140 20.705 74.470 20.905 ;
        RECT 70.945 19.715 71.115 20.325 ;
        RECT 71.285 19.935 71.615 20.370 ;
        RECT 71.835 19.885 72.175 20.515 ;
        RECT 72.345 19.715 72.595 20.515 ;
        RECT 72.785 20.365 74.010 20.535 ;
        RECT 72.785 19.885 73.115 20.365 ;
        RECT 73.285 19.715 73.510 20.175 ;
        RECT 73.680 19.885 74.010 20.365 ;
        RECT 74.640 20.495 74.810 21.125 ;
        RECT 76.435 21.100 76.725 22.265 ;
        RECT 77.560 21.295 77.890 22.095 ;
        RECT 78.060 21.465 78.390 22.265 ;
        RECT 78.690 21.295 79.020 22.095 ;
        RECT 79.665 21.465 79.915 22.265 ;
        RECT 77.560 21.125 79.995 21.295 ;
        RECT 80.185 21.125 80.355 22.265 ;
        RECT 80.525 21.125 80.865 22.095 ;
        RECT 81.240 21.295 81.570 22.095 ;
        RECT 81.740 21.465 82.070 22.265 ;
        RECT 82.370 21.295 82.700 22.095 ;
        RECT 83.345 21.465 83.595 22.265 ;
        RECT 81.240 21.125 83.675 21.295 ;
        RECT 83.865 21.125 84.035 22.265 ;
        RECT 84.205 21.125 84.545 22.095 ;
        RECT 84.805 21.335 84.975 22.095 ;
        RECT 85.190 21.505 85.520 22.265 ;
        RECT 84.805 21.165 85.520 21.335 ;
        RECT 85.690 21.190 85.945 22.095 ;
        RECT 74.995 20.705 75.345 20.955 ;
        RECT 77.355 20.705 77.705 20.955 ;
        RECT 77.890 20.495 78.060 21.125 ;
        RECT 78.230 20.705 78.560 20.905 ;
        RECT 78.730 20.705 79.060 20.905 ;
        RECT 79.230 20.705 79.650 20.905 ;
        RECT 79.825 20.875 79.995 21.125 ;
        RECT 79.825 20.705 80.520 20.875 ;
        RECT 74.640 19.885 75.140 20.495 ;
        RECT 76.435 19.715 76.725 20.440 ;
        RECT 77.560 19.885 78.060 20.495 ;
        RECT 78.690 20.365 79.915 20.535 ;
        RECT 80.690 20.515 80.865 21.125 ;
        RECT 81.035 20.705 81.385 20.955 ;
        RECT 78.690 19.885 79.020 20.365 ;
        RECT 79.190 19.715 79.415 20.175 ;
        RECT 79.585 19.885 79.915 20.365 ;
        RECT 80.105 19.715 80.355 20.515 ;
        RECT 80.525 19.885 80.865 20.515 ;
        RECT 81.570 20.495 81.740 21.125 ;
        RECT 81.910 20.705 82.240 20.905 ;
        RECT 82.410 20.705 82.740 20.905 ;
        RECT 82.910 20.705 83.330 20.905 ;
        RECT 83.505 20.875 83.675 21.125 ;
        RECT 83.505 20.705 84.200 20.875 ;
        RECT 81.240 19.885 81.740 20.495 ;
        RECT 82.370 20.365 83.595 20.535 ;
        RECT 84.370 20.515 84.545 21.125 ;
        RECT 84.715 20.615 85.070 20.985 ;
        RECT 85.350 20.955 85.520 21.165 ;
        RECT 85.350 20.625 85.605 20.955 ;
        RECT 82.370 19.885 82.700 20.365 ;
        RECT 82.870 19.715 83.095 20.175 ;
        RECT 83.265 19.885 83.595 20.365 ;
        RECT 83.785 19.715 84.035 20.515 ;
        RECT 84.205 19.885 84.545 20.515 ;
        RECT 85.350 20.435 85.520 20.625 ;
        RECT 85.775 20.460 85.945 21.190 ;
        RECT 86.120 21.115 86.380 22.265 ;
        RECT 86.645 21.335 86.815 22.095 ;
        RECT 87.030 21.505 87.360 22.265 ;
        RECT 86.645 21.165 87.360 21.335 ;
        RECT 87.530 21.190 87.785 22.095 ;
        RECT 86.555 20.615 86.910 20.985 ;
        RECT 87.190 20.955 87.360 21.165 ;
        RECT 87.190 20.625 87.445 20.955 ;
        RECT 84.805 20.265 85.520 20.435 ;
        RECT 84.805 19.885 84.975 20.265 ;
        RECT 85.190 19.715 85.520 20.095 ;
        RECT 85.690 19.885 85.945 20.460 ;
        RECT 86.120 19.715 86.380 20.555 ;
        RECT 87.190 20.435 87.360 20.625 ;
        RECT 87.615 20.460 87.785 21.190 ;
        RECT 87.960 21.115 88.220 22.265 ;
        RECT 89.315 21.175 90.525 22.265 ;
        RECT 89.315 20.635 89.835 21.175 ;
        RECT 86.645 20.265 87.360 20.435 ;
        RECT 86.645 19.885 86.815 20.265 ;
        RECT 87.030 19.715 87.360 20.095 ;
        RECT 87.530 19.885 87.785 20.460 ;
        RECT 87.960 19.715 88.220 20.555 ;
        RECT 90.005 20.465 90.525 21.005 ;
        RECT 89.315 19.715 90.525 20.465 ;
        RECT 11.950 19.545 90.610 19.715 ;
        RECT 12.035 18.795 13.245 19.545 ;
        RECT 14.500 19.035 14.740 19.545 ;
        RECT 14.920 19.035 15.200 19.365 ;
        RECT 15.430 19.035 15.645 19.545 ;
        RECT 12.035 18.255 12.555 18.795 ;
        RECT 12.725 18.085 13.245 18.625 ;
        RECT 14.395 18.305 14.750 18.865 ;
        RECT 14.920 18.135 15.090 19.035 ;
        RECT 15.260 18.305 15.525 18.865 ;
        RECT 15.815 18.805 16.430 19.375 ;
        RECT 15.775 18.135 15.945 18.635 ;
        RECT 12.035 16.995 13.245 18.085 ;
        RECT 14.520 17.965 15.945 18.135 ;
        RECT 14.520 17.790 14.910 17.965 ;
        RECT 15.395 16.995 15.725 17.795 ;
        RECT 16.115 17.785 16.430 18.805 ;
        RECT 16.635 18.795 17.845 19.545 ;
        RECT 18.105 18.995 18.275 19.285 ;
        RECT 18.445 19.165 18.775 19.545 ;
        RECT 18.105 18.825 18.770 18.995 ;
        RECT 16.635 18.255 17.155 18.795 ;
        RECT 17.325 18.085 17.845 18.625 ;
        RECT 15.895 17.165 16.430 17.785 ;
        RECT 16.635 16.995 17.845 18.085 ;
        RECT 18.020 18.005 18.370 18.655 ;
        RECT 18.540 17.835 18.770 18.825 ;
        RECT 18.105 17.665 18.770 17.835 ;
        RECT 18.105 17.165 18.275 17.665 ;
        RECT 18.445 16.995 18.775 17.495 ;
        RECT 18.945 17.165 19.130 19.285 ;
        RECT 19.385 19.085 19.635 19.545 ;
        RECT 19.805 19.095 20.140 19.265 ;
        RECT 20.335 19.095 21.010 19.265 ;
        RECT 19.805 18.955 19.975 19.095 ;
        RECT 19.300 17.965 19.580 18.915 ;
        RECT 19.750 18.825 19.975 18.955 ;
        RECT 19.750 17.720 19.920 18.825 ;
        RECT 20.145 18.675 20.670 18.895 ;
        RECT 20.090 17.910 20.330 18.505 ;
        RECT 20.500 17.975 20.670 18.675 ;
        RECT 20.840 18.315 21.010 19.095 ;
        RECT 21.330 19.045 21.700 19.545 ;
        RECT 21.880 19.095 22.285 19.265 ;
        RECT 22.455 19.095 23.240 19.265 ;
        RECT 21.880 18.865 22.050 19.095 ;
        RECT 21.220 18.565 22.050 18.865 ;
        RECT 22.435 18.595 22.900 18.925 ;
        RECT 21.220 18.535 21.420 18.565 ;
        RECT 21.540 18.315 21.710 18.385 ;
        RECT 20.840 18.145 21.710 18.315 ;
        RECT 21.200 18.055 21.710 18.145 ;
        RECT 19.750 17.590 20.055 17.720 ;
        RECT 20.500 17.610 21.030 17.975 ;
        RECT 19.370 16.995 19.635 17.455 ;
        RECT 19.805 17.165 20.055 17.590 ;
        RECT 21.200 17.440 21.370 18.055 ;
        RECT 20.265 17.270 21.370 17.440 ;
        RECT 21.540 16.995 21.710 17.795 ;
        RECT 21.880 17.495 22.050 18.565 ;
        RECT 22.220 17.665 22.410 18.385 ;
        RECT 22.580 17.635 22.900 18.595 ;
        RECT 23.070 18.635 23.240 19.095 ;
        RECT 23.515 19.015 23.725 19.545 ;
        RECT 23.985 18.805 24.315 19.330 ;
        RECT 24.485 18.935 24.655 19.545 ;
        RECT 24.825 18.890 25.155 19.325 ;
        RECT 25.540 19.035 25.780 19.545 ;
        RECT 25.960 19.035 26.240 19.365 ;
        RECT 26.470 19.035 26.685 19.545 ;
        RECT 24.825 18.805 25.205 18.890 ;
        RECT 24.115 18.635 24.315 18.805 ;
        RECT 24.980 18.765 25.205 18.805 ;
        RECT 23.070 18.305 23.945 18.635 ;
        RECT 24.115 18.305 24.865 18.635 ;
        RECT 21.880 17.165 22.130 17.495 ;
        RECT 23.070 17.465 23.240 18.305 ;
        RECT 24.115 18.100 24.305 18.305 ;
        RECT 25.035 18.185 25.205 18.765 ;
        RECT 25.435 18.305 25.790 18.865 ;
        RECT 24.990 18.135 25.205 18.185 ;
        RECT 25.960 18.135 26.130 19.035 ;
        RECT 26.300 18.305 26.565 18.865 ;
        RECT 26.855 18.805 27.470 19.375 ;
        RECT 27.765 18.995 27.935 19.285 ;
        RECT 28.105 19.165 28.435 19.545 ;
        RECT 27.765 18.825 28.430 18.995 ;
        RECT 26.815 18.135 26.985 18.635 ;
        RECT 23.410 17.725 24.305 18.100 ;
        RECT 24.815 18.055 25.205 18.135 ;
        RECT 22.355 17.295 23.240 17.465 ;
        RECT 23.420 16.995 23.735 17.495 ;
        RECT 23.965 17.165 24.305 17.725 ;
        RECT 24.475 16.995 24.645 18.005 ;
        RECT 24.815 17.210 25.145 18.055 ;
        RECT 25.560 17.965 26.985 18.135 ;
        RECT 25.560 17.790 25.950 17.965 ;
        RECT 26.435 16.995 26.765 17.795 ;
        RECT 27.155 17.785 27.470 18.805 ;
        RECT 27.680 18.005 28.030 18.655 ;
        RECT 28.200 17.835 28.430 18.825 ;
        RECT 26.935 17.165 27.470 17.785 ;
        RECT 27.765 17.665 28.430 17.835 ;
        RECT 27.765 17.165 27.935 17.665 ;
        RECT 28.105 16.995 28.435 17.495 ;
        RECT 28.605 17.165 28.790 19.285 ;
        RECT 29.045 19.085 29.295 19.545 ;
        RECT 29.465 19.095 29.800 19.265 ;
        RECT 29.995 19.095 30.670 19.265 ;
        RECT 29.465 18.955 29.635 19.095 ;
        RECT 28.960 17.965 29.240 18.915 ;
        RECT 29.410 18.825 29.635 18.955 ;
        RECT 29.410 17.720 29.580 18.825 ;
        RECT 29.805 18.675 30.330 18.895 ;
        RECT 29.750 17.910 29.990 18.505 ;
        RECT 30.160 17.975 30.330 18.675 ;
        RECT 30.500 18.315 30.670 19.095 ;
        RECT 30.990 19.045 31.360 19.545 ;
        RECT 31.540 19.095 31.945 19.265 ;
        RECT 32.115 19.095 32.900 19.265 ;
        RECT 31.540 18.865 31.710 19.095 ;
        RECT 30.880 18.565 31.710 18.865 ;
        RECT 32.095 18.595 32.560 18.925 ;
        RECT 30.880 18.535 31.080 18.565 ;
        RECT 31.200 18.315 31.370 18.385 ;
        RECT 30.500 18.145 31.370 18.315 ;
        RECT 30.860 18.055 31.370 18.145 ;
        RECT 29.410 17.590 29.715 17.720 ;
        RECT 30.160 17.610 30.690 17.975 ;
        RECT 29.030 16.995 29.295 17.455 ;
        RECT 29.465 17.165 29.715 17.590 ;
        RECT 30.860 17.440 31.030 18.055 ;
        RECT 29.925 17.270 31.030 17.440 ;
        RECT 31.200 16.995 31.370 17.795 ;
        RECT 31.540 17.495 31.710 18.565 ;
        RECT 31.880 17.665 32.070 18.385 ;
        RECT 32.240 17.635 32.560 18.595 ;
        RECT 32.730 18.635 32.900 19.095 ;
        RECT 33.175 19.015 33.385 19.545 ;
        RECT 33.645 18.805 33.975 19.330 ;
        RECT 34.145 18.935 34.315 19.545 ;
        RECT 34.485 18.890 34.815 19.325 ;
        RECT 34.485 18.805 34.865 18.890 ;
        RECT 33.775 18.635 33.975 18.805 ;
        RECT 34.640 18.765 34.865 18.805 ;
        RECT 32.730 18.305 33.605 18.635 ;
        RECT 33.775 18.305 34.525 18.635 ;
        RECT 31.540 17.165 31.790 17.495 ;
        RECT 32.730 17.465 32.900 18.305 ;
        RECT 33.775 18.100 33.965 18.305 ;
        RECT 34.695 18.185 34.865 18.765 ;
        RECT 34.650 18.135 34.865 18.185 ;
        RECT 33.070 17.725 33.965 18.100 ;
        RECT 34.475 18.055 34.865 18.135 ;
        RECT 35.070 18.805 35.685 19.375 ;
        RECT 35.855 19.035 36.070 19.545 ;
        RECT 36.300 19.035 36.580 19.365 ;
        RECT 36.760 19.035 37.000 19.545 ;
        RECT 32.015 17.295 32.900 17.465 ;
        RECT 33.080 16.995 33.395 17.495 ;
        RECT 33.625 17.165 33.965 17.725 ;
        RECT 34.135 16.995 34.305 18.005 ;
        RECT 34.475 17.210 34.805 18.055 ;
        RECT 35.070 17.785 35.385 18.805 ;
        RECT 35.555 18.135 35.725 18.635 ;
        RECT 35.975 18.305 36.240 18.865 ;
        RECT 36.410 18.135 36.580 19.035 ;
        RECT 36.750 18.305 37.105 18.865 ;
        RECT 37.795 18.820 38.085 19.545 ;
        RECT 38.765 18.890 39.095 19.325 ;
        RECT 39.265 18.935 39.435 19.545 ;
        RECT 38.715 18.805 39.095 18.890 ;
        RECT 39.605 18.805 39.935 19.330 ;
        RECT 40.195 19.015 40.405 19.545 ;
        RECT 40.680 19.095 41.465 19.265 ;
        RECT 41.635 19.095 42.040 19.265 ;
        RECT 38.715 18.765 38.940 18.805 ;
        RECT 38.715 18.185 38.885 18.765 ;
        RECT 39.605 18.635 39.805 18.805 ;
        RECT 40.680 18.635 40.850 19.095 ;
        RECT 39.055 18.305 39.805 18.635 ;
        RECT 39.975 18.305 40.850 18.635 ;
        RECT 35.555 17.965 36.980 18.135 ;
        RECT 35.070 17.165 35.605 17.785 ;
        RECT 35.775 16.995 36.105 17.795 ;
        RECT 36.590 17.790 36.980 17.965 ;
        RECT 37.795 16.995 38.085 18.160 ;
        RECT 38.715 18.135 38.930 18.185 ;
        RECT 38.715 18.055 39.105 18.135 ;
        RECT 38.775 17.210 39.105 18.055 ;
        RECT 39.615 18.100 39.805 18.305 ;
        RECT 39.275 16.995 39.445 18.005 ;
        RECT 39.615 17.725 40.510 18.100 ;
        RECT 39.615 17.165 39.955 17.725 ;
        RECT 40.185 16.995 40.500 17.495 ;
        RECT 40.680 17.465 40.850 18.305 ;
        RECT 41.020 18.595 41.485 18.925 ;
        RECT 41.870 18.865 42.040 19.095 ;
        RECT 42.220 19.045 42.590 19.545 ;
        RECT 42.910 19.095 43.585 19.265 ;
        RECT 43.780 19.095 44.115 19.265 ;
        RECT 41.020 17.635 41.340 18.595 ;
        RECT 41.870 18.565 42.700 18.865 ;
        RECT 41.510 17.665 41.700 18.385 ;
        RECT 41.870 17.495 42.040 18.565 ;
        RECT 42.500 18.535 42.700 18.565 ;
        RECT 42.210 18.315 42.380 18.385 ;
        RECT 42.910 18.315 43.080 19.095 ;
        RECT 43.945 18.955 44.115 19.095 ;
        RECT 44.285 19.085 44.535 19.545 ;
        RECT 42.210 18.145 43.080 18.315 ;
        RECT 43.250 18.675 43.775 18.895 ;
        RECT 43.945 18.825 44.170 18.955 ;
        RECT 42.210 18.055 42.720 18.145 ;
        RECT 40.680 17.295 41.565 17.465 ;
        RECT 41.790 17.165 42.040 17.495 ;
        RECT 42.210 16.995 42.380 17.795 ;
        RECT 42.550 17.440 42.720 18.055 ;
        RECT 43.250 17.975 43.420 18.675 ;
        RECT 42.890 17.610 43.420 17.975 ;
        RECT 43.590 17.910 43.830 18.505 ;
        RECT 44.000 17.720 44.170 18.825 ;
        RECT 44.340 17.965 44.620 18.915 ;
        RECT 43.865 17.590 44.170 17.720 ;
        RECT 42.550 17.270 43.655 17.440 ;
        RECT 43.865 17.165 44.115 17.590 ;
        RECT 44.285 16.995 44.550 17.455 ;
        RECT 44.790 17.165 44.975 19.285 ;
        RECT 45.145 19.165 45.475 19.545 ;
        RECT 45.645 18.995 45.815 19.285 ;
        RECT 45.150 18.825 45.815 18.995 ;
        RECT 46.625 18.995 46.795 19.285 ;
        RECT 46.965 19.165 47.295 19.545 ;
        RECT 46.625 18.825 47.290 18.995 ;
        RECT 45.150 17.835 45.380 18.825 ;
        RECT 45.550 18.005 45.900 18.655 ;
        RECT 46.540 18.005 46.890 18.655 ;
        RECT 47.060 17.835 47.290 18.825 ;
        RECT 45.150 17.665 45.815 17.835 ;
        RECT 45.145 16.995 45.475 17.495 ;
        RECT 45.645 17.165 45.815 17.665 ;
        RECT 46.625 17.665 47.290 17.835 ;
        RECT 46.625 17.165 46.795 17.665 ;
        RECT 46.965 16.995 47.295 17.495 ;
        RECT 47.465 17.165 47.650 19.285 ;
        RECT 47.905 19.085 48.155 19.545 ;
        RECT 48.325 19.095 48.660 19.265 ;
        RECT 48.855 19.095 49.530 19.265 ;
        RECT 48.325 18.955 48.495 19.095 ;
        RECT 47.820 17.965 48.100 18.915 ;
        RECT 48.270 18.825 48.495 18.955 ;
        RECT 48.270 17.720 48.440 18.825 ;
        RECT 48.665 18.675 49.190 18.895 ;
        RECT 48.610 17.910 48.850 18.505 ;
        RECT 49.020 17.975 49.190 18.675 ;
        RECT 49.360 18.315 49.530 19.095 ;
        RECT 49.850 19.045 50.220 19.545 ;
        RECT 50.400 19.095 50.805 19.265 ;
        RECT 50.975 19.095 51.760 19.265 ;
        RECT 50.400 18.865 50.570 19.095 ;
        RECT 49.740 18.565 50.570 18.865 ;
        RECT 50.955 18.595 51.420 18.925 ;
        RECT 49.740 18.535 49.940 18.565 ;
        RECT 50.060 18.315 50.230 18.385 ;
        RECT 49.360 18.145 50.230 18.315 ;
        RECT 49.720 18.055 50.230 18.145 ;
        RECT 48.270 17.590 48.575 17.720 ;
        RECT 49.020 17.610 49.550 17.975 ;
        RECT 47.890 16.995 48.155 17.455 ;
        RECT 48.325 17.165 48.575 17.590 ;
        RECT 49.720 17.440 49.890 18.055 ;
        RECT 48.785 17.270 49.890 17.440 ;
        RECT 50.060 16.995 50.230 17.795 ;
        RECT 50.400 17.495 50.570 18.565 ;
        RECT 50.740 17.665 50.930 18.385 ;
        RECT 51.100 17.635 51.420 18.595 ;
        RECT 51.590 18.635 51.760 19.095 ;
        RECT 52.035 19.015 52.245 19.545 ;
        RECT 52.505 18.805 52.835 19.330 ;
        RECT 53.005 18.935 53.175 19.545 ;
        RECT 53.345 18.890 53.675 19.325 ;
        RECT 53.985 18.995 54.155 19.285 ;
        RECT 54.325 19.165 54.655 19.545 ;
        RECT 53.345 18.805 53.725 18.890 ;
        RECT 53.985 18.825 54.650 18.995 ;
        RECT 52.635 18.635 52.835 18.805 ;
        RECT 53.500 18.765 53.725 18.805 ;
        RECT 51.590 18.305 52.465 18.635 ;
        RECT 52.635 18.305 53.385 18.635 ;
        RECT 50.400 17.165 50.650 17.495 ;
        RECT 51.590 17.465 51.760 18.305 ;
        RECT 52.635 18.100 52.825 18.305 ;
        RECT 53.555 18.185 53.725 18.765 ;
        RECT 53.510 18.135 53.725 18.185 ;
        RECT 51.930 17.725 52.825 18.100 ;
        RECT 53.335 18.055 53.725 18.135 ;
        RECT 50.875 17.295 51.760 17.465 ;
        RECT 51.940 16.995 52.255 17.495 ;
        RECT 52.485 17.165 52.825 17.725 ;
        RECT 52.995 16.995 53.165 18.005 ;
        RECT 53.335 17.210 53.665 18.055 ;
        RECT 53.900 18.005 54.250 18.655 ;
        RECT 54.420 17.835 54.650 18.825 ;
        RECT 53.985 17.665 54.650 17.835 ;
        RECT 53.985 17.165 54.155 17.665 ;
        RECT 54.325 16.995 54.655 17.495 ;
        RECT 54.825 17.165 55.010 19.285 ;
        RECT 55.265 19.085 55.515 19.545 ;
        RECT 55.685 19.095 56.020 19.265 ;
        RECT 56.215 19.095 56.890 19.265 ;
        RECT 55.685 18.955 55.855 19.095 ;
        RECT 55.180 17.965 55.460 18.915 ;
        RECT 55.630 18.825 55.855 18.955 ;
        RECT 55.630 17.720 55.800 18.825 ;
        RECT 56.025 18.675 56.550 18.895 ;
        RECT 55.970 17.910 56.210 18.505 ;
        RECT 56.380 17.975 56.550 18.675 ;
        RECT 56.720 18.315 56.890 19.095 ;
        RECT 57.210 19.045 57.580 19.545 ;
        RECT 57.760 19.095 58.165 19.265 ;
        RECT 58.335 19.095 59.120 19.265 ;
        RECT 57.760 18.865 57.930 19.095 ;
        RECT 57.100 18.565 57.930 18.865 ;
        RECT 58.315 18.595 58.780 18.925 ;
        RECT 57.100 18.535 57.300 18.565 ;
        RECT 57.420 18.315 57.590 18.385 ;
        RECT 56.720 18.145 57.590 18.315 ;
        RECT 57.080 18.055 57.590 18.145 ;
        RECT 55.630 17.590 55.935 17.720 ;
        RECT 56.380 17.610 56.910 17.975 ;
        RECT 55.250 16.995 55.515 17.455 ;
        RECT 55.685 17.165 55.935 17.590 ;
        RECT 57.080 17.440 57.250 18.055 ;
        RECT 56.145 17.270 57.250 17.440 ;
        RECT 57.420 16.995 57.590 17.795 ;
        RECT 57.760 17.495 57.930 18.565 ;
        RECT 58.100 17.665 58.290 18.385 ;
        RECT 58.460 17.635 58.780 18.595 ;
        RECT 58.950 18.635 59.120 19.095 ;
        RECT 59.395 19.015 59.605 19.545 ;
        RECT 59.865 18.805 60.195 19.330 ;
        RECT 60.365 18.935 60.535 19.545 ;
        RECT 60.705 18.890 61.035 19.325 ;
        RECT 60.705 18.805 61.085 18.890 ;
        RECT 59.995 18.635 60.195 18.805 ;
        RECT 60.860 18.765 61.085 18.805 ;
        RECT 58.950 18.305 59.825 18.635 ;
        RECT 59.995 18.305 60.745 18.635 ;
        RECT 57.760 17.165 58.010 17.495 ;
        RECT 58.950 17.465 59.120 18.305 ;
        RECT 59.995 18.100 60.185 18.305 ;
        RECT 60.915 18.185 61.085 18.765 ;
        RECT 60.870 18.135 61.085 18.185 ;
        RECT 59.290 17.725 60.185 18.100 ;
        RECT 60.695 18.055 61.085 18.135 ;
        RECT 61.290 18.805 61.905 19.375 ;
        RECT 62.075 19.035 62.290 19.545 ;
        RECT 62.520 19.035 62.800 19.365 ;
        RECT 62.980 19.035 63.220 19.545 ;
        RECT 58.235 17.295 59.120 17.465 ;
        RECT 59.300 16.995 59.615 17.495 ;
        RECT 59.845 17.165 60.185 17.725 ;
        RECT 60.355 16.995 60.525 18.005 ;
        RECT 60.695 17.210 61.025 18.055 ;
        RECT 61.290 17.785 61.605 18.805 ;
        RECT 61.775 18.135 61.945 18.635 ;
        RECT 62.195 18.305 62.460 18.865 ;
        RECT 62.630 18.135 62.800 19.035 ;
        RECT 62.970 18.305 63.325 18.865 ;
        RECT 63.555 18.820 63.845 19.545 ;
        RECT 64.015 19.045 64.275 19.375 ;
        RECT 64.445 19.185 64.775 19.545 ;
        RECT 65.030 19.165 66.330 19.375 ;
        RECT 61.775 17.965 63.200 18.135 ;
        RECT 61.290 17.165 61.825 17.785 ;
        RECT 61.995 16.995 62.325 17.795 ;
        RECT 62.810 17.790 63.200 17.965 ;
        RECT 63.555 16.995 63.845 18.160 ;
        RECT 64.015 17.845 64.185 19.045 ;
        RECT 65.030 19.015 65.200 19.165 ;
        RECT 64.445 18.890 65.200 19.015 ;
        RECT 64.355 18.845 65.200 18.890 ;
        RECT 64.355 18.725 64.625 18.845 ;
        RECT 64.355 18.150 64.525 18.725 ;
        RECT 64.755 18.285 65.165 18.590 ;
        RECT 65.455 18.555 65.665 18.955 ;
        RECT 65.335 18.345 65.665 18.555 ;
        RECT 65.910 18.555 66.130 18.955 ;
        RECT 66.605 18.780 67.060 19.545 ;
        RECT 67.235 18.795 68.445 19.545 ;
        RECT 68.705 18.995 68.875 19.285 ;
        RECT 69.045 19.165 69.375 19.545 ;
        RECT 68.705 18.825 69.370 18.995 ;
        RECT 65.910 18.345 66.385 18.555 ;
        RECT 66.575 18.355 67.065 18.555 ;
        RECT 67.235 18.255 67.755 18.795 ;
        RECT 64.355 18.115 64.555 18.150 ;
        RECT 65.885 18.115 67.060 18.175 ;
        RECT 64.355 18.005 67.060 18.115 ;
        RECT 67.925 18.085 68.445 18.625 ;
        RECT 64.415 17.945 66.215 18.005 ;
        RECT 65.885 17.915 66.215 17.945 ;
        RECT 64.015 17.165 64.275 17.845 ;
        RECT 64.445 16.995 64.695 17.775 ;
        RECT 64.945 17.745 65.780 17.755 ;
        RECT 66.370 17.745 66.555 17.835 ;
        RECT 64.945 17.545 66.555 17.745 ;
        RECT 64.945 17.165 65.195 17.545 ;
        RECT 66.325 17.505 66.555 17.545 ;
        RECT 66.805 17.385 67.060 18.005 ;
        RECT 65.365 16.995 65.720 17.375 ;
        RECT 66.725 17.165 67.060 17.385 ;
        RECT 67.235 16.995 68.445 18.085 ;
        RECT 68.620 18.005 68.970 18.655 ;
        RECT 69.140 17.835 69.370 18.825 ;
        RECT 68.705 17.665 69.370 17.835 ;
        RECT 68.705 17.165 68.875 17.665 ;
        RECT 69.045 16.995 69.375 17.495 ;
        RECT 69.545 17.165 69.730 19.285 ;
        RECT 69.985 19.085 70.235 19.545 ;
        RECT 70.405 19.095 70.740 19.265 ;
        RECT 70.935 19.095 71.610 19.265 ;
        RECT 70.405 18.955 70.575 19.095 ;
        RECT 69.900 17.965 70.180 18.915 ;
        RECT 70.350 18.825 70.575 18.955 ;
        RECT 70.350 17.720 70.520 18.825 ;
        RECT 70.745 18.675 71.270 18.895 ;
        RECT 70.690 17.910 70.930 18.505 ;
        RECT 71.100 17.975 71.270 18.675 ;
        RECT 71.440 18.315 71.610 19.095 ;
        RECT 71.930 19.045 72.300 19.545 ;
        RECT 72.480 19.095 72.885 19.265 ;
        RECT 73.055 19.095 73.840 19.265 ;
        RECT 72.480 18.865 72.650 19.095 ;
        RECT 71.820 18.565 72.650 18.865 ;
        RECT 73.035 18.595 73.500 18.925 ;
        RECT 71.820 18.535 72.020 18.565 ;
        RECT 72.140 18.315 72.310 18.385 ;
        RECT 71.440 18.145 72.310 18.315 ;
        RECT 71.800 18.055 72.310 18.145 ;
        RECT 70.350 17.590 70.655 17.720 ;
        RECT 71.100 17.610 71.630 17.975 ;
        RECT 69.970 16.995 70.235 17.455 ;
        RECT 70.405 17.165 70.655 17.590 ;
        RECT 71.800 17.440 71.970 18.055 ;
        RECT 70.865 17.270 71.970 17.440 ;
        RECT 72.140 16.995 72.310 17.795 ;
        RECT 72.480 17.495 72.650 18.565 ;
        RECT 72.820 17.665 73.010 18.385 ;
        RECT 73.180 17.635 73.500 18.595 ;
        RECT 73.670 18.635 73.840 19.095 ;
        RECT 74.115 19.015 74.325 19.545 ;
        RECT 74.585 18.805 74.915 19.330 ;
        RECT 75.085 18.935 75.255 19.545 ;
        RECT 75.425 18.890 75.755 19.325 ;
        RECT 76.140 19.035 76.380 19.545 ;
        RECT 76.560 19.035 76.840 19.365 ;
        RECT 77.070 19.035 77.285 19.545 ;
        RECT 75.425 18.805 75.805 18.890 ;
        RECT 74.715 18.635 74.915 18.805 ;
        RECT 75.580 18.765 75.805 18.805 ;
        RECT 73.670 18.305 74.545 18.635 ;
        RECT 74.715 18.305 75.465 18.635 ;
        RECT 72.480 17.165 72.730 17.495 ;
        RECT 73.670 17.465 73.840 18.305 ;
        RECT 74.715 18.100 74.905 18.305 ;
        RECT 75.635 18.185 75.805 18.765 ;
        RECT 76.035 18.305 76.390 18.865 ;
        RECT 75.590 18.135 75.805 18.185 ;
        RECT 76.560 18.135 76.730 19.035 ;
        RECT 76.900 18.305 77.165 18.865 ;
        RECT 77.455 18.805 78.070 19.375 ;
        RECT 77.415 18.135 77.585 18.635 ;
        RECT 74.010 17.725 74.905 18.100 ;
        RECT 75.415 18.055 75.805 18.135 ;
        RECT 72.955 17.295 73.840 17.465 ;
        RECT 74.020 16.995 74.335 17.495 ;
        RECT 74.565 17.165 74.905 17.725 ;
        RECT 75.075 16.995 75.245 18.005 ;
        RECT 75.415 17.210 75.745 18.055 ;
        RECT 76.160 17.965 77.585 18.135 ;
        RECT 76.160 17.790 76.550 17.965 ;
        RECT 77.035 16.995 77.365 17.795 ;
        RECT 77.755 17.785 78.070 18.805 ;
        RECT 78.275 18.795 79.485 19.545 ;
        RECT 79.745 18.995 79.915 19.285 ;
        RECT 80.085 19.165 80.415 19.545 ;
        RECT 79.745 18.825 80.410 18.995 ;
        RECT 78.275 18.255 78.795 18.795 ;
        RECT 78.965 18.085 79.485 18.625 ;
        RECT 77.535 17.165 78.070 17.785 ;
        RECT 78.275 16.995 79.485 18.085 ;
        RECT 79.660 18.005 80.010 18.655 ;
        RECT 80.180 17.835 80.410 18.825 ;
        RECT 79.745 17.665 80.410 17.835 ;
        RECT 79.745 17.165 79.915 17.665 ;
        RECT 80.085 16.995 80.415 17.495 ;
        RECT 80.585 17.165 80.770 19.285 ;
        RECT 81.025 19.085 81.275 19.545 ;
        RECT 81.445 19.095 81.780 19.265 ;
        RECT 81.975 19.095 82.650 19.265 ;
        RECT 81.445 18.955 81.615 19.095 ;
        RECT 80.940 17.965 81.220 18.915 ;
        RECT 81.390 18.825 81.615 18.955 ;
        RECT 81.390 17.720 81.560 18.825 ;
        RECT 81.785 18.675 82.310 18.895 ;
        RECT 81.730 17.910 81.970 18.505 ;
        RECT 82.140 17.975 82.310 18.675 ;
        RECT 82.480 18.315 82.650 19.095 ;
        RECT 82.970 19.045 83.340 19.545 ;
        RECT 83.520 19.095 83.925 19.265 ;
        RECT 84.095 19.095 84.880 19.265 ;
        RECT 83.520 18.865 83.690 19.095 ;
        RECT 82.860 18.565 83.690 18.865 ;
        RECT 84.075 18.595 84.540 18.925 ;
        RECT 82.860 18.535 83.060 18.565 ;
        RECT 83.180 18.315 83.350 18.385 ;
        RECT 82.480 18.145 83.350 18.315 ;
        RECT 82.840 18.055 83.350 18.145 ;
        RECT 81.390 17.590 81.695 17.720 ;
        RECT 82.140 17.610 82.670 17.975 ;
        RECT 81.010 16.995 81.275 17.455 ;
        RECT 81.445 17.165 81.695 17.590 ;
        RECT 82.840 17.440 83.010 18.055 ;
        RECT 81.905 17.270 83.010 17.440 ;
        RECT 83.180 16.995 83.350 17.795 ;
        RECT 83.520 17.495 83.690 18.565 ;
        RECT 83.860 17.665 84.050 18.385 ;
        RECT 84.220 17.635 84.540 18.595 ;
        RECT 84.710 18.635 84.880 19.095 ;
        RECT 85.155 19.015 85.365 19.545 ;
        RECT 85.625 18.805 85.955 19.330 ;
        RECT 86.125 18.935 86.295 19.545 ;
        RECT 86.465 18.890 86.795 19.325 ;
        RECT 87.105 18.995 87.275 19.375 ;
        RECT 87.490 19.165 87.820 19.545 ;
        RECT 86.465 18.805 86.845 18.890 ;
        RECT 87.105 18.825 87.820 18.995 ;
        RECT 85.755 18.635 85.955 18.805 ;
        RECT 86.620 18.765 86.845 18.805 ;
        RECT 84.710 18.305 85.585 18.635 ;
        RECT 85.755 18.305 86.505 18.635 ;
        RECT 83.520 17.165 83.770 17.495 ;
        RECT 84.710 17.465 84.880 18.305 ;
        RECT 85.755 18.100 85.945 18.305 ;
        RECT 86.675 18.185 86.845 18.765 ;
        RECT 87.015 18.275 87.370 18.645 ;
        RECT 87.650 18.635 87.820 18.825 ;
        RECT 87.990 18.800 88.245 19.375 ;
        RECT 87.650 18.305 87.905 18.635 ;
        RECT 86.630 18.135 86.845 18.185 ;
        RECT 85.050 17.725 85.945 18.100 ;
        RECT 86.455 18.055 86.845 18.135 ;
        RECT 87.650 18.095 87.820 18.305 ;
        RECT 83.995 17.295 84.880 17.465 ;
        RECT 85.060 16.995 85.375 17.495 ;
        RECT 85.605 17.165 85.945 17.725 ;
        RECT 86.115 16.995 86.285 18.005 ;
        RECT 86.455 17.210 86.785 18.055 ;
        RECT 87.105 17.925 87.820 18.095 ;
        RECT 88.075 18.070 88.245 18.800 ;
        RECT 88.420 18.705 88.680 19.545 ;
        RECT 89.315 18.795 90.525 19.545 ;
        RECT 87.105 17.165 87.275 17.925 ;
        RECT 87.490 16.995 87.820 17.755 ;
        RECT 87.990 17.165 88.245 18.070 ;
        RECT 88.420 16.995 88.680 18.145 ;
        RECT 89.315 18.085 89.835 18.625 ;
        RECT 90.005 18.255 90.525 18.795 ;
        RECT 89.315 16.995 90.525 18.085 ;
        RECT 11.950 16.825 90.610 16.995 ;
        RECT 12.035 15.735 13.245 16.825 ;
        RECT 13.505 16.155 13.675 16.655 ;
        RECT 13.845 16.325 14.175 16.825 ;
        RECT 13.505 15.985 14.170 16.155 ;
        RECT 12.035 15.025 12.555 15.565 ;
        RECT 12.725 15.195 13.245 15.735 ;
        RECT 13.420 15.165 13.770 15.815 ;
        RECT 12.035 14.275 13.245 15.025 ;
        RECT 13.940 14.995 14.170 15.985 ;
        RECT 13.505 14.825 14.170 14.995 ;
        RECT 13.505 14.535 13.675 14.825 ;
        RECT 13.845 14.275 14.175 14.655 ;
        RECT 14.345 14.535 14.530 16.655 ;
        RECT 14.770 16.365 15.035 16.825 ;
        RECT 15.205 16.230 15.455 16.655 ;
        RECT 15.665 16.380 16.770 16.550 ;
        RECT 15.150 16.100 15.455 16.230 ;
        RECT 14.700 14.905 14.980 15.855 ;
        RECT 15.150 14.995 15.320 16.100 ;
        RECT 15.490 15.315 15.730 15.910 ;
        RECT 15.900 15.845 16.430 16.210 ;
        RECT 15.900 15.145 16.070 15.845 ;
        RECT 16.600 15.765 16.770 16.380 ;
        RECT 16.940 16.025 17.110 16.825 ;
        RECT 17.280 16.325 17.530 16.655 ;
        RECT 17.755 16.355 18.640 16.525 ;
        RECT 16.600 15.675 17.110 15.765 ;
        RECT 15.150 14.865 15.375 14.995 ;
        RECT 15.545 14.925 16.070 15.145 ;
        RECT 16.240 15.505 17.110 15.675 ;
        RECT 14.785 14.275 15.035 14.735 ;
        RECT 15.205 14.725 15.375 14.865 ;
        RECT 16.240 14.725 16.410 15.505 ;
        RECT 16.940 15.435 17.110 15.505 ;
        RECT 16.620 15.255 16.820 15.285 ;
        RECT 17.280 15.255 17.450 16.325 ;
        RECT 17.620 15.435 17.810 16.155 ;
        RECT 16.620 14.955 17.450 15.255 ;
        RECT 17.980 15.225 18.300 16.185 ;
        RECT 15.205 14.555 15.540 14.725 ;
        RECT 15.735 14.555 16.410 14.725 ;
        RECT 16.730 14.275 17.100 14.775 ;
        RECT 17.280 14.725 17.450 14.955 ;
        RECT 17.835 14.895 18.300 15.225 ;
        RECT 18.470 15.515 18.640 16.355 ;
        RECT 18.820 16.325 19.135 16.825 ;
        RECT 19.365 16.095 19.705 16.655 ;
        RECT 18.810 15.720 19.705 16.095 ;
        RECT 19.875 15.815 20.045 16.825 ;
        RECT 19.515 15.515 19.705 15.720 ;
        RECT 20.215 15.765 20.545 16.610 ;
        RECT 21.730 16.035 22.265 16.655 ;
        RECT 20.215 15.685 20.605 15.765 ;
        RECT 20.390 15.635 20.605 15.685 ;
        RECT 18.470 15.185 19.345 15.515 ;
        RECT 19.515 15.185 20.265 15.515 ;
        RECT 18.470 14.725 18.640 15.185 ;
        RECT 19.515 15.015 19.715 15.185 ;
        RECT 20.435 15.055 20.605 15.635 ;
        RECT 20.380 15.015 20.605 15.055 ;
        RECT 17.280 14.555 17.685 14.725 ;
        RECT 17.855 14.555 18.640 14.725 ;
        RECT 18.915 14.275 19.125 14.805 ;
        RECT 19.385 14.490 19.715 15.015 ;
        RECT 20.225 14.930 20.605 15.015 ;
        RECT 21.730 15.015 22.045 16.035 ;
        RECT 22.435 16.025 22.765 16.825 ;
        RECT 23.250 15.855 23.640 16.030 ;
        RECT 22.215 15.685 23.640 15.855 ;
        RECT 22.215 15.185 22.385 15.685 ;
        RECT 19.885 14.275 20.055 14.885 ;
        RECT 20.225 14.495 20.555 14.930 ;
        RECT 21.730 14.445 22.345 15.015 ;
        RECT 22.635 14.955 22.900 15.515 ;
        RECT 23.070 14.785 23.240 15.685 ;
        RECT 24.915 15.660 25.205 16.825 ;
        RECT 26.300 15.675 26.560 16.825 ;
        RECT 26.735 15.750 26.990 16.655 ;
        RECT 27.160 16.065 27.490 16.825 ;
        RECT 27.705 15.895 27.875 16.655 ;
        RECT 23.410 14.955 23.765 15.515 ;
        RECT 22.515 14.275 22.730 14.785 ;
        RECT 22.960 14.455 23.240 14.785 ;
        RECT 23.420 14.275 23.660 14.785 ;
        RECT 24.915 14.275 25.205 15.000 ;
        RECT 26.300 14.275 26.560 15.115 ;
        RECT 26.735 15.020 26.905 15.750 ;
        RECT 27.160 15.725 27.875 15.895 ;
        RECT 27.160 15.515 27.330 15.725 ;
        RECT 28.600 15.675 28.860 16.825 ;
        RECT 29.035 15.750 29.290 16.655 ;
        RECT 29.460 16.065 29.790 16.825 ;
        RECT 30.005 15.895 30.175 16.655 ;
        RECT 27.075 15.185 27.330 15.515 ;
        RECT 26.735 14.445 26.990 15.020 ;
        RECT 27.160 14.995 27.330 15.185 ;
        RECT 27.610 15.175 27.965 15.545 ;
        RECT 27.160 14.825 27.875 14.995 ;
        RECT 27.160 14.275 27.490 14.655 ;
        RECT 27.705 14.445 27.875 14.825 ;
        RECT 28.600 14.275 28.860 15.115 ;
        RECT 29.035 15.020 29.205 15.750 ;
        RECT 29.460 15.725 30.175 15.895 ;
        RECT 29.460 15.515 29.630 15.725 ;
        RECT 30.440 15.675 30.700 16.825 ;
        RECT 30.875 15.750 31.130 16.655 ;
        RECT 31.300 16.065 31.630 16.825 ;
        RECT 31.845 15.895 32.015 16.655 ;
        RECT 29.375 15.185 29.630 15.515 ;
        RECT 29.035 14.445 29.290 15.020 ;
        RECT 29.460 14.995 29.630 15.185 ;
        RECT 29.910 15.175 30.265 15.545 ;
        RECT 29.460 14.825 30.175 14.995 ;
        RECT 29.460 14.275 29.790 14.655 ;
        RECT 30.005 14.445 30.175 14.825 ;
        RECT 30.440 14.275 30.700 15.115 ;
        RECT 30.875 15.020 31.045 15.750 ;
        RECT 31.300 15.725 32.015 15.895 ;
        RECT 31.300 15.515 31.470 15.725 ;
        RECT 32.280 15.675 32.540 16.825 ;
        RECT 32.715 15.750 32.970 16.655 ;
        RECT 33.140 16.065 33.470 16.825 ;
        RECT 33.685 15.895 33.855 16.655 ;
        RECT 31.215 15.185 31.470 15.515 ;
        RECT 30.875 14.445 31.130 15.020 ;
        RECT 31.300 14.995 31.470 15.185 ;
        RECT 31.750 15.175 32.105 15.545 ;
        RECT 31.300 14.825 32.015 14.995 ;
        RECT 31.300 14.275 31.630 14.655 ;
        RECT 31.845 14.445 32.015 14.825 ;
        RECT 32.280 14.275 32.540 15.115 ;
        RECT 32.715 15.020 32.885 15.750 ;
        RECT 33.140 15.725 33.855 15.895 ;
        RECT 33.140 15.515 33.310 15.725 ;
        RECT 34.120 15.675 34.380 16.825 ;
        RECT 34.555 15.750 34.810 16.655 ;
        RECT 34.980 16.065 35.310 16.825 ;
        RECT 35.525 15.895 35.695 16.655 ;
        RECT 33.055 15.185 33.310 15.515 ;
        RECT 32.715 14.445 32.970 15.020 ;
        RECT 33.140 14.995 33.310 15.185 ;
        RECT 33.590 15.175 33.945 15.545 ;
        RECT 33.140 14.825 33.855 14.995 ;
        RECT 33.140 14.275 33.470 14.655 ;
        RECT 33.685 14.445 33.855 14.825 ;
        RECT 34.120 14.275 34.380 15.115 ;
        RECT 34.555 15.020 34.725 15.750 ;
        RECT 34.980 15.725 35.695 15.895 ;
        RECT 34.980 15.515 35.150 15.725 ;
        RECT 35.960 15.675 36.220 16.825 ;
        RECT 36.395 15.750 36.650 16.655 ;
        RECT 36.820 16.065 37.150 16.825 ;
        RECT 37.365 15.895 37.535 16.655 ;
        RECT 34.895 15.185 35.150 15.515 ;
        RECT 34.555 14.445 34.810 15.020 ;
        RECT 34.980 14.995 35.150 15.185 ;
        RECT 35.430 15.175 35.785 15.545 ;
        RECT 34.980 14.825 35.695 14.995 ;
        RECT 34.980 14.275 35.310 14.655 ;
        RECT 35.525 14.445 35.695 14.825 ;
        RECT 35.960 14.275 36.220 15.115 ;
        RECT 36.395 15.020 36.565 15.750 ;
        RECT 36.820 15.725 37.535 15.895 ;
        RECT 36.820 15.515 36.990 15.725 ;
        RECT 37.795 15.660 38.085 16.825 ;
        RECT 39.180 16.435 39.515 16.655 ;
        RECT 40.520 16.445 40.875 16.825 ;
        RECT 39.180 15.815 39.435 16.435 ;
        RECT 39.685 16.275 39.915 16.315 ;
        RECT 41.045 16.275 41.295 16.655 ;
        RECT 39.685 16.075 41.295 16.275 ;
        RECT 39.685 15.985 39.870 16.075 ;
        RECT 40.460 16.065 41.295 16.075 ;
        RECT 41.545 16.045 41.795 16.825 ;
        RECT 41.965 15.975 42.225 16.655 ;
        RECT 40.025 15.875 40.355 15.905 ;
        RECT 40.025 15.815 41.825 15.875 ;
        RECT 39.180 15.705 41.885 15.815 ;
        RECT 39.180 15.645 40.355 15.705 ;
        RECT 41.685 15.670 41.885 15.705 ;
        RECT 36.735 15.185 36.990 15.515 ;
        RECT 36.395 14.445 36.650 15.020 ;
        RECT 36.820 14.995 36.990 15.185 ;
        RECT 37.270 15.175 37.625 15.545 ;
        RECT 39.175 15.265 39.665 15.465 ;
        RECT 39.855 15.265 40.330 15.475 ;
        RECT 36.820 14.825 37.535 14.995 ;
        RECT 36.820 14.275 37.150 14.655 ;
        RECT 37.365 14.445 37.535 14.825 ;
        RECT 37.795 14.275 38.085 15.000 ;
        RECT 39.180 14.275 39.635 15.040 ;
        RECT 40.110 14.865 40.330 15.265 ;
        RECT 40.575 15.265 40.905 15.475 ;
        RECT 40.575 14.865 40.785 15.265 ;
        RECT 41.075 15.230 41.485 15.535 ;
        RECT 41.715 15.095 41.885 15.670 ;
        RECT 41.615 14.975 41.885 15.095 ;
        RECT 41.040 14.930 41.885 14.975 ;
        RECT 41.040 14.805 41.795 14.930 ;
        RECT 41.040 14.655 41.210 14.805 ;
        RECT 42.055 14.775 42.225 15.975 ;
        RECT 42.580 15.855 42.970 16.030 ;
        RECT 43.455 16.025 43.785 16.825 ;
        RECT 43.955 16.035 44.490 16.655 ;
        RECT 42.580 15.685 44.005 15.855 ;
        RECT 42.455 14.955 42.810 15.515 ;
        RECT 42.980 14.785 43.150 15.685 ;
        RECT 43.320 14.955 43.585 15.515 ;
        RECT 43.835 15.185 44.005 15.685 ;
        RECT 44.175 15.015 44.490 16.035 ;
        RECT 44.700 15.675 44.960 16.825 ;
        RECT 45.135 15.750 45.390 16.655 ;
        RECT 45.560 16.065 45.890 16.825 ;
        RECT 46.105 15.895 46.275 16.655 ;
        RECT 39.910 14.445 41.210 14.655 ;
        RECT 41.465 14.275 41.795 14.635 ;
        RECT 41.965 14.445 42.225 14.775 ;
        RECT 42.560 14.275 42.800 14.785 ;
        RECT 42.980 14.455 43.260 14.785 ;
        RECT 43.490 14.275 43.705 14.785 ;
        RECT 43.875 14.445 44.490 15.015 ;
        RECT 44.700 14.275 44.960 15.115 ;
        RECT 45.135 15.020 45.305 15.750 ;
        RECT 45.560 15.725 46.275 15.895 ;
        RECT 46.625 15.895 46.795 16.655 ;
        RECT 47.010 16.065 47.340 16.825 ;
        RECT 46.625 15.725 47.340 15.895 ;
        RECT 47.510 15.750 47.765 16.655 ;
        RECT 45.560 15.515 45.730 15.725 ;
        RECT 45.475 15.185 45.730 15.515 ;
        RECT 45.135 14.445 45.390 15.020 ;
        RECT 45.560 14.995 45.730 15.185 ;
        RECT 46.010 15.175 46.365 15.545 ;
        RECT 46.535 15.175 46.890 15.545 ;
        RECT 47.170 15.515 47.340 15.725 ;
        RECT 47.170 15.185 47.425 15.515 ;
        RECT 47.170 14.995 47.340 15.185 ;
        RECT 47.595 15.020 47.765 15.750 ;
        RECT 47.940 15.675 48.200 16.825 ;
        RECT 48.560 15.855 48.950 16.030 ;
        RECT 49.435 16.025 49.765 16.825 ;
        RECT 49.935 16.035 50.470 16.655 ;
        RECT 48.560 15.685 49.985 15.855 ;
        RECT 45.560 14.825 46.275 14.995 ;
        RECT 45.560 14.275 45.890 14.655 ;
        RECT 46.105 14.445 46.275 14.825 ;
        RECT 46.625 14.825 47.340 14.995 ;
        RECT 46.625 14.445 46.795 14.825 ;
        RECT 47.010 14.275 47.340 14.655 ;
        RECT 47.510 14.445 47.765 15.020 ;
        RECT 47.940 14.275 48.200 15.115 ;
        RECT 48.435 14.955 48.790 15.515 ;
        RECT 48.960 14.785 49.130 15.685 ;
        RECT 49.300 14.955 49.565 15.515 ;
        RECT 49.815 15.185 49.985 15.685 ;
        RECT 50.155 15.015 50.470 16.035 ;
        RECT 50.675 15.660 50.965 16.825 ;
        RECT 52.060 15.675 52.320 16.825 ;
        RECT 52.495 15.750 52.750 16.655 ;
        RECT 52.920 16.065 53.250 16.825 ;
        RECT 53.465 15.895 53.635 16.655 ;
        RECT 48.540 14.275 48.780 14.785 ;
        RECT 48.960 14.455 49.240 14.785 ;
        RECT 49.470 14.275 49.685 14.785 ;
        RECT 49.855 14.445 50.470 15.015 ;
        RECT 50.675 14.275 50.965 15.000 ;
        RECT 52.060 14.275 52.320 15.115 ;
        RECT 52.495 15.020 52.665 15.750 ;
        RECT 52.920 15.725 53.635 15.895 ;
        RECT 53.895 15.735 55.105 16.825 ;
        RECT 52.920 15.515 53.090 15.725 ;
        RECT 52.835 15.185 53.090 15.515 ;
        RECT 52.495 14.445 52.750 15.020 ;
        RECT 52.920 14.995 53.090 15.185 ;
        RECT 53.370 15.175 53.725 15.545 ;
        RECT 53.895 15.025 54.415 15.565 ;
        RECT 54.585 15.195 55.105 15.735 ;
        RECT 55.280 15.675 55.540 16.825 ;
        RECT 55.715 15.750 55.970 16.655 ;
        RECT 56.140 16.065 56.470 16.825 ;
        RECT 56.685 15.895 56.855 16.655 ;
        RECT 52.920 14.825 53.635 14.995 ;
        RECT 52.920 14.275 53.250 14.655 ;
        RECT 53.465 14.445 53.635 14.825 ;
        RECT 53.895 14.275 55.105 15.025 ;
        RECT 55.280 14.275 55.540 15.115 ;
        RECT 55.715 15.020 55.885 15.750 ;
        RECT 56.140 15.725 56.855 15.895 ;
        RECT 57.115 15.735 58.325 16.825 ;
        RECT 56.140 15.515 56.310 15.725 ;
        RECT 56.055 15.185 56.310 15.515 ;
        RECT 55.715 14.445 55.970 15.020 ;
        RECT 56.140 14.995 56.310 15.185 ;
        RECT 56.590 15.175 56.945 15.545 ;
        RECT 57.115 15.025 57.635 15.565 ;
        RECT 57.805 15.195 58.325 15.735 ;
        RECT 58.585 15.895 58.755 16.655 ;
        RECT 58.970 16.065 59.300 16.825 ;
        RECT 58.585 15.725 59.300 15.895 ;
        RECT 59.470 15.750 59.725 16.655 ;
        RECT 58.495 15.175 58.850 15.545 ;
        RECT 59.130 15.515 59.300 15.725 ;
        RECT 59.130 15.185 59.385 15.515 ;
        RECT 56.140 14.825 56.855 14.995 ;
        RECT 56.140 14.275 56.470 14.655 ;
        RECT 56.685 14.445 56.855 14.825 ;
        RECT 57.115 14.275 58.325 15.025 ;
        RECT 59.130 14.995 59.300 15.185 ;
        RECT 59.555 15.020 59.725 15.750 ;
        RECT 59.900 15.675 60.160 16.825 ;
        RECT 60.335 15.735 61.545 16.825 ;
        RECT 58.585 14.825 59.300 14.995 ;
        RECT 58.585 14.445 58.755 14.825 ;
        RECT 58.970 14.275 59.300 14.655 ;
        RECT 59.470 14.445 59.725 15.020 ;
        RECT 59.900 14.275 60.160 15.115 ;
        RECT 60.335 15.025 60.855 15.565 ;
        RECT 61.025 15.195 61.545 15.735 ;
        RECT 61.720 15.675 61.980 16.825 ;
        RECT 62.155 15.750 62.410 16.655 ;
        RECT 62.580 16.065 62.910 16.825 ;
        RECT 63.125 15.895 63.295 16.655 ;
        RECT 60.335 14.275 61.545 15.025 ;
        RECT 61.720 14.275 61.980 15.115 ;
        RECT 62.155 15.020 62.325 15.750 ;
        RECT 62.580 15.725 63.295 15.895 ;
        RECT 62.580 15.515 62.750 15.725 ;
        RECT 63.555 15.660 63.845 16.825 ;
        RECT 64.940 15.675 65.200 16.825 ;
        RECT 65.375 15.750 65.630 16.655 ;
        RECT 65.800 16.065 66.130 16.825 ;
        RECT 66.345 15.895 66.515 16.655 ;
        RECT 62.495 15.185 62.750 15.515 ;
        RECT 62.155 14.445 62.410 15.020 ;
        RECT 62.580 14.995 62.750 15.185 ;
        RECT 63.030 15.175 63.385 15.545 ;
        RECT 62.580 14.825 63.295 14.995 ;
        RECT 62.580 14.275 62.910 14.655 ;
        RECT 63.125 14.445 63.295 14.825 ;
        RECT 63.555 14.275 63.845 15.000 ;
        RECT 64.940 14.275 65.200 15.115 ;
        RECT 65.375 15.020 65.545 15.750 ;
        RECT 65.800 15.725 66.515 15.895 ;
        RECT 66.775 15.735 67.985 16.825 ;
        RECT 65.800 15.515 65.970 15.725 ;
        RECT 65.715 15.185 65.970 15.515 ;
        RECT 65.375 14.445 65.630 15.020 ;
        RECT 65.800 14.995 65.970 15.185 ;
        RECT 66.250 15.175 66.605 15.545 ;
        RECT 66.775 15.025 67.295 15.565 ;
        RECT 67.465 15.195 67.985 15.735 ;
        RECT 68.160 15.675 68.420 16.825 ;
        RECT 68.595 15.750 68.850 16.655 ;
        RECT 69.020 16.065 69.350 16.825 ;
        RECT 69.565 15.895 69.735 16.655 ;
        RECT 65.800 14.825 66.515 14.995 ;
        RECT 65.800 14.275 66.130 14.655 ;
        RECT 66.345 14.445 66.515 14.825 ;
        RECT 66.775 14.275 67.985 15.025 ;
        RECT 68.160 14.275 68.420 15.115 ;
        RECT 68.595 15.020 68.765 15.750 ;
        RECT 69.020 15.725 69.735 15.895 ;
        RECT 69.995 15.735 71.205 16.825 ;
        RECT 69.020 15.515 69.190 15.725 ;
        RECT 68.935 15.185 69.190 15.515 ;
        RECT 68.595 14.445 68.850 15.020 ;
        RECT 69.020 14.995 69.190 15.185 ;
        RECT 69.470 15.175 69.825 15.545 ;
        RECT 69.995 15.025 70.515 15.565 ;
        RECT 70.685 15.195 71.205 15.735 ;
        RECT 71.465 15.895 71.635 16.655 ;
        RECT 71.850 16.065 72.180 16.825 ;
        RECT 71.465 15.725 72.180 15.895 ;
        RECT 72.350 15.750 72.605 16.655 ;
        RECT 71.375 15.175 71.730 15.545 ;
        RECT 72.010 15.515 72.180 15.725 ;
        RECT 72.010 15.185 72.265 15.515 ;
        RECT 69.020 14.825 69.735 14.995 ;
        RECT 69.020 14.275 69.350 14.655 ;
        RECT 69.565 14.445 69.735 14.825 ;
        RECT 69.995 14.275 71.205 15.025 ;
        RECT 72.010 14.995 72.180 15.185 ;
        RECT 72.435 15.020 72.605 15.750 ;
        RECT 72.780 15.675 73.040 16.825 ;
        RECT 73.215 15.735 74.425 16.825 ;
        RECT 71.465 14.825 72.180 14.995 ;
        RECT 71.465 14.445 71.635 14.825 ;
        RECT 71.850 14.275 72.180 14.655 ;
        RECT 72.350 14.445 72.605 15.020 ;
        RECT 72.780 14.275 73.040 15.115 ;
        RECT 73.215 15.025 73.735 15.565 ;
        RECT 73.905 15.195 74.425 15.735 ;
        RECT 74.600 15.675 74.860 16.825 ;
        RECT 75.035 15.750 75.290 16.655 ;
        RECT 75.460 16.065 75.790 16.825 ;
        RECT 76.005 15.895 76.175 16.655 ;
        RECT 73.215 14.275 74.425 15.025 ;
        RECT 74.600 14.275 74.860 15.115 ;
        RECT 75.035 15.020 75.205 15.750 ;
        RECT 75.460 15.725 76.175 15.895 ;
        RECT 75.460 15.515 75.630 15.725 ;
        RECT 76.435 15.660 76.725 16.825 ;
        RECT 77.080 15.855 77.470 16.030 ;
        RECT 77.955 16.025 78.285 16.825 ;
        RECT 78.455 16.035 78.990 16.655 ;
        RECT 77.080 15.685 78.505 15.855 ;
        RECT 75.375 15.185 75.630 15.515 ;
        RECT 75.035 14.445 75.290 15.020 ;
        RECT 75.460 14.995 75.630 15.185 ;
        RECT 75.910 15.175 76.265 15.545 ;
        RECT 75.460 14.825 76.175 14.995 ;
        RECT 75.460 14.275 75.790 14.655 ;
        RECT 76.005 14.445 76.175 14.825 ;
        RECT 76.435 14.275 76.725 15.000 ;
        RECT 76.955 14.955 77.310 15.515 ;
        RECT 77.480 14.785 77.650 15.685 ;
        RECT 77.820 14.955 78.085 15.515 ;
        RECT 78.335 15.185 78.505 15.685 ;
        RECT 78.675 15.015 78.990 16.035 ;
        RECT 79.380 15.855 79.770 16.030 ;
        RECT 80.255 16.025 80.585 16.825 ;
        RECT 80.755 16.035 81.290 16.655 ;
        RECT 79.380 15.685 80.805 15.855 ;
        RECT 77.060 14.275 77.300 14.785 ;
        RECT 77.480 14.455 77.760 14.785 ;
        RECT 77.990 14.275 78.205 14.785 ;
        RECT 78.375 14.445 78.990 15.015 ;
        RECT 79.255 14.955 79.610 15.515 ;
        RECT 79.780 14.785 79.950 15.685 ;
        RECT 80.120 14.955 80.385 15.515 ;
        RECT 80.635 15.185 80.805 15.685 ;
        RECT 80.975 15.015 81.290 16.035 ;
        RECT 82.045 16.155 82.215 16.655 ;
        RECT 82.385 16.325 82.715 16.825 ;
        RECT 82.045 15.985 82.710 16.155 ;
        RECT 81.960 15.165 82.310 15.815 ;
        RECT 79.360 14.275 79.600 14.785 ;
        RECT 79.780 14.455 80.060 14.785 ;
        RECT 80.290 14.275 80.505 14.785 ;
        RECT 80.675 14.445 81.290 15.015 ;
        RECT 82.480 14.995 82.710 15.985 ;
        RECT 82.045 14.825 82.710 14.995 ;
        RECT 82.045 14.535 82.215 14.825 ;
        RECT 82.385 14.275 82.715 14.655 ;
        RECT 82.885 14.535 83.070 16.655 ;
        RECT 83.310 16.365 83.575 16.825 ;
        RECT 83.745 16.230 83.995 16.655 ;
        RECT 84.205 16.380 85.310 16.550 ;
        RECT 83.690 16.100 83.995 16.230 ;
        RECT 83.240 14.905 83.520 15.855 ;
        RECT 83.690 14.995 83.860 16.100 ;
        RECT 84.030 15.315 84.270 15.910 ;
        RECT 84.440 15.845 84.970 16.210 ;
        RECT 84.440 15.145 84.610 15.845 ;
        RECT 85.140 15.765 85.310 16.380 ;
        RECT 85.480 16.025 85.650 16.825 ;
        RECT 85.820 16.325 86.070 16.655 ;
        RECT 86.295 16.355 87.180 16.525 ;
        RECT 85.140 15.675 85.650 15.765 ;
        RECT 83.690 14.865 83.915 14.995 ;
        RECT 84.085 14.925 84.610 15.145 ;
        RECT 84.780 15.505 85.650 15.675 ;
        RECT 83.325 14.275 83.575 14.735 ;
        RECT 83.745 14.725 83.915 14.865 ;
        RECT 84.780 14.725 84.950 15.505 ;
        RECT 85.480 15.435 85.650 15.505 ;
        RECT 85.160 15.255 85.360 15.285 ;
        RECT 85.820 15.255 85.990 16.325 ;
        RECT 86.160 15.435 86.350 16.155 ;
        RECT 85.160 14.955 85.990 15.255 ;
        RECT 86.520 15.225 86.840 16.185 ;
        RECT 83.745 14.555 84.080 14.725 ;
        RECT 84.275 14.555 84.950 14.725 ;
        RECT 85.270 14.275 85.640 14.775 ;
        RECT 85.820 14.725 85.990 14.955 ;
        RECT 86.375 14.895 86.840 15.225 ;
        RECT 87.010 15.515 87.180 16.355 ;
        RECT 87.360 16.325 87.675 16.825 ;
        RECT 87.905 16.095 88.245 16.655 ;
        RECT 87.350 15.720 88.245 16.095 ;
        RECT 88.415 15.815 88.585 16.825 ;
        RECT 88.055 15.515 88.245 15.720 ;
        RECT 88.755 15.765 89.085 16.610 ;
        RECT 88.755 15.685 89.145 15.765 ;
        RECT 88.930 15.635 89.145 15.685 ;
        RECT 87.010 15.185 87.885 15.515 ;
        RECT 88.055 15.185 88.805 15.515 ;
        RECT 87.010 14.725 87.180 15.185 ;
        RECT 88.055 15.015 88.255 15.185 ;
        RECT 88.975 15.055 89.145 15.635 ;
        RECT 89.315 15.735 90.525 16.825 ;
        RECT 89.315 15.195 89.835 15.735 ;
        RECT 88.920 15.015 89.145 15.055 ;
        RECT 90.005 15.025 90.525 15.565 ;
        RECT 85.820 14.555 86.225 14.725 ;
        RECT 86.395 14.555 87.180 14.725 ;
        RECT 87.455 14.275 87.665 14.805 ;
        RECT 87.925 14.490 88.255 15.015 ;
        RECT 88.765 14.930 89.145 15.015 ;
        RECT 88.425 14.275 88.595 14.885 ;
        RECT 88.765 14.495 89.095 14.930 ;
        RECT 89.315 14.275 90.525 15.025 ;
        RECT 11.950 14.105 90.610 14.275 ;
      LAYER met1 ;
        RECT 149.710 221.830 149.970 222.150 ;
        RECT 149.150 220.770 149.410 221.090 ;
        RECT 115.800 220.285 116.060 220.605 ;
        RECT 110.950 206.310 111.210 206.630 ;
        RECT 109.950 205.860 110.210 206.180 ;
        RECT 11.950 201.630 90.610 202.110 ;
        RECT 49.740 201.430 50.060 201.490 ;
        RECT 57.575 201.430 57.865 201.475 ;
        RECT 49.740 201.290 57.865 201.430 ;
        RECT 49.740 201.230 50.060 201.290 ;
        RECT 57.575 201.245 57.865 201.290 ;
        RECT 61.240 200.410 61.560 200.470 ;
        RECT 61.715 200.410 62.005 200.455 ;
        RECT 61.240 200.270 62.005 200.410 ;
        RECT 61.240 200.210 61.560 200.270 ;
        RECT 61.715 200.225 62.005 200.270 ;
        RECT 70.900 200.410 71.220 200.470 ;
        RECT 72.295 200.410 72.585 200.455 ;
        RECT 70.900 200.270 72.585 200.410 ;
        RECT 70.900 200.210 71.220 200.270 ;
        RECT 72.295 200.225 72.585 200.270 ;
        RECT 47.440 200.070 47.760 200.130 ;
        RECT 58.495 200.070 58.785 200.115 ;
        RECT 47.440 199.930 58.785 200.070 ;
        RECT 47.440 199.870 47.760 199.930 ;
        RECT 58.495 199.885 58.785 199.930 ;
        RECT 56.640 199.530 56.960 199.790 ;
        RECT 57.495 199.730 57.785 199.775 ;
        RECT 60.320 199.730 60.640 199.790 ;
        RECT 57.495 199.590 60.640 199.730 ;
        RECT 57.495 199.545 57.785 199.590 ;
        RECT 60.320 199.530 60.640 199.590 ;
        RECT 62.635 199.730 62.925 199.775 ;
        RECT 63.080 199.730 63.400 199.790 ;
        RECT 62.635 199.590 63.400 199.730 ;
        RECT 62.635 199.545 62.925 199.590 ;
        RECT 63.080 199.530 63.400 199.590 ;
        RECT 69.520 199.730 69.840 199.790 ;
        RECT 71.375 199.730 71.665 199.775 ;
        RECT 69.520 199.590 71.665 199.730 ;
        RECT 69.520 199.530 69.840 199.590 ;
        RECT 71.375 199.545 71.665 199.590 ;
        RECT 11.950 198.910 90.610 199.390 ;
        RECT 44.235 198.525 44.525 198.755 ;
        RECT 56.640 198.710 56.960 198.770 ;
        RECT 56.640 198.570 57.330 198.710 ;
        RECT 41.460 198.370 41.780 198.430 ;
        RECT 43.300 198.415 43.620 198.430 ;
        RECT 42.395 198.370 42.685 198.415 ;
        RECT 41.460 198.230 42.685 198.370 ;
        RECT 41.460 198.170 41.780 198.230 ;
        RECT 42.395 198.185 42.685 198.230 ;
        RECT 43.300 198.185 43.685 198.415 ;
        RECT 44.310 198.370 44.450 198.525 ;
        RECT 56.640 198.510 56.960 198.570 ;
        RECT 57.190 198.415 57.330 198.570 ;
        RECT 45.920 198.370 46.210 198.415 ;
        RECT 44.310 198.230 46.210 198.370 ;
        RECT 45.920 198.185 46.210 198.230 ;
        RECT 57.070 198.185 57.360 198.415 ;
        RECT 41.000 197.830 41.320 198.090 ;
        RECT 41.920 197.830 42.240 198.090 ;
        RECT 42.470 198.030 42.610 198.185 ;
        RECT 43.300 198.170 43.620 198.185 ;
        RECT 47.440 198.030 47.760 198.090 ;
        RECT 42.470 197.890 47.760 198.030 ;
        RECT 47.440 197.830 47.760 197.890 ;
        RECT 69.980 198.030 70.300 198.090 ;
        RECT 71.880 198.030 72.170 198.075 ;
        RECT 69.980 197.890 72.170 198.030 ;
        RECT 69.980 197.830 70.300 197.890 ;
        RECT 71.880 197.845 72.170 197.890 ;
        RECT 36.860 197.690 37.180 197.750 ;
        RECT 44.695 197.690 44.985 197.735 ;
        RECT 36.860 197.550 44.985 197.690 ;
        RECT 36.860 197.490 37.180 197.550 ;
        RECT 44.695 197.505 44.985 197.550 ;
        RECT 45.575 197.690 45.865 197.735 ;
        RECT 46.765 197.690 47.055 197.735 ;
        RECT 49.285 197.690 49.575 197.735 ;
        RECT 45.575 197.550 49.575 197.690 ;
        RECT 45.575 197.505 45.865 197.550 ;
        RECT 46.765 197.505 47.055 197.550 ;
        RECT 49.285 197.505 49.575 197.550 ;
        RECT 55.260 197.690 55.580 197.750 ;
        RECT 55.735 197.690 56.025 197.735 ;
        RECT 55.260 197.550 56.025 197.690 ;
        RECT 55.260 197.490 55.580 197.550 ;
        RECT 55.735 197.505 56.025 197.550 ;
        RECT 56.615 197.690 56.905 197.735 ;
        RECT 57.805 197.690 58.095 197.735 ;
        RECT 60.325 197.690 60.615 197.735 ;
        RECT 56.615 197.550 60.615 197.690 ;
        RECT 56.615 197.505 56.905 197.550 ;
        RECT 57.805 197.505 58.095 197.550 ;
        RECT 60.325 197.505 60.615 197.550 ;
        RECT 68.625 197.690 68.915 197.735 ;
        RECT 71.145 197.690 71.435 197.735 ;
        RECT 72.335 197.690 72.625 197.735 ;
        RECT 68.625 197.550 72.625 197.690 ;
        RECT 68.625 197.505 68.915 197.550 ;
        RECT 71.145 197.505 71.435 197.550 ;
        RECT 72.335 197.505 72.625 197.550 ;
        RECT 73.215 197.690 73.505 197.735 ;
        RECT 75.960 197.690 76.280 197.750 ;
        RECT 73.215 197.550 76.280 197.690 ;
        RECT 73.215 197.505 73.505 197.550 ;
        RECT 75.960 197.490 76.280 197.550 ;
        RECT 45.180 197.350 45.470 197.395 ;
        RECT 47.280 197.350 47.570 197.395 ;
        RECT 48.850 197.350 49.140 197.395 ;
        RECT 45.180 197.210 49.140 197.350 ;
        RECT 45.180 197.165 45.470 197.210 ;
        RECT 47.280 197.165 47.570 197.210 ;
        RECT 48.850 197.165 49.140 197.210 ;
        RECT 56.220 197.350 56.510 197.395 ;
        RECT 58.320 197.350 58.610 197.395 ;
        RECT 59.890 197.350 60.180 197.395 ;
        RECT 56.220 197.210 60.180 197.350 ;
        RECT 56.220 197.165 56.510 197.210 ;
        RECT 58.320 197.165 58.610 197.210 ;
        RECT 59.890 197.165 60.180 197.210 ;
        RECT 69.060 197.350 69.350 197.395 ;
        RECT 70.630 197.350 70.920 197.395 ;
        RECT 72.730 197.350 73.020 197.395 ;
        RECT 69.060 197.210 73.020 197.350 ;
        RECT 69.060 197.165 69.350 197.210 ;
        RECT 70.630 197.165 70.920 197.210 ;
        RECT 72.730 197.165 73.020 197.210 ;
        RECT 41.920 196.810 42.240 197.070 ;
        RECT 43.315 197.010 43.605 197.055 ;
        RECT 46.060 197.010 46.380 197.070 ;
        RECT 43.315 196.870 46.380 197.010 ;
        RECT 43.315 196.825 43.605 196.870 ;
        RECT 46.060 196.810 46.380 196.870 ;
        RECT 47.900 197.010 48.220 197.070 ;
        RECT 51.595 197.010 51.885 197.055 ;
        RECT 47.900 196.870 51.885 197.010 ;
        RECT 47.900 196.810 48.220 196.870 ;
        RECT 51.595 196.825 51.885 196.870 ;
        RECT 61.700 197.010 62.020 197.070 ;
        RECT 62.635 197.010 62.925 197.055 ;
        RECT 61.700 196.870 62.925 197.010 ;
        RECT 61.700 196.810 62.020 196.870 ;
        RECT 62.635 196.825 62.925 196.870 ;
        RECT 66.315 197.010 66.605 197.055 ;
        RECT 66.760 197.010 67.080 197.070 ;
        RECT 66.315 196.870 67.080 197.010 ;
        RECT 66.315 196.825 66.605 196.870 ;
        RECT 66.760 196.810 67.080 196.870 ;
        RECT 11.950 196.190 90.610 196.670 ;
        RECT 45.140 195.990 45.460 196.050 ;
        RECT 45.615 195.990 45.905 196.035 ;
        RECT 45.140 195.850 45.905 195.990 ;
        RECT 45.140 195.790 45.460 195.850 ;
        RECT 45.615 195.805 45.905 195.850 ;
        RECT 46.060 195.990 46.380 196.050 ;
        RECT 49.295 195.990 49.585 196.035 ;
        RECT 49.740 195.990 50.060 196.050 ;
        RECT 46.060 195.850 50.060 195.990 ;
        RECT 46.060 195.790 46.380 195.850 ;
        RECT 49.295 195.805 49.585 195.850 ;
        RECT 49.740 195.790 50.060 195.850 ;
        RECT 60.320 195.790 60.640 196.050 ;
        RECT 66.775 195.990 67.065 196.035 ;
        RECT 67.220 195.990 67.540 196.050 ;
        RECT 66.775 195.850 67.540 195.990 ;
        RECT 66.775 195.805 67.065 195.850 ;
        RECT 67.220 195.790 67.540 195.850 ;
        RECT 67.695 195.990 67.985 196.035 ;
        RECT 69.980 195.990 70.300 196.050 ;
        RECT 67.695 195.850 70.300 195.990 ;
        RECT 67.695 195.805 67.985 195.850 ;
        RECT 69.980 195.790 70.300 195.850 ;
        RECT 37.360 195.650 37.650 195.695 ;
        RECT 39.460 195.650 39.750 195.695 ;
        RECT 41.030 195.650 41.320 195.695 ;
        RECT 37.360 195.510 41.320 195.650 ;
        RECT 37.360 195.465 37.650 195.510 ;
        RECT 39.460 195.465 39.750 195.510 ;
        RECT 41.030 195.465 41.320 195.510 ;
        RECT 43.300 195.650 43.620 195.710 ;
        RECT 46.995 195.650 47.285 195.695 ;
        RECT 43.300 195.510 47.285 195.650 ;
        RECT 43.300 195.450 43.620 195.510 ;
        RECT 46.995 195.465 47.285 195.510 ;
        RECT 51.620 195.650 51.910 195.695 ;
        RECT 53.720 195.650 54.010 195.695 ;
        RECT 55.290 195.650 55.580 195.695 ;
        RECT 51.620 195.510 55.580 195.650 ;
        RECT 51.620 195.465 51.910 195.510 ;
        RECT 53.720 195.465 54.010 195.510 ;
        RECT 55.290 195.465 55.580 195.510 ;
        RECT 71.820 195.650 72.110 195.695 ;
        RECT 73.390 195.650 73.680 195.695 ;
        RECT 75.490 195.650 75.780 195.695 ;
        RECT 71.820 195.510 75.780 195.650 ;
        RECT 71.820 195.465 72.110 195.510 ;
        RECT 73.390 195.465 73.680 195.510 ;
        RECT 75.490 195.465 75.780 195.510 ;
        RECT 36.860 195.110 37.180 195.370 ;
        RECT 37.755 195.310 38.045 195.355 ;
        RECT 38.945 195.310 39.235 195.355 ;
        RECT 41.465 195.310 41.755 195.355 ;
        RECT 52.015 195.310 52.305 195.355 ;
        RECT 53.205 195.310 53.495 195.355 ;
        RECT 55.725 195.310 56.015 195.355 ;
        RECT 62.175 195.310 62.465 195.355 ;
        RECT 37.755 195.170 41.755 195.310 ;
        RECT 37.755 195.125 38.045 195.170 ;
        RECT 38.945 195.125 39.235 195.170 ;
        RECT 41.465 195.125 41.755 195.170 ;
        RECT 44.770 195.170 48.130 195.310 ;
        RECT 38.210 194.630 38.500 194.675 ;
        RECT 39.620 194.630 39.940 194.690 ;
        RECT 38.210 194.490 39.940 194.630 ;
        RECT 38.210 194.445 38.500 194.490 ;
        RECT 39.620 194.430 39.940 194.490 ;
        RECT 44.770 194.350 44.910 195.170 ;
        RECT 46.980 194.770 47.300 195.030 ;
        RECT 47.990 195.015 48.130 195.170 ;
        RECT 52.015 195.170 56.015 195.310 ;
        RECT 52.015 195.125 52.305 195.170 ;
        RECT 53.205 195.125 53.495 195.170 ;
        RECT 55.725 195.125 56.015 195.170 ;
        RECT 60.410 195.170 62.465 195.310 ;
        RECT 47.915 194.785 48.205 195.015 ;
        RECT 48.820 194.970 49.140 195.030 ;
        RECT 51.135 194.970 51.425 195.015 ;
        RECT 55.260 194.970 55.580 195.030 ;
        RECT 48.820 194.830 55.580 194.970 ;
        RECT 48.820 194.770 49.140 194.830 ;
        RECT 51.135 194.785 51.425 194.830 ;
        RECT 55.260 194.770 55.580 194.830 ;
        RECT 59.400 194.770 59.720 195.030 ;
        RECT 60.410 195.015 60.550 195.170 ;
        RECT 62.175 195.125 62.465 195.170 ;
        RECT 71.385 195.310 71.675 195.355 ;
        RECT 73.905 195.310 74.195 195.355 ;
        RECT 75.095 195.310 75.385 195.355 ;
        RECT 71.385 195.170 75.385 195.310 ;
        RECT 71.385 195.125 71.675 195.170 ;
        RECT 73.905 195.125 74.195 195.170 ;
        RECT 75.095 195.125 75.385 195.170 ;
        RECT 75.960 195.110 76.280 195.370 ;
        RECT 60.335 194.785 60.625 195.015 ;
        RECT 61.700 194.770 62.020 195.030 ;
        RECT 62.635 194.970 62.925 195.015 ;
        RECT 64.000 194.970 64.320 195.030 ;
        RECT 64.475 194.970 64.765 195.015 ;
        RECT 62.635 194.830 64.765 194.970 ;
        RECT 62.635 194.785 62.925 194.830 ;
        RECT 64.000 194.770 64.320 194.830 ;
        RECT 64.475 194.785 64.765 194.830 ;
        RECT 65.395 194.970 65.685 195.015 ;
        RECT 67.220 194.970 67.540 195.030 ;
        RECT 65.395 194.830 67.540 194.970 ;
        RECT 65.395 194.785 65.685 194.830 ;
        RECT 67.220 194.770 67.540 194.830 ;
        RECT 46.535 194.445 46.825 194.675 ;
        RECT 47.440 194.630 47.760 194.690 ;
        RECT 48.375 194.630 48.665 194.675 ;
        RECT 52.360 194.630 52.650 194.675 ;
        RECT 47.440 194.490 48.665 194.630 ;
        RECT 43.775 194.290 44.065 194.335 ;
        RECT 44.220 194.290 44.540 194.350 ;
        RECT 43.775 194.150 44.540 194.290 ;
        RECT 43.775 194.105 44.065 194.150 ;
        RECT 44.220 194.090 44.540 194.150 ;
        RECT 44.680 194.090 45.000 194.350 ;
        RECT 45.600 194.335 45.920 194.350 ;
        RECT 45.535 194.105 45.920 194.335 ;
        RECT 46.610 194.290 46.750 194.445 ;
        RECT 47.440 194.430 47.760 194.490 ;
        RECT 48.375 194.445 48.665 194.490 ;
        RECT 50.290 194.490 52.650 194.630 ;
        RECT 47.900 194.290 48.220 194.350 ;
        RECT 46.610 194.150 48.220 194.290 ;
        RECT 45.600 194.090 45.920 194.105 ;
        RECT 47.900 194.090 48.220 194.150 ;
        RECT 49.280 194.335 49.600 194.350 ;
        RECT 50.290 194.335 50.430 194.490 ;
        RECT 52.360 194.445 52.650 194.490 ;
        RECT 65.840 194.430 66.160 194.690 ;
        RECT 71.820 194.630 72.140 194.690 ;
        RECT 74.640 194.630 74.930 194.675 ;
        RECT 71.820 194.490 74.930 194.630 ;
        RECT 71.820 194.430 72.140 194.490 ;
        RECT 74.640 194.445 74.930 194.490 ;
        RECT 49.280 194.105 49.665 194.335 ;
        RECT 50.215 194.105 50.505 194.335 ;
        RECT 49.280 194.090 49.600 194.105 ;
        RECT 58.020 194.090 58.340 194.350 ;
        RECT 64.935 194.290 65.225 194.335 ;
        RECT 66.855 194.290 67.145 194.335 ;
        RECT 64.935 194.150 67.145 194.290 ;
        RECT 64.935 194.105 65.225 194.150 ;
        RECT 66.855 194.105 67.145 194.150 ;
        RECT 68.140 194.290 68.460 194.350 ;
        RECT 69.075 194.290 69.365 194.335 ;
        RECT 68.140 194.150 69.365 194.290 ;
        RECT 68.140 194.090 68.460 194.150 ;
        RECT 69.075 194.105 69.365 194.150 ;
        RECT 11.950 193.470 90.610 193.950 ;
        RECT 39.620 193.070 39.940 193.330 ;
        RECT 40.475 193.270 40.765 193.315 ;
        RECT 41.920 193.270 42.240 193.330 ;
        RECT 40.475 193.130 42.240 193.270 ;
        RECT 40.475 193.085 40.765 193.130 ;
        RECT 41.920 193.070 42.240 193.130 ;
        RECT 42.380 193.070 42.700 193.330 ;
        RECT 44.680 193.070 45.000 193.330 ;
        RECT 46.980 193.315 47.300 193.330 ;
        RECT 46.980 193.270 47.315 193.315 ;
        RECT 46.815 193.130 47.315 193.270 ;
        RECT 46.980 193.085 47.315 193.130 ;
        RECT 47.455 193.270 47.745 193.315 ;
        RECT 50.200 193.270 50.520 193.330 ;
        RECT 56.180 193.270 56.500 193.330 ;
        RECT 58.020 193.270 58.340 193.330 ;
        RECT 47.455 193.130 58.340 193.270 ;
        RECT 47.455 193.085 47.745 193.130 ;
        RECT 46.980 193.070 47.300 193.085 ;
        RECT 50.200 193.070 50.520 193.130 ;
        RECT 56.180 193.070 56.500 193.130 ;
        RECT 58.020 193.070 58.340 193.130 ;
        RECT 59.400 193.270 59.720 193.330 ;
        RECT 66.775 193.270 67.065 193.315 ;
        RECT 59.400 193.130 67.065 193.270 ;
        RECT 59.400 193.070 59.720 193.130 ;
        RECT 66.775 193.085 67.065 193.130 ;
        RECT 67.680 193.270 68.000 193.330 ;
        RECT 69.995 193.270 70.285 193.315 ;
        RECT 67.680 193.130 70.285 193.270 ;
        RECT 67.680 193.070 68.000 193.130 ;
        RECT 69.995 193.085 70.285 193.130 ;
        RECT 71.820 193.070 72.140 193.330 ;
        RECT 41.460 192.730 41.780 192.990 ;
        RECT 44.770 192.930 44.910 193.070 ;
        RECT 42.010 192.790 44.910 192.930 ;
        RECT 45.155 192.930 45.445 192.975 ;
        RECT 45.600 192.930 45.920 192.990 ;
        RECT 45.155 192.790 48.130 192.930 ;
        RECT 42.010 192.635 42.150 192.790 ;
        RECT 45.155 192.745 45.445 192.790 ;
        RECT 45.600 192.730 45.920 192.790 ;
        RECT 41.935 192.405 42.225 192.635 ;
        RECT 42.855 192.590 43.145 192.635 ;
        RECT 44.220 192.590 44.540 192.650 ;
        RECT 42.855 192.450 44.540 192.590 ;
        RECT 42.855 192.405 43.145 192.450 ;
        RECT 44.220 192.390 44.540 192.450 ;
        RECT 44.680 192.390 45.000 192.650 ;
        RECT 47.990 192.635 48.130 192.790 ;
        RECT 50.200 192.635 50.520 192.650 ;
        RECT 46.535 192.590 46.825 192.635 ;
        RECT 47.915 192.590 48.205 192.635 ;
        RECT 50.200 192.590 50.540 192.635 ;
        RECT 46.535 192.450 47.210 192.590 ;
        RECT 46.535 192.405 46.825 192.450 ;
        RECT 43.315 191.910 43.605 191.955 ;
        RECT 47.070 191.910 47.210 192.450 ;
        RECT 47.915 192.450 49.925 192.590 ;
        RECT 47.915 192.405 48.205 192.450 ;
        RECT 48.375 192.250 48.665 192.295 ;
        RECT 49.280 192.250 49.600 192.310 ;
        RECT 48.375 192.110 49.600 192.250 ;
        RECT 49.785 192.250 49.925 192.450 ;
        RECT 50.200 192.450 50.715 192.590 ;
        RECT 50.200 192.405 50.540 192.450 ;
        RECT 50.200 192.390 50.520 192.405 ;
        RECT 50.675 192.250 50.965 192.295 ;
        RECT 59.490 192.250 59.630 193.070 ;
        RECT 62.635 192.930 62.925 192.975 ;
        RECT 69.520 192.930 69.840 192.990 ;
        RECT 62.635 192.790 69.840 192.930 ;
        RECT 62.635 192.745 62.925 192.790 ;
        RECT 69.520 192.730 69.840 192.790 ;
        RECT 70.915 192.930 71.205 192.975 ;
        RECT 74.135 192.930 74.425 192.975 ;
        RECT 70.915 192.790 74.425 192.930 ;
        RECT 70.915 192.745 71.205 192.790 ;
        RECT 74.135 192.745 74.425 192.790 ;
        RECT 61.700 192.590 62.020 192.650 ;
        RECT 64.015 192.590 64.305 192.635 ;
        RECT 64.935 192.590 65.225 192.635 ;
        RECT 61.700 192.450 64.305 192.590 ;
        RECT 61.700 192.390 62.020 192.450 ;
        RECT 64.015 192.405 64.305 192.450 ;
        RECT 64.550 192.450 65.225 192.590 ;
        RECT 49.785 192.110 59.630 192.250 ;
        RECT 62.620 192.250 62.940 192.310 ;
        RECT 64.550 192.250 64.690 192.450 ;
        RECT 64.935 192.405 65.225 192.450 ;
        RECT 65.395 192.405 65.685 192.635 ;
        RECT 65.855 192.405 66.145 192.635 ;
        RECT 66.760 192.590 67.080 192.650 ;
        RECT 67.235 192.590 67.525 192.635 ;
        RECT 66.760 192.450 67.525 192.590 ;
        RECT 65.470 192.250 65.610 192.405 ;
        RECT 62.620 192.110 64.690 192.250 ;
        RECT 65.010 192.110 65.610 192.250 ;
        RECT 65.930 192.250 66.070 192.405 ;
        RECT 66.760 192.390 67.080 192.450 ;
        RECT 67.235 192.405 67.525 192.450 ;
        RECT 68.140 192.390 68.460 192.650 ;
        RECT 68.615 192.590 68.905 192.635 ;
        RECT 68.615 192.450 69.290 192.590 ;
        RECT 68.615 192.405 68.905 192.450 ;
        RECT 69.150 192.250 69.290 192.450 ;
        RECT 70.440 192.390 70.760 192.650 ;
        RECT 72.295 192.405 72.585 192.635 ;
        RECT 69.520 192.250 69.840 192.310 ;
        RECT 72.370 192.250 72.510 192.405 ;
        RECT 73.200 192.390 73.520 192.650 ;
        RECT 110.010 192.545 110.150 205.860 ;
        RECT 111.010 201.530 111.150 206.310 ;
        RECT 111.360 205.830 111.620 206.150 ;
        RECT 111.420 202.635 111.560 205.830 ;
        RECT 111.330 202.375 111.650 202.635 ;
        RECT 111.010 201.390 111.640 201.530 ;
        RECT 111.500 198.530 111.640 201.390 ;
        RECT 111.410 198.200 111.740 198.530 ;
        RECT 65.930 192.110 72.510 192.250 ;
        RECT 109.950 192.225 110.210 192.545 ;
        RECT 48.375 192.065 48.665 192.110 ;
        RECT 49.280 192.050 49.600 192.110 ;
        RECT 50.675 192.065 50.965 192.110 ;
        RECT 62.620 192.050 62.940 192.110 ;
        RECT 65.010 191.970 65.150 192.110 ;
        RECT 69.520 192.050 69.840 192.110 ;
        RECT 47.900 191.910 48.220 191.970 ;
        RECT 43.315 191.770 48.220 191.910 ;
        RECT 43.315 191.725 43.605 191.770 ;
        RECT 47.900 191.710 48.220 191.770 ;
        RECT 64.920 191.710 65.240 191.970 ;
        RECT 67.220 191.710 67.540 191.970 ;
        RECT 69.075 191.910 69.365 191.955 ;
        RECT 68.460 191.770 69.365 191.910 ;
        RECT 40.540 191.370 40.860 191.630 ;
        RECT 41.000 191.570 41.320 191.630 ;
        RECT 46.075 191.570 46.365 191.615 ;
        RECT 41.000 191.430 46.365 191.570 ;
        RECT 41.000 191.370 41.320 191.430 ;
        RECT 46.075 191.385 46.365 191.430 ;
        RECT 60.780 191.570 61.100 191.630 ;
        RECT 61.255 191.570 61.545 191.615 ;
        RECT 60.780 191.430 61.545 191.570 ;
        RECT 60.780 191.370 61.100 191.430 ;
        RECT 61.255 191.385 61.545 191.430 ;
        RECT 62.160 191.570 62.480 191.630 ;
        RECT 65.840 191.570 66.160 191.630 ;
        RECT 68.460 191.570 68.600 191.770 ;
        RECT 69.075 191.725 69.365 191.770 ;
        RECT 62.160 191.430 68.600 191.570 ;
        RECT 62.160 191.370 62.480 191.430 ;
        RECT 65.840 191.370 66.160 191.430 ;
        RECT 11.950 190.750 90.610 191.230 ;
        RECT 40.540 190.550 40.860 190.610 ;
        RECT 41.015 190.550 41.305 190.595 ;
        RECT 49.740 190.550 50.060 190.610 ;
        RECT 40.540 190.410 50.060 190.550 ;
        RECT 40.540 190.350 40.860 190.410 ;
        RECT 41.015 190.365 41.305 190.410 ;
        RECT 49.740 190.350 50.060 190.410 ;
        RECT 64.000 190.350 64.320 190.610 ;
        RECT 64.920 190.350 65.240 190.610 ;
        RECT 69.995 190.550 70.285 190.595 ;
        RECT 70.440 190.550 70.760 190.610 ;
        RECT 69.995 190.410 70.760 190.550 ;
        RECT 69.995 190.365 70.285 190.410 ;
        RECT 70.440 190.350 70.760 190.410 ;
        RECT 57.115 190.210 57.405 190.255 ;
        RECT 59.400 190.210 59.720 190.270 ;
        RECT 57.115 190.070 59.720 190.210 ;
        RECT 57.115 190.025 57.405 190.070 ;
        RECT 59.400 190.010 59.720 190.070 ;
        RECT 60.780 190.210 61.100 190.270 ;
        RECT 60.780 190.070 63.310 190.210 ;
        RECT 60.780 190.010 61.100 190.070 ;
        RECT 63.170 189.915 63.310 190.070 ;
        RECT 59.875 189.870 60.165 189.915 ;
        RECT 56.270 189.730 59.170 189.870 ;
        RECT 56.270 189.590 56.410 189.730 ;
        RECT 41.460 189.330 41.780 189.590 ;
        RECT 55.720 189.330 56.040 189.590 ;
        RECT 56.180 189.330 56.500 189.590 ;
        RECT 59.030 189.575 59.170 189.730 ;
        RECT 59.875 189.730 61.930 189.870 ;
        RECT 59.875 189.685 60.165 189.730 ;
        RECT 61.790 189.590 61.930 189.730 ;
        RECT 63.095 189.685 63.385 189.915 ;
        RECT 64.920 189.870 65.240 189.930 ;
        RECT 68.140 189.870 68.460 189.930 ;
        RECT 64.920 189.730 70.670 189.870 ;
        RECT 64.920 189.670 65.240 189.730 ;
        RECT 68.140 189.670 68.460 189.730 ;
        RECT 58.495 189.530 58.785 189.575 ;
        RECT 56.730 189.390 58.785 189.530 ;
        RECT 41.550 189.190 41.690 189.330 ;
        RECT 41.935 189.190 42.225 189.235 ;
        RECT 41.550 189.050 42.225 189.190 ;
        RECT 55.810 189.190 55.950 189.330 ;
        RECT 56.730 189.190 56.870 189.390 ;
        RECT 58.495 189.345 58.785 189.390 ;
        RECT 58.955 189.345 59.245 189.575 ;
        RECT 60.320 189.330 60.640 189.590 ;
        RECT 61.700 189.330 62.020 189.590 ;
        RECT 62.620 189.330 62.940 189.590 ;
        RECT 69.520 189.530 69.840 189.590 ;
        RECT 70.530 189.575 70.670 189.730 ;
        RECT 65.470 189.390 69.840 189.530 ;
        RECT 55.810 189.050 56.870 189.190 ;
        RECT 57.115 189.190 57.405 189.235 ;
        RECT 60.795 189.190 61.085 189.235 ;
        RECT 57.115 189.050 61.085 189.190 ;
        RECT 41.935 189.005 42.225 189.050 ;
        RECT 57.115 189.005 57.405 189.050 ;
        RECT 60.795 189.005 61.085 189.050 ;
        RECT 64.855 189.190 65.145 189.235 ;
        RECT 65.470 189.190 65.610 189.390 ;
        RECT 69.520 189.330 69.840 189.390 ;
        RECT 70.455 189.530 70.745 189.575 ;
        RECT 73.200 189.530 73.520 189.590 ;
        RECT 70.455 189.390 73.520 189.530 ;
        RECT 70.455 189.345 70.745 189.390 ;
        RECT 73.200 189.330 73.520 189.390 ;
        RECT 64.855 189.050 65.610 189.190 ;
        RECT 65.855 189.190 66.145 189.235 ;
        RECT 66.760 189.190 67.080 189.250 ;
        RECT 65.855 189.050 67.080 189.190 ;
        RECT 69.610 189.190 69.750 189.330 ;
        RECT 71.360 189.190 71.680 189.250 ;
        RECT 69.610 189.050 71.680 189.190 ;
        RECT 64.855 189.005 65.145 189.050 ;
        RECT 65.855 189.005 66.145 189.050 ;
        RECT 40.080 188.650 40.400 188.910 ;
        RECT 40.935 188.850 41.225 188.895 ;
        RECT 41.460 188.850 41.780 188.910 ;
        RECT 40.935 188.710 41.780 188.850 ;
        RECT 40.935 188.665 41.225 188.710 ;
        RECT 41.460 188.650 41.780 188.710 ;
        RECT 56.640 188.850 56.960 188.910 ;
        RECT 57.575 188.850 57.865 188.895 ;
        RECT 56.640 188.710 57.865 188.850 ;
        RECT 56.640 188.650 56.960 188.710 ;
        RECT 57.575 188.665 57.865 188.710 ;
        RECT 62.620 188.850 62.940 188.910 ;
        RECT 65.930 188.850 66.070 189.005 ;
        RECT 66.760 188.990 67.080 189.050 ;
        RECT 71.360 188.990 71.680 189.050 ;
        RECT 62.620 188.710 66.070 188.850 ;
        RECT 62.620 188.650 62.940 188.710 ;
        RECT 11.950 188.030 90.610 188.510 ;
        RECT 55.735 187.830 56.025 187.875 ;
        RECT 56.180 187.830 56.500 187.890 ;
        RECT 55.735 187.690 56.500 187.830 ;
        RECT 55.735 187.645 56.025 187.690 ;
        RECT 56.180 187.630 56.500 187.690 ;
        RECT 21.220 187.535 21.540 187.550 ;
        RECT 21.155 187.305 21.540 187.535 ;
        RECT 22.155 187.305 22.445 187.535 ;
        RECT 39.590 187.490 39.880 187.535 ;
        RECT 40.080 187.490 40.400 187.550 ;
        RECT 39.590 187.350 40.400 187.490 ;
        RECT 39.590 187.305 39.880 187.350 ;
        RECT 21.220 187.290 21.540 187.305 ;
        RECT 16.620 186.810 16.940 186.870 ;
        RECT 22.230 186.810 22.370 187.305 ;
        RECT 40.080 187.290 40.400 187.350 ;
        RECT 51.580 187.490 51.900 187.550 ;
        RECT 62.160 187.490 62.480 187.550 ;
        RECT 51.580 187.350 62.480 187.490 ;
        RECT 51.580 187.290 51.900 187.350 ;
        RECT 62.160 187.290 62.480 187.350 ;
        RECT 26.740 187.150 27.060 187.210 ;
        RECT 27.575 187.150 27.865 187.195 ;
        RECT 26.740 187.010 27.865 187.150 ;
        RECT 26.740 186.950 27.060 187.010 ;
        RECT 27.575 186.965 27.865 187.010 ;
        RECT 36.860 187.150 37.180 187.210 ;
        RECT 38.255 187.150 38.545 187.195 ;
        RECT 36.860 187.010 38.545 187.150 ;
        RECT 36.860 186.950 37.180 187.010 ;
        RECT 38.255 186.965 38.545 187.010 ;
        RECT 55.275 186.965 55.565 187.195 ;
        RECT 16.620 186.670 22.370 186.810 ;
        RECT 24.440 186.810 24.760 186.870 ;
        RECT 26.295 186.810 26.585 186.855 ;
        RECT 24.440 186.670 26.585 186.810 ;
        RECT 16.620 186.610 16.940 186.670 ;
        RECT 24.440 186.610 24.760 186.670 ;
        RECT 26.295 186.625 26.585 186.670 ;
        RECT 27.175 186.810 27.465 186.855 ;
        RECT 28.365 186.810 28.655 186.855 ;
        RECT 30.885 186.810 31.175 186.855 ;
        RECT 27.175 186.670 31.175 186.810 ;
        RECT 27.175 186.625 27.465 186.670 ;
        RECT 28.365 186.625 28.655 186.670 ;
        RECT 30.885 186.625 31.175 186.670 ;
        RECT 39.135 186.810 39.425 186.855 ;
        RECT 40.325 186.810 40.615 186.855 ;
        RECT 42.845 186.810 43.135 186.855 ;
        RECT 39.135 186.670 43.135 186.810 ;
        RECT 55.350 186.810 55.490 186.965 ;
        RECT 56.640 186.950 56.960 187.210 ;
        RECT 58.480 187.150 58.800 187.210 ;
        RECT 59.415 187.150 59.705 187.195 ;
        RECT 58.480 187.010 59.705 187.150 ;
        RECT 58.480 186.950 58.800 187.010 ;
        RECT 59.415 186.965 59.705 187.010 ;
        RECT 59.875 187.150 60.165 187.195 ;
        RECT 62.620 187.150 62.940 187.210 ;
        RECT 59.875 187.010 62.940 187.150 ;
        RECT 59.875 186.965 60.165 187.010 ;
        RECT 62.620 186.950 62.940 187.010 ;
        RECT 55.720 186.810 56.040 186.870 ;
        RECT 57.560 186.810 57.880 186.870 ;
        RECT 55.350 186.670 57.880 186.810 ;
        RECT 39.135 186.625 39.425 186.670 ;
        RECT 40.325 186.625 40.615 186.670 ;
        RECT 42.845 186.625 43.135 186.670 ;
        RECT 55.720 186.610 56.040 186.670 ;
        RECT 57.560 186.610 57.880 186.670 ;
        RECT 60.795 186.810 61.085 186.855 ;
        RECT 64.920 186.810 65.240 186.870 ;
        RECT 60.795 186.670 65.240 186.810 ;
        RECT 60.795 186.625 61.085 186.670 ;
        RECT 64.920 186.610 65.240 186.670 ;
        RECT 26.780 186.470 27.070 186.515 ;
        RECT 28.880 186.470 29.170 186.515 ;
        RECT 30.450 186.470 30.740 186.515 ;
        RECT 26.780 186.330 30.740 186.470 ;
        RECT 26.780 186.285 27.070 186.330 ;
        RECT 28.880 186.285 29.170 186.330 ;
        RECT 30.450 186.285 30.740 186.330 ;
        RECT 38.740 186.470 39.030 186.515 ;
        RECT 40.840 186.470 41.130 186.515 ;
        RECT 42.410 186.470 42.700 186.515 ;
        RECT 38.740 186.330 42.700 186.470 ;
        RECT 38.740 186.285 39.030 186.330 ;
        RECT 40.840 186.285 41.130 186.330 ;
        RECT 42.410 186.285 42.700 186.330 ;
        RECT 46.060 186.470 46.380 186.530 ;
        RECT 47.440 186.470 47.760 186.530 ;
        RECT 67.220 186.470 67.540 186.530 ;
        RECT 46.060 186.330 67.540 186.470 ;
        RECT 46.060 186.270 46.380 186.330 ;
        RECT 47.440 186.270 47.760 186.330 ;
        RECT 67.220 186.270 67.540 186.330 ;
        RECT 20.300 185.930 20.620 186.190 ;
        RECT 21.235 186.130 21.525 186.175 ;
        RECT 26.280 186.130 26.600 186.190 ;
        RECT 21.235 185.990 26.600 186.130 ;
        RECT 21.235 185.945 21.525 185.990 ;
        RECT 26.280 185.930 26.600 185.990 ;
        RECT 33.180 185.930 33.500 186.190 ;
        RECT 42.840 186.130 43.160 186.190 ;
        RECT 45.155 186.130 45.445 186.175 ;
        RECT 42.840 185.990 45.445 186.130 ;
        RECT 42.840 185.930 43.160 185.990 ;
        RECT 45.155 185.945 45.445 185.990 ;
        RECT 56.655 186.130 56.945 186.175 ;
        RECT 58.940 186.130 59.260 186.190 ;
        RECT 56.655 185.990 59.260 186.130 ;
        RECT 56.655 185.945 56.945 185.990 ;
        RECT 58.940 185.930 59.260 185.990 ;
        RECT 60.320 185.930 60.640 186.190 ;
        RECT 11.950 185.310 90.610 185.790 ;
        RECT 16.620 184.910 16.940 185.170 ;
        RECT 26.295 185.110 26.585 185.155 ;
        RECT 26.740 185.110 27.060 185.170 ;
        RECT 26.295 184.970 27.060 185.110 ;
        RECT 26.295 184.925 26.585 184.970 ;
        RECT 26.740 184.910 27.060 184.970 ;
        RECT 27.200 184.910 27.520 185.170 ;
        RECT 36.875 185.110 37.165 185.155 ;
        RECT 27.750 184.970 37.165 185.110 ;
        RECT 20.300 184.770 20.590 184.815 ;
        RECT 21.870 184.770 22.160 184.815 ;
        RECT 23.970 184.770 24.260 184.815 ;
        RECT 20.300 184.630 24.260 184.770 ;
        RECT 20.300 184.585 20.590 184.630 ;
        RECT 21.870 184.585 22.160 184.630 ;
        RECT 23.970 184.585 24.260 184.630 ;
        RECT 19.865 184.430 20.155 184.475 ;
        RECT 22.385 184.430 22.675 184.475 ;
        RECT 23.575 184.430 23.865 184.475 ;
        RECT 19.865 184.290 23.865 184.430 ;
        RECT 19.865 184.245 20.155 184.290 ;
        RECT 22.385 184.245 22.675 184.290 ;
        RECT 23.575 184.245 23.865 184.290 ;
        RECT 16.175 183.905 16.465 184.135 ;
        RECT 16.250 183.750 16.390 183.905 ;
        RECT 17.080 183.890 17.400 184.150 ;
        RECT 20.300 184.090 20.620 184.150 ;
        RECT 23.120 184.090 23.410 184.135 ;
        RECT 20.300 183.950 23.410 184.090 ;
        RECT 20.300 183.890 20.620 183.950 ;
        RECT 23.120 183.905 23.410 183.950 ;
        RECT 24.440 183.890 24.760 184.150 ;
        RECT 27.135 183.750 27.425 183.795 ;
        RECT 27.750 183.750 27.890 184.970 ;
        RECT 36.875 184.925 37.165 184.970 ;
        RECT 41.460 184.910 41.780 185.170 ;
        RECT 56.640 185.110 56.960 185.170 ;
        RECT 63.540 185.110 63.860 185.170 ;
        RECT 56.640 184.970 63.860 185.110 ;
        RECT 56.640 184.910 56.960 184.970 ;
        RECT 29.590 184.630 35.250 184.770 ;
        RECT 29.040 184.090 29.360 184.150 ;
        RECT 29.590 184.135 29.730 184.630 ;
        RECT 29.960 184.430 30.280 184.490 ;
        RECT 29.960 184.290 32.950 184.430 ;
        RECT 29.960 184.230 30.280 184.290 ;
        RECT 29.515 184.090 29.805 184.135 ;
        RECT 29.040 183.950 29.805 184.090 ;
        RECT 29.040 183.890 29.360 183.950 ;
        RECT 29.515 183.905 29.805 183.950 ;
        RECT 30.420 183.890 30.740 184.150 ;
        RECT 30.880 183.890 31.200 184.150 ;
        RECT 32.810 184.135 32.950 184.290 ;
        RECT 32.735 184.090 33.025 184.135 ;
        RECT 33.180 184.090 33.500 184.150 ;
        RECT 32.735 183.950 33.500 184.090 ;
        RECT 33.730 184.100 33.870 184.630 ;
        RECT 35.110 184.430 35.250 184.630 ;
        RECT 40.095 184.430 40.385 184.475 ;
        RECT 41.000 184.430 41.320 184.490 ;
        RECT 35.110 184.290 38.470 184.430 ;
        RECT 34.115 184.100 34.405 184.135 ;
        RECT 33.730 183.960 34.405 184.100 ;
        RECT 32.735 183.905 33.025 183.950 ;
        RECT 33.180 183.890 33.500 183.950 ;
        RECT 34.115 183.905 34.405 183.960 ;
        RECT 34.560 183.890 34.880 184.150 ;
        RECT 35.110 184.090 35.250 184.290 ;
        RECT 35.495 184.090 35.785 184.135 ;
        RECT 35.110 183.950 35.785 184.090 ;
        RECT 35.495 183.905 35.785 183.950 ;
        RECT 35.940 183.890 36.260 184.150 ;
        RECT 38.330 184.135 38.470 184.290 ;
        RECT 40.095 184.290 41.320 184.430 ;
        RECT 40.095 184.245 40.385 184.290 ;
        RECT 41.000 184.230 41.320 184.290 ;
        RECT 36.875 184.090 37.165 184.135 ;
        RECT 36.875 183.950 38.010 184.090 ;
        RECT 36.875 183.905 37.165 183.950 ;
        RECT 16.250 183.610 17.770 183.750 ;
        RECT 17.630 183.455 17.770 183.610 ;
        RECT 27.135 183.610 27.890 183.750 ;
        RECT 28.135 183.750 28.425 183.795 ;
        RECT 31.815 183.750 32.105 183.795 ;
        RECT 32.260 183.750 32.580 183.810 ;
        RECT 28.135 183.610 32.580 183.750 ;
        RECT 33.270 183.750 33.410 183.890 ;
        RECT 37.335 183.750 37.625 183.795 ;
        RECT 33.270 183.610 37.625 183.750 ;
        RECT 27.135 183.565 27.425 183.610 ;
        RECT 28.135 183.565 28.425 183.610 ;
        RECT 31.815 183.565 32.105 183.610 ;
        RECT 32.260 183.550 32.580 183.610 ;
        RECT 37.335 183.565 37.625 183.610 ;
        RECT 17.555 183.410 17.845 183.455 ;
        RECT 22.600 183.410 22.920 183.470 ;
        RECT 17.555 183.270 22.920 183.410 ;
        RECT 17.555 183.225 17.845 183.270 ;
        RECT 22.600 183.210 22.920 183.270 ;
        RECT 28.595 183.410 28.885 183.455 ;
        RECT 29.500 183.410 29.820 183.470 ;
        RECT 28.595 183.270 29.820 183.410 ;
        RECT 28.595 183.225 28.885 183.270 ;
        RECT 29.500 183.210 29.820 183.270 ;
        RECT 31.340 183.410 31.660 183.470 ;
        RECT 33.180 183.410 33.500 183.470 ;
        RECT 33.655 183.410 33.945 183.455 ;
        RECT 37.870 183.410 38.010 183.950 ;
        RECT 38.255 183.905 38.545 184.135 ;
        RECT 39.635 184.090 39.925 184.135 ;
        RECT 42.380 184.090 42.700 184.150 ;
        RECT 39.635 183.950 42.700 184.090 ;
        RECT 39.635 183.905 39.925 183.950 ;
        RECT 42.380 183.890 42.700 183.950 ;
        RECT 52.040 183.890 52.360 184.150 ;
        RECT 53.435 184.090 53.725 184.135 ;
        RECT 56.180 184.090 56.500 184.150 ;
        RECT 58.110 184.135 58.250 184.970 ;
        RECT 63.540 184.910 63.860 184.970 ;
        RECT 67.220 185.110 67.540 185.170 ;
        RECT 67.695 185.110 67.985 185.155 ;
        RECT 67.220 184.970 67.985 185.110 ;
        RECT 67.220 184.910 67.540 184.970 ;
        RECT 67.695 184.925 67.985 184.970 ;
        RECT 59.415 184.770 59.705 184.815 ;
        RECT 60.320 184.770 60.640 184.830 ;
        RECT 59.415 184.630 60.640 184.770 ;
        RECT 59.415 184.585 59.705 184.630 ;
        RECT 60.320 184.570 60.640 184.630 ;
        RECT 66.760 184.770 67.080 184.830 ;
        RECT 69.075 184.770 69.365 184.815 ;
        RECT 66.760 184.630 69.365 184.770 ;
        RECT 66.760 184.570 67.080 184.630 ;
        RECT 69.075 184.585 69.365 184.630 ;
        RECT 71.820 184.770 72.110 184.815 ;
        RECT 73.390 184.770 73.680 184.815 ;
        RECT 75.490 184.770 75.780 184.815 ;
        RECT 71.820 184.630 75.780 184.770 ;
        RECT 71.820 184.585 72.110 184.630 ;
        RECT 73.390 184.585 73.680 184.630 ;
        RECT 75.490 184.585 75.780 184.630 ;
        RECT 61.330 184.290 63.310 184.430 ;
        RECT 53.435 183.950 56.500 184.090 ;
        RECT 53.435 183.905 53.725 183.950 ;
        RECT 56.180 183.890 56.500 183.950 ;
        RECT 58.035 183.905 58.325 184.135 ;
        RECT 58.955 184.090 59.245 184.135 ;
        RECT 59.400 184.090 59.720 184.150 ;
        RECT 58.955 183.950 59.720 184.090 ;
        RECT 58.955 183.905 59.245 183.950 ;
        RECT 59.400 183.890 59.720 183.950 ;
        RECT 59.875 183.905 60.165 184.135 ;
        RECT 60.335 184.100 60.625 184.135 ;
        RECT 61.330 184.100 61.470 184.290 ;
        RECT 60.335 183.960 61.470 184.100 ;
        RECT 62.160 184.090 62.480 184.150 ;
        RECT 62.635 184.090 62.925 184.135 ;
        RECT 60.335 183.905 60.625 183.960 ;
        RECT 62.160 183.950 62.925 184.090 ;
        RECT 63.170 184.090 63.310 184.290 ;
        RECT 63.540 184.230 63.860 184.490 ;
        RECT 71.385 184.430 71.675 184.475 ;
        RECT 73.905 184.430 74.195 184.475 ;
        RECT 75.095 184.430 75.385 184.475 ;
        RECT 71.385 184.290 75.385 184.430 ;
        RECT 71.385 184.245 71.675 184.290 ;
        RECT 73.905 184.245 74.195 184.290 ;
        RECT 75.095 184.245 75.385 184.290 ;
        RECT 75.960 184.230 76.280 184.490 ;
        RECT 63.170 183.950 63.770 184.090 ;
        RECT 41.920 183.750 42.240 183.810 ;
        RECT 46.535 183.750 46.825 183.795 ;
        RECT 41.920 183.610 46.825 183.750 ;
        RECT 41.920 183.550 42.240 183.610 ;
        RECT 46.535 183.565 46.825 183.610 ;
        RECT 49.280 183.750 49.600 183.810 ;
        RECT 52.975 183.750 53.265 183.795 ;
        RECT 49.280 183.610 53.265 183.750 ;
        RECT 59.950 183.750 60.090 183.905 ;
        RECT 62.160 183.890 62.480 183.950 ;
        RECT 62.635 183.905 62.925 183.950 ;
        RECT 63.080 183.750 63.400 183.810 ;
        RECT 59.950 183.610 63.400 183.750 ;
        RECT 63.630 183.750 63.770 183.950 ;
        RECT 64.000 183.890 64.320 184.150 ;
        RECT 65.855 184.090 66.145 184.135 ;
        RECT 71.820 184.090 72.140 184.150 ;
        RECT 65.855 183.950 72.140 184.090 ;
        RECT 65.855 183.905 66.145 183.950 ;
        RECT 71.820 183.890 72.140 183.950 ;
        RECT 64.475 183.750 64.765 183.795 ;
        RECT 63.630 183.610 64.765 183.750 ;
        RECT 49.280 183.550 49.600 183.610 ;
        RECT 52.975 183.565 53.265 183.610 ;
        RECT 63.080 183.550 63.400 183.610 ;
        RECT 64.475 183.565 64.765 183.610 ;
        RECT 70.440 183.750 70.760 183.810 ;
        RECT 74.640 183.750 74.930 183.795 ;
        RECT 70.440 183.610 74.930 183.750 ;
        RECT 70.440 183.550 70.760 183.610 ;
        RECT 74.640 183.565 74.930 183.610 ;
        RECT 31.340 183.270 38.010 183.410 ;
        RECT 43.760 183.410 44.080 183.470 ;
        RECT 46.075 183.410 46.365 183.455 ;
        RECT 47.440 183.410 47.760 183.470 ;
        RECT 43.760 183.270 47.760 183.410 ;
        RECT 31.340 183.210 31.660 183.270 ;
        RECT 33.180 183.210 33.500 183.270 ;
        RECT 33.655 183.225 33.945 183.270 ;
        RECT 43.760 183.210 44.080 183.270 ;
        RECT 46.075 183.225 46.365 183.270 ;
        RECT 47.440 183.210 47.760 183.270 ;
        RECT 51.135 183.410 51.425 183.455 ;
        RECT 51.580 183.410 51.900 183.470 ;
        RECT 51.135 183.270 51.900 183.410 ;
        RECT 51.135 183.225 51.425 183.270 ;
        RECT 51.580 183.210 51.900 183.270 ;
        RECT 59.400 183.410 59.720 183.470 ;
        RECT 61.255 183.410 61.545 183.455 ;
        RECT 59.400 183.270 61.545 183.410 ;
        RECT 59.400 183.210 59.720 183.270 ;
        RECT 61.255 183.225 61.545 183.270 ;
        RECT 61.700 183.210 62.020 183.470 ;
        RECT 67.680 183.210 68.000 183.470 ;
        RECT 68.600 183.210 68.920 183.470 ;
        RECT 11.950 182.590 90.610 183.070 ;
        RECT 20.775 182.390 21.065 182.435 ;
        RECT 21.220 182.390 21.540 182.450 ;
        RECT 20.775 182.250 21.540 182.390 ;
        RECT 20.775 182.205 21.065 182.250 ;
        RECT 21.220 182.190 21.540 182.250 ;
        RECT 30.420 182.390 30.740 182.450 ;
        RECT 32.720 182.390 33.040 182.450 ;
        RECT 34.100 182.390 34.420 182.450 ;
        RECT 30.420 182.250 31.110 182.390 ;
        RECT 30.420 182.190 30.740 182.250 ;
        RECT 22.600 182.050 22.920 182.110 ;
        RECT 29.040 182.050 29.360 182.110 ;
        RECT 30.970 182.095 31.110 182.250 ;
        RECT 32.720 182.250 34.420 182.390 ;
        RECT 32.720 182.190 33.040 182.250 ;
        RECT 34.100 182.190 34.420 182.250 ;
        RECT 41.935 182.390 42.225 182.435 ;
        RECT 47.915 182.390 48.205 182.435 ;
        RECT 41.935 182.250 48.205 182.390 ;
        RECT 41.935 182.205 42.225 182.250 ;
        RECT 47.915 182.205 48.205 182.250 ;
        RECT 49.280 182.190 49.600 182.450 ;
        RECT 51.135 182.390 51.425 182.435 ;
        RECT 52.040 182.390 52.360 182.450 ;
        RECT 51.135 182.250 52.360 182.390 ;
        RECT 51.135 182.205 51.425 182.250 ;
        RECT 52.040 182.190 52.360 182.250 ;
        RECT 56.180 182.190 56.500 182.450 ;
        RECT 57.560 182.390 57.880 182.450 ;
        RECT 63.095 182.390 63.385 182.435 ;
        RECT 64.000 182.390 64.320 182.450 ;
        RECT 57.560 182.250 62.390 182.390 ;
        RECT 57.560 182.190 57.880 182.250 ;
        RECT 29.975 182.050 30.265 182.095 ;
        RECT 22.600 181.910 30.265 182.050 ;
        RECT 22.600 181.850 22.920 181.910 ;
        RECT 29.040 181.850 29.360 181.910 ;
        RECT 29.975 181.865 30.265 181.910 ;
        RECT 30.895 182.050 31.185 182.095 ;
        RECT 42.855 182.050 43.145 182.095 ;
        RECT 48.500 182.050 48.790 182.095 ;
        RECT 30.895 181.910 35.250 182.050 ;
        RECT 30.895 181.865 31.185 181.910 ;
        RECT 35.110 181.770 35.250 181.910 ;
        RECT 42.855 181.910 48.790 182.050 ;
        RECT 49.370 182.050 49.510 182.190 ;
        RECT 58.020 182.050 58.340 182.110 ;
        RECT 61.700 182.050 62.020 182.110 ;
        RECT 49.370 181.910 54.570 182.050 ;
        RECT 42.855 181.865 43.145 181.910 ;
        RECT 48.500 181.865 48.790 181.910 ;
        RECT 17.080 181.710 17.400 181.770 ;
        RECT 21.695 181.710 21.985 181.755 ;
        RECT 17.080 181.570 21.985 181.710 ;
        RECT 17.080 181.510 17.400 181.570 ;
        RECT 21.695 181.525 21.985 181.570 ;
        RECT 21.770 181.370 21.910 181.525 ;
        RECT 30.420 181.510 30.740 181.770 ;
        RECT 33.655 181.525 33.945 181.755 ;
        RECT 31.815 181.370 32.105 181.415 ;
        RECT 33.180 181.370 33.500 181.430 ;
        RECT 21.770 181.230 33.500 181.370 ;
        RECT 33.730 181.370 33.870 181.525 ;
        RECT 34.100 181.510 34.420 181.770 ;
        RECT 34.560 181.510 34.880 181.770 ;
        RECT 35.020 181.510 35.340 181.770 ;
        RECT 40.080 181.510 40.400 181.770 ;
        RECT 42.380 181.510 42.700 181.770 ;
        RECT 43.315 181.710 43.605 181.755 ;
        RECT 43.760 181.710 44.080 181.770 ;
        RECT 43.315 181.570 44.080 181.710 ;
        RECT 43.315 181.525 43.605 181.570 ;
        RECT 43.760 181.510 44.080 181.570 ;
        RECT 44.695 181.525 44.985 181.755 ;
        RECT 45.615 181.710 45.905 181.755 ;
        RECT 47.455 181.710 47.745 181.755 ;
        RECT 45.615 181.570 47.745 181.710 ;
        RECT 45.615 181.525 45.905 181.570 ;
        RECT 47.455 181.525 47.745 181.570 ;
        RECT 49.755 181.710 50.045 181.755 ;
        RECT 49.755 181.570 50.890 181.710 ;
        RECT 49.755 181.525 50.045 181.570 ;
        RECT 36.400 181.370 36.720 181.430 ;
        RECT 39.635 181.370 39.925 181.415 ;
        RECT 33.730 181.230 39.925 181.370 ;
        RECT 42.470 181.370 42.610 181.510 ;
        RECT 44.770 181.370 44.910 181.525 ;
        RECT 42.470 181.230 44.910 181.370 ;
        RECT 31.815 181.185 32.105 181.230 ;
        RECT 33.180 181.170 33.500 181.230 ;
        RECT 36.400 181.170 36.720 181.230 ;
        RECT 39.635 181.185 39.925 181.230 ;
        RECT 27.200 180.690 27.520 180.750 ;
        RECT 29.055 180.690 29.345 180.735 ;
        RECT 29.960 180.690 30.280 180.750 ;
        RECT 27.200 180.550 30.280 180.690 ;
        RECT 27.200 180.490 27.520 180.550 ;
        RECT 29.055 180.505 29.345 180.550 ;
        RECT 29.960 180.490 30.280 180.550 ;
        RECT 32.735 180.690 33.025 180.735 ;
        RECT 33.180 180.690 33.500 180.750 ;
        RECT 32.735 180.550 33.500 180.690 ;
        RECT 44.770 180.690 44.910 181.230 ;
        RECT 46.075 181.370 46.365 181.415 ;
        RECT 46.520 181.370 46.840 181.430 ;
        RECT 46.075 181.230 46.840 181.370 ;
        RECT 47.530 181.370 47.670 181.525 ;
        RECT 50.215 181.370 50.505 181.415 ;
        RECT 47.530 181.230 50.505 181.370 ;
        RECT 46.075 181.185 46.365 181.230 ;
        RECT 46.520 181.170 46.840 181.230 ;
        RECT 50.215 181.185 50.505 181.230 ;
        RECT 45.600 181.030 45.920 181.090 ;
        RECT 50.750 181.030 50.890 181.570 ;
        RECT 52.515 181.525 52.805 181.755 ;
        RECT 53.435 181.710 53.725 181.755 ;
        RECT 53.880 181.710 54.200 181.770 ;
        RECT 54.430 181.755 54.570 181.910 ;
        RECT 58.020 181.910 62.020 182.050 ;
        RECT 62.250 182.050 62.390 182.250 ;
        RECT 63.095 182.250 64.320 182.390 ;
        RECT 63.095 182.205 63.385 182.250 ;
        RECT 64.000 182.190 64.320 182.250 ;
        RECT 71.820 182.390 72.140 182.450 ;
        RECT 76.435 182.390 76.725 182.435 ;
        RECT 100.970 182.410 102.630 184.070 ;
        RECT 112.120 183.415 112.600 219.295 ;
        RECT 113.420 207.865 113.680 208.185 ;
        RECT 112.755 206.960 112.985 207.250 ;
        RECT 112.800 205.425 112.940 206.960 ;
        RECT 112.740 205.105 113.000 205.425 ;
        RECT 112.755 204.660 112.985 204.950 ;
        RECT 112.800 202.665 112.940 204.660 ;
        RECT 113.435 203.955 113.665 204.030 ;
        RECT 113.435 203.815 114.640 203.955 ;
        RECT 113.435 203.740 113.665 203.815 ;
        RECT 113.435 203.280 113.665 203.570 ;
        RECT 113.480 203.125 113.620 203.280 ;
        RECT 113.420 202.805 113.680 203.125 ;
        RECT 114.115 202.795 114.345 203.085 ;
        RECT 112.740 202.345 113.000 202.665 ;
        RECT 113.775 202.400 114.005 202.690 ;
        RECT 113.095 201.945 113.325 202.235 ;
        RECT 113.140 200.825 113.280 201.945 ;
        RECT 113.820 201.500 113.960 202.400 ;
        RECT 113.775 201.210 114.005 201.500 ;
        RECT 113.080 200.505 113.340 200.825 ;
        RECT 113.820 198.980 113.960 201.210 ;
        RECT 114.160 200.985 114.300 202.795 ;
        RECT 114.115 200.695 114.345 200.985 ;
        RECT 114.160 199.415 114.300 200.695 ;
        RECT 114.115 199.125 114.345 199.415 ;
        RECT 113.775 198.690 114.005 198.980 ;
        RECT 112.740 198.435 113.000 198.525 ;
        RECT 112.740 198.295 113.280 198.435 ;
        RECT 112.740 198.205 113.000 198.295 ;
        RECT 112.755 195.675 112.985 195.750 ;
        RECT 113.140 195.675 113.280 198.295 ;
        RECT 114.500 198.065 114.640 203.815 ;
        RECT 114.440 197.745 114.700 198.065 ;
        RECT 114.115 196.380 114.345 196.670 ;
        RECT 112.755 195.535 113.280 195.675 ;
        RECT 112.755 195.460 112.985 195.535 ;
        RECT 114.160 194.845 114.300 196.380 ;
        RECT 113.420 194.525 113.680 194.845 ;
        RECT 114.100 194.525 114.360 194.845 ;
        RECT 112.740 192.225 113.000 192.545 ;
        RECT 112.800 191.150 112.940 192.225 ;
        RECT 113.420 191.765 113.680 192.085 ;
        RECT 112.755 190.860 112.985 191.150 ;
        RECT 114.455 189.940 114.685 190.230 ;
        RECT 113.760 189.465 114.020 189.785 ;
        RECT 113.420 189.005 113.680 189.325 ;
        RECT 113.820 187.930 113.960 189.465 ;
        RECT 114.100 188.545 114.360 188.865 ;
        RECT 113.775 187.640 114.005 187.930 ;
        RECT 114.160 186.550 114.300 188.545 ;
        RECT 114.500 188.405 114.640 189.940 ;
        RECT 114.440 188.085 114.700 188.405 ;
        RECT 114.115 186.260 114.345 186.550 ;
        RECT 114.440 185.785 114.700 186.105 ;
        RECT 114.500 185.630 114.640 185.785 ;
        RECT 114.455 185.340 114.685 185.630 ;
        RECT 114.840 183.415 115.320 219.295 ;
        RECT 115.860 217.370 116.000 220.285 ;
        RECT 148.630 220.050 148.950 220.310 ;
        RECT 148.140 219.570 148.400 219.890 ;
        RECT 116.480 217.525 116.740 217.845 ;
        RECT 115.815 217.080 116.045 217.370 ;
        RECT 116.540 216.450 116.680 217.525 ;
        RECT 116.495 216.160 116.725 216.450 ;
        RECT 117.160 214.765 117.420 215.085 ;
        RECT 117.160 212.925 117.420 213.245 ;
        RECT 117.160 212.465 117.420 212.785 ;
        RECT 116.155 211.560 116.385 211.850 ;
        RECT 116.200 206.345 116.340 211.560 ;
        RECT 117.160 210.165 117.420 210.485 ;
        RECT 117.220 208.185 117.360 210.165 ;
        RECT 117.160 207.865 117.420 208.185 ;
        RECT 116.140 206.025 116.400 206.345 ;
        RECT 117.220 205.870 117.360 207.865 ;
        RECT 117.175 205.580 117.405 205.870 ;
        RECT 116.155 203.270 116.385 203.560 ;
        RECT 115.815 202.835 116.045 203.125 ;
        RECT 115.860 201.555 116.000 202.835 ;
        RECT 115.815 201.265 116.045 201.555 ;
        RECT 115.460 200.505 115.720 200.825 ;
        RECT 115.520 198.510 115.660 200.505 ;
        RECT 115.860 199.455 116.000 201.265 ;
        RECT 116.200 201.040 116.340 203.270 ;
        RECT 117.160 201.655 117.420 201.745 ;
        RECT 116.540 201.515 117.420 201.655 ;
        RECT 116.155 200.750 116.385 201.040 ;
        RECT 116.200 199.850 116.340 200.750 ;
        RECT 116.540 200.305 116.680 201.515 ;
        RECT 117.160 201.425 117.420 201.515 ;
        RECT 116.820 200.505 117.080 200.825 ;
        RECT 116.495 200.015 116.725 200.305 ;
        RECT 116.155 199.560 116.385 199.850 ;
        RECT 115.815 199.165 116.045 199.455 ;
        RECT 116.495 198.895 116.725 198.970 ;
        RECT 116.880 198.895 117.020 200.505 ;
        RECT 116.495 198.755 117.020 198.895 ;
        RECT 116.495 198.680 116.725 198.755 ;
        RECT 115.475 198.220 115.705 198.510 ;
        RECT 116.495 196.380 116.725 196.670 ;
        RECT 116.140 194.985 116.400 195.305 ;
        RECT 116.140 194.525 116.400 194.845 ;
        RECT 116.200 190.230 116.340 194.525 ;
        RECT 116.540 192.990 116.680 196.380 ;
        RECT 117.160 195.905 117.420 196.225 ;
        RECT 116.495 192.700 116.725 192.990 ;
        RECT 116.155 189.940 116.385 190.230 ;
        RECT 116.140 189.465 116.400 189.785 ;
        RECT 116.200 188.390 116.340 189.465 ;
        RECT 116.480 189.005 116.740 189.325 ;
        RECT 116.155 188.100 116.385 188.390 ;
        RECT 116.155 187.640 116.385 187.930 ;
        RECT 116.200 185.185 116.340 187.640 ;
        RECT 116.540 187.010 116.680 189.005 ;
        RECT 116.495 186.720 116.725 187.010 ;
        RECT 117.160 186.245 117.420 186.565 ;
        RECT 117.220 186.090 117.360 186.245 ;
        RECT 117.175 185.800 117.405 186.090 ;
        RECT 116.140 184.865 116.400 185.185 ;
        RECT 117.560 183.415 118.040 219.295 ;
        RECT 119.880 217.525 120.140 217.845 ;
        RECT 119.215 215.230 119.445 215.520 ;
        RECT 118.520 214.765 118.780 215.085 ;
        RECT 118.580 212.265 118.720 214.765 ;
        RECT 119.260 213.000 119.400 215.230 ;
        RECT 119.555 214.795 119.785 215.085 ;
        RECT 119.600 213.515 119.740 214.795 ;
        RECT 119.555 213.225 119.785 213.515 ;
        RECT 119.215 212.710 119.445 213.000 ;
        RECT 118.535 211.975 118.765 212.265 ;
        RECT 119.260 211.810 119.400 212.710 ;
        RECT 119.215 211.520 119.445 211.810 ;
        RECT 119.600 211.415 119.740 213.225 ;
        RECT 119.555 211.125 119.785 211.415 ;
        RECT 119.200 210.625 119.460 210.945 ;
        RECT 118.875 205.580 119.105 205.870 ;
        RECT 118.920 201.285 119.060 205.580 ;
        RECT 118.860 200.965 119.120 201.285 ;
        RECT 119.880 200.505 120.140 200.825 ;
        RECT 119.940 199.430 120.080 200.505 ;
        RECT 119.895 199.140 120.125 199.430 ;
        RECT 118.875 195.215 119.105 195.290 ;
        RECT 118.875 195.075 119.400 195.215 ;
        RECT 118.875 195.000 119.105 195.075 ;
        RECT 118.860 193.605 119.120 193.925 ;
        RECT 118.195 192.915 118.425 192.990 ;
        RECT 118.195 192.775 118.720 192.915 ;
        RECT 118.195 192.700 118.425 192.775 ;
        RECT 118.195 189.940 118.425 190.230 ;
        RECT 118.240 189.785 118.380 189.940 ;
        RECT 118.180 189.465 118.440 189.785 ;
        RECT 118.580 189.695 118.720 192.775 ;
        RECT 118.860 192.225 119.120 192.545 ;
        RECT 118.860 190.845 119.120 191.165 ;
        RECT 118.875 189.695 119.105 189.770 ;
        RECT 118.580 189.555 119.105 189.695 ;
        RECT 118.180 189.005 118.440 189.325 ;
        RECT 118.580 187.395 118.720 189.555 ;
        RECT 118.875 189.480 119.105 189.555 ;
        RECT 118.875 188.560 119.105 188.850 ;
        RECT 118.920 188.405 119.060 188.560 ;
        RECT 118.860 188.085 119.120 188.405 ;
        RECT 118.860 187.395 119.120 187.485 ;
        RECT 118.580 187.255 119.120 187.395 ;
        RECT 118.860 187.165 119.120 187.255 ;
        RECT 118.860 185.785 119.120 186.105 ;
        RECT 119.260 185.645 119.400 195.075 ;
        RECT 119.555 194.080 119.785 194.370 ;
        RECT 119.600 188.865 119.740 194.080 ;
        RECT 119.895 191.320 120.125 191.610 ;
        RECT 119.940 189.325 120.080 191.320 ;
        RECT 119.880 189.005 120.140 189.325 ;
        RECT 119.540 188.545 119.800 188.865 ;
        RECT 119.895 188.100 120.125 188.390 ;
        RECT 119.940 187.945 120.080 188.100 ;
        RECT 119.880 187.625 120.140 187.945 ;
        RECT 119.200 185.325 119.460 185.645 ;
        RECT 118.860 184.865 119.120 185.185 ;
        RECT 120.280 183.415 120.760 219.295 ;
        RECT 121.240 217.985 121.500 218.305 ;
        RECT 121.300 217.370 121.440 217.985 ;
        RECT 121.580 217.525 121.840 217.845 ;
        RECT 121.255 217.080 121.485 217.370 ;
        RECT 121.640 215.070 121.780 217.525 ;
        RECT 121.935 216.160 122.165 216.450 ;
        RECT 121.595 214.780 121.825 215.070 ;
        RECT 120.900 212.925 121.160 213.245 ;
        RECT 120.960 211.850 121.100 212.925 ;
        RECT 121.240 212.465 121.500 212.785 ;
        RECT 120.915 211.560 121.145 211.850 ;
        RECT 120.915 202.820 121.145 203.110 ;
        RECT 120.960 201.745 121.100 202.820 ;
        RECT 120.900 201.425 121.160 201.745 ;
        RECT 121.300 200.735 121.440 212.465 ;
        RECT 121.580 210.165 121.840 210.485 ;
        RECT 121.980 210.025 122.120 216.160 ;
        RECT 121.920 209.705 122.180 210.025 ;
        RECT 121.935 206.960 122.165 207.250 ;
        RECT 121.580 206.025 121.840 206.345 ;
        RECT 121.595 205.120 121.825 205.410 ;
        RECT 121.640 201.195 121.780 205.120 ;
        RECT 121.980 204.950 122.120 206.960 ;
        RECT 121.935 204.660 122.165 204.950 ;
        RECT 121.640 201.055 122.460 201.195 ;
        RECT 120.960 200.595 121.440 200.735 ;
        RECT 120.960 194.385 121.100 200.595 ;
        RECT 121.920 200.505 122.180 200.825 ;
        RECT 121.255 200.035 121.485 200.325 ;
        RECT 121.300 198.225 121.440 200.035 ;
        RECT 121.595 199.640 121.825 199.930 ;
        RECT 121.640 198.740 121.780 199.640 ;
        RECT 121.935 199.185 122.165 199.475 ;
        RECT 121.595 198.450 121.825 198.740 ;
        RECT 121.255 197.935 121.485 198.225 ;
        RECT 121.300 196.655 121.440 197.935 ;
        RECT 121.255 196.365 121.485 196.655 ;
        RECT 121.640 196.220 121.780 198.450 ;
        RECT 121.595 195.930 121.825 196.220 ;
        RECT 121.980 195.675 122.120 199.185 ;
        RECT 122.320 196.225 122.460 201.055 ;
        RECT 122.260 195.905 122.520 196.225 ;
        RECT 121.300 195.535 122.120 195.675 ;
        RECT 120.900 194.065 121.160 194.385 ;
        RECT 120.915 193.620 121.145 193.910 ;
        RECT 120.960 192.085 121.100 193.620 ;
        RECT 121.300 192.990 121.440 195.535 ;
        RECT 121.920 194.985 122.180 195.305 ;
        RECT 121.580 194.065 121.840 194.385 ;
        RECT 121.255 192.700 121.485 192.990 ;
        RECT 120.900 191.765 121.160 192.085 ;
        RECT 121.640 190.690 121.780 194.065 ;
        RECT 121.595 190.400 121.825 190.690 ;
        RECT 121.595 190.155 121.825 190.230 ;
        RECT 121.980 190.155 122.120 194.985 ;
        RECT 122.600 190.845 122.860 191.165 ;
        RECT 121.595 190.015 122.120 190.155 ;
        RECT 121.595 189.940 121.825 190.015 ;
        RECT 121.580 189.005 121.840 189.325 ;
        RECT 120.900 188.085 121.160 188.405 ;
        RECT 120.960 186.550 121.100 188.085 ;
        RECT 121.255 187.640 121.485 187.930 ;
        RECT 120.915 186.260 121.145 186.550 ;
        RECT 121.300 185.185 121.440 187.640 ;
        RECT 121.640 186.105 121.780 189.005 ;
        RECT 121.920 188.545 122.180 188.865 ;
        RECT 121.920 187.165 122.180 187.485 ;
        RECT 122.600 187.165 122.860 187.485 ;
        RECT 121.980 186.550 122.120 187.165 ;
        RECT 122.260 186.705 122.520 187.025 ;
        RECT 121.935 186.260 122.165 186.550 ;
        RECT 121.580 185.785 121.840 186.105 ;
        RECT 121.240 184.865 121.500 185.185 ;
        RECT 122.320 185.170 122.460 186.705 ;
        RECT 122.275 184.880 122.505 185.170 ;
        RECT 123.000 183.415 123.480 219.295 ;
        RECT 124.640 217.755 124.900 217.845 ;
        RECT 124.360 217.615 124.900 217.755 ;
        RECT 123.975 216.205 124.205 216.495 ;
        RECT 124.020 215.545 124.160 216.205 ;
        RECT 123.960 215.225 124.220 215.545 ;
        RECT 124.360 210.945 124.500 217.615 ;
        RECT 124.640 217.525 124.900 217.615 ;
        RECT 124.995 217.055 125.225 217.345 ;
        RECT 124.655 216.660 124.885 216.950 ;
        RECT 124.700 215.760 124.840 216.660 ;
        RECT 124.655 215.470 124.885 215.760 ;
        RECT 124.700 213.240 124.840 215.470 ;
        RECT 125.040 215.245 125.180 217.055 ;
        RECT 124.995 214.955 125.225 215.245 ;
        RECT 125.040 213.675 125.180 214.955 ;
        RECT 124.995 213.385 125.225 213.675 ;
        RECT 124.655 212.950 124.885 213.240 ;
        RECT 124.300 210.625 124.560 210.945 ;
        RECT 125.335 210.640 125.565 210.930 ;
        RECT 124.360 205.870 124.500 210.625 ;
        RECT 125.380 210.025 125.520 210.640 ;
        RECT 125.320 209.705 125.580 210.025 ;
        RECT 124.315 205.795 124.545 205.870 ;
        RECT 123.680 205.655 124.545 205.795 ;
        RECT 123.680 200.825 123.820 205.655 ;
        RECT 124.315 205.580 124.545 205.655 ;
        RECT 124.995 205.095 125.225 205.385 ;
        RECT 123.960 204.645 124.220 204.965 ;
        RECT 124.655 204.700 124.885 204.990 ;
        RECT 124.020 204.415 124.160 204.645 ;
        RECT 124.315 204.415 124.545 204.535 ;
        RECT 124.020 204.275 124.545 204.415 ;
        RECT 124.315 204.245 124.545 204.275 ;
        RECT 124.700 203.800 124.840 204.700 ;
        RECT 124.655 203.510 124.885 203.800 ;
        RECT 124.700 201.280 124.840 203.510 ;
        RECT 125.040 203.285 125.180 205.095 ;
        RECT 124.995 202.995 125.225 203.285 ;
        RECT 125.040 201.715 125.180 202.995 ;
        RECT 124.995 201.425 125.225 201.715 ;
        RECT 124.655 200.990 124.885 201.280 ;
        RECT 123.620 200.505 123.880 200.825 ;
        RECT 123.635 198.680 123.865 198.970 ;
        RECT 123.680 198.065 123.820 198.680 ;
        RECT 124.655 198.220 124.885 198.510 ;
        RECT 123.620 197.745 123.880 198.065 ;
        RECT 124.700 197.605 124.840 198.220 ;
        RECT 124.640 197.285 124.900 197.605 ;
        RECT 124.980 196.365 125.240 196.685 ;
        RECT 125.335 195.920 125.565 196.210 ;
        RECT 125.380 195.305 125.520 195.920 ;
        RECT 125.320 194.985 125.580 195.305 ;
        RECT 124.300 191.765 124.560 192.085 ;
        RECT 123.620 190.845 123.880 191.165 ;
        RECT 123.680 188.850 123.820 190.845 ;
        RECT 124.640 189.465 124.900 189.785 ;
        RECT 124.300 189.005 124.560 189.325 ;
        RECT 123.635 188.560 123.865 188.850 ;
        RECT 124.360 187.470 124.500 189.005 ;
        RECT 124.315 187.180 124.545 187.470 ;
        RECT 124.300 186.705 124.560 187.025 ;
        RECT 124.300 186.245 124.560 186.565 ;
        RECT 124.315 186.015 124.545 186.090 ;
        RECT 124.700 186.015 124.840 189.465 ;
        RECT 125.320 189.005 125.580 189.325 ;
        RECT 125.380 188.390 125.520 189.005 ;
        RECT 125.335 188.100 125.565 188.390 ;
        RECT 124.315 185.875 124.840 186.015 ;
        RECT 124.315 185.800 124.545 185.875 ;
        RECT 125.720 183.415 126.200 219.295 ;
        RECT 128.040 217.985 128.300 218.305 ;
        RECT 126.680 217.525 126.940 217.845 ;
        RECT 127.360 217.525 127.620 217.845 ;
        RECT 126.340 215.225 126.600 215.545 ;
        RECT 126.740 211.315 126.880 217.525 ;
        RECT 127.420 216.450 127.560 217.525 ;
        RECT 128.100 217.370 128.240 217.985 ;
        RECT 128.055 217.080 128.285 217.370 ;
        RECT 127.375 216.160 127.605 216.450 ;
        RECT 128.055 213.400 128.285 213.690 ;
        RECT 127.035 212.940 127.265 213.230 ;
        RECT 127.080 212.785 127.220 212.940 ;
        RECT 128.100 212.785 128.240 213.400 ;
        RECT 127.020 212.465 127.280 212.785 ;
        RECT 128.040 212.465 128.300 212.785 ;
        RECT 127.020 212.005 127.280 212.325 ;
        RECT 127.035 211.315 127.265 211.390 ;
        RECT 126.740 211.175 127.265 211.315 ;
        RECT 127.035 211.100 127.265 211.175 ;
        RECT 126.695 210.615 126.925 210.905 ;
        RECT 126.740 208.805 126.880 210.615 ;
        RECT 127.035 210.220 127.265 210.510 ;
        RECT 127.080 209.320 127.220 210.220 ;
        RECT 127.715 209.765 127.945 210.055 ;
        RECT 127.035 209.030 127.265 209.320 ;
        RECT 126.695 208.515 126.925 208.805 ;
        RECT 126.740 207.235 126.880 208.515 ;
        RECT 126.695 206.945 126.925 207.235 ;
        RECT 127.080 206.800 127.220 209.030 ;
        RECT 127.035 206.510 127.265 206.800 ;
        RECT 127.760 206.345 127.900 209.765 ;
        RECT 127.700 206.025 127.960 206.345 ;
        RECT 127.760 204.965 127.900 206.025 ;
        RECT 126.680 204.645 126.940 204.965 ;
        RECT 127.700 204.645 127.960 204.965 ;
        RECT 126.740 204.030 126.880 204.645 ;
        RECT 128.040 204.185 128.300 204.505 ;
        RECT 126.695 203.740 126.925 204.030 ;
        RECT 127.375 201.900 127.605 202.190 ;
        RECT 127.035 201.655 127.265 201.730 ;
        RECT 126.740 201.515 127.265 201.655 ;
        RECT 126.740 196.225 126.880 201.515 ;
        RECT 127.035 201.440 127.265 201.515 ;
        RECT 127.035 200.520 127.265 200.810 ;
        RECT 127.080 198.525 127.220 200.520 ;
        RECT 127.420 199.890 127.560 201.900 ;
        RECT 127.375 199.600 127.605 199.890 ;
        RECT 127.020 198.205 127.280 198.525 ;
        RECT 127.020 197.745 127.280 198.065 ;
        RECT 127.080 197.130 127.220 197.745 ;
        RECT 128.100 197.605 128.240 204.185 ;
        RECT 128.040 197.285 128.300 197.605 ;
        RECT 127.035 196.840 127.265 197.130 ;
        RECT 126.680 195.905 126.940 196.225 ;
        RECT 126.740 190.230 126.880 195.905 ;
        RECT 127.360 193.605 127.620 193.925 ;
        RECT 127.420 192.530 127.560 193.605 ;
        RECT 127.375 192.240 127.605 192.530 ;
        RECT 127.375 191.995 127.605 192.070 ;
        RECT 127.375 191.855 127.900 191.995 ;
        RECT 127.375 191.780 127.605 191.855 ;
        RECT 127.360 191.305 127.620 191.625 ;
        RECT 127.035 190.860 127.265 191.150 ;
        RECT 126.695 189.940 126.925 190.230 ;
        RECT 127.080 187.485 127.220 190.860 ;
        RECT 127.760 189.785 127.900 191.855 ;
        RECT 127.700 189.465 127.960 189.785 ;
        RECT 127.375 188.560 127.605 188.850 ;
        RECT 127.420 188.405 127.560 188.560 ;
        RECT 127.360 188.085 127.620 188.405 ;
        RECT 127.360 187.625 127.620 187.945 ;
        RECT 128.040 187.625 128.300 187.945 ;
        RECT 127.020 187.165 127.280 187.485 ;
        RECT 127.375 186.260 127.605 186.550 ;
        RECT 127.420 186.105 127.560 186.260 ;
        RECT 127.360 185.785 127.620 186.105 ;
        RECT 128.100 185.630 128.240 187.625 ;
        RECT 128.055 185.340 128.285 185.630 ;
        RECT 128.440 183.415 128.920 219.295 ;
        RECT 130.080 217.525 130.340 217.845 ;
        RECT 130.140 216.450 130.280 217.525 ;
        RECT 130.095 216.160 130.325 216.450 ;
        RECT 130.760 212.925 131.020 213.245 ;
        RECT 129.060 212.465 129.320 212.785 ;
        RECT 129.740 209.705 130.000 210.025 ;
        RECT 129.755 205.795 129.985 205.870 ;
        RECT 129.460 205.655 129.985 205.795 ;
        RECT 129.460 200.350 129.600 205.655 ;
        RECT 129.755 205.580 129.985 205.655 ;
        RECT 129.755 204.875 129.985 204.950 ;
        RECT 129.755 204.735 130.280 204.875 ;
        RECT 129.755 204.660 129.985 204.735 ;
        RECT 129.740 204.185 130.000 204.505 ;
        RECT 130.140 203.495 130.280 204.735 ;
        RECT 130.760 204.645 131.020 204.965 ;
        RECT 130.760 204.185 131.020 204.505 ;
        RECT 130.435 203.495 130.665 203.570 ;
        RECT 130.140 203.355 130.665 203.495 ;
        RECT 130.435 203.280 130.665 203.355 ;
        RECT 130.095 202.820 130.325 203.110 ;
        RECT 129.755 201.900 129.985 202.190 ;
        RECT 129.800 201.745 129.940 201.900 ;
        RECT 129.740 201.425 130.000 201.745 ;
        RECT 129.740 200.505 130.000 200.825 ;
        RECT 129.415 200.060 129.645 200.350 ;
        RECT 130.140 197.515 130.280 202.820 ;
        RECT 130.480 200.365 130.620 203.280 ;
        RECT 130.820 202.650 130.960 204.185 ;
        RECT 130.775 202.360 131.005 202.650 ;
        RECT 130.420 200.045 130.680 200.365 ;
        RECT 130.140 197.375 130.620 197.515 ;
        RECT 130.080 196.825 130.340 197.145 ;
        RECT 130.480 196.225 130.620 197.375 ;
        RECT 130.420 195.905 130.680 196.225 ;
        RECT 129.075 195.000 129.305 195.290 ;
        RECT 129.120 194.385 129.260 195.000 ;
        RECT 129.060 194.065 129.320 194.385 ;
        RECT 129.755 194.295 129.985 194.370 ;
        RECT 129.755 194.155 130.280 194.295 ;
        RECT 129.755 194.080 129.985 194.155 ;
        RECT 129.755 193.160 129.985 193.450 ;
        RECT 129.415 191.780 129.645 192.070 ;
        RECT 129.060 191.305 129.320 191.625 ;
        RECT 129.120 191.150 129.260 191.305 ;
        RECT 129.075 190.860 129.305 191.150 ;
        RECT 129.460 189.785 129.600 191.780 ;
        RECT 129.800 191.610 129.940 193.160 ;
        RECT 129.755 191.320 129.985 191.610 ;
        RECT 129.800 191.165 129.940 191.320 ;
        RECT 129.740 190.845 130.000 191.165 ;
        RECT 129.755 190.615 129.985 190.690 ;
        RECT 130.140 190.615 130.280 194.155 ;
        RECT 130.760 193.605 131.020 193.925 ;
        RECT 129.755 190.475 130.280 190.615 ;
        RECT 129.755 190.400 129.985 190.475 ;
        RECT 129.740 189.925 130.000 190.245 ;
        RECT 129.400 189.465 129.660 189.785 ;
        RECT 129.075 189.235 129.305 189.310 ;
        RECT 129.075 189.095 129.600 189.235 ;
        RECT 129.075 189.020 129.305 189.095 ;
        RECT 129.460 188.775 129.600 189.095 ;
        RECT 129.755 188.775 129.985 188.850 ;
        RECT 129.460 188.635 129.985 188.775 ;
        RECT 129.460 187.025 129.600 188.635 ;
        RECT 129.755 188.560 129.985 188.635 ;
        RECT 129.740 187.625 130.000 187.945 ;
        RECT 130.140 187.855 130.280 190.475 ;
        RECT 130.420 187.855 130.680 187.945 ;
        RECT 130.140 187.715 130.680 187.855 ;
        RECT 130.420 187.625 130.680 187.715 ;
        RECT 129.740 187.165 130.000 187.485 ;
        RECT 129.400 186.705 129.660 187.025 ;
        RECT 129.800 186.550 129.940 187.165 ;
        RECT 129.755 186.260 129.985 186.550 ;
        RECT 130.760 186.245 131.020 186.565 ;
        RECT 130.820 185.630 130.960 186.245 ;
        RECT 130.775 185.340 131.005 185.630 ;
        RECT 131.160 183.415 131.640 219.295 ;
        RECT 131.780 217.525 132.040 217.845 ;
        RECT 133.140 217.525 133.400 217.845 ;
        RECT 132.475 215.230 132.705 215.520 ;
        RECT 132.135 214.795 132.365 215.085 ;
        RECT 132.180 213.515 132.320 214.795 ;
        RECT 132.135 213.225 132.365 213.515 ;
        RECT 132.180 211.415 132.320 213.225 ;
        RECT 132.520 213.000 132.660 215.230 ;
        RECT 132.475 212.710 132.705 213.000 ;
        RECT 132.520 211.810 132.660 212.710 ;
        RECT 133.200 212.265 133.340 217.525 ;
        RECT 133.155 211.975 133.385 212.265 ;
        RECT 132.475 211.520 132.705 211.810 ;
        RECT 132.135 211.125 132.365 211.415 ;
        RECT 132.800 210.625 133.060 210.945 ;
        RECT 133.140 206.945 133.400 207.265 ;
        RECT 131.780 200.965 132.040 201.285 ;
        RECT 131.840 200.810 131.980 200.965 ;
        RECT 131.795 200.520 132.025 200.810 ;
        RECT 132.460 200.505 132.720 200.825 ;
        RECT 131.780 195.905 132.040 196.225 ;
        RECT 131.840 192.990 131.980 195.905 ;
        RECT 132.520 195.290 132.660 200.505 ;
        RECT 133.480 197.745 133.740 198.065 ;
        RECT 133.480 195.445 133.740 195.765 ;
        RECT 132.475 195.000 132.705 195.290 ;
        RECT 131.795 192.700 132.025 192.990 ;
        RECT 132.800 192.685 133.060 193.005 ;
        RECT 132.800 191.765 133.060 192.085 ;
        RECT 133.540 191.150 133.680 195.445 ;
        RECT 133.495 190.860 133.725 191.150 ;
        RECT 131.780 189.465 132.040 189.785 ;
        RECT 131.840 186.550 131.980 189.465 ;
        RECT 132.800 187.395 133.060 187.485 ;
        RECT 132.800 187.255 133.340 187.395 ;
        RECT 132.800 187.165 133.060 187.255 ;
        RECT 131.795 186.260 132.025 186.550 ;
        RECT 132.815 186.260 133.045 186.550 ;
        RECT 132.860 186.105 133.000 186.260 ;
        RECT 132.800 185.785 133.060 186.105 ;
        RECT 133.200 186.015 133.340 187.255 ;
        RECT 133.495 186.015 133.725 186.090 ;
        RECT 133.200 185.875 133.725 186.015 ;
        RECT 133.495 185.800 133.725 185.875 ;
        RECT 132.800 184.865 133.060 185.185 ;
        RECT 133.880 183.415 134.360 219.295 ;
        RECT 134.500 217.525 134.760 217.845 ;
        RECT 134.515 215.700 134.745 215.990 ;
        RECT 134.560 213.245 134.700 215.700 ;
        RECT 135.520 215.225 135.780 215.545 ;
        RECT 135.535 214.320 135.765 214.610 ;
        RECT 135.195 213.400 135.425 213.690 ;
        RECT 135.580 213.615 135.720 214.320 ;
        RECT 135.580 213.475 136.400 213.615 ;
        RECT 134.500 212.925 134.760 213.245 ;
        RECT 134.900 212.355 135.040 212.760 ;
        RECT 134.855 212.325 135.085 212.355 ;
        RECT 134.840 212.005 135.100 212.325 ;
        RECT 134.900 204.875 135.040 212.005 ;
        RECT 135.240 210.945 135.380 213.400 ;
        RECT 135.875 212.915 136.105 213.205 ;
        RECT 135.535 212.520 135.765 212.810 ;
        RECT 135.580 211.620 135.720 212.520 ;
        RECT 135.535 211.330 135.765 211.620 ;
        RECT 135.180 210.625 135.440 210.945 ;
        RECT 135.240 208.185 135.380 210.625 ;
        RECT 135.580 209.100 135.720 211.330 ;
        RECT 135.920 211.105 136.060 212.915 ;
        RECT 135.875 210.815 136.105 211.105 ;
        RECT 135.920 209.535 136.060 210.815 ;
        RECT 135.875 209.245 136.105 209.535 ;
        RECT 135.535 208.810 135.765 209.100 ;
        RECT 135.180 207.865 135.440 208.185 ;
        RECT 135.875 206.715 136.105 206.790 ;
        RECT 134.560 204.735 135.040 204.875 ;
        RECT 135.240 206.575 136.105 206.715 ;
        RECT 134.560 198.525 134.700 204.735 ;
        RECT 134.855 204.245 135.085 204.535 ;
        RECT 134.500 198.205 134.760 198.525 ;
        RECT 134.560 197.590 134.700 198.205 ;
        RECT 134.900 198.065 135.040 204.245 ;
        RECT 134.840 197.745 135.100 198.065 ;
        RECT 135.240 197.605 135.380 206.575 ;
        RECT 135.875 206.500 136.105 206.575 ;
        RECT 135.520 205.565 135.780 205.885 ;
        RECT 135.875 205.095 136.105 205.385 ;
        RECT 135.535 204.700 135.765 204.990 ;
        RECT 135.580 203.800 135.720 204.700 ;
        RECT 135.535 203.510 135.765 203.800 ;
        RECT 135.580 201.280 135.720 203.510 ;
        RECT 135.920 203.285 136.060 205.095 ;
        RECT 136.260 204.965 136.400 213.475 ;
        RECT 136.200 204.645 136.460 204.965 ;
        RECT 135.875 202.995 136.105 203.285 ;
        RECT 135.920 201.715 136.060 202.995 ;
        RECT 135.875 201.425 136.105 201.715 ;
        RECT 135.535 200.990 135.765 201.280 ;
        RECT 136.215 198.680 136.445 198.970 ;
        RECT 136.260 198.525 136.400 198.680 ;
        RECT 136.200 198.205 136.460 198.525 ;
        RECT 134.515 197.300 134.745 197.590 ;
        RECT 135.180 197.285 135.440 197.605 ;
        RECT 134.840 196.595 135.100 196.685 ;
        RECT 135.240 196.595 135.380 197.285 ;
        RECT 135.860 196.825 136.120 197.145 ;
        RECT 134.840 196.455 135.380 196.595 ;
        RECT 134.840 196.365 135.100 196.455 ;
        RECT 134.900 195.290 135.040 196.365 ;
        RECT 134.855 195.000 135.085 195.290 ;
        RECT 134.515 193.620 134.745 193.910 ;
        RECT 134.560 193.005 134.700 193.620 ;
        RECT 134.500 192.685 134.760 193.005 ;
        RECT 135.195 192.915 135.425 192.990 ;
        RECT 134.900 192.775 135.425 192.915 ;
        RECT 134.900 192.455 135.040 192.775 ;
        RECT 135.195 192.700 135.425 192.775 ;
        RECT 134.560 192.315 135.040 192.455 ;
        RECT 135.535 192.455 135.765 192.530 ;
        RECT 135.535 192.315 136.060 192.455 ;
        RECT 134.560 187.855 134.700 192.315 ;
        RECT 135.535 192.240 135.765 192.315 ;
        RECT 135.535 191.780 135.765 192.070 ;
        RECT 135.195 191.535 135.425 191.610 ;
        RECT 134.900 191.395 135.425 191.535 ;
        RECT 134.900 190.230 135.040 191.395 ;
        RECT 135.195 191.320 135.425 191.395 ;
        RECT 135.180 190.845 135.440 191.165 ;
        RECT 135.240 190.690 135.380 190.845 ;
        RECT 135.195 190.400 135.425 190.690 ;
        RECT 134.855 189.940 135.085 190.230 ;
        RECT 135.195 189.480 135.425 189.770 ;
        RECT 135.240 188.405 135.380 189.480 ;
        RECT 135.580 189.325 135.720 191.780 ;
        RECT 135.920 190.245 136.060 192.315 ;
        RECT 135.860 189.925 136.120 190.245 ;
        RECT 135.520 189.005 135.780 189.325 ;
        RECT 135.180 188.085 135.440 188.405 ;
        RECT 135.180 187.855 135.440 187.945 ;
        RECT 134.560 187.715 135.440 187.855 ;
        RECT 135.180 187.625 135.440 187.715 ;
        RECT 135.180 186.245 135.440 186.565 ;
        RECT 135.180 185.785 135.440 186.105 ;
        RECT 135.240 185.630 135.380 185.785 ;
        RECT 135.920 185.645 136.060 189.925 ;
        RECT 136.215 188.560 136.445 188.850 ;
        RECT 136.260 187.025 136.400 188.560 ;
        RECT 136.200 186.705 136.460 187.025 ;
        RECT 135.195 185.340 135.425 185.630 ;
        RECT 135.860 185.325 136.120 185.645 ;
        RECT 136.600 183.415 137.080 219.295 ;
        RECT 138.920 217.985 139.180 218.305 ;
        RECT 138.980 217.370 139.120 217.985 ;
        RECT 138.935 217.080 139.165 217.370 ;
        RECT 138.255 216.160 138.485 216.450 ;
        RECT 137.560 215.225 137.820 215.545 ;
        RECT 137.620 213.615 137.760 215.225 ;
        RECT 137.915 213.615 138.145 213.690 ;
        RECT 137.620 213.475 138.145 213.615 ;
        RECT 137.235 200.980 137.465 201.270 ;
        RECT 137.280 200.825 137.420 200.980 ;
        RECT 137.220 200.505 137.480 200.825 ;
        RECT 137.620 195.765 137.760 213.475 ;
        RECT 137.915 213.400 138.145 213.475 ;
        RECT 137.915 212.480 138.145 212.770 ;
        RECT 137.960 212.325 138.100 212.480 ;
        RECT 137.900 212.005 138.160 212.325 ;
        RECT 138.300 210.945 138.440 216.160 ;
        RECT 138.920 215.685 139.180 216.005 ;
        RECT 138.935 213.860 139.165 214.150 ;
        RECT 138.240 210.625 138.500 210.945 ;
        RECT 138.980 210.485 139.120 213.860 ;
        RECT 138.920 210.165 139.180 210.485 ;
        RECT 138.920 207.865 139.180 208.185 ;
        RECT 138.980 205.885 139.120 207.865 ;
        RECT 138.920 205.565 139.180 205.885 ;
        RECT 138.920 204.645 139.180 204.965 ;
        RECT 138.255 201.440 138.485 201.730 ;
        RECT 138.300 201.285 138.440 201.440 ;
        RECT 138.980 201.285 139.120 204.645 ;
        RECT 138.240 200.965 138.500 201.285 ;
        RECT 138.920 200.965 139.180 201.285 ;
        RECT 137.915 197.760 138.145 198.050 ;
        RECT 137.960 197.605 138.100 197.760 ;
        RECT 137.900 197.285 138.160 197.605 ;
        RECT 138.580 195.905 138.840 196.225 ;
        RECT 137.560 195.445 137.820 195.765 ;
        RECT 137.915 195.000 138.145 195.290 ;
        RECT 137.235 194.755 137.465 194.830 ;
        RECT 137.235 194.615 137.760 194.755 ;
        RECT 137.235 194.540 137.465 194.615 ;
        RECT 137.220 193.605 137.480 193.925 ;
        RECT 137.620 191.165 137.760 194.615 ;
        RECT 137.960 191.995 138.100 195.000 ;
        RECT 138.255 194.755 138.485 194.830 ;
        RECT 138.255 194.615 139.120 194.755 ;
        RECT 138.255 194.540 138.485 194.615 ;
        RECT 138.595 192.700 138.825 192.990 ;
        RECT 138.240 191.995 138.500 192.085 ;
        RECT 137.960 191.855 138.500 191.995 ;
        RECT 138.240 191.765 138.500 191.855 ;
        RECT 138.640 191.625 138.780 192.700 ;
        RECT 138.580 191.305 138.840 191.625 ;
        RECT 137.560 190.845 137.820 191.165 ;
        RECT 138.580 190.845 138.840 191.165 ;
        RECT 138.255 190.615 138.485 190.690 ;
        RECT 137.960 190.475 138.485 190.615 ;
        RECT 137.960 189.310 138.100 190.475 ;
        RECT 138.255 190.400 138.485 190.475 ;
        RECT 138.255 189.695 138.485 189.770 ;
        RECT 138.640 189.695 138.780 190.845 ;
        RECT 138.255 189.555 138.780 189.695 ;
        RECT 138.255 189.480 138.485 189.555 ;
        RECT 137.915 189.020 138.145 189.310 ;
        RECT 138.240 188.085 138.500 188.405 ;
        RECT 138.240 186.705 138.500 187.025 ;
        RECT 138.255 185.800 138.485 186.090 ;
        RECT 138.640 186.015 138.780 189.555 ;
        RECT 138.980 188.405 139.120 194.615 ;
        RECT 138.920 188.085 139.180 188.405 ;
        RECT 138.920 186.015 139.180 186.105 ;
        RECT 138.640 185.875 139.180 186.015 ;
        RECT 138.300 185.645 138.440 185.800 ;
        RECT 138.920 185.785 139.180 185.875 ;
        RECT 138.240 185.325 138.500 185.645 ;
        RECT 139.320 183.415 139.800 219.295 ;
        RECT 140.635 217.540 140.865 217.830 ;
        RECT 140.295 216.205 140.525 216.495 ;
        RECT 140.340 216.005 140.480 216.205 ;
        RECT 140.280 215.685 140.540 216.005 ;
        RECT 139.940 210.855 140.200 210.945 ;
        RECT 139.940 210.715 140.480 210.855 ;
        RECT 139.940 210.625 140.200 210.715 ;
        RECT 139.940 210.165 140.200 210.485 ;
        RECT 140.340 207.635 140.480 210.715 ;
        RECT 140.680 208.185 140.820 217.540 ;
        RECT 141.315 217.055 141.545 217.345 ;
        RECT 140.975 216.660 141.205 216.950 ;
        RECT 141.020 215.760 141.160 216.660 ;
        RECT 140.975 215.470 141.205 215.760 ;
        RECT 141.020 213.240 141.160 215.470 ;
        RECT 141.360 215.245 141.500 217.055 ;
        RECT 141.315 214.955 141.545 215.245 ;
        RECT 141.360 213.675 141.500 214.955 ;
        RECT 141.315 213.385 141.545 213.675 ;
        RECT 140.975 212.950 141.205 213.240 ;
        RECT 140.620 207.865 140.880 208.185 ;
        RECT 140.635 207.635 140.865 207.710 ;
        RECT 140.340 207.495 140.865 207.635 ;
        RECT 140.635 207.420 140.865 207.495 ;
        RECT 141.640 205.565 141.900 205.885 ;
        RECT 140.635 203.740 140.865 204.030 ;
        RECT 140.295 203.280 140.525 203.570 ;
        RECT 139.940 201.425 140.200 201.745 ;
        RECT 140.000 199.430 140.140 201.425 ;
        RECT 139.955 199.140 140.185 199.430 ;
        RECT 140.340 195.765 140.480 203.280 ;
        RECT 140.680 201.745 140.820 203.740 ;
        RECT 140.975 202.575 141.205 202.650 ;
        RECT 140.975 202.435 141.500 202.575 ;
        RECT 140.975 202.360 141.205 202.435 ;
        RECT 140.620 201.425 140.880 201.745 ;
        RECT 140.620 200.965 140.880 201.285 ;
        RECT 140.620 200.045 140.880 200.365 ;
        RECT 140.680 198.525 140.820 200.045 ;
        RECT 140.620 198.205 140.880 198.525 ;
        RECT 140.620 197.745 140.880 198.065 ;
        RECT 140.680 197.145 140.820 197.745 ;
        RECT 140.960 197.285 141.220 197.605 ;
        RECT 141.360 197.515 141.500 202.435 ;
        RECT 141.640 200.505 141.900 200.825 ;
        RECT 141.700 198.510 141.840 200.505 ;
        RECT 141.655 198.220 141.885 198.510 ;
        RECT 141.360 197.375 141.840 197.515 ;
        RECT 140.620 196.825 140.880 197.145 ;
        RECT 141.315 196.815 141.545 197.105 ;
        RECT 140.975 196.420 141.205 196.710 ;
        RECT 140.635 195.965 140.865 196.255 ;
        RECT 140.280 195.445 140.540 195.765 ;
        RECT 140.680 194.845 140.820 195.965 ;
        RECT 141.020 195.520 141.160 196.420 ;
        RECT 140.975 195.230 141.205 195.520 ;
        RECT 140.620 194.525 140.880 194.845 ;
        RECT 141.020 193.000 141.160 195.230 ;
        RECT 141.360 195.005 141.500 196.815 ;
        RECT 141.700 195.765 141.840 197.375 ;
        RECT 141.640 195.445 141.900 195.765 ;
        RECT 141.315 194.715 141.545 195.005 ;
        RECT 141.360 193.435 141.500 194.715 ;
        RECT 141.315 193.145 141.545 193.435 ;
        RECT 140.975 192.710 141.205 193.000 ;
        RECT 141.700 192.455 141.840 195.445 ;
        RECT 140.680 192.315 141.840 192.455 ;
        RECT 140.680 189.770 140.820 192.315 ;
        RECT 141.640 190.385 141.900 190.705 ;
        RECT 140.635 189.480 140.865 189.770 ;
        RECT 140.620 188.545 140.880 188.865 ;
        RECT 141.640 187.625 141.900 187.945 ;
        RECT 140.620 187.165 140.880 187.485 ;
        RECT 139.940 186.245 140.200 186.565 ;
        RECT 139.940 185.785 140.200 186.105 ;
        RECT 140.620 184.865 140.880 185.185 ;
        RECT 142.040 183.415 142.520 219.295 ;
        RECT 144.360 213.385 144.620 213.705 ;
        RECT 143.355 211.090 143.585 211.380 ;
        RECT 143.015 210.655 143.245 210.945 ;
        RECT 143.060 209.375 143.200 210.655 ;
        RECT 143.015 209.085 143.245 209.375 ;
        RECT 142.660 207.865 142.920 208.185 ;
        RECT 142.720 206.255 142.860 207.865 ;
        RECT 143.060 207.275 143.200 209.085 ;
        RECT 143.400 208.860 143.540 211.090 ;
        RECT 143.355 208.570 143.585 208.860 ;
        RECT 144.360 208.785 144.620 209.105 ;
        RECT 143.400 207.670 143.540 208.570 ;
        RECT 143.695 207.780 143.925 208.070 ;
        RECT 143.355 207.380 143.585 207.670 ;
        RECT 143.015 206.985 143.245 207.275 ;
        RECT 143.355 206.500 143.585 206.790 ;
        RECT 143.400 206.330 143.540 206.500 ;
        RECT 143.355 206.255 143.585 206.330 ;
        RECT 142.720 206.115 143.585 206.255 ;
        RECT 142.720 197.605 142.860 206.115 ;
        RECT 143.355 206.040 143.585 206.115 ;
        RECT 143.740 205.885 143.880 207.780 ;
        RECT 144.020 206.485 144.280 206.805 ;
        RECT 143.015 205.555 143.245 205.845 ;
        RECT 143.680 205.565 143.940 205.885 ;
        RECT 143.060 203.745 143.200 205.555 ;
        RECT 143.355 205.160 143.585 205.450 ;
        RECT 143.400 204.260 143.540 205.160 ;
        RECT 144.080 205.105 144.220 206.485 ;
        RECT 144.035 204.815 144.265 205.105 ;
        RECT 143.355 203.970 143.585 204.260 ;
        RECT 143.015 203.455 143.245 203.745 ;
        RECT 143.060 202.175 143.200 203.455 ;
        RECT 143.015 201.885 143.245 202.175 ;
        RECT 143.400 201.740 143.540 203.970 ;
        RECT 144.420 203.955 144.560 208.785 ;
        RECT 144.080 203.815 144.560 203.955 ;
        RECT 143.355 201.450 143.585 201.740 ;
        RECT 143.000 200.965 143.260 201.285 ;
        RECT 142.660 197.285 142.920 197.605 ;
        RECT 143.060 195.750 143.200 200.965 ;
        RECT 143.340 200.045 143.600 200.365 ;
        RECT 143.400 196.595 143.540 200.045 ;
        RECT 144.080 198.970 144.220 203.815 ;
        RECT 144.375 199.140 144.605 199.430 ;
        RECT 144.035 198.680 144.265 198.970 ;
        RECT 144.420 198.525 144.560 199.140 ;
        RECT 144.360 198.205 144.620 198.525 ;
        RECT 144.020 197.745 144.280 198.065 ;
        RECT 143.680 196.825 143.940 197.145 ;
        RECT 143.695 196.595 143.925 196.670 ;
        RECT 143.400 196.455 143.925 196.595 ;
        RECT 143.695 196.380 143.925 196.455 ;
        RECT 143.340 195.905 143.600 196.225 ;
        RECT 143.015 195.460 143.245 195.750 ;
        RECT 142.660 194.525 142.920 194.845 ;
        RECT 142.720 192.990 142.860 194.525 ;
        RECT 143.015 194.080 143.245 194.370 ;
        RECT 142.675 192.700 142.905 192.990 ;
        RECT 143.060 191.610 143.200 194.080 ;
        RECT 143.400 193.835 143.540 195.905 ;
        RECT 143.680 195.445 143.940 195.765 ;
        RECT 143.740 194.830 143.880 195.445 ;
        RECT 143.695 194.540 143.925 194.830 ;
        RECT 143.680 193.835 143.940 193.925 ;
        RECT 143.400 193.695 143.940 193.835 ;
        RECT 143.680 193.605 143.940 193.695 ;
        RECT 143.740 192.070 143.880 193.605 ;
        RECT 143.695 191.780 143.925 192.070 ;
        RECT 143.015 191.320 143.245 191.610 ;
        RECT 143.680 190.845 143.940 191.165 ;
        RECT 143.000 190.385 143.260 190.705 ;
        RECT 143.695 190.400 143.925 190.690 ;
        RECT 143.060 189.695 143.200 190.385 ;
        RECT 143.355 189.695 143.585 189.770 ;
        RECT 143.060 189.555 143.585 189.695 ;
        RECT 143.355 189.480 143.585 189.555 ;
        RECT 142.660 188.545 142.920 188.865 ;
        RECT 142.720 186.550 142.860 188.545 ;
        RECT 143.740 187.945 143.880 190.400 ;
        RECT 143.680 187.625 143.940 187.945 ;
        RECT 143.000 187.165 143.260 187.485 ;
        RECT 142.675 186.260 142.905 186.550 ;
        RECT 143.060 186.090 143.200 187.165 ;
        RECT 143.015 185.800 143.245 186.090 ;
        RECT 143.680 184.865 143.940 185.185 ;
        RECT 144.760 183.415 145.240 219.295 ;
        RECT 146.060 213.385 146.320 213.705 ;
        RECT 146.120 211.390 146.260 213.385 ;
        RECT 146.075 211.315 146.305 211.390 ;
        RECT 146.075 211.175 146.600 211.315 ;
        RECT 146.075 211.100 146.305 211.175 ;
        RECT 146.060 208.785 146.320 209.105 ;
        RECT 146.060 208.325 146.320 208.645 ;
        RECT 146.075 207.420 146.305 207.710 ;
        RECT 145.380 206.485 145.640 206.805 ;
        RECT 145.380 201.425 145.640 201.745 ;
        RECT 146.120 199.355 146.260 207.420 ;
        RECT 146.460 204.950 146.600 211.175 ;
        RECT 147.095 210.180 147.325 210.470 ;
        RECT 146.755 207.880 146.985 208.170 ;
        RECT 146.415 204.660 146.645 204.950 ;
        RECT 146.800 200.825 146.940 207.880 ;
        RECT 147.140 205.425 147.280 210.180 ;
        RECT 147.080 205.105 147.340 205.425 ;
        RECT 146.740 200.505 147.000 200.825 ;
        RECT 147.095 199.600 147.325 199.890 ;
        RECT 146.120 199.215 146.940 199.355 ;
        RECT 146.075 198.680 146.305 198.970 ;
        RECT 146.120 198.525 146.260 198.680 ;
        RECT 146.060 198.205 146.320 198.525 ;
        RECT 145.380 197.745 145.640 198.065 ;
        RECT 145.440 195.290 145.580 197.745 ;
        RECT 146.060 195.445 146.320 195.765 ;
        RECT 145.395 195.000 145.625 195.290 ;
        RECT 146.120 194.830 146.260 195.445 ;
        RECT 146.075 194.540 146.305 194.830 ;
        RECT 146.800 193.925 146.940 199.215 ;
        RECT 147.140 198.985 147.280 199.600 ;
        RECT 147.080 198.665 147.340 198.985 ;
        RECT 146.740 193.605 147.000 193.925 ;
        RECT 147.080 192.225 147.340 192.545 ;
        RECT 145.380 191.765 145.640 192.085 ;
        RECT 145.440 188.850 145.580 191.765 ;
        RECT 147.140 191.610 147.280 192.225 ;
        RECT 147.095 191.320 147.325 191.610 ;
        RECT 146.060 190.385 146.320 190.705 ;
        RECT 145.395 188.560 145.625 188.850 ;
        RECT 145.380 188.085 145.640 188.405 ;
        RECT 145.440 187.470 145.580 188.085 ;
        RECT 146.060 187.625 146.320 187.945 ;
        RECT 145.395 187.180 145.625 187.470 ;
        RECT 146.060 186.245 146.320 186.565 ;
        RECT 145.395 185.800 145.625 186.090 ;
        RECT 145.440 185.645 145.580 185.800 ;
        RECT 145.380 185.325 145.640 185.645 ;
        RECT 146.060 184.865 146.320 185.185 ;
        RECT 147.480 183.415 147.960 219.295 ;
        RECT 148.200 201.290 148.340 219.570 ;
        RECT 148.110 200.960 148.440 201.290 ;
        RECT 148.720 198.955 148.860 220.050 ;
        RECT 148.630 198.695 148.950 198.955 ;
        RECT 149.210 198.060 149.350 220.770 ;
        RECT 149.770 205.430 149.910 221.830 ;
        RECT 149.680 205.100 150.000 205.430 ;
        RECT 148.670 197.920 149.350 198.060 ;
        RECT 148.670 192.550 148.810 197.920 ;
        RECT 148.570 192.220 148.900 192.550 ;
        RECT 71.820 182.250 76.725 182.390 ;
        RECT 71.820 182.190 72.140 182.250 ;
        RECT 76.435 182.205 76.725 182.250 ;
        RECT 63.540 182.050 63.860 182.110 ;
        RECT 64.935 182.050 65.225 182.095 ;
        RECT 62.250 181.910 65.225 182.050 ;
        RECT 58.020 181.850 58.340 181.910 ;
        RECT 61.700 181.850 62.020 181.910 ;
        RECT 63.540 181.850 63.860 181.910 ;
        RECT 64.935 181.865 65.225 181.910 ;
        RECT 67.220 181.850 67.540 182.110 ;
        RECT 68.140 182.095 68.460 182.110 ;
        RECT 68.140 181.865 68.525 182.095 ;
        RECT 69.060 182.050 69.380 182.110 ;
        RECT 70.760 182.050 71.050 182.095 ;
        RECT 69.060 181.910 71.050 182.050 ;
        RECT 68.140 181.850 68.460 181.865 ;
        RECT 69.060 181.850 69.380 181.910 ;
        RECT 70.760 181.865 71.050 181.910 ;
        RECT 53.435 181.570 54.200 181.710 ;
        RECT 53.435 181.525 53.725 181.570 ;
        RECT 51.120 181.170 51.440 181.430 ;
        RECT 52.590 181.370 52.730 181.525 ;
        RECT 53.880 181.510 54.200 181.570 ;
        RECT 54.355 181.525 54.645 181.755 ;
        RECT 55.735 181.710 56.025 181.755 ;
        RECT 56.180 181.710 56.500 181.770 ;
        RECT 55.735 181.570 56.500 181.710 ;
        RECT 55.735 181.525 56.025 181.570 ;
        RECT 56.180 181.510 56.500 181.570 ;
        RECT 57.115 181.525 57.405 181.755 ;
        RECT 54.800 181.370 55.120 181.430 ;
        RECT 52.590 181.230 55.120 181.370 ;
        RECT 45.600 180.890 50.890 181.030 ;
        RECT 45.600 180.830 45.920 180.890 ;
        RECT 46.980 180.690 47.300 180.750 ;
        RECT 44.770 180.550 47.300 180.690 ;
        RECT 32.735 180.505 33.025 180.550 ;
        RECT 33.180 180.490 33.500 180.550 ;
        RECT 46.980 180.490 47.300 180.550 ;
        RECT 47.440 180.690 47.760 180.750 ;
        RECT 52.590 180.690 52.730 181.230 ;
        RECT 54.800 181.170 55.120 181.230 ;
        RECT 55.260 181.370 55.580 181.430 ;
        RECT 57.190 181.370 57.330 181.525 ;
        RECT 57.560 181.510 57.880 181.770 ;
        RECT 58.940 181.510 59.260 181.770 ;
        RECT 59.400 181.510 59.720 181.770 ;
        RECT 60.335 181.710 60.625 181.755 ;
        RECT 66.760 181.710 67.080 181.770 ;
        RECT 60.335 181.570 61.470 181.710 ;
        RECT 60.335 181.525 60.625 181.570 ;
        RECT 61.330 181.430 61.470 181.570 ;
        RECT 62.250 181.570 67.080 181.710 ;
        RECT 55.260 181.230 57.330 181.370 ;
        RECT 55.260 181.170 55.580 181.230 ;
        RECT 61.240 181.170 61.560 181.430 ;
        RECT 61.715 181.185 62.005 181.415 ;
        RECT 60.780 181.030 61.100 181.090 ;
        RECT 61.790 181.030 61.930 181.185 ;
        RECT 60.780 180.890 61.930 181.030 ;
        RECT 60.780 180.830 61.100 180.890 ;
        RECT 47.440 180.550 52.730 180.690 ;
        RECT 47.440 180.490 47.760 180.550 ;
        RECT 55.720 180.490 56.040 180.750 ;
        RECT 62.250 180.735 62.390 181.570 ;
        RECT 66.760 181.510 67.080 181.570 ;
        RECT 68.600 181.370 68.920 181.430 ;
        RECT 65.010 181.230 68.920 181.370 ;
        RECT 63.080 181.030 63.400 181.090 ;
        RECT 64.015 181.030 64.305 181.075 ;
        RECT 63.080 180.890 64.305 181.030 ;
        RECT 63.080 180.830 63.400 180.890 ;
        RECT 64.015 180.845 64.305 180.890 ;
        RECT 65.010 180.735 65.150 181.230 ;
        RECT 68.600 181.170 68.920 181.230 ;
        RECT 69.520 181.170 69.840 181.430 ;
        RECT 70.415 181.370 70.705 181.415 ;
        RECT 71.605 181.370 71.895 181.415 ;
        RECT 74.125 181.370 74.415 181.415 ;
        RECT 70.415 181.230 74.415 181.370 ;
        RECT 70.415 181.185 70.705 181.230 ;
        RECT 71.605 181.185 71.895 181.230 ;
        RECT 74.125 181.185 74.415 181.230 ;
        RECT 70.020 181.030 70.310 181.075 ;
        RECT 72.120 181.030 72.410 181.075 ;
        RECT 73.690 181.030 73.980 181.075 ;
        RECT 70.020 180.890 73.980 181.030 ;
        RECT 70.020 180.845 70.310 180.890 ;
        RECT 72.120 180.845 72.410 180.890 ;
        RECT 73.690 180.845 73.980 180.890 ;
        RECT 62.175 180.505 62.465 180.735 ;
        RECT 64.935 180.505 65.225 180.735 ;
        RECT 67.680 180.690 68.000 180.750 ;
        RECT 68.155 180.690 68.445 180.735 ;
        RECT 67.680 180.550 68.445 180.690 ;
        RECT 67.680 180.490 68.000 180.550 ;
        RECT 68.155 180.505 68.445 180.550 ;
        RECT 69.075 180.690 69.365 180.735 ;
        RECT 70.440 180.690 70.760 180.750 ;
        RECT 69.075 180.550 70.760 180.690 ;
        RECT 69.075 180.505 69.365 180.550 ;
        RECT 70.440 180.490 70.760 180.550 ;
        RECT 11.950 179.870 90.610 180.350 ;
        RECT 17.080 179.670 17.400 179.730 ;
        RECT 17.555 179.670 17.845 179.715 ;
        RECT 17.080 179.530 17.845 179.670 ;
        RECT 17.080 179.470 17.400 179.530 ;
        RECT 17.555 179.485 17.845 179.530 ;
        RECT 27.215 179.670 27.505 179.715 ;
        RECT 29.500 179.670 29.820 179.730 ;
        RECT 27.215 179.530 29.820 179.670 ;
        RECT 27.215 179.485 27.505 179.530 ;
        RECT 29.500 179.470 29.820 179.530 ;
        RECT 35.020 179.670 35.340 179.730 ;
        RECT 35.495 179.670 35.785 179.715 ;
        RECT 35.020 179.530 35.785 179.670 ;
        RECT 35.020 179.470 35.340 179.530 ;
        RECT 35.495 179.485 35.785 179.530 ;
        RECT 36.400 179.470 36.720 179.730 ;
        RECT 46.520 179.470 46.840 179.730 ;
        RECT 48.360 179.470 48.680 179.730 ;
        RECT 49.370 179.530 50.430 179.670 ;
        RECT 20.300 179.330 20.590 179.375 ;
        RECT 21.870 179.330 22.160 179.375 ;
        RECT 23.970 179.330 24.260 179.375 ;
        RECT 20.300 179.190 24.260 179.330 ;
        RECT 20.300 179.145 20.590 179.190 ;
        RECT 21.870 179.145 22.160 179.190 ;
        RECT 23.970 179.145 24.260 179.190 ;
        RECT 25.375 179.330 25.665 179.375 ;
        RECT 26.740 179.330 27.060 179.390 ;
        RECT 25.375 179.190 27.060 179.330 ;
        RECT 25.375 179.145 25.665 179.190 ;
        RECT 26.740 179.130 27.060 179.190 ;
        RECT 29.080 179.330 29.370 179.375 ;
        RECT 31.180 179.330 31.470 179.375 ;
        RECT 32.750 179.330 33.040 179.375 ;
        RECT 29.080 179.190 33.040 179.330 ;
        RECT 29.080 179.145 29.370 179.190 ;
        RECT 31.180 179.145 31.470 179.190 ;
        RECT 32.750 179.145 33.040 179.190 ;
        RECT 35.940 179.330 36.260 179.390 ;
        RECT 37.335 179.330 37.625 179.375 ;
        RECT 40.540 179.330 40.860 179.390 ;
        RECT 35.940 179.190 40.860 179.330 ;
        RECT 35.940 179.130 36.260 179.190 ;
        RECT 37.335 179.145 37.625 179.190 ;
        RECT 40.540 179.130 40.860 179.190 ;
        RECT 19.865 178.990 20.155 179.035 ;
        RECT 22.385 178.990 22.675 179.035 ;
        RECT 23.575 178.990 23.865 179.035 ;
        RECT 19.865 178.850 23.865 178.990 ;
        RECT 19.865 178.805 20.155 178.850 ;
        RECT 22.385 178.805 22.675 178.850 ;
        RECT 23.575 178.805 23.865 178.850 ;
        RECT 29.475 178.990 29.765 179.035 ;
        RECT 30.665 178.990 30.955 179.035 ;
        RECT 33.185 178.990 33.475 179.035 ;
        RECT 29.475 178.850 33.475 178.990 ;
        RECT 29.475 178.805 29.765 178.850 ;
        RECT 30.665 178.805 30.955 178.850 ;
        RECT 33.185 178.805 33.475 178.850 ;
        RECT 24.440 178.450 24.760 178.710 ;
        RECT 28.595 178.650 28.885 178.695 ;
        RECT 36.860 178.650 37.180 178.710 ;
        RECT 28.595 178.510 37.180 178.650 ;
        RECT 28.595 178.465 28.885 178.510 ;
        RECT 36.860 178.450 37.180 178.510 ;
        RECT 44.220 178.650 44.540 178.710 ;
        RECT 44.695 178.650 44.985 178.695 ;
        RECT 44.220 178.510 44.985 178.650 ;
        RECT 44.220 178.450 44.540 178.510 ;
        RECT 44.695 178.465 44.985 178.510 ;
        RECT 45.600 178.450 45.920 178.710 ;
        RECT 46.610 178.650 46.750 179.470 ;
        RECT 46.980 178.990 47.300 179.050 ;
        RECT 47.915 178.990 48.205 179.035 ;
        RECT 46.980 178.850 48.205 178.990 ;
        RECT 46.980 178.790 47.300 178.850 ;
        RECT 47.915 178.805 48.205 178.850 ;
        RECT 47.455 178.650 47.745 178.695 ;
        RECT 46.610 178.510 47.745 178.650 ;
        RECT 47.455 178.465 47.745 178.510 ;
        RECT 48.835 178.650 49.125 178.695 ;
        RECT 49.370 178.650 49.510 179.530 ;
        RECT 49.755 179.145 50.045 179.375 ;
        RECT 50.290 179.330 50.430 179.530 ;
        RECT 51.120 179.470 51.440 179.730 ;
        RECT 55.260 179.470 55.580 179.730 ;
        RECT 56.180 179.470 56.500 179.730 ;
        RECT 57.115 179.670 57.405 179.715 ;
        RECT 57.560 179.670 57.880 179.730 ;
        RECT 61.255 179.670 61.545 179.715 ;
        RECT 57.115 179.530 61.545 179.670 ;
        RECT 57.115 179.485 57.405 179.530 ;
        RECT 57.560 179.470 57.880 179.530 ;
        RECT 61.255 179.485 61.545 179.530 ;
        RECT 68.140 179.670 68.460 179.730 ;
        RECT 68.140 179.530 70.670 179.670 ;
        RECT 68.140 179.470 68.460 179.530 ;
        RECT 52.960 179.330 53.280 179.390 ;
        RECT 58.480 179.330 58.800 179.390 ;
        RECT 50.290 179.190 58.800 179.330 ;
        RECT 48.835 178.510 49.510 178.650 ;
        RECT 49.830 178.650 49.970 179.145 ;
        RECT 52.960 179.130 53.280 179.190 ;
        RECT 58.480 179.130 58.800 179.190 ;
        RECT 59.415 179.330 59.705 179.375 ;
        RECT 60.320 179.330 60.640 179.390 ;
        RECT 59.415 179.190 60.640 179.330 ;
        RECT 59.415 179.145 59.705 179.190 ;
        RECT 60.320 179.130 60.640 179.190 ;
        RECT 53.435 178.990 53.725 179.035 ;
        RECT 56.180 178.990 56.500 179.050 ;
        RECT 67.680 178.990 68.000 179.050 ;
        RECT 70.530 179.035 70.670 179.530 ;
        RECT 53.435 178.850 54.800 178.990 ;
        RECT 53.435 178.805 53.725 178.850 ;
        RECT 54.660 178.710 54.800 178.850 ;
        RECT 56.180 178.850 68.000 178.990 ;
        RECT 56.180 178.790 56.500 178.850 ;
        RECT 67.680 178.790 68.000 178.850 ;
        RECT 69.075 178.990 69.365 179.035 ;
        RECT 69.075 178.850 70.210 178.990 ;
        RECT 69.075 178.805 69.365 178.850 ;
        RECT 52.055 178.650 52.345 178.695 ;
        RECT 49.830 178.510 52.345 178.650 ;
        RECT 48.835 178.465 49.125 178.510 ;
        RECT 52.055 178.465 52.345 178.510 ;
        RECT 52.515 178.465 52.805 178.695 ;
        RECT 21.680 178.310 22.000 178.370 ;
        RECT 23.120 178.310 23.410 178.355 ;
        RECT 29.820 178.310 30.110 178.355 ;
        RECT 21.680 178.170 23.410 178.310 ;
        RECT 21.680 178.110 22.000 178.170 ;
        RECT 23.120 178.125 23.410 178.170 ;
        RECT 28.210 178.170 30.110 178.310 ;
        RECT 27.200 177.770 27.520 178.030 ;
        RECT 28.210 178.015 28.350 178.170 ;
        RECT 29.820 178.125 30.110 178.170 ;
        RECT 34.100 178.310 34.420 178.370 ;
        RECT 38.715 178.310 39.005 178.355 ;
        RECT 34.100 178.170 39.005 178.310 ;
        RECT 34.100 178.110 34.420 178.170 ;
        RECT 38.715 178.125 39.005 178.170 ;
        RECT 40.080 178.310 40.400 178.370 ;
        RECT 47.900 178.310 48.220 178.370 ;
        RECT 52.590 178.310 52.730 178.465 ;
        RECT 53.880 178.450 54.200 178.710 ;
        RECT 54.660 178.510 55.120 178.710 ;
        RECT 54.800 178.450 55.120 178.510 ;
        RECT 55.735 178.650 56.025 178.695 ;
        RECT 58.940 178.650 59.260 178.710 ;
        RECT 59.875 178.650 60.165 178.695 ;
        RECT 55.735 178.510 58.710 178.650 ;
        RECT 55.735 178.465 56.025 178.510 ;
        RECT 40.080 178.170 52.730 178.310 ;
        RECT 54.890 178.310 55.030 178.450 ;
        RECT 58.570 178.370 58.710 178.510 ;
        RECT 58.940 178.510 60.165 178.650 ;
        RECT 58.940 178.450 59.260 178.510 ;
        RECT 59.875 178.465 60.165 178.510 ;
        RECT 62.635 178.465 62.925 178.695 ;
        RECT 57.560 178.310 57.880 178.370 ;
        RECT 54.890 178.170 57.880 178.310 ;
        RECT 40.080 178.110 40.400 178.170 ;
        RECT 47.900 178.110 48.220 178.170 ;
        RECT 57.560 178.110 57.880 178.170 ;
        RECT 58.020 178.110 58.340 178.370 ;
        RECT 58.480 178.110 58.800 178.370 ;
        RECT 28.135 177.785 28.425 178.015 ;
        RECT 57.035 177.970 57.325 178.015 ;
        RECT 59.875 177.970 60.165 178.015 ;
        RECT 57.035 177.830 60.165 177.970 ;
        RECT 62.710 177.970 62.850 178.465 ;
        RECT 63.080 178.450 63.400 178.710 ;
        RECT 63.555 178.650 63.845 178.695 ;
        RECT 64.000 178.650 64.320 178.710 ;
        RECT 63.555 178.510 64.320 178.650 ;
        RECT 63.555 178.465 63.845 178.510 ;
        RECT 64.000 178.450 64.320 178.510 ;
        RECT 64.460 178.450 64.780 178.710 ;
        RECT 70.070 178.695 70.210 178.850 ;
        RECT 70.455 178.805 70.745 179.035 ;
        RECT 68.645 178.465 68.935 178.695 ;
        RECT 69.535 178.465 69.825 178.695 ;
        RECT 69.995 178.465 70.285 178.695 ;
        RECT 70.915 178.650 71.205 178.695 ;
        RECT 71.360 178.650 71.680 178.710 ;
        RECT 70.915 178.510 71.680 178.650 ;
        RECT 70.915 178.465 71.205 178.510 ;
        RECT 66.760 178.310 67.080 178.370 ;
        RECT 68.690 178.310 68.830 178.465 ;
        RECT 66.760 178.170 68.830 178.310 ;
        RECT 66.760 178.110 67.080 178.170 ;
        RECT 68.600 177.970 68.920 178.030 ;
        RECT 62.710 177.830 68.920 177.970 ;
        RECT 69.610 177.970 69.750 178.465 ;
        RECT 71.360 178.450 71.680 178.510 ;
        RECT 101.005 178.120 102.595 182.410 ;
        RECT 100.100 178.100 140.370 178.120 ;
        RECT 100.100 178.080 140.860 178.100 ;
        RECT 69.980 177.970 70.300 178.030 ;
        RECT 69.610 177.830 70.300 177.970 ;
        RECT 57.035 177.785 57.325 177.830 ;
        RECT 59.875 177.785 60.165 177.830 ;
        RECT 68.600 177.770 68.920 177.830 ;
        RECT 69.980 177.770 70.300 177.830 ;
        RECT 11.950 177.150 90.610 177.630 ;
        RECT 99.990 177.050 140.860 178.080 ;
        RECT 21.680 176.750 22.000 177.010 ;
        RECT 48.360 176.950 48.680 177.010 ;
        RECT 62.160 176.950 62.480 177.010 ;
        RECT 48.360 176.810 62.480 176.950 ;
        RECT 48.360 176.750 48.680 176.810 ;
        RECT 62.160 176.750 62.480 176.810 ;
        RECT 99.990 176.770 100.770 177.050 ;
        RECT 17.080 176.610 17.400 176.670 ;
        RECT 19.395 176.610 19.685 176.655 ;
        RECT 17.080 176.470 19.685 176.610 ;
        RECT 17.080 176.410 17.400 176.470 ;
        RECT 19.395 176.425 19.685 176.470 ;
        RECT 59.860 176.610 60.180 176.670 ;
        RECT 63.080 176.610 63.400 176.670 ;
        RECT 70.915 176.610 71.205 176.655 ;
        RECT 72.280 176.610 72.600 176.670 ;
        RECT 59.860 176.470 63.400 176.610 ;
        RECT 59.860 176.410 60.180 176.470 ;
        RECT 63.080 176.410 63.400 176.470 ;
        RECT 70.070 176.470 71.205 176.610 ;
        RECT 70.070 176.330 70.210 176.470 ;
        RECT 70.915 176.425 71.205 176.470 ;
        RECT 71.450 176.470 72.600 176.610 ;
        RECT 43.315 176.270 43.605 176.315 ;
        RECT 43.760 176.270 44.080 176.330 ;
        RECT 43.315 176.130 44.080 176.270 ;
        RECT 43.315 176.085 43.605 176.130 ;
        RECT 43.760 176.070 44.080 176.130 ;
        RECT 44.235 176.270 44.525 176.315 ;
        RECT 47.440 176.270 47.760 176.330 ;
        RECT 44.235 176.130 47.760 176.270 ;
        RECT 44.235 176.085 44.525 176.130 ;
        RECT 47.440 176.070 47.760 176.130 ;
        RECT 67.680 176.070 68.000 176.330 ;
        RECT 69.060 176.070 69.380 176.330 ;
        RECT 69.980 176.070 70.300 176.330 ;
        RECT 70.440 176.070 70.760 176.330 ;
        RECT 71.450 176.315 71.590 176.470 ;
        RECT 72.280 176.410 72.600 176.470 ;
        RECT 71.375 176.085 71.665 176.315 ;
        RECT 71.820 176.070 72.140 176.330 ;
        RECT 72.755 176.270 73.045 176.315 ;
        RECT 73.200 176.270 73.520 176.330 ;
        RECT 72.755 176.130 73.520 176.270 ;
        RECT 72.755 176.085 73.045 176.130 ;
        RECT 73.200 176.070 73.520 176.130 ;
        RECT 67.235 175.930 67.525 175.975 ;
        RECT 68.600 175.930 68.920 175.990 ;
        RECT 67.235 175.790 68.920 175.930 ;
        RECT 67.235 175.745 67.525 175.790 ;
        RECT 20.760 175.590 21.080 175.650 ;
        RECT 27.200 175.590 27.520 175.650 ;
        RECT 20.760 175.450 27.520 175.590 ;
        RECT 20.760 175.390 21.080 175.450 ;
        RECT 27.200 175.390 27.520 175.450 ;
        RECT 42.840 175.590 43.160 175.650 ;
        RECT 49.740 175.590 50.060 175.650 ;
        RECT 52.500 175.590 52.820 175.650 ;
        RECT 42.840 175.450 52.820 175.590 ;
        RECT 68.230 175.590 68.370 175.790 ;
        RECT 68.600 175.730 68.920 175.790 ;
        RECT 69.535 175.930 69.825 175.975 ;
        RECT 70.900 175.930 71.220 175.990 ;
        RECT 69.535 175.790 71.220 175.930 ;
        RECT 69.535 175.745 69.825 175.790 ;
        RECT 70.900 175.730 71.220 175.790 ;
        RECT 70.440 175.590 70.760 175.650 ;
        RECT 68.230 175.450 70.760 175.590 ;
        RECT 42.840 175.390 43.160 175.450 ;
        RECT 49.740 175.390 50.060 175.450 ;
        RECT 52.500 175.390 52.820 175.450 ;
        RECT 70.440 175.390 70.760 175.450 ;
        RECT 42.380 175.250 42.700 175.310 ;
        RECT 43.315 175.250 43.605 175.295 ;
        RECT 42.380 175.110 43.605 175.250 ;
        RECT 42.380 175.050 42.700 175.110 ;
        RECT 43.315 175.065 43.605 175.110 ;
        RECT 51.580 175.250 51.900 175.310 ;
        RECT 68.140 175.250 68.460 175.310 ;
        RECT 51.580 175.110 68.460 175.250 ;
        RECT 51.580 175.050 51.900 175.110 ;
        RECT 68.140 175.050 68.460 175.110 ;
        RECT 69.980 175.250 70.300 175.310 ;
        RECT 71.360 175.250 71.680 175.310 ;
        RECT 99.990 175.260 100.880 176.770 ;
        RECT 106.550 176.380 107.800 176.820 ;
        RECT 117.640 176.640 118.600 176.800 ;
        RECT 120.030 176.750 120.810 177.050 ;
        RECT 140.080 176.800 140.860 177.050 ;
        RECT 104.490 176.370 109.730 176.380 ;
        RECT 101.540 176.270 116.840 176.370 ;
        RECT 101.540 176.260 116.875 176.270 ;
        RECT 101.500 176.140 116.875 176.260 ;
        RECT 101.500 176.030 105.500 176.140 ;
        RECT 106.550 176.060 108.290 176.140 ;
        RECT 108.870 176.060 116.875 176.140 ;
        RECT 106.550 175.980 107.800 176.060 ;
        RECT 108.875 176.040 116.875 176.060 ;
        RECT 69.980 175.110 71.680 175.250 ;
        RECT 69.980 175.050 70.300 175.110 ;
        RECT 71.360 175.050 71.680 175.110 ;
        RECT 11.950 174.430 90.610 174.910 ;
        RECT 100.050 174.670 100.880 175.260 ;
        RECT 101.110 175.730 101.340 175.980 ;
        RECT 105.660 175.840 105.890 175.980 ;
        RECT 108.440 175.840 108.670 175.990 ;
        RECT 105.660 175.730 108.670 175.840 ;
        RECT 117.080 175.730 117.310 175.990 ;
        RECT 101.110 175.290 117.310 175.730 ;
        RECT 101.110 175.020 101.340 175.290 ;
        RECT 105.660 175.260 117.310 175.290 ;
        RECT 105.660 175.170 108.670 175.260 ;
        RECT 105.660 175.020 105.890 175.170 ;
        RECT 108.440 175.030 108.670 175.170 ;
        RECT 117.080 175.030 117.310 175.260 ;
        RECT 101.500 174.740 105.500 174.970 ;
        RECT 108.875 174.760 116.875 174.980 ;
        RECT 117.640 174.760 118.880 176.640 ;
        RECT 108.875 174.750 118.880 174.760 ;
        RECT 101.500 174.670 105.490 174.740 ;
        RECT 100.050 174.560 105.490 174.670 ;
        RECT 108.930 174.620 118.880 174.750 ;
        RECT 119.930 175.260 120.810 176.750 ;
        RECT 126.430 176.330 127.680 176.770 ;
        RECT 137.520 176.620 138.480 176.750 ;
        RECT 124.370 176.320 129.610 176.330 ;
        RECT 121.420 176.220 136.720 176.320 ;
        RECT 121.420 176.210 136.755 176.220 ;
        RECT 121.380 176.090 136.755 176.210 ;
        RECT 121.380 175.980 125.380 176.090 ;
        RECT 126.430 176.010 128.170 176.090 ;
        RECT 128.750 176.010 136.755 176.090 ;
        RECT 126.430 175.930 127.680 176.010 ;
        RECT 128.755 175.990 136.755 176.010 ;
        RECT 120.990 175.680 121.220 175.930 ;
        RECT 125.540 175.790 125.770 175.930 ;
        RECT 128.320 175.790 128.550 175.940 ;
        RECT 125.540 175.680 128.550 175.790 ;
        RECT 136.960 175.680 137.190 175.940 ;
        RECT 119.930 174.620 120.760 175.260 ;
        RECT 120.990 175.240 137.190 175.680 ;
        RECT 120.990 174.970 121.220 175.240 ;
        RECT 125.540 175.210 137.190 175.240 ;
        RECT 125.540 175.120 128.550 175.210 ;
        RECT 125.540 174.970 125.770 175.120 ;
        RECT 128.320 174.980 128.550 175.120 ;
        RECT 136.960 174.980 137.190 175.210 ;
        RECT 121.380 174.690 125.380 174.920 ;
        RECT 128.755 174.710 136.755 174.930 ;
        RECT 137.520 174.710 138.700 176.620 ;
        RECT 128.755 174.700 138.700 174.710 ;
        RECT 121.380 174.620 125.370 174.690 ;
        RECT 108.930 174.590 118.600 174.620 ;
        RECT 100.050 174.470 103.180 174.560 ;
        RECT 116.670 174.540 118.600 174.590 ;
        RECT 29.040 174.230 29.360 174.290 ;
        RECT 29.515 174.230 29.805 174.275 ;
        RECT 29.040 174.090 29.805 174.230 ;
        RECT 29.040 174.030 29.360 174.090 ;
        RECT 29.515 174.045 29.805 174.090 ;
        RECT 31.815 174.230 32.105 174.275 ;
        RECT 35.940 174.230 36.260 174.290 ;
        RECT 31.815 174.090 36.260 174.230 ;
        RECT 31.815 174.045 32.105 174.090 ;
        RECT 27.200 173.890 27.520 173.950 ;
        RECT 30.895 173.890 31.185 173.935 ;
        RECT 27.200 173.750 31.185 173.890 ;
        RECT 27.200 173.690 27.520 173.750 ;
        RECT 30.895 173.705 31.185 173.750 ;
        RECT 28.580 173.550 28.900 173.610 ;
        RECT 31.890 173.550 32.030 174.045 ;
        RECT 35.940 174.030 36.260 174.090 ;
        RECT 42.395 174.230 42.685 174.275 ;
        RECT 42.840 174.230 43.160 174.290 ;
        RECT 42.395 174.090 43.160 174.230 ;
        RECT 42.395 174.045 42.685 174.090 ;
        RECT 42.840 174.030 43.160 174.090 ;
        RECT 44.695 174.230 44.985 174.275 ;
        RECT 45.600 174.230 45.920 174.290 ;
        RECT 44.695 174.090 45.920 174.230 ;
        RECT 44.695 174.045 44.985 174.090 ;
        RECT 45.600 174.030 45.920 174.090 ;
        RECT 47.440 174.030 47.760 174.290 ;
        RECT 57.575 174.230 57.865 174.275 ;
        RECT 58.480 174.230 58.800 174.290 ;
        RECT 57.575 174.090 58.800 174.230 ;
        RECT 57.575 174.045 57.865 174.090 ;
        RECT 58.480 174.030 58.800 174.090 ;
        RECT 68.615 174.230 68.905 174.275 ;
        RECT 69.060 174.230 69.380 174.290 ;
        RECT 68.615 174.090 69.380 174.230 ;
        RECT 68.615 174.045 68.905 174.090 ;
        RECT 69.060 174.030 69.380 174.090 ;
        RECT 71.820 174.230 72.140 174.290 ;
        RECT 75.040 174.230 75.360 174.290 ;
        RECT 71.820 174.090 75.360 174.230 ;
        RECT 71.820 174.030 72.140 174.090 ;
        RECT 75.040 174.030 75.360 174.090 ;
        RECT 43.300 173.890 43.620 173.950 ;
        RECT 46.060 173.890 46.380 173.950 ;
        RECT 52.515 173.890 52.805 173.935 ;
        RECT 43.300 173.750 52.805 173.890 ;
        RECT 43.300 173.690 43.620 173.750 ;
        RECT 46.060 173.690 46.380 173.750 ;
        RECT 52.515 173.705 52.805 173.750 ;
        RECT 57.115 173.705 57.405 173.935 ;
        RECT 65.395 173.890 65.685 173.935 ;
        RECT 69.980 173.890 70.300 173.950 ;
        RECT 65.395 173.750 70.300 173.890 ;
        RECT 65.395 173.705 65.685 173.750 ;
        RECT 28.580 173.410 32.030 173.550 ;
        RECT 28.580 173.350 28.900 173.410 ;
        RECT 36.860 173.350 37.180 173.610 ;
        RECT 56.640 173.550 56.960 173.610 ;
        RECT 41.090 173.410 56.960 173.550 ;
        RECT 57.190 173.550 57.330 173.705 ;
        RECT 69.980 173.690 70.300 173.750 ;
        RECT 71.360 173.890 71.680 173.950 ;
        RECT 73.200 173.890 73.520 173.950 ;
        RECT 71.360 173.750 73.520 173.890 ;
        RECT 71.360 173.690 71.680 173.750 ;
        RECT 73.200 173.690 73.520 173.750 ;
        RECT 77.380 173.890 77.670 173.935 ;
        RECT 79.480 173.890 79.770 173.935 ;
        RECT 81.050 173.890 81.340 173.935 ;
        RECT 77.380 173.750 81.340 173.890 ;
        RECT 77.380 173.705 77.670 173.750 ;
        RECT 79.480 173.705 79.770 173.750 ;
        RECT 81.050 173.705 81.340 173.750 ;
        RECT 68.155 173.550 68.445 173.595 ;
        RECT 68.600 173.550 68.920 173.610 ;
        RECT 75.960 173.550 76.280 173.610 ;
        RECT 76.895 173.550 77.185 173.595 ;
        RECT 57.190 173.410 60.550 173.550 ;
        RECT 28.120 173.210 28.440 173.270 ;
        RECT 29.960 173.210 30.280 173.270 ;
        RECT 41.090 173.255 41.230 173.410 ;
        RECT 56.640 173.350 56.960 173.410 ;
        RECT 28.120 173.070 30.280 173.210 ;
        RECT 28.120 173.010 28.440 173.070 ;
        RECT 29.960 173.010 30.280 173.070 ;
        RECT 41.015 173.025 41.305 173.255 ;
        RECT 41.460 173.210 41.780 173.270 ;
        RECT 46.075 173.210 46.365 173.255 ;
        RECT 41.460 173.070 46.365 173.210 ;
        RECT 41.460 173.010 41.780 173.070 ;
        RECT 26.280 172.870 26.600 172.930 ;
        RECT 28.595 172.870 28.885 172.915 ;
        RECT 26.280 172.730 28.885 172.870 ;
        RECT 30.050 172.870 30.190 173.010 ;
        RECT 31.655 172.870 31.945 172.915 ;
        RECT 30.050 172.730 31.945 172.870 ;
        RECT 26.280 172.670 26.600 172.730 ;
        RECT 28.595 172.685 28.885 172.730 ;
        RECT 31.655 172.685 31.945 172.730 ;
        RECT 32.735 172.870 33.025 172.915 ;
        RECT 33.640 172.870 33.960 172.930 ;
        RECT 42.380 172.915 42.700 172.930 ;
        RECT 32.735 172.730 33.960 172.870 ;
        RECT 32.735 172.685 33.025 172.730 ;
        RECT 33.640 172.670 33.960 172.730 ;
        RECT 42.315 172.685 42.700 172.915 ;
        RECT 42.380 172.670 42.700 172.685 ;
        RECT 43.300 172.670 43.620 172.930 ;
        RECT 44.770 172.915 44.910 173.070 ;
        RECT 46.075 173.025 46.365 173.070 ;
        RECT 46.520 173.210 46.840 173.270 ;
        RECT 47.455 173.210 47.745 173.255 ;
        RECT 46.520 173.070 47.745 173.210 ;
        RECT 46.520 173.010 46.840 173.070 ;
        RECT 47.455 173.025 47.745 173.070 ;
        RECT 51.580 173.010 51.900 173.270 ;
        RECT 53.895 173.210 54.185 173.255 ;
        RECT 55.720 173.210 56.040 173.270 ;
        RECT 53.895 173.070 56.040 173.210 ;
        RECT 53.895 173.025 54.185 173.070 ;
        RECT 55.720 173.010 56.040 173.070 ;
        RECT 56.180 173.010 56.500 173.270 ;
        RECT 57.115 173.025 57.405 173.255 ;
        RECT 44.615 172.730 44.910 172.915 ;
        RECT 44.615 172.685 44.905 172.730 ;
        RECT 45.615 172.685 45.905 172.915 ;
        RECT 52.500 172.870 52.820 172.930 ;
        RECT 52.975 172.870 53.265 172.915 ;
        RECT 52.500 172.730 53.265 172.870 ;
        RECT 57.190 172.870 57.330 173.025 ;
        RECT 58.480 173.010 58.800 173.270 ;
        RECT 60.410 173.255 60.550 173.410 ;
        RECT 62.710 173.410 68.920 173.550 ;
        RECT 62.710 173.270 62.850 173.410 ;
        RECT 68.155 173.365 68.445 173.410 ;
        RECT 68.600 173.350 68.920 173.410 ;
        RECT 69.610 173.410 72.510 173.550 ;
        RECT 60.335 173.025 60.625 173.255 ;
        RECT 62.160 173.210 62.480 173.270 ;
        RECT 61.965 173.070 62.480 173.210 ;
        RECT 62.160 173.010 62.480 173.070 ;
        RECT 62.620 173.010 62.940 173.270 ;
        RECT 66.775 173.210 67.065 173.255 ;
        RECT 67.680 173.210 68.000 173.270 ;
        RECT 69.610 173.255 69.750 173.410 ;
        RECT 72.370 173.270 72.510 173.410 ;
        RECT 75.960 173.410 77.185 173.550 ;
        RECT 75.960 173.350 76.280 173.410 ;
        RECT 76.895 173.365 77.185 173.410 ;
        RECT 77.775 173.550 78.065 173.595 ;
        RECT 78.965 173.550 79.255 173.595 ;
        RECT 81.485 173.550 81.775 173.595 ;
        RECT 77.775 173.410 81.775 173.550 ;
        RECT 77.775 173.365 78.065 173.410 ;
        RECT 78.965 173.365 79.255 173.410 ;
        RECT 81.485 173.365 81.775 173.410 ;
        RECT 66.775 173.070 68.000 173.210 ;
        RECT 66.775 173.025 67.065 173.070 ;
        RECT 67.680 173.010 68.000 173.070 ;
        RECT 69.535 173.025 69.825 173.255 ;
        RECT 70.440 173.010 70.760 173.270 ;
        RECT 72.280 173.010 72.600 173.270 ;
        RECT 73.675 173.210 73.965 173.255 ;
        RECT 78.175 173.210 78.465 173.255 ;
        RECT 73.675 173.070 78.465 173.210 ;
        RECT 73.675 173.025 73.965 173.070 ;
        RECT 78.175 173.025 78.465 173.070 ;
        RECT 58.955 172.870 59.245 172.915 ;
        RECT 57.190 172.730 59.245 172.870 ;
        RECT 29.500 172.575 29.820 172.590 ;
        RECT 29.500 172.345 29.885 172.575 ;
        RECT 29.500 172.330 29.820 172.345 ;
        RECT 30.420 172.330 30.740 172.590 ;
        RECT 41.000 172.530 41.320 172.590 ;
        RECT 41.475 172.530 41.765 172.575 ;
        RECT 41.000 172.390 41.765 172.530 ;
        RECT 41.000 172.330 41.320 172.390 ;
        RECT 41.475 172.345 41.765 172.390 ;
        RECT 43.760 172.330 44.080 172.590 ;
        RECT 45.690 172.530 45.830 172.685 ;
        RECT 52.500 172.670 52.820 172.730 ;
        RECT 52.975 172.685 53.265 172.730 ;
        RECT 58.955 172.685 59.245 172.730 ;
        RECT 59.415 172.870 59.705 172.915 ;
        RECT 60.795 172.870 61.085 172.915 ;
        RECT 59.415 172.730 61.085 172.870 ;
        RECT 59.415 172.685 59.705 172.730 ;
        RECT 60.795 172.685 61.085 172.730 ;
        RECT 66.315 172.870 66.605 172.915 ;
        RECT 68.140 172.870 68.460 172.930 ;
        RECT 70.915 172.870 71.205 172.915 ;
        RECT 72.755 172.870 73.045 172.915 ;
        RECT 74.135 172.870 74.425 172.915 ;
        RECT 66.315 172.730 67.910 172.870 ;
        RECT 66.315 172.685 66.605 172.730 ;
        RECT 46.535 172.530 46.825 172.575 ;
        RECT 46.980 172.530 47.300 172.590 ;
        RECT 45.690 172.390 47.300 172.530 ;
        RECT 59.030 172.530 59.170 172.685 ;
        RECT 66.390 172.530 66.530 172.685 ;
        RECT 59.030 172.390 66.530 172.530 ;
        RECT 66.760 172.530 67.080 172.590 ;
        RECT 67.235 172.530 67.525 172.575 ;
        RECT 66.760 172.390 67.525 172.530 ;
        RECT 67.770 172.530 67.910 172.730 ;
        RECT 68.140 172.730 72.510 172.870 ;
        RECT 68.140 172.670 68.460 172.730 ;
        RECT 70.915 172.685 71.205 172.730 ;
        RECT 72.370 172.590 72.510 172.730 ;
        RECT 72.755 172.730 74.425 172.870 ;
        RECT 72.755 172.685 73.045 172.730 ;
        RECT 74.135 172.685 74.425 172.730 ;
        RECT 75.040 172.670 75.360 172.930 ;
        RECT 75.975 172.685 76.265 172.915 ;
        RECT 71.360 172.530 71.680 172.590 ;
        RECT 67.770 172.390 71.680 172.530 ;
        RECT 46.535 172.345 46.825 172.390 ;
        RECT 46.980 172.330 47.300 172.390 ;
        RECT 66.760 172.330 67.080 172.390 ;
        RECT 67.235 172.345 67.525 172.390 ;
        RECT 71.360 172.330 71.680 172.390 ;
        RECT 71.820 172.330 72.140 172.590 ;
        RECT 72.280 172.330 72.600 172.590 ;
        RECT 73.200 172.530 73.520 172.590 ;
        RECT 76.050 172.530 76.190 172.685 ;
        RECT 83.795 172.530 84.085 172.575 ;
        RECT 73.200 172.390 84.085 172.530 ;
        RECT 73.200 172.330 73.520 172.390 ;
        RECT 83.795 172.345 84.085 172.390 ;
        RECT 11.950 171.710 90.610 172.190 ;
        RECT 29.040 171.310 29.360 171.570 ;
        RECT 56.180 171.510 56.500 171.570 ;
        RECT 60.320 171.510 60.640 171.570 ;
        RECT 41.090 171.370 60.640 171.510 ;
        RECT 24.440 171.170 24.760 171.230 ;
        RECT 29.500 171.170 29.820 171.230 ;
        RECT 36.860 171.170 37.180 171.230 ;
        RECT 20.850 171.030 29.820 171.170 ;
        RECT 20.850 170.875 20.990 171.030 ;
        RECT 24.440 170.970 24.760 171.030 ;
        RECT 29.500 170.970 29.820 171.030 ;
        RECT 30.510 171.030 37.180 171.170 ;
        RECT 20.775 170.645 21.065 170.875 ;
        RECT 21.220 170.830 21.540 170.890 ;
        RECT 22.055 170.830 22.345 170.875 ;
        RECT 21.220 170.690 22.345 170.830 ;
        RECT 21.220 170.630 21.540 170.690 ;
        RECT 22.055 170.645 22.345 170.690 ;
        RECT 28.120 170.630 28.440 170.890 ;
        RECT 28.580 170.830 28.900 170.890 ;
        RECT 29.055 170.830 29.345 170.875 ;
        RECT 30.510 170.830 30.650 171.030 ;
        RECT 36.860 170.970 37.180 171.030 ;
        RECT 30.880 170.875 31.200 170.890 ;
        RECT 28.580 170.690 29.345 170.830 ;
        RECT 28.580 170.630 28.900 170.690 ;
        RECT 29.055 170.645 29.345 170.690 ;
        RECT 29.590 170.690 30.650 170.830 ;
        RECT 30.850 170.830 31.200 170.875 ;
        RECT 40.540 170.830 40.860 170.890 ;
        RECT 41.090 170.875 41.230 171.370 ;
        RECT 56.180 171.310 56.500 171.370 ;
        RECT 60.320 171.310 60.640 171.370 ;
        RECT 64.015 171.510 64.305 171.555 ;
        RECT 64.460 171.510 64.780 171.570 ;
        RECT 64.015 171.370 64.780 171.510 ;
        RECT 64.015 171.325 64.305 171.370 ;
        RECT 64.460 171.310 64.780 171.370 ;
        RECT 64.920 171.310 65.240 171.570 ;
        RECT 57.100 171.170 57.420 171.230 ;
        RECT 69.520 171.170 69.840 171.230 ;
        RECT 48.910 171.030 69.840 171.170 ;
        RECT 48.910 170.890 49.050 171.030 ;
        RECT 57.100 170.970 57.420 171.030 ;
        RECT 69.520 170.970 69.840 171.030 ;
        RECT 100.050 171.200 100.880 174.470 ;
        RECT 104.530 174.010 109.780 174.020 ;
        RECT 104.530 173.900 116.840 174.010 ;
        RECT 101.560 173.840 116.840 173.900 ;
        RECT 101.560 173.830 116.875 173.840 ;
        RECT 101.500 173.700 116.875 173.830 ;
        RECT 101.500 173.690 106.660 173.700 ;
        RECT 101.500 173.600 105.500 173.690 ;
        RECT 108.875 173.610 116.875 173.700 ;
        RECT 108.960 173.600 116.850 173.610 ;
        RECT 101.110 173.240 101.340 173.550 ;
        RECT 101.560 173.240 105.460 173.600 ;
        RECT 105.660 173.240 105.890 173.550 ;
        RECT 101.110 171.900 105.890 173.240 ;
        RECT 101.110 171.590 101.340 171.900 ;
        RECT 105.660 171.590 105.890 171.900 ;
        RECT 108.440 173.020 108.670 173.560 ;
        RECT 109.480 173.020 110.490 173.050 ;
        RECT 117.080 173.020 117.310 173.560 ;
        RECT 108.440 172.120 117.310 173.020 ;
        RECT 108.440 171.600 108.670 172.120 ;
        RECT 109.480 172.050 110.490 172.120 ;
        RECT 117.080 171.600 117.310 172.120 ;
        RECT 101.500 171.310 105.500 171.540 ;
        RECT 108.875 171.320 116.875 171.550 ;
        RECT 100.050 171.160 101.180 171.200 ;
        RECT 100.050 171.080 101.420 171.160 ;
        RECT 101.790 171.090 105.450 171.310 ;
        RECT 101.790 171.080 103.230 171.090 ;
        RECT 100.050 171.040 103.230 171.080 ;
        RECT 100.050 170.950 102.740 171.040 ;
        RECT 108.940 171.030 116.830 171.320 ;
        RECT 100.050 170.890 102.070 170.950 ;
        RECT 41.015 170.830 41.305 170.875 ;
        RECT 30.850 170.690 31.350 170.830 ;
        RECT 40.540 170.690 41.305 170.830 ;
        RECT 29.590 170.535 29.730 170.690 ;
        RECT 30.850 170.645 31.200 170.690 ;
        RECT 30.880 170.630 31.200 170.645 ;
        RECT 40.540 170.630 40.860 170.690 ;
        RECT 41.015 170.645 41.305 170.690 ;
        RECT 45.155 170.830 45.445 170.875 ;
        RECT 47.900 170.830 48.220 170.890 ;
        RECT 45.155 170.690 48.220 170.830 ;
        RECT 45.155 170.645 45.445 170.690 ;
        RECT 47.900 170.630 48.220 170.690 ;
        RECT 48.375 170.830 48.665 170.875 ;
        RECT 48.820 170.830 49.140 170.890 ;
        RECT 49.740 170.875 50.060 170.890 ;
        RECT 48.375 170.690 49.140 170.830 ;
        RECT 48.375 170.645 48.665 170.690 ;
        RECT 48.820 170.630 49.140 170.690 ;
        RECT 49.710 170.645 50.060 170.875 ;
        RECT 55.735 170.830 56.025 170.875 ;
        RECT 49.740 170.630 50.060 170.645 ;
        RECT 55.350 170.690 56.025 170.830 ;
        RECT 21.655 170.490 21.945 170.535 ;
        RECT 22.845 170.490 23.135 170.535 ;
        RECT 25.365 170.490 25.655 170.535 ;
        RECT 21.655 170.350 25.655 170.490 ;
        RECT 21.655 170.305 21.945 170.350 ;
        RECT 22.845 170.305 23.135 170.350 ;
        RECT 25.365 170.305 25.655 170.350 ;
        RECT 29.515 170.305 29.805 170.535 ;
        RECT 30.395 170.490 30.685 170.535 ;
        RECT 31.585 170.490 31.875 170.535 ;
        RECT 34.105 170.490 34.395 170.535 ;
        RECT 30.395 170.350 34.395 170.490 ;
        RECT 30.395 170.305 30.685 170.350 ;
        RECT 31.585 170.305 31.875 170.350 ;
        RECT 34.105 170.305 34.395 170.350 ;
        RECT 39.175 170.490 39.465 170.535 ;
        RECT 44.235 170.490 44.525 170.535 ;
        RECT 39.175 170.350 44.525 170.490 ;
        RECT 39.175 170.305 39.465 170.350 ;
        RECT 44.235 170.305 44.525 170.350 ;
        RECT 49.255 170.490 49.545 170.535 ;
        RECT 50.445 170.490 50.735 170.535 ;
        RECT 52.965 170.490 53.255 170.535 ;
        RECT 49.255 170.350 53.255 170.490 ;
        RECT 49.255 170.305 49.545 170.350 ;
        RECT 50.445 170.305 50.735 170.350 ;
        RECT 52.965 170.305 53.255 170.350 ;
        RECT 21.260 170.150 21.550 170.195 ;
        RECT 23.360 170.150 23.650 170.195 ;
        RECT 24.930 170.150 25.220 170.195 ;
        RECT 21.260 170.010 25.220 170.150 ;
        RECT 21.260 169.965 21.550 170.010 ;
        RECT 23.360 169.965 23.650 170.010 ;
        RECT 24.930 169.965 25.220 170.010 ;
        RECT 30.000 170.150 30.290 170.195 ;
        RECT 32.100 170.150 32.390 170.195 ;
        RECT 33.670 170.150 33.960 170.195 ;
        RECT 30.000 170.010 33.960 170.150 ;
        RECT 30.000 169.965 30.290 170.010 ;
        RECT 32.100 169.965 32.390 170.010 ;
        RECT 33.670 169.965 33.960 170.010 ;
        RECT 44.680 169.950 45.000 170.210 ;
        RECT 48.860 170.150 49.150 170.195 ;
        RECT 50.960 170.150 51.250 170.195 ;
        RECT 52.530 170.150 52.820 170.195 ;
        RECT 48.860 170.010 52.820 170.150 ;
        RECT 48.860 169.965 49.150 170.010 ;
        RECT 50.960 169.965 51.250 170.010 ;
        RECT 52.530 169.965 52.820 170.010 ;
        RECT 25.820 169.810 26.140 169.870 ;
        RECT 27.675 169.810 27.965 169.855 ;
        RECT 25.820 169.670 27.965 169.810 ;
        RECT 25.820 169.610 26.140 169.670 ;
        RECT 27.675 169.625 27.965 169.670 ;
        RECT 28.120 169.810 28.440 169.870 ;
        RECT 30.420 169.810 30.740 169.870 ;
        RECT 28.120 169.670 30.740 169.810 ;
        RECT 28.120 169.610 28.440 169.670 ;
        RECT 30.420 169.610 30.740 169.670 ;
        RECT 35.940 169.810 36.260 169.870 ;
        RECT 36.415 169.810 36.705 169.855 ;
        RECT 35.940 169.670 36.705 169.810 ;
        RECT 35.940 169.610 36.260 169.670 ;
        RECT 36.415 169.625 36.705 169.670 ;
        RECT 50.200 169.810 50.520 169.870 ;
        RECT 53.880 169.810 54.200 169.870 ;
        RECT 55.350 169.855 55.490 170.690 ;
        RECT 55.735 170.645 56.025 170.690 ;
        RECT 56.180 170.830 56.500 170.890 ;
        RECT 57.575 170.830 57.865 170.875 ;
        RECT 56.180 170.690 57.865 170.830 ;
        RECT 56.180 170.630 56.500 170.690 ;
        RECT 57.575 170.645 57.865 170.690 ;
        RECT 60.320 170.630 60.640 170.890 ;
        RECT 64.920 170.830 65.210 170.875 ;
        RECT 66.300 170.830 66.620 170.890 ;
        RECT 64.920 170.690 66.620 170.830 ;
        RECT 64.920 170.645 65.210 170.690 ;
        RECT 66.300 170.630 66.620 170.690 ;
        RECT 66.775 170.830 67.065 170.875 ;
        RECT 67.680 170.830 68.000 170.890 ;
        RECT 70.440 170.830 70.760 170.890 ;
        RECT 75.100 170.830 75.390 170.875 ;
        RECT 66.775 170.690 68.600 170.830 ;
        RECT 66.775 170.645 67.065 170.690 ;
        RECT 67.680 170.630 68.000 170.690 ;
        RECT 56.655 170.490 56.945 170.535 ;
        RECT 62.620 170.490 62.940 170.550 ;
        RECT 56.655 170.350 62.940 170.490 ;
        RECT 56.655 170.305 56.945 170.350 ;
        RECT 62.620 170.290 62.940 170.350 ;
        RECT 67.220 170.290 67.540 170.550 ;
        RECT 56.195 170.150 56.485 170.195 ;
        RECT 58.480 170.150 58.800 170.210 ;
        RECT 56.195 170.010 58.800 170.150 ;
        RECT 68.460 170.150 68.600 170.690 ;
        RECT 70.440 170.690 75.390 170.830 ;
        RECT 70.440 170.630 70.760 170.690 ;
        RECT 75.100 170.645 75.390 170.690 ;
        RECT 75.960 170.830 76.280 170.890 ;
        RECT 76.435 170.830 76.725 170.875 ;
        RECT 75.960 170.690 76.725 170.830 ;
        RECT 75.960 170.630 76.280 170.690 ;
        RECT 76.435 170.645 76.725 170.690 ;
        RECT 100.050 170.840 101.820 170.890 ;
        RECT 71.845 170.490 72.135 170.535 ;
        RECT 74.365 170.490 74.655 170.535 ;
        RECT 75.555 170.490 75.845 170.535 ;
        RECT 71.845 170.350 75.845 170.490 ;
        RECT 71.845 170.305 72.135 170.350 ;
        RECT 74.365 170.305 74.655 170.350 ;
        RECT 75.555 170.305 75.845 170.350 ;
        RECT 69.535 170.150 69.825 170.195 ;
        RECT 68.460 170.010 69.825 170.150 ;
        RECT 56.195 169.965 56.485 170.010 ;
        RECT 58.480 169.950 58.800 170.010 ;
        RECT 69.535 169.965 69.825 170.010 ;
        RECT 72.280 170.150 72.570 170.195 ;
        RECT 73.850 170.150 74.140 170.195 ;
        RECT 75.950 170.150 76.240 170.195 ;
        RECT 72.280 170.010 76.240 170.150 ;
        RECT 72.280 169.965 72.570 170.010 ;
        RECT 73.850 169.965 74.140 170.010 ;
        RECT 75.950 169.965 76.240 170.010 ;
        RECT 55.275 169.810 55.565 169.855 ;
        RECT 50.200 169.670 55.565 169.810 ;
        RECT 50.200 169.610 50.520 169.670 ;
        RECT 53.880 169.610 54.200 169.670 ;
        RECT 55.275 169.625 55.565 169.670 ;
        RECT 56.655 169.810 56.945 169.855 ;
        RECT 58.940 169.810 59.260 169.870 ;
        RECT 56.655 169.670 59.260 169.810 ;
        RECT 56.655 169.625 56.945 169.670 ;
        RECT 58.940 169.610 59.260 169.670 ;
        RECT 59.400 169.610 59.720 169.870 ;
        RECT 60.320 169.810 60.640 169.870 ;
        RECT 69.980 169.810 70.300 169.870 ;
        RECT 60.320 169.670 70.300 169.810 ;
        RECT 60.320 169.610 60.640 169.670 ;
        RECT 69.980 169.610 70.300 169.670 ;
        RECT 11.950 168.990 90.610 169.470 ;
        RECT 21.220 168.590 21.540 168.850 ;
        RECT 22.155 168.790 22.445 168.835 ;
        RECT 25.375 168.790 25.665 168.835 ;
        RECT 40.540 168.790 40.860 168.850 ;
        RECT 22.155 168.650 25.665 168.790 ;
        RECT 22.155 168.605 22.445 168.650 ;
        RECT 25.375 168.605 25.665 168.650 ;
        RECT 35.110 168.650 40.860 168.790 ;
        RECT 23.995 168.450 24.285 168.495 ;
        RECT 26.740 168.450 27.060 168.510 ;
        RECT 23.995 168.310 27.060 168.450 ;
        RECT 23.995 168.265 24.285 168.310 ;
        RECT 26.740 168.250 27.060 168.310 ;
        RECT 30.420 168.110 30.740 168.170 ;
        RECT 27.750 167.970 30.740 168.110 ;
        RECT 27.750 167.830 27.890 167.970 ;
        RECT 30.420 167.910 30.740 167.970 ;
        RECT 25.820 167.770 26.140 167.830 ;
        RECT 26.295 167.770 26.585 167.815 ;
        RECT 25.820 167.630 26.585 167.770 ;
        RECT 25.820 167.570 26.140 167.630 ;
        RECT 26.295 167.585 26.585 167.630 ;
        RECT 26.370 167.430 26.510 167.585 ;
        RECT 27.660 167.570 27.980 167.830 ;
        RECT 29.500 167.570 29.820 167.830 ;
        RECT 34.100 167.570 34.420 167.830 ;
        RECT 35.110 167.815 35.250 168.650 ;
        RECT 40.540 168.590 40.860 168.650 ;
        RECT 46.520 168.590 46.840 168.850 ;
        RECT 49.740 168.790 50.060 168.850 ;
        RECT 50.215 168.790 50.505 168.835 ;
        RECT 49.740 168.650 50.505 168.790 ;
        RECT 49.740 168.590 50.060 168.650 ;
        RECT 50.215 168.605 50.505 168.650 ;
        RECT 52.960 168.790 53.280 168.850 ;
        RECT 55.720 168.790 56.040 168.850 ;
        RECT 52.960 168.650 56.040 168.790 ;
        RECT 52.960 168.590 53.280 168.650 ;
        RECT 55.720 168.590 56.040 168.650 ;
        RECT 70.440 168.590 70.760 168.850 ;
        RECT 71.375 168.790 71.665 168.835 ;
        RECT 71.820 168.790 72.140 168.850 ;
        RECT 71.375 168.650 72.140 168.790 ;
        RECT 71.375 168.605 71.665 168.650 ;
        RECT 40.120 168.450 40.410 168.495 ;
        RECT 42.220 168.450 42.510 168.495 ;
        RECT 43.790 168.450 44.080 168.495 ;
        RECT 40.120 168.310 44.080 168.450 ;
        RECT 40.120 168.265 40.410 168.310 ;
        RECT 42.220 168.265 42.510 168.310 ;
        RECT 43.790 168.265 44.080 168.310 ;
        RECT 47.900 168.450 48.220 168.510 ;
        RECT 53.420 168.450 53.740 168.510 ;
        RECT 55.275 168.450 55.565 168.495 ;
        RECT 47.900 168.310 62.390 168.450 ;
        RECT 47.900 168.250 48.220 168.310 ;
        RECT 53.420 168.250 53.740 168.310 ;
        RECT 55.275 168.265 55.565 168.310 ;
        RECT 62.250 168.170 62.390 168.310 ;
        RECT 40.515 168.110 40.805 168.155 ;
        RECT 41.705 168.110 41.995 168.155 ;
        RECT 44.225 168.110 44.515 168.155 ;
        RECT 40.515 167.970 44.515 168.110 ;
        RECT 40.515 167.925 40.805 167.970 ;
        RECT 41.705 167.925 41.995 167.970 ;
        RECT 44.225 167.925 44.515 167.970 ;
        RECT 47.070 167.970 52.270 168.110 ;
        RECT 35.035 167.585 35.325 167.815 ;
        RECT 36.415 167.770 36.705 167.815 ;
        RECT 36.860 167.770 37.180 167.830 ;
        RECT 38.700 167.770 39.020 167.830 ;
        RECT 41.000 167.815 41.320 167.830 ;
        RECT 39.635 167.770 39.925 167.815 ;
        RECT 40.970 167.770 41.320 167.815 ;
        RECT 36.415 167.630 39.925 167.770 ;
        RECT 40.805 167.630 41.320 167.770 ;
        RECT 36.415 167.585 36.705 167.630 ;
        RECT 36.860 167.570 37.180 167.630 ;
        RECT 38.700 167.570 39.020 167.630 ;
        RECT 39.635 167.585 39.925 167.630 ;
        RECT 40.970 167.585 41.320 167.630 ;
        RECT 41.000 167.570 41.320 167.585 ;
        RECT 43.300 167.770 43.620 167.830 ;
        RECT 47.070 167.815 47.210 167.970 ;
        RECT 46.995 167.770 47.285 167.815 ;
        RECT 43.300 167.630 47.285 167.770 ;
        RECT 43.300 167.570 43.620 167.630 ;
        RECT 46.995 167.585 47.285 167.630 ;
        RECT 47.900 167.570 48.220 167.830 ;
        RECT 48.375 167.585 48.665 167.815 ;
        RECT 48.835 167.770 49.125 167.815 ;
        RECT 50.200 167.770 50.520 167.830 ;
        RECT 48.835 167.630 50.520 167.770 ;
        RECT 48.835 167.585 49.125 167.630 ;
        RECT 28.120 167.430 28.440 167.490 ;
        RECT 26.370 167.290 28.440 167.430 ;
        RECT 28.120 167.230 28.440 167.290 ;
        RECT 35.955 167.430 36.245 167.475 ;
        RECT 41.460 167.430 41.780 167.490 ;
        RECT 35.955 167.290 41.780 167.430 ;
        RECT 35.955 167.245 36.245 167.290 ;
        RECT 41.460 167.230 41.780 167.290 ;
        RECT 43.760 167.430 44.080 167.490 ;
        RECT 48.450 167.430 48.590 167.585 ;
        RECT 50.200 167.570 50.520 167.630 ;
        RECT 51.135 167.770 51.425 167.815 ;
        RECT 51.580 167.770 51.900 167.830 ;
        RECT 52.130 167.815 52.270 167.970 ;
        RECT 56.180 167.910 56.500 168.170 ;
        RECT 57.100 168.110 57.420 168.170 ;
        RECT 60.335 168.110 60.625 168.155 ;
        RECT 60.780 168.110 61.100 168.170 ;
        RECT 57.100 167.970 61.100 168.110 ;
        RECT 57.100 167.910 57.420 167.970 ;
        RECT 60.335 167.925 60.625 167.970 ;
        RECT 60.780 167.910 61.100 167.970 ;
        RECT 62.160 167.910 62.480 168.170 ;
        RECT 64.475 168.110 64.765 168.155 ;
        RECT 67.220 168.110 67.540 168.170 ;
        RECT 71.450 168.110 71.590 168.605 ;
        RECT 71.820 168.590 72.140 168.650 ;
        RECT 64.475 167.970 67.540 168.110 ;
        RECT 64.475 167.925 64.765 167.970 ;
        RECT 67.220 167.910 67.540 167.970 ;
        RECT 68.460 167.970 71.590 168.110 ;
        RECT 51.135 167.630 51.900 167.770 ;
        RECT 51.135 167.585 51.425 167.630 ;
        RECT 43.760 167.290 48.590 167.430 ;
        RECT 49.280 167.430 49.600 167.490 ;
        RECT 51.210 167.430 51.350 167.585 ;
        RECT 51.580 167.570 51.900 167.630 ;
        RECT 52.055 167.585 52.345 167.815 ;
        RECT 52.515 167.585 52.805 167.815 ;
        RECT 52.590 167.430 52.730 167.585 ;
        RECT 56.640 167.570 56.960 167.830 ;
        RECT 59.400 167.770 59.720 167.830 ;
        RECT 62.635 167.770 62.925 167.815 ;
        RECT 57.650 167.630 62.925 167.770 ;
        RECT 57.650 167.490 57.790 167.630 ;
        RECT 59.400 167.570 59.720 167.630 ;
        RECT 62.635 167.585 62.925 167.630 ;
        RECT 53.895 167.430 54.185 167.475 ;
        RECT 57.560 167.430 57.880 167.490 ;
        RECT 49.280 167.290 51.350 167.430 ;
        RECT 51.670 167.290 57.880 167.430 ;
        RECT 43.760 167.230 44.080 167.290 ;
        RECT 49.280 167.230 49.600 167.290 ;
        RECT 22.155 167.090 22.445 167.135 ;
        RECT 23.980 167.090 24.300 167.150 ;
        RECT 26.280 167.090 26.600 167.150 ;
        RECT 22.155 166.950 26.600 167.090 ;
        RECT 22.155 166.905 22.445 166.950 ;
        RECT 23.980 166.890 24.300 166.950 ;
        RECT 26.280 166.890 26.600 166.950 ;
        RECT 26.740 167.090 27.060 167.150 ;
        RECT 27.215 167.090 27.505 167.135 ;
        RECT 35.480 167.090 35.800 167.150 ;
        RECT 26.740 166.950 35.800 167.090 ;
        RECT 26.740 166.890 27.060 166.950 ;
        RECT 27.215 166.905 27.505 166.950 ;
        RECT 35.480 166.890 35.800 166.950 ;
        RECT 37.780 167.090 38.100 167.150 ;
        RECT 51.670 167.090 51.810 167.290 ;
        RECT 53.895 167.245 54.185 167.290 ;
        RECT 57.560 167.230 57.880 167.290 ;
        RECT 37.780 166.950 51.810 167.090 ;
        RECT 37.780 166.890 38.100 166.950 ;
        RECT 52.040 166.890 52.360 167.150 ;
        RECT 52.500 167.090 52.820 167.150 ;
        RECT 68.460 167.090 68.600 167.970 ;
        RECT 69.535 167.770 69.825 167.815 ;
        RECT 75.960 167.770 76.280 167.830 ;
        RECT 69.535 167.630 76.280 167.770 ;
        RECT 69.535 167.585 69.825 167.630 ;
        RECT 75.960 167.570 76.280 167.630 ;
        RECT 100.050 167.500 100.880 170.840 ;
        RECT 108.930 170.540 116.850 170.550 ;
        RECT 105.160 170.530 116.850 170.540 ;
        RECT 101.540 170.410 116.850 170.530 ;
        RECT 101.540 170.400 116.875 170.410 ;
        RECT 101.500 170.280 116.875 170.400 ;
        RECT 101.500 170.170 105.500 170.280 ;
        RECT 101.110 169.830 101.340 170.120 ;
        RECT 101.560 169.830 105.450 170.170 ;
        RECT 105.660 169.830 105.890 170.120 ;
        RECT 101.110 168.460 105.890 169.830 ;
        RECT 101.110 168.160 101.340 168.460 ;
        RECT 105.660 168.160 105.890 168.460 ;
        RECT 101.500 167.880 105.500 168.110 ;
        RECT 101.750 167.650 105.320 167.880 ;
        RECT 101.750 167.500 105.440 167.650 ;
        RECT 70.900 167.475 71.220 167.490 ;
        RECT 70.900 167.245 71.505 167.475 ;
        RECT 70.900 167.230 71.220 167.245 ;
        RECT 72.280 167.230 72.600 167.490 ;
        RECT 100.050 167.240 105.440 167.500 ;
        RECT 106.690 167.330 107.310 170.280 ;
        RECT 108.875 170.180 116.875 170.280 ;
        RECT 108.930 170.170 116.850 170.180 ;
        RECT 108.440 169.470 108.670 170.130 ;
        RECT 109.450 169.470 110.450 169.560 ;
        RECT 117.080 169.470 117.310 170.130 ;
        RECT 108.440 168.650 117.310 169.470 ;
        RECT 108.440 168.170 108.670 168.650 ;
        RECT 109.450 168.560 110.450 168.650 ;
        RECT 117.080 168.170 117.310 168.650 ;
        RECT 108.875 167.890 116.875 168.120 ;
        RECT 52.500 166.950 68.600 167.090 ;
        RECT 100.010 167.220 105.440 167.240 ;
        RECT 52.500 166.890 52.820 166.950 ;
        RECT 100.010 166.760 105.450 167.220 ;
        RECT 11.950 166.270 90.610 166.750 ;
        RECT 25.835 166.070 26.125 166.115 ;
        RECT 27.660 166.070 27.980 166.130 ;
        RECT 25.835 165.930 27.980 166.070 ;
        RECT 25.835 165.885 26.125 165.930 ;
        RECT 27.660 165.870 27.980 165.930 ;
        RECT 32.260 166.070 32.580 166.130 ;
        RECT 44.680 166.070 45.000 166.130 ;
        RECT 58.940 166.070 59.260 166.130 ;
        RECT 32.260 165.930 59.260 166.070 ;
        RECT 32.260 165.870 32.580 165.930 ;
        RECT 44.680 165.870 45.000 165.930 ;
        RECT 58.940 165.870 59.260 165.930 ;
        RECT 63.095 166.070 63.385 166.115 ;
        RECT 64.920 166.070 65.240 166.130 ;
        RECT 63.095 165.930 65.240 166.070 ;
        RECT 63.095 165.885 63.385 165.930 ;
        RECT 64.920 165.870 65.240 165.930 ;
        RECT 22.615 165.730 22.905 165.775 ;
        RECT 27.200 165.730 27.520 165.790 ;
        RECT 22.615 165.590 27.520 165.730 ;
        RECT 22.615 165.545 22.905 165.590 ;
        RECT 27.200 165.530 27.520 165.590 ;
        RECT 35.035 165.730 35.325 165.775 ;
        RECT 37.780 165.730 38.100 165.790 ;
        RECT 35.035 165.590 38.100 165.730 ;
        RECT 35.035 165.545 35.325 165.590 ;
        RECT 37.780 165.530 38.100 165.590 ;
        RECT 56.640 165.730 56.960 165.790 ;
        RECT 65.840 165.730 66.160 165.790 ;
        RECT 67.235 165.730 67.525 165.775 ;
        RECT 56.640 165.590 67.525 165.730 ;
        RECT 56.640 165.530 56.960 165.590 ;
        RECT 65.840 165.530 66.160 165.590 ;
        RECT 67.235 165.545 67.525 165.590 ;
        RECT 71.375 165.730 71.665 165.775 ;
        RECT 75.960 165.730 76.280 165.790 ;
        RECT 71.375 165.590 76.280 165.730 ;
        RECT 71.375 165.545 71.665 165.590 ;
        RECT 75.960 165.530 76.280 165.590 ;
        RECT 23.535 165.205 23.825 165.435 ;
        RECT 23.610 165.050 23.750 165.205 ;
        RECT 26.280 165.190 26.600 165.450 ;
        RECT 26.755 165.390 27.045 165.435 ;
        RECT 28.120 165.390 28.440 165.450 ;
        RECT 26.755 165.250 30.650 165.390 ;
        RECT 26.755 165.205 27.045 165.250 ;
        RECT 28.120 165.190 28.440 165.250 ;
        RECT 29.055 165.050 29.345 165.095 ;
        RECT 29.500 165.050 29.820 165.110 ;
        RECT 23.610 164.910 27.890 165.050 ;
        RECT 27.750 164.755 27.890 164.910 ;
        RECT 29.055 164.910 29.820 165.050 ;
        RECT 30.510 165.050 30.650 165.250 ;
        RECT 32.720 165.190 33.040 165.450 ;
        RECT 34.115 165.205 34.405 165.435 ;
        RECT 35.495 165.390 35.785 165.435 ;
        RECT 35.940 165.390 36.260 165.450 ;
        RECT 35.495 165.250 36.260 165.390 ;
        RECT 35.495 165.205 35.785 165.250 ;
        RECT 33.640 165.050 33.960 165.110 ;
        RECT 34.190 165.050 34.330 165.205 ;
        RECT 35.940 165.190 36.260 165.250 ;
        RECT 57.100 165.190 57.420 165.450 ;
        RECT 57.560 165.390 57.880 165.450 ;
        RECT 62.160 165.435 62.480 165.450 ;
        RECT 61.255 165.390 61.545 165.435 ;
        RECT 57.560 165.250 61.545 165.390 ;
        RECT 57.560 165.190 57.880 165.250 ;
        RECT 61.255 165.205 61.545 165.250 ;
        RECT 62.025 165.205 62.480 165.435 ;
        RECT 62.160 165.190 62.480 165.205 ;
        RECT 62.620 165.390 62.940 165.450 ;
        RECT 64.475 165.390 64.765 165.435 ;
        RECT 62.620 165.250 64.765 165.390 ;
        RECT 62.620 165.190 62.940 165.250 ;
        RECT 64.475 165.205 64.765 165.250 ;
        RECT 100.010 165.410 102.050 166.760 ;
        RECT 103.800 166.750 105.450 166.760 ;
        RECT 102.490 165.480 103.490 166.200 ;
        RECT 103.800 165.940 104.110 166.750 ;
        RECT 104.570 166.470 105.450 166.750 ;
        RECT 105.690 166.930 107.310 167.330 ;
        RECT 108.960 166.980 116.830 167.890 ;
        RECT 104.510 166.240 105.510 166.470 ;
        RECT 105.690 166.280 106.040 166.930 ;
        RECT 106.690 166.920 107.310 166.930 ;
        RECT 108.875 166.750 116.875 166.980 ;
        RECT 108.960 166.740 116.830 166.750 ;
        RECT 104.570 166.030 105.450 166.050 ;
        RECT 103.840 165.650 104.110 165.940 ;
        RECT 104.510 165.800 105.510 166.030 ;
        RECT 105.670 165.990 106.040 166.280 ;
        RECT 105.700 165.930 106.040 165.990 ;
        RECT 106.800 166.600 107.560 166.650 ;
        RECT 108.440 166.600 108.670 166.700 ;
        RECT 106.800 166.390 108.670 166.600 ;
        RECT 117.080 166.390 117.310 166.700 ;
        RECT 106.800 165.970 109.340 166.390 ;
        RECT 116.710 165.970 117.310 166.390 ;
        RECT 104.570 165.650 105.450 165.800 ;
        RECT 104.580 165.480 105.310 165.650 ;
        RECT 36.400 165.050 36.720 165.110 ;
        RECT 30.510 164.910 36.720 165.050 ;
        RECT 29.055 164.865 29.345 164.910 ;
        RECT 29.500 164.850 29.820 164.910 ;
        RECT 33.640 164.850 33.960 164.910 ;
        RECT 36.400 164.850 36.720 164.910 ;
        RECT 27.675 164.710 27.965 164.755 ;
        RECT 30.420 164.710 30.740 164.770 ;
        RECT 27.675 164.570 30.740 164.710 ;
        RECT 27.675 164.525 27.965 164.570 ;
        RECT 30.420 164.510 30.740 164.570 ;
        RECT 24.440 164.170 24.760 164.430 ;
        RECT 24.900 164.170 25.220 164.430 ;
        RECT 31.340 164.370 31.660 164.430 ;
        RECT 33.195 164.370 33.485 164.415 ;
        RECT 31.340 164.230 33.485 164.370 ;
        RECT 62.250 164.370 62.390 165.190 ;
        RECT 63.540 164.370 63.860 164.430 ;
        RECT 64.935 164.370 65.225 164.415 ;
        RECT 62.250 164.230 65.225 164.370 ;
        RECT 31.340 164.170 31.660 164.230 ;
        RECT 33.195 164.185 33.485 164.230 ;
        RECT 63.540 164.170 63.860 164.230 ;
        RECT 64.935 164.185 65.225 164.230 ;
        RECT 11.950 163.550 90.610 164.030 ;
        RECT 24.440 163.350 24.760 163.410 ;
        RECT 27.215 163.350 27.505 163.395 ;
        RECT 24.440 163.210 27.505 163.350 ;
        RECT 24.440 163.150 24.760 163.210 ;
        RECT 27.215 163.165 27.505 163.210 ;
        RECT 29.960 163.350 30.280 163.410 ;
        RECT 30.435 163.350 30.725 163.395 ;
        RECT 35.940 163.350 36.260 163.410 ;
        RECT 29.960 163.210 30.725 163.350 ;
        RECT 29.960 163.150 30.280 163.210 ;
        RECT 30.435 163.165 30.725 163.210 ;
        RECT 30.970 163.210 36.260 163.350 ;
        RECT 24.900 163.010 25.220 163.070 ;
        RECT 25.375 163.010 25.665 163.055 ;
        RECT 24.900 162.870 25.665 163.010 ;
        RECT 24.900 162.810 25.220 162.870 ;
        RECT 25.375 162.825 25.665 162.870 ;
        RECT 30.970 162.670 31.110 163.210 ;
        RECT 35.940 163.150 36.260 163.210 ;
        RECT 41.460 163.350 41.780 163.410 ;
        RECT 41.460 163.210 55.030 163.350 ;
        RECT 41.460 163.150 41.780 163.210 ;
        RECT 32.260 163.010 32.580 163.070 ;
        RECT 33.640 163.010 33.960 163.070 ;
        RECT 35.035 163.010 35.325 163.055 ;
        RECT 32.260 162.870 32.950 163.010 ;
        RECT 32.260 162.810 32.580 162.870 ;
        RECT 28.210 162.530 31.110 162.670 ;
        RECT 21.220 162.330 21.540 162.390 ;
        RECT 21.220 162.190 26.050 162.330 ;
        RECT 21.220 162.130 21.540 162.190 ;
        RECT 25.910 161.990 26.050 162.190 ;
        RECT 27.215 161.990 27.505 162.035 ;
        RECT 25.910 161.850 27.505 161.990 ;
        RECT 28.210 161.990 28.350 162.530 ;
        RECT 28.595 162.330 28.885 162.375 ;
        RECT 30.880 162.330 31.200 162.390 ;
        RECT 28.595 162.190 31.200 162.330 ;
        RECT 28.595 162.145 28.885 162.190 ;
        RECT 30.880 162.130 31.200 162.190 ;
        RECT 31.340 162.130 31.660 162.390 ;
        RECT 32.810 162.375 32.950 162.870 ;
        RECT 33.640 162.870 35.325 163.010 ;
        RECT 33.640 162.810 33.960 162.870 ;
        RECT 35.035 162.825 35.325 162.870 ;
        RECT 37.320 163.010 37.640 163.070 ;
        RECT 37.320 162.870 49.510 163.010 ;
        RECT 37.320 162.810 37.640 162.870 ;
        RECT 33.180 162.470 33.500 162.730 ;
        RECT 35.495 162.670 35.785 162.715 ;
        RECT 34.190 162.530 35.785 162.670 ;
        RECT 34.190 162.375 34.330 162.530 ;
        RECT 35.495 162.485 35.785 162.530 ;
        RECT 35.940 162.670 36.260 162.730 ;
        RECT 35.940 162.530 37.550 162.670 ;
        RECT 35.940 162.470 36.260 162.530 ;
        RECT 32.275 162.330 32.565 162.375 ;
        RECT 32.165 162.190 32.565 162.330 ;
        RECT 32.275 162.145 32.565 162.190 ;
        RECT 32.735 162.330 33.025 162.375 ;
        RECT 32.735 162.190 33.135 162.330 ;
        RECT 32.735 162.145 33.025 162.190 ;
        RECT 34.115 162.145 34.405 162.375 ;
        RECT 29.515 161.990 29.805 162.035 ;
        RECT 28.210 161.850 29.805 161.990 ;
        RECT 27.215 161.805 27.505 161.850 ;
        RECT 29.515 161.805 29.805 161.850 ;
        RECT 30.420 161.990 30.740 162.050 ;
        RECT 32.350 161.990 32.490 162.145 ;
        RECT 30.420 161.850 32.490 161.990 ;
        RECT 32.810 161.990 32.950 162.145 ;
        RECT 36.400 162.130 36.720 162.390 ;
        RECT 37.410 162.375 37.550 162.530 ;
        RECT 41.460 162.470 41.780 162.730 ;
        RECT 49.370 162.715 49.510 162.870 ;
        RECT 49.295 162.485 49.585 162.715 ;
        RECT 37.335 162.145 37.625 162.375 ;
        RECT 37.780 162.130 38.100 162.390 ;
        RECT 41.000 162.130 41.320 162.390 ;
        RECT 48.375 162.330 48.665 162.375 ;
        RECT 41.550 162.190 48.665 162.330 ;
        RECT 33.180 161.990 33.500 162.050 ;
        RECT 32.810 161.850 33.500 161.990 ;
        RECT 30.420 161.790 30.740 161.850 ;
        RECT 33.180 161.790 33.500 161.850 ;
        RECT 40.540 161.990 40.860 162.050 ;
        RECT 41.550 161.990 41.690 162.190 ;
        RECT 48.375 162.145 48.665 162.190 ;
        RECT 48.820 162.130 49.140 162.390 ;
        RECT 49.755 162.330 50.045 162.375 ;
        RECT 52.960 162.330 53.280 162.390 ;
        RECT 54.890 162.375 55.030 163.210 ;
        RECT 59.490 162.870 67.450 163.010 ;
        RECT 58.035 162.670 58.325 162.715 ;
        RECT 58.035 162.530 59.170 162.670 ;
        RECT 58.035 162.485 58.325 162.530 ;
        RECT 53.435 162.330 53.725 162.375 ;
        RECT 49.755 162.190 53.725 162.330 ;
        RECT 49.755 162.145 50.045 162.190 ;
        RECT 52.960 162.130 53.280 162.190 ;
        RECT 53.435 162.145 53.725 162.190 ;
        RECT 54.815 162.145 55.105 162.375 ;
        RECT 57.560 162.130 57.880 162.390 ;
        RECT 59.030 162.375 59.170 162.530 ;
        RECT 58.495 162.330 58.785 162.375 ;
        RECT 58.385 162.190 58.785 162.330 ;
        RECT 59.030 162.190 59.345 162.375 ;
        RECT 58.495 162.145 58.785 162.190 ;
        RECT 59.055 162.145 59.345 162.190 ;
        RECT 40.540 161.850 41.690 161.990 ;
        RECT 46.535 161.990 46.825 162.035 ;
        RECT 46.535 161.850 53.650 161.990 ;
        RECT 40.540 161.790 40.860 161.850 ;
        RECT 46.535 161.805 46.825 161.850 ;
        RECT 53.510 161.710 53.650 161.850 ;
        RECT 54.355 161.805 54.645 162.035 ;
        RECT 58.570 161.990 58.710 162.145 ;
        RECT 59.490 161.990 59.630 162.870 ;
        RECT 62.175 162.670 62.465 162.715 ;
        RECT 59.950 162.530 62.465 162.670 ;
        RECT 59.950 162.375 60.090 162.530 ;
        RECT 62.175 162.485 62.465 162.530 ;
        RECT 66.775 162.485 67.065 162.715 ;
        RECT 59.875 162.145 60.165 162.375 ;
        RECT 60.335 162.145 60.625 162.375 ;
        RECT 60.915 162.330 61.205 162.375 ;
        RECT 63.540 162.330 63.860 162.390 ;
        RECT 60.870 162.145 61.205 162.330 ;
        RECT 63.345 162.190 63.860 162.330 ;
        RECT 60.410 161.990 60.550 162.145 ;
        RECT 58.570 161.850 60.550 161.990 ;
        RECT 28.120 161.450 28.440 161.710 ;
        RECT 39.160 161.450 39.480 161.710 ;
        RECT 46.060 161.450 46.380 161.710 ;
        RECT 46.980 161.650 47.300 161.710 ;
        RECT 47.455 161.650 47.745 161.695 ;
        RECT 46.980 161.510 47.745 161.650 ;
        RECT 46.980 161.450 47.300 161.510 ;
        RECT 47.455 161.465 47.745 161.510 ;
        RECT 52.040 161.650 52.360 161.710 ;
        RECT 52.515 161.650 52.805 161.695 ;
        RECT 52.040 161.510 52.805 161.650 ;
        RECT 52.040 161.450 52.360 161.510 ;
        RECT 52.515 161.465 52.805 161.510 ;
        RECT 53.420 161.450 53.740 161.710 ;
        RECT 53.880 161.650 54.200 161.710 ;
        RECT 54.430 161.650 54.570 161.805 ;
        RECT 55.735 161.650 56.025 161.695 ;
        RECT 60.870 161.650 61.010 162.145 ;
        RECT 63.540 162.130 63.860 162.190 ;
        RECT 64.000 162.330 64.320 162.390 ;
        RECT 66.850 162.330 66.990 162.485 ;
        RECT 67.310 162.375 67.450 162.870 ;
        RECT 69.075 162.670 69.365 162.715 ;
        RECT 71.960 162.670 72.250 162.715 ;
        RECT 69.075 162.530 72.250 162.670 ;
        RECT 69.075 162.485 69.365 162.530 ;
        RECT 71.960 162.485 72.250 162.530 ;
        RECT 64.000 162.190 66.990 162.330 ;
        RECT 67.235 162.330 67.525 162.375 ;
        RECT 68.600 162.330 68.920 162.390 ;
        RECT 67.235 162.190 68.920 162.330 ;
        RECT 64.000 162.130 64.320 162.190 ;
        RECT 67.235 162.145 67.525 162.190 ;
        RECT 68.600 162.130 68.920 162.190 ;
        RECT 69.520 162.130 69.840 162.390 ;
        RECT 70.900 162.130 71.220 162.390 ;
        RECT 71.360 162.130 71.680 162.390 ;
        RECT 100.010 161.770 100.780 165.410 ;
        RECT 102.460 164.360 105.310 165.480 ;
        RECT 105.700 165.180 106.050 165.930 ;
        RECT 106.800 165.810 108.670 165.970 ;
        RECT 106.800 165.760 107.560 165.810 ;
        RECT 108.440 165.740 108.670 165.810 ;
        RECT 117.080 165.740 117.310 165.970 ;
        RECT 108.875 165.460 116.875 165.690 ;
        RECT 105.700 165.120 105.990 165.180 ;
        RECT 105.610 165.000 105.990 165.120 ;
        RECT 108.970 165.060 116.830 165.460 ;
        RECT 117.640 165.060 118.600 174.540 ;
        RECT 119.930 174.510 125.370 174.620 ;
        RECT 128.810 174.600 138.700 174.700 ;
        RECT 139.960 175.280 140.860 176.800 ;
        RECT 146.460 176.380 147.710 176.820 ;
        RECT 144.400 176.370 149.640 176.380 ;
        RECT 141.450 176.270 156.750 176.370 ;
        RECT 141.450 176.260 156.785 176.270 ;
        RECT 141.410 176.140 156.785 176.260 ;
        RECT 141.410 176.030 145.410 176.140 ;
        RECT 146.460 176.060 148.200 176.140 ;
        RECT 148.780 176.060 156.785 176.140 ;
        RECT 146.460 175.980 147.710 176.060 ;
        RECT 148.785 176.040 156.785 176.060 ;
        RECT 141.020 175.730 141.250 175.980 ;
        RECT 145.570 175.840 145.800 175.980 ;
        RECT 148.350 175.840 148.580 175.990 ;
        RECT 145.570 175.730 148.580 175.840 ;
        RECT 156.990 175.730 157.220 175.990 ;
        RECT 141.020 175.290 157.220 175.730 ;
        RECT 139.960 174.670 140.790 175.280 ;
        RECT 141.020 175.020 141.250 175.290 ;
        RECT 145.570 175.260 157.220 175.290 ;
        RECT 145.570 175.170 148.580 175.260 ;
        RECT 145.570 175.020 145.800 175.170 ;
        RECT 148.350 175.030 148.580 175.170 ;
        RECT 156.990 175.030 157.220 175.260 ;
        RECT 141.410 174.740 145.410 174.970 ;
        RECT 148.785 174.760 156.785 174.980 ;
        RECT 157.550 174.760 158.510 176.800 ;
        RECT 148.785 174.750 158.510 174.760 ;
        RECT 141.410 174.670 145.400 174.740 ;
        RECT 128.810 174.540 138.480 174.600 ;
        RECT 119.930 174.420 123.060 174.510 ;
        RECT 136.550 174.490 138.480 174.540 ;
        RECT 119.930 171.150 120.760 174.420 ;
        RECT 124.410 173.960 129.660 173.970 ;
        RECT 124.410 173.850 136.720 173.960 ;
        RECT 121.440 173.790 136.720 173.850 ;
        RECT 121.440 173.780 136.755 173.790 ;
        RECT 121.380 173.650 136.755 173.780 ;
        RECT 121.380 173.640 126.540 173.650 ;
        RECT 121.380 173.550 125.380 173.640 ;
        RECT 128.755 173.560 136.755 173.650 ;
        RECT 128.840 173.550 136.730 173.560 ;
        RECT 120.990 173.190 121.220 173.500 ;
        RECT 121.440 173.190 125.340 173.550 ;
        RECT 125.540 173.190 125.770 173.500 ;
        RECT 120.990 171.850 125.770 173.190 ;
        RECT 120.990 171.540 121.220 171.850 ;
        RECT 125.540 171.540 125.770 171.850 ;
        RECT 128.320 172.970 128.550 173.510 ;
        RECT 129.360 172.970 130.370 173.000 ;
        RECT 136.960 172.970 137.190 173.510 ;
        RECT 128.320 172.070 137.190 172.970 ;
        RECT 128.320 171.550 128.550 172.070 ;
        RECT 129.360 172.000 130.370 172.070 ;
        RECT 136.960 171.550 137.190 172.070 ;
        RECT 121.380 171.260 125.380 171.490 ;
        RECT 128.755 171.270 136.755 171.500 ;
        RECT 119.930 171.110 121.060 171.150 ;
        RECT 119.930 171.030 121.300 171.110 ;
        RECT 121.670 171.040 125.330 171.260 ;
        RECT 121.670 171.030 123.110 171.040 ;
        RECT 119.930 170.990 123.110 171.030 ;
        RECT 119.930 170.900 122.620 170.990 ;
        RECT 128.820 170.980 136.710 171.270 ;
        RECT 119.930 170.840 121.950 170.900 ;
        RECT 119.930 170.790 121.700 170.840 ;
        RECT 119.930 167.450 120.760 170.790 ;
        RECT 128.810 170.490 136.730 170.500 ;
        RECT 125.040 170.480 136.730 170.490 ;
        RECT 121.420 170.360 136.730 170.480 ;
        RECT 121.420 170.350 136.755 170.360 ;
        RECT 121.380 170.230 136.755 170.350 ;
        RECT 121.380 170.120 125.380 170.230 ;
        RECT 120.990 169.780 121.220 170.070 ;
        RECT 121.440 169.780 125.330 170.120 ;
        RECT 125.540 169.780 125.770 170.070 ;
        RECT 120.990 168.410 125.770 169.780 ;
        RECT 120.990 168.110 121.220 168.410 ;
        RECT 125.540 168.110 125.770 168.410 ;
        RECT 121.380 167.830 125.380 168.060 ;
        RECT 121.630 167.600 125.200 167.830 ;
        RECT 121.630 167.450 125.320 167.600 ;
        RECT 119.930 167.170 125.320 167.450 ;
        RECT 126.570 167.280 127.190 170.230 ;
        RECT 128.755 170.130 136.755 170.230 ;
        RECT 128.810 170.120 136.730 170.130 ;
        RECT 128.320 169.420 128.550 170.080 ;
        RECT 129.330 169.420 130.330 169.510 ;
        RECT 136.960 169.420 137.190 170.080 ;
        RECT 128.320 168.600 137.190 169.420 ;
        RECT 128.320 168.120 128.550 168.600 ;
        RECT 129.330 168.510 130.330 168.600 ;
        RECT 136.960 168.120 137.190 168.600 ;
        RECT 128.755 167.840 136.755 168.070 ;
        RECT 119.930 166.710 125.330 167.170 ;
        RECT 119.930 165.370 121.930 166.710 ;
        RECT 123.680 166.700 125.330 166.710 ;
        RECT 122.370 165.430 123.370 166.150 ;
        RECT 123.680 165.890 123.990 166.700 ;
        RECT 124.450 166.420 125.330 166.700 ;
        RECT 125.570 166.880 127.190 167.280 ;
        RECT 128.840 166.930 136.710 167.840 ;
        RECT 124.390 166.190 125.390 166.420 ;
        RECT 125.570 166.230 125.920 166.880 ;
        RECT 126.570 166.870 127.190 166.880 ;
        RECT 128.755 166.700 136.755 166.930 ;
        RECT 128.840 166.690 136.710 166.700 ;
        RECT 124.450 165.980 125.330 166.000 ;
        RECT 123.720 165.600 123.990 165.890 ;
        RECT 124.390 165.750 125.390 165.980 ;
        RECT 125.550 165.940 125.920 166.230 ;
        RECT 125.580 165.880 125.920 165.940 ;
        RECT 126.680 166.550 127.440 166.600 ;
        RECT 128.320 166.550 128.550 166.650 ;
        RECT 126.680 166.340 128.550 166.550 ;
        RECT 136.960 166.340 137.190 166.650 ;
        RECT 126.680 165.920 129.220 166.340 ;
        RECT 136.590 165.920 137.190 166.340 ;
        RECT 124.450 165.600 125.330 165.750 ;
        RECT 124.460 165.430 125.190 165.600 ;
        RECT 102.400 164.130 105.400 164.360 ;
        RECT 105.610 164.170 105.950 165.000 ;
        RECT 107.960 164.990 118.600 165.060 ;
        RECT 102.450 164.100 105.310 164.130 ;
        RECT 102.450 164.080 103.620 164.100 ;
        RECT 104.580 164.090 105.310 164.100 ;
        RECT 102.400 163.690 105.400 163.920 ;
        RECT 105.605 163.880 105.950 164.170 ;
        RECT 106.140 163.950 118.600 164.990 ;
        RECT 120.000 165.360 121.930 165.370 ;
        RECT 106.140 163.930 118.560 163.950 ;
        RECT 105.610 163.770 105.950 163.880 ;
        RECT 106.180 163.920 111.850 163.930 ;
        RECT 112.850 163.920 118.560 163.930 ;
        RECT 102.490 163.520 105.350 163.690 ;
        RECT 106.180 163.520 106.610 163.920 ;
        RECT 102.460 163.150 106.610 163.520 ;
        RECT 53.880 161.510 61.010 161.650 ;
        RECT 53.880 161.450 54.200 161.510 ;
        RECT 55.735 161.465 56.025 161.510 ;
        RECT 61.700 161.450 62.020 161.710 ;
        RECT 72.755 161.650 73.045 161.695 ;
        RECT 73.200 161.650 73.520 161.710 ;
        RECT 72.755 161.510 73.520 161.650 ;
        RECT 72.755 161.465 73.045 161.510 ;
        RECT 73.200 161.450 73.520 161.510 ;
        RECT 11.950 160.830 90.610 161.310 ;
        RECT 23.075 160.445 23.365 160.675 ;
        RECT 23.150 159.950 23.290 160.445 ;
        RECT 29.960 160.430 30.280 160.690 ;
        RECT 30.420 160.630 30.740 160.690 ;
        RECT 31.355 160.630 31.645 160.675 ;
        RECT 30.420 160.490 31.645 160.630 ;
        RECT 30.420 160.430 30.740 160.490 ;
        RECT 31.355 160.445 31.645 160.490 ;
        RECT 37.335 160.630 37.625 160.675 ;
        RECT 41.460 160.630 41.780 160.690 ;
        RECT 45.615 160.630 45.905 160.675 ;
        RECT 48.820 160.630 49.140 160.690 ;
        RECT 37.335 160.490 41.780 160.630 ;
        RECT 45.405 160.490 49.140 160.630 ;
        RECT 37.335 160.445 37.625 160.490 ;
        RECT 41.460 160.430 41.780 160.490 ;
        RECT 45.615 160.445 45.905 160.490 ;
        RECT 28.120 160.290 28.440 160.350 ;
        RECT 28.640 160.290 28.930 160.335 ;
        RECT 28.120 160.150 28.930 160.290 ;
        RECT 28.120 160.090 28.440 160.150 ;
        RECT 28.640 160.105 28.930 160.150 ;
        RECT 30.050 159.950 30.190 160.430 ;
        RECT 40.540 160.290 40.860 160.350 ;
        RECT 36.490 160.150 40.860 160.290 ;
        RECT 32.260 159.950 32.580 160.010 ;
        RECT 36.490 159.995 36.630 160.150 ;
        RECT 40.540 160.090 40.860 160.150 ;
        RECT 41.000 160.290 41.320 160.350 ;
        RECT 45.690 160.290 45.830 160.445 ;
        RECT 48.820 160.430 49.140 160.490 ;
        RECT 52.960 160.430 53.280 160.690 ;
        RECT 60.780 160.290 61.100 160.350 ;
        RECT 72.280 160.290 72.600 160.350 ;
        RECT 73.200 160.335 73.520 160.350 ;
        RECT 41.000 160.150 45.830 160.290 ;
        RECT 46.150 160.150 61.100 160.290 ;
        RECT 41.000 160.090 41.320 160.150 ;
        RECT 23.150 159.810 32.580 159.950 ;
        RECT 32.260 159.750 32.580 159.810 ;
        RECT 36.415 159.765 36.705 159.995 ;
        RECT 37.320 159.950 37.640 160.010 ;
        RECT 38.240 159.950 38.560 160.010 ;
        RECT 37.320 159.810 38.560 159.950 ;
        RECT 37.320 159.750 37.640 159.810 ;
        RECT 38.240 159.750 38.560 159.810 ;
        RECT 38.700 159.750 39.020 160.010 ;
        RECT 40.080 159.995 40.400 160.010 ;
        RECT 46.150 159.995 46.290 160.150 ;
        RECT 60.780 160.090 61.100 160.150 ;
        RECT 68.460 160.150 72.600 160.290 ;
        RECT 47.440 159.995 47.760 160.010 ;
        RECT 40.050 159.765 40.400 159.995 ;
        RECT 46.075 159.765 46.365 159.995 ;
        RECT 47.410 159.765 47.760 159.995 ;
        RECT 40.080 159.750 40.400 159.765 ;
        RECT 47.440 159.750 47.760 159.765 ;
        RECT 52.040 159.950 52.360 160.010 ;
        RECT 55.735 159.950 56.025 159.995 ;
        RECT 52.040 159.810 56.025 159.950 ;
        RECT 52.040 159.750 52.360 159.810 ;
        RECT 55.735 159.765 56.025 159.810 ;
        RECT 56.180 159.950 56.500 160.010 ;
        RECT 56.655 159.950 56.945 159.995 ;
        RECT 56.180 159.810 56.945 159.950 ;
        RECT 56.180 159.750 56.500 159.810 ;
        RECT 56.655 159.765 56.945 159.810 ;
        RECT 57.115 159.950 57.405 159.995 ;
        RECT 64.000 159.950 64.320 160.010 ;
        RECT 68.460 159.950 68.600 160.150 ;
        RECT 72.280 160.090 72.600 160.150 ;
        RECT 73.170 160.105 73.520 160.335 ;
        RECT 73.200 160.090 73.520 160.105 ;
        RECT 74.120 160.090 74.440 160.350 ;
        RECT 74.210 159.950 74.350 160.090 ;
        RECT 57.115 159.810 68.600 159.950 ;
        RECT 71.450 159.810 74.350 159.950 ;
        RECT 57.115 159.765 57.405 159.810 ;
        RECT 64.000 159.750 64.320 159.810 ;
        RECT 71.450 159.670 71.590 159.810 ;
        RECT 100.010 159.670 100.880 161.770 ;
        RECT 106.550 161.380 107.800 161.820 ;
        RECT 117.700 161.800 118.560 163.920 ;
        RECT 120.000 161.800 120.770 165.360 ;
        RECT 122.340 164.310 125.190 165.430 ;
        RECT 125.580 165.130 125.930 165.880 ;
        RECT 126.680 165.760 128.550 165.920 ;
        RECT 126.680 165.710 127.440 165.760 ;
        RECT 128.320 165.690 128.550 165.760 ;
        RECT 136.960 165.690 137.190 165.920 ;
        RECT 128.755 165.410 136.755 165.640 ;
        RECT 125.580 165.070 125.870 165.130 ;
        RECT 125.490 164.950 125.870 165.070 ;
        RECT 128.850 165.010 136.710 165.410 ;
        RECT 137.520 165.010 138.480 174.490 ;
        RECT 139.960 174.560 145.400 174.670 ;
        RECT 148.840 174.590 158.510 174.750 ;
        RECT 139.960 174.470 143.090 174.560 ;
        RECT 156.580 174.540 158.510 174.590 ;
        RECT 139.960 171.200 140.790 174.470 ;
        RECT 144.440 174.010 149.690 174.020 ;
        RECT 144.440 173.900 156.750 174.010 ;
        RECT 141.470 173.840 156.750 173.900 ;
        RECT 141.470 173.830 156.785 173.840 ;
        RECT 141.410 173.700 156.785 173.830 ;
        RECT 141.410 173.690 146.570 173.700 ;
        RECT 141.410 173.600 145.410 173.690 ;
        RECT 148.785 173.610 156.785 173.700 ;
        RECT 148.870 173.600 156.760 173.610 ;
        RECT 141.020 173.240 141.250 173.550 ;
        RECT 141.470 173.240 145.370 173.600 ;
        RECT 145.570 173.240 145.800 173.550 ;
        RECT 141.020 171.900 145.800 173.240 ;
        RECT 141.020 171.590 141.250 171.900 ;
        RECT 145.570 171.590 145.800 171.900 ;
        RECT 148.350 173.020 148.580 173.560 ;
        RECT 149.390 173.020 150.400 173.050 ;
        RECT 156.990 173.020 157.220 173.560 ;
        RECT 148.350 172.120 157.220 173.020 ;
        RECT 148.350 171.600 148.580 172.120 ;
        RECT 149.390 172.050 150.400 172.120 ;
        RECT 156.990 171.600 157.220 172.120 ;
        RECT 141.410 171.310 145.410 171.540 ;
        RECT 148.785 171.320 156.785 171.550 ;
        RECT 139.960 171.160 141.090 171.200 ;
        RECT 139.960 171.080 141.330 171.160 ;
        RECT 141.700 171.090 145.360 171.310 ;
        RECT 141.700 171.080 143.140 171.090 ;
        RECT 139.960 171.040 143.140 171.080 ;
        RECT 139.960 170.950 142.650 171.040 ;
        RECT 148.850 171.030 156.740 171.320 ;
        RECT 139.960 170.890 141.980 170.950 ;
        RECT 139.960 170.840 141.730 170.890 ;
        RECT 139.960 167.500 140.790 170.840 ;
        RECT 148.840 170.540 156.760 170.550 ;
        RECT 145.070 170.530 156.760 170.540 ;
        RECT 141.450 170.410 156.760 170.530 ;
        RECT 141.450 170.400 156.785 170.410 ;
        RECT 141.410 170.280 156.785 170.400 ;
        RECT 141.410 170.170 145.410 170.280 ;
        RECT 141.020 169.830 141.250 170.120 ;
        RECT 141.470 169.830 145.360 170.170 ;
        RECT 145.570 169.830 145.800 170.120 ;
        RECT 141.020 168.460 145.800 169.830 ;
        RECT 141.020 168.160 141.250 168.460 ;
        RECT 145.570 168.160 145.800 168.460 ;
        RECT 141.410 167.880 145.410 168.110 ;
        RECT 141.660 167.650 145.230 167.880 ;
        RECT 141.660 167.500 145.350 167.650 ;
        RECT 139.960 167.270 145.350 167.500 ;
        RECT 146.600 167.330 147.220 170.280 ;
        RECT 148.785 170.180 156.785 170.280 ;
        RECT 148.840 170.170 156.760 170.180 ;
        RECT 148.350 169.470 148.580 170.130 ;
        RECT 149.360 169.470 150.360 169.560 ;
        RECT 156.990 169.470 157.220 170.130 ;
        RECT 148.350 168.650 157.220 169.470 ;
        RECT 148.350 168.170 148.580 168.650 ;
        RECT 149.360 168.560 150.360 168.650 ;
        RECT 156.990 168.170 157.220 168.650 ;
        RECT 148.785 167.890 156.785 168.120 ;
        RECT 122.280 164.080 125.280 164.310 ;
        RECT 125.490 164.120 125.830 164.950 ;
        RECT 127.840 164.940 138.480 165.010 ;
        RECT 122.330 164.050 125.190 164.080 ;
        RECT 122.330 164.030 123.500 164.050 ;
        RECT 124.460 164.040 125.190 164.050 ;
        RECT 122.280 163.640 125.280 163.870 ;
        RECT 125.485 163.830 125.830 164.120 ;
        RECT 126.020 163.900 138.480 164.940 ;
        RECT 139.930 167.220 145.350 167.270 ;
        RECT 139.930 166.760 145.360 167.220 ;
        RECT 139.930 165.410 141.960 166.760 ;
        RECT 143.710 166.750 145.360 166.760 ;
        RECT 142.400 165.480 143.400 166.200 ;
        RECT 143.710 165.940 144.020 166.750 ;
        RECT 144.480 166.470 145.360 166.750 ;
        RECT 145.600 166.930 147.220 167.330 ;
        RECT 148.870 166.980 156.740 167.890 ;
        RECT 144.420 166.240 145.420 166.470 ;
        RECT 145.600 166.280 145.950 166.930 ;
        RECT 146.600 166.920 147.220 166.930 ;
        RECT 148.785 166.750 156.785 166.980 ;
        RECT 148.870 166.740 156.740 166.750 ;
        RECT 144.480 166.030 145.360 166.050 ;
        RECT 143.750 165.650 144.020 165.940 ;
        RECT 144.420 165.800 145.420 166.030 ;
        RECT 145.580 165.990 145.950 166.280 ;
        RECT 145.610 165.930 145.950 165.990 ;
        RECT 146.710 166.600 147.470 166.650 ;
        RECT 148.350 166.600 148.580 166.700 ;
        RECT 146.710 166.390 148.580 166.600 ;
        RECT 156.990 166.390 157.220 166.700 ;
        RECT 146.710 165.970 149.250 166.390 ;
        RECT 156.620 165.970 157.220 166.390 ;
        RECT 144.480 165.650 145.360 165.800 ;
        RECT 144.490 165.480 145.220 165.650 ;
        RECT 126.020 163.880 138.460 163.900 ;
        RECT 125.490 163.720 125.830 163.830 ;
        RECT 126.060 163.870 131.730 163.880 ;
        RECT 132.730 163.870 138.460 163.880 ;
        RECT 122.370 163.470 125.230 163.640 ;
        RECT 126.060 163.470 126.490 163.870 ;
        RECT 122.340 163.100 126.490 163.470 ;
        RECT 104.490 161.370 109.730 161.380 ;
        RECT 101.540 161.270 116.840 161.370 ;
        RECT 101.540 161.260 116.875 161.270 ;
        RECT 101.500 161.140 116.875 161.260 ;
        RECT 101.500 161.030 105.500 161.140 ;
        RECT 106.550 161.060 108.290 161.140 ;
        RECT 108.870 161.060 116.875 161.140 ;
        RECT 106.550 160.980 107.800 161.060 ;
        RECT 108.875 161.040 116.875 161.060 ;
        RECT 101.110 160.730 101.340 160.980 ;
        RECT 105.660 160.840 105.890 160.980 ;
        RECT 108.440 160.840 108.670 160.990 ;
        RECT 105.660 160.730 108.670 160.840 ;
        RECT 117.080 160.730 117.310 160.990 ;
        RECT 101.110 160.290 117.310 160.730 ;
        RECT 101.110 160.020 101.340 160.290 ;
        RECT 105.660 160.260 117.310 160.290 ;
        RECT 105.660 160.170 108.670 160.260 ;
        RECT 105.660 160.020 105.890 160.170 ;
        RECT 108.440 160.030 108.670 160.170 ;
        RECT 117.080 160.030 117.310 160.260 ;
        RECT 101.500 159.740 105.500 159.970 ;
        RECT 108.875 159.760 116.875 159.980 ;
        RECT 117.640 159.760 118.600 161.800 ;
        RECT 108.875 159.750 118.600 159.760 ;
        RECT 101.500 159.670 105.490 159.740 ;
        RECT 25.385 159.610 25.675 159.655 ;
        RECT 27.905 159.610 28.195 159.655 ;
        RECT 29.095 159.610 29.385 159.655 ;
        RECT 25.385 159.470 29.385 159.610 ;
        RECT 25.385 159.425 25.675 159.470 ;
        RECT 27.905 159.425 28.195 159.470 ;
        RECT 29.095 159.425 29.385 159.470 ;
        RECT 29.960 159.410 30.280 159.670 ;
        RECT 33.655 159.610 33.945 159.655 ;
        RECT 34.560 159.610 34.880 159.670 ;
        RECT 33.655 159.470 34.880 159.610 ;
        RECT 33.655 159.425 33.945 159.470 ;
        RECT 34.560 159.410 34.880 159.470 ;
        RECT 39.595 159.610 39.885 159.655 ;
        RECT 40.785 159.610 41.075 159.655 ;
        RECT 43.305 159.610 43.595 159.655 ;
        RECT 39.595 159.470 43.595 159.610 ;
        RECT 39.595 159.425 39.885 159.470 ;
        RECT 40.785 159.425 41.075 159.470 ;
        RECT 43.305 159.425 43.595 159.470 ;
        RECT 46.955 159.610 47.245 159.655 ;
        RECT 48.145 159.610 48.435 159.655 ;
        RECT 50.665 159.610 50.955 159.655 ;
        RECT 46.955 159.470 50.955 159.610 ;
        RECT 46.955 159.425 47.245 159.470 ;
        RECT 48.145 159.425 48.435 159.470 ;
        RECT 50.665 159.425 50.955 159.470 ;
        RECT 53.420 159.610 53.740 159.670 ;
        RECT 71.360 159.610 71.680 159.670 ;
        RECT 53.420 159.470 71.680 159.610 ;
        RECT 53.420 159.410 53.740 159.470 ;
        RECT 71.360 159.410 71.680 159.470 ;
        RECT 71.835 159.610 72.125 159.655 ;
        RECT 72.715 159.610 73.005 159.655 ;
        RECT 73.905 159.610 74.195 159.655 ;
        RECT 76.425 159.610 76.715 159.655 ;
        RECT 71.835 159.425 72.175 159.610 ;
        RECT 72.715 159.470 76.715 159.610 ;
        RECT 72.715 159.425 73.005 159.470 ;
        RECT 73.905 159.425 74.195 159.470 ;
        RECT 76.425 159.425 76.715 159.470 ;
        RECT 100.010 159.560 105.490 159.670 ;
        RECT 108.930 159.590 118.600 159.750 ;
        RECT 100.010 159.470 103.180 159.560 ;
        RECT 116.670 159.540 118.600 159.590 ;
        RECT 25.820 159.270 26.110 159.315 ;
        RECT 27.390 159.270 27.680 159.315 ;
        RECT 29.490 159.270 29.780 159.315 ;
        RECT 25.820 159.130 29.780 159.270 ;
        RECT 25.820 159.085 26.110 159.130 ;
        RECT 27.390 159.085 27.680 159.130 ;
        RECT 29.490 159.085 29.780 159.130 ;
        RECT 39.200 159.270 39.490 159.315 ;
        RECT 41.300 159.270 41.590 159.315 ;
        RECT 42.870 159.270 43.160 159.315 ;
        RECT 39.200 159.130 43.160 159.270 ;
        RECT 39.200 159.085 39.490 159.130 ;
        RECT 41.300 159.085 41.590 159.130 ;
        RECT 42.870 159.085 43.160 159.130 ;
        RECT 46.560 159.270 46.850 159.315 ;
        RECT 48.660 159.270 48.950 159.315 ;
        RECT 50.230 159.270 50.520 159.315 ;
        RECT 46.560 159.130 50.520 159.270 ;
        RECT 46.560 159.085 46.850 159.130 ;
        RECT 48.660 159.085 48.950 159.130 ;
        RECT 50.230 159.085 50.520 159.130 ;
        RECT 51.120 159.270 51.440 159.330 ;
        RECT 69.520 159.270 69.840 159.330 ;
        RECT 70.440 159.270 70.760 159.330 ;
        RECT 51.120 159.130 70.760 159.270 ;
        RECT 51.120 159.070 51.440 159.130 ;
        RECT 69.520 159.070 69.840 159.130 ;
        RECT 70.440 159.070 70.760 159.130 ;
        RECT 33.195 158.930 33.485 158.975 ;
        RECT 34.100 158.930 34.420 158.990 ;
        RECT 33.195 158.790 34.420 158.930 ;
        RECT 33.195 158.745 33.485 158.790 ;
        RECT 34.100 158.730 34.420 158.790 ;
        RECT 54.815 158.930 55.105 158.975 ;
        RECT 59.860 158.930 60.180 158.990 ;
        RECT 54.815 158.790 60.180 158.930 ;
        RECT 54.815 158.745 55.105 158.790 ;
        RECT 59.860 158.730 60.180 158.790 ;
        RECT 60.320 158.930 60.640 158.990 ;
        RECT 71.360 158.930 71.680 158.990 ;
        RECT 60.320 158.790 71.680 158.930 ;
        RECT 72.035 158.930 72.175 159.425 ;
        RECT 72.320 159.270 72.610 159.315 ;
        RECT 74.420 159.270 74.710 159.315 ;
        RECT 75.990 159.270 76.280 159.315 ;
        RECT 72.320 159.130 76.280 159.270 ;
        RECT 72.320 159.085 72.610 159.130 ;
        RECT 74.420 159.085 74.710 159.130 ;
        RECT 75.990 159.085 76.280 159.130 ;
        RECT 76.880 158.930 77.200 158.990 ;
        RECT 72.035 158.790 77.200 158.930 ;
        RECT 60.320 158.730 60.640 158.790 ;
        RECT 71.360 158.730 71.680 158.790 ;
        RECT 76.880 158.730 77.200 158.790 ;
        RECT 78.720 158.730 79.040 158.990 ;
        RECT 11.950 158.110 90.610 158.590 ;
        RECT 39.175 157.910 39.465 157.955 ;
        RECT 40.080 157.910 40.400 157.970 ;
        RECT 39.175 157.770 40.400 157.910 ;
        RECT 39.175 157.725 39.465 157.770 ;
        RECT 40.080 157.710 40.400 157.770 ;
        RECT 47.440 157.710 47.760 157.970 ;
        RECT 52.975 157.910 53.265 157.955 ;
        RECT 53.420 157.910 53.740 157.970 ;
        RECT 52.975 157.770 53.740 157.910 ;
        RECT 52.975 157.725 53.265 157.770 ;
        RECT 53.420 157.710 53.740 157.770 ;
        RECT 59.415 157.910 59.705 157.955 ;
        RECT 61.700 157.910 62.020 157.970 ;
        RECT 59.415 157.770 62.020 157.910 ;
        RECT 59.415 157.725 59.705 157.770 ;
        RECT 61.700 157.710 62.020 157.770 ;
        RECT 70.440 157.910 70.760 157.970 ;
        RECT 72.740 157.910 73.060 157.970 ;
        RECT 70.440 157.770 73.060 157.910 ;
        RECT 70.440 157.710 70.760 157.770 ;
        RECT 72.740 157.710 73.060 157.770 ;
        RECT 51.120 157.570 51.440 157.630 ;
        RECT 44.310 157.430 51.440 157.570 ;
        RECT 24.900 157.230 25.220 157.290 ;
        RECT 32.260 157.230 32.580 157.290 ;
        RECT 33.655 157.230 33.945 157.275 ;
        RECT 24.900 157.090 26.510 157.230 ;
        RECT 24.900 157.030 25.220 157.090 ;
        RECT 25.375 156.890 25.665 156.935 ;
        RECT 25.820 156.890 26.140 156.950 ;
        RECT 26.370 156.935 26.510 157.090 ;
        RECT 32.260 157.090 33.945 157.230 ;
        RECT 32.260 157.030 32.580 157.090 ;
        RECT 33.655 157.045 33.945 157.090 ;
        RECT 39.160 157.230 39.480 157.290 ;
        RECT 44.310 157.275 44.450 157.430 ;
        RECT 51.120 157.370 51.440 157.430 ;
        RECT 55.735 157.570 56.025 157.615 ;
        RECT 56.655 157.570 56.945 157.615 ;
        RECT 60.320 157.570 60.640 157.630 ;
        RECT 66.775 157.570 67.065 157.615 ;
        RECT 55.735 157.430 56.945 157.570 ;
        RECT 55.735 157.385 56.025 157.430 ;
        RECT 56.655 157.385 56.945 157.430 ;
        RECT 57.190 157.430 60.640 157.570 ;
        RECT 39.970 157.230 40.260 157.275 ;
        RECT 39.160 157.090 40.260 157.230 ;
        RECT 39.160 157.030 39.480 157.090 ;
        RECT 39.970 157.045 40.260 157.090 ;
        RECT 42.395 157.230 42.685 157.275 ;
        RECT 44.235 157.230 44.525 157.275 ;
        RECT 57.190 157.230 57.330 157.430 ;
        RECT 60.320 157.370 60.640 157.430 ;
        RECT 63.170 157.430 67.065 157.570 ;
        RECT 42.395 157.090 44.525 157.230 ;
        RECT 42.395 157.045 42.685 157.090 ;
        RECT 44.235 157.045 44.525 157.090 ;
        RECT 49.830 157.090 57.330 157.230 ;
        RECT 58.495 157.230 58.785 157.275 ;
        RECT 62.160 157.230 62.480 157.290 ;
        RECT 58.495 157.090 62.480 157.230 ;
        RECT 25.375 156.750 26.140 156.890 ;
        RECT 25.375 156.705 25.665 156.750 ;
        RECT 25.820 156.690 26.140 156.750 ;
        RECT 26.295 156.705 26.585 156.935 ;
        RECT 32.735 156.890 33.025 156.935 ;
        RECT 33.180 156.890 33.500 156.950 ;
        RECT 32.735 156.750 33.500 156.890 ;
        RECT 32.735 156.705 33.025 156.750 ;
        RECT 33.180 156.690 33.500 156.750 ;
        RECT 46.520 156.935 46.840 156.950 ;
        RECT 46.520 156.705 46.950 156.935 ;
        RECT 46.520 156.690 46.840 156.705 ;
        RECT 41.015 156.550 41.305 156.595 ;
        RECT 45.615 156.550 45.905 156.595 ;
        RECT 48.360 156.550 48.680 156.610 ;
        RECT 41.015 156.410 48.680 156.550 ;
        RECT 41.015 156.365 41.305 156.410 ;
        RECT 45.615 156.365 45.905 156.410 ;
        RECT 48.360 156.350 48.680 156.410 ;
        RECT 22.140 156.210 22.460 156.270 ;
        RECT 25.375 156.210 25.665 156.255 ;
        RECT 22.140 156.070 25.665 156.210 ;
        RECT 22.140 156.010 22.460 156.070 ;
        RECT 25.375 156.025 25.665 156.070 ;
        RECT 30.420 156.210 30.740 156.270 ;
        RECT 31.815 156.210 32.105 156.255 ;
        RECT 30.420 156.070 32.105 156.210 ;
        RECT 30.420 156.010 30.740 156.070 ;
        RECT 31.815 156.025 32.105 156.070 ;
        RECT 40.555 156.210 40.845 156.255 ;
        RECT 41.460 156.210 41.780 156.270 ;
        RECT 46.060 156.210 46.380 156.270 ;
        RECT 49.830 156.210 49.970 157.090 ;
        RECT 58.495 157.045 58.785 157.090 ;
        RECT 62.160 157.030 62.480 157.090 ;
        RECT 63.170 156.950 63.310 157.430 ;
        RECT 66.775 157.385 67.065 157.430 ;
        RECT 71.360 157.570 71.680 157.630 ;
        RECT 73.660 157.570 73.980 157.630 ;
        RECT 71.360 157.430 73.980 157.570 ;
        RECT 71.360 157.370 71.680 157.430 ;
        RECT 73.660 157.370 73.980 157.430 ;
        RECT 77.380 157.570 77.670 157.615 ;
        RECT 79.480 157.570 79.770 157.615 ;
        RECT 81.050 157.570 81.340 157.615 ;
        RECT 77.380 157.430 81.340 157.570 ;
        RECT 77.380 157.385 77.670 157.430 ;
        RECT 79.480 157.385 79.770 157.430 ;
        RECT 81.050 157.385 81.340 157.430 ;
        RECT 64.920 157.030 65.240 157.290 ;
        RECT 67.220 157.230 67.540 157.290 ;
        RECT 69.075 157.230 69.365 157.275 ;
        RECT 76.420 157.230 76.740 157.290 ;
        RECT 67.220 157.090 69.365 157.230 ;
        RECT 67.220 157.030 67.540 157.090 ;
        RECT 69.075 157.045 69.365 157.090 ;
        RECT 71.450 157.090 76.740 157.230 ;
        RECT 52.960 156.890 53.280 156.950 ;
        RECT 53.600 156.890 53.890 156.935 ;
        RECT 52.960 156.750 53.890 156.890 ;
        RECT 52.960 156.690 53.280 156.750 ;
        RECT 53.600 156.705 53.890 156.750 ;
        RECT 56.180 156.690 56.500 156.950 ;
        RECT 57.560 156.690 57.880 156.950 ;
        RECT 59.860 156.690 60.180 156.950 ;
        RECT 61.240 156.690 61.560 156.950 ;
        RECT 61.715 156.705 62.005 156.935 ;
        RECT 62.635 156.890 62.925 156.935 ;
        RECT 62.250 156.750 62.925 156.890 ;
        RECT 61.790 156.550 61.930 156.705 ;
        RECT 54.660 156.410 61.930 156.550 ;
        RECT 40.555 156.070 49.970 156.210 ;
        RECT 52.960 156.210 53.280 156.270 ;
        RECT 53.880 156.210 54.200 156.270 ;
        RECT 54.660 156.210 54.800 156.410 ;
        RECT 52.960 156.070 54.800 156.210 ;
        RECT 40.555 156.025 40.845 156.070 ;
        RECT 41.460 156.010 41.780 156.070 ;
        RECT 46.060 156.010 46.380 156.070 ;
        RECT 52.960 156.010 53.280 156.070 ;
        RECT 53.880 156.010 54.200 156.070 ;
        RECT 60.320 156.010 60.640 156.270 ;
        RECT 62.250 156.210 62.390 156.750 ;
        RECT 62.635 156.705 62.925 156.750 ;
        RECT 63.080 156.690 63.400 156.950 ;
        RECT 65.380 156.690 65.700 156.950 ;
        RECT 68.600 156.690 68.920 156.950 ;
        RECT 70.440 156.690 70.760 156.950 ;
        RECT 71.450 156.935 71.590 157.090 ;
        RECT 76.420 157.030 76.740 157.090 ;
        RECT 76.880 157.030 77.200 157.290 ;
        RECT 77.775 157.230 78.065 157.275 ;
        RECT 78.965 157.230 79.255 157.275 ;
        RECT 81.485 157.230 81.775 157.275 ;
        RECT 77.775 157.090 81.775 157.230 ;
        RECT 77.775 157.045 78.065 157.090 ;
        RECT 78.965 157.045 79.255 157.090 ;
        RECT 81.485 157.045 81.775 157.090 ;
        RECT 71.375 156.705 71.665 156.935 ;
        RECT 71.835 156.890 72.125 156.935 ;
        RECT 72.740 156.890 73.060 156.950 ;
        RECT 71.835 156.750 73.060 156.890 ;
        RECT 71.835 156.705 72.125 156.750 ;
        RECT 72.740 156.690 73.060 156.750 ;
        RECT 73.660 156.690 73.980 156.950 ;
        RECT 70.915 156.550 71.205 156.595 ;
        RECT 74.260 156.550 74.550 156.595 ;
        RECT 78.120 156.550 78.410 156.595 ;
        RECT 70.915 156.410 74.550 156.550 ;
        RECT 70.915 156.365 71.205 156.410 ;
        RECT 74.260 156.365 74.550 156.410 ;
        RECT 75.130 156.410 78.410 156.550 ;
        RECT 62.620 156.210 62.940 156.270 ;
        RECT 63.555 156.210 63.845 156.255 ;
        RECT 62.250 156.070 63.845 156.210 ;
        RECT 62.620 156.010 62.940 156.070 ;
        RECT 63.555 156.025 63.845 156.070 ;
        RECT 71.820 156.210 72.140 156.270 ;
        RECT 75.130 156.255 75.270 156.410 ;
        RECT 78.120 156.365 78.410 156.410 ;
        RECT 73.215 156.210 73.505 156.255 ;
        RECT 71.820 156.070 73.505 156.210 ;
        RECT 71.820 156.010 72.140 156.070 ;
        RECT 73.215 156.025 73.505 156.070 ;
        RECT 75.055 156.025 75.345 156.255 ;
        RECT 76.880 156.210 77.200 156.270 ;
        RECT 83.795 156.210 84.085 156.255 ;
        RECT 76.880 156.070 84.085 156.210 ;
        RECT 76.880 156.010 77.200 156.070 ;
        RECT 83.795 156.025 84.085 156.070 ;
        RECT 100.010 156.200 100.880 159.470 ;
        RECT 104.530 159.010 109.780 159.020 ;
        RECT 104.530 158.900 116.840 159.010 ;
        RECT 101.560 158.840 116.840 158.900 ;
        RECT 101.560 158.830 116.875 158.840 ;
        RECT 101.500 158.700 116.875 158.830 ;
        RECT 101.500 158.690 106.660 158.700 ;
        RECT 101.500 158.600 105.500 158.690 ;
        RECT 108.875 158.610 116.875 158.700 ;
        RECT 108.960 158.600 116.850 158.610 ;
        RECT 101.110 158.240 101.340 158.550 ;
        RECT 101.560 158.240 105.460 158.600 ;
        RECT 105.660 158.240 105.890 158.550 ;
        RECT 101.110 156.900 105.890 158.240 ;
        RECT 101.110 156.590 101.340 156.900 ;
        RECT 105.660 156.590 105.890 156.900 ;
        RECT 108.440 158.020 108.670 158.560 ;
        RECT 109.480 158.020 110.490 158.050 ;
        RECT 117.080 158.020 117.310 158.560 ;
        RECT 108.440 157.120 117.310 158.020 ;
        RECT 108.440 156.600 108.670 157.120 ;
        RECT 109.480 157.050 110.490 157.120 ;
        RECT 117.080 156.600 117.310 157.120 ;
        RECT 101.500 156.310 105.500 156.540 ;
        RECT 108.875 156.320 116.875 156.550 ;
        RECT 100.010 156.160 101.180 156.200 ;
        RECT 100.010 156.080 101.420 156.160 ;
        RECT 101.790 156.090 105.450 156.310 ;
        RECT 101.790 156.080 103.230 156.090 ;
        RECT 100.010 156.040 103.230 156.080 ;
        RECT 100.010 155.950 102.740 156.040 ;
        RECT 108.940 156.030 116.830 156.320 ;
        RECT 100.010 155.890 102.070 155.950 ;
        RECT 11.950 155.390 90.610 155.870 ;
        RECT 100.010 155.840 101.820 155.890 ;
        RECT 25.820 155.190 26.140 155.250 ;
        RECT 24.530 155.050 26.140 155.190 ;
        RECT 21.220 154.650 21.540 154.910 ;
        RECT 24.530 154.895 24.670 155.050 ;
        RECT 25.820 154.990 26.140 155.050 ;
        RECT 32.735 155.190 33.025 155.235 ;
        RECT 33.180 155.190 33.500 155.250 ;
        RECT 34.100 155.190 34.420 155.250 ;
        RECT 32.735 155.050 34.420 155.190 ;
        RECT 32.735 155.005 33.025 155.050 ;
        RECT 33.180 154.990 33.500 155.050 ;
        RECT 34.100 154.990 34.420 155.050 ;
        RECT 48.820 155.190 49.140 155.250 ;
        RECT 56.180 155.190 56.500 155.250 ;
        RECT 60.795 155.190 61.085 155.235 ;
        RECT 70.440 155.190 70.760 155.250 ;
        RECT 73.200 155.190 73.520 155.250 ;
        RECT 48.820 155.050 51.810 155.190 ;
        RECT 48.820 154.990 49.140 155.050 ;
        RECT 22.315 154.850 22.605 154.895 ;
        RECT 23.535 154.850 23.825 154.895 ;
        RECT 22.315 154.710 23.825 154.850 ;
        RECT 22.315 154.665 22.605 154.710 ;
        RECT 23.535 154.665 23.825 154.710 ;
        RECT 24.455 154.665 24.745 154.895 ;
        RECT 24.900 154.850 25.220 154.910 ;
        RECT 25.375 154.850 25.665 154.895 ;
        RECT 29.960 154.850 30.280 154.910 ;
        RECT 24.900 154.710 25.665 154.850 ;
        RECT 24.900 154.650 25.220 154.710 ;
        RECT 25.375 154.665 25.665 154.710 ;
        RECT 25.910 154.710 30.280 154.850 ;
        RECT 25.910 154.555 26.050 154.710 ;
        RECT 29.960 154.650 30.280 154.710 ;
        RECT 38.240 154.850 38.560 154.910 ;
        RECT 38.240 154.710 49.970 154.850 ;
        RECT 38.240 154.650 38.560 154.710 ;
        RECT 25.835 154.325 26.125 154.555 ;
        RECT 27.115 154.510 27.405 154.555 ;
        RECT 26.370 154.370 27.405 154.510 ;
        RECT 26.370 154.170 26.510 154.370 ;
        RECT 27.115 154.325 27.405 154.370 ;
        RECT 47.900 154.510 48.220 154.570 ;
        RECT 49.830 154.555 49.970 154.710 ;
        RECT 51.670 154.555 51.810 155.050 ;
        RECT 56.180 155.050 61.085 155.190 ;
        RECT 56.180 154.990 56.500 155.050 ;
        RECT 60.795 155.005 61.085 155.050 ;
        RECT 69.150 155.050 70.210 155.190 ;
        RECT 69.150 154.895 69.290 155.050 ;
        RECT 69.075 154.665 69.365 154.895 ;
        RECT 69.520 154.650 69.840 154.910 ;
        RECT 70.070 154.850 70.210 155.050 ;
        RECT 70.440 155.050 73.520 155.190 ;
        RECT 70.440 154.990 70.760 155.050 ;
        RECT 73.200 154.990 73.520 155.050 ;
        RECT 72.280 154.850 72.600 154.910 ;
        RECT 73.975 154.850 74.265 154.895 ;
        RECT 70.070 154.710 74.265 154.850 ;
        RECT 72.280 154.650 72.600 154.710 ;
        RECT 73.975 154.665 74.265 154.710 ;
        RECT 75.055 154.850 75.345 154.895 ;
        RECT 76.880 154.850 77.200 154.910 ;
        RECT 75.055 154.710 77.200 154.850 ;
        RECT 75.055 154.665 75.345 154.710 ;
        RECT 48.835 154.510 49.125 154.555 ;
        RECT 47.900 154.370 49.125 154.510 ;
        RECT 47.900 154.310 48.220 154.370 ;
        RECT 48.835 154.325 49.125 154.370 ;
        RECT 49.755 154.510 50.045 154.555 ;
        RECT 51.135 154.510 51.425 154.555 ;
        RECT 49.755 154.370 51.425 154.510 ;
        RECT 49.755 154.325 50.045 154.370 ;
        RECT 51.135 154.325 51.425 154.370 ;
        RECT 51.595 154.325 51.885 154.555 ;
        RECT 52.040 154.510 52.360 154.570 ;
        RECT 52.515 154.510 52.805 154.555 ;
        RECT 52.040 154.370 52.805 154.510 ;
        RECT 23.150 154.030 26.510 154.170 ;
        RECT 26.715 154.170 27.005 154.215 ;
        RECT 27.905 154.170 28.195 154.215 ;
        RECT 30.425 154.170 30.715 154.215 ;
        RECT 26.715 154.030 30.715 154.170 ;
        RECT 48.910 154.170 49.050 154.325 ;
        RECT 51.670 154.170 51.810 154.325 ;
        RECT 52.040 154.310 52.360 154.370 ;
        RECT 52.515 154.325 52.805 154.370 ;
        RECT 53.420 154.310 53.740 154.570 ;
        RECT 54.815 154.510 55.105 154.555 ;
        RECT 55.720 154.510 56.040 154.570 ;
        RECT 54.815 154.370 56.040 154.510 ;
        RECT 54.815 154.325 55.105 154.370 ;
        RECT 55.720 154.310 56.040 154.370 ;
        RECT 61.700 154.310 62.020 154.570 ;
        RECT 62.635 154.510 62.925 154.555 ;
        RECT 63.080 154.510 63.400 154.570 ;
        RECT 62.635 154.370 63.400 154.510 ;
        RECT 62.635 154.325 62.925 154.370 ;
        RECT 63.080 154.310 63.400 154.370 ;
        RECT 65.380 154.510 65.700 154.570 ;
        RECT 65.855 154.510 66.145 154.555 ;
        RECT 65.380 154.370 66.145 154.510 ;
        RECT 65.380 154.310 65.700 154.370 ;
        RECT 65.855 154.325 66.145 154.370 ;
        RECT 66.775 154.510 67.065 154.555 ;
        RECT 67.220 154.510 67.540 154.570 ;
        RECT 66.775 154.370 67.540 154.510 ;
        RECT 66.775 154.325 67.065 154.370 ;
        RECT 53.895 154.170 54.185 154.215 ;
        RECT 48.910 154.030 51.350 154.170 ;
        RECT 51.670 154.030 54.185 154.170 ;
        RECT 65.930 154.170 66.070 154.325 ;
        RECT 67.220 154.310 67.540 154.370 ;
        RECT 68.600 154.510 68.920 154.570 ;
        RECT 69.995 154.510 70.285 154.555 ;
        RECT 75.130 154.510 75.270 154.665 ;
        RECT 76.880 154.650 77.200 154.710 ;
        RECT 68.600 154.370 75.270 154.510 ;
        RECT 68.600 154.310 68.920 154.370 ;
        RECT 69.995 154.325 70.285 154.370 ;
        RECT 75.515 154.325 75.805 154.555 ;
        RECT 75.975 154.510 76.265 154.555 ;
        RECT 78.720 154.510 79.040 154.570 ;
        RECT 75.975 154.370 79.040 154.510 ;
        RECT 75.975 154.325 76.265 154.370 ;
        RECT 72.280 154.170 72.600 154.230 ;
        RECT 75.040 154.170 75.360 154.230 ;
        RECT 75.590 154.170 75.730 154.325 ;
        RECT 65.930 154.030 71.130 154.170 ;
        RECT 23.150 153.875 23.290 154.030 ;
        RECT 26.715 153.985 27.005 154.030 ;
        RECT 27.905 153.985 28.195 154.030 ;
        RECT 30.425 153.985 30.715 154.030 ;
        RECT 23.075 153.645 23.365 153.875 ;
        RECT 26.320 153.830 26.610 153.875 ;
        RECT 28.420 153.830 28.710 153.875 ;
        RECT 29.990 153.830 30.280 153.875 ;
        RECT 26.320 153.690 30.280 153.830 ;
        RECT 26.320 153.645 26.610 153.690 ;
        RECT 28.420 153.645 28.710 153.690 ;
        RECT 29.990 153.645 30.280 153.690 ;
        RECT 34.560 153.830 34.880 153.890 ;
        RECT 37.780 153.830 38.100 153.890 ;
        RECT 51.210 153.830 51.350 154.030 ;
        RECT 53.895 153.985 54.185 154.030 ;
        RECT 52.055 153.830 52.345 153.875 ;
        RECT 52.960 153.830 53.280 153.890 ;
        RECT 54.340 153.830 54.660 153.890 ;
        RECT 68.600 153.830 68.920 153.890 ;
        RECT 70.990 153.875 71.130 154.030 ;
        RECT 72.280 154.030 75.730 154.170 ;
        RECT 72.280 153.970 72.600 154.030 ;
        RECT 75.040 153.970 75.360 154.030 ;
        RECT 34.560 153.690 50.890 153.830 ;
        RECT 51.210 153.690 53.280 153.830 ;
        RECT 34.560 153.630 34.880 153.690 ;
        RECT 37.780 153.630 38.100 153.690 ;
        RECT 22.140 153.290 22.460 153.550 ;
        RECT 48.820 153.290 49.140 153.550 ;
        RECT 50.200 153.290 50.520 153.550 ;
        RECT 50.750 153.490 50.890 153.690 ;
        RECT 52.055 153.645 52.345 153.690 ;
        RECT 52.960 153.630 53.280 153.690 ;
        RECT 53.510 153.690 54.660 153.830 ;
        RECT 53.510 153.535 53.650 153.690 ;
        RECT 54.340 153.630 54.660 153.690 ;
        RECT 66.850 153.690 68.920 153.830 ;
        RECT 53.435 153.490 53.725 153.535 ;
        RECT 50.750 153.350 53.725 153.490 ;
        RECT 53.435 153.305 53.725 153.350 ;
        RECT 53.880 153.490 54.200 153.550 ;
        RECT 55.735 153.490 56.025 153.535 ;
        RECT 53.880 153.350 56.025 153.490 ;
        RECT 53.880 153.290 54.200 153.350 ;
        RECT 55.735 153.305 56.025 153.350 ;
        RECT 62.620 153.290 62.940 153.550 ;
        RECT 63.540 153.490 63.860 153.550 ;
        RECT 66.850 153.535 66.990 153.690 ;
        RECT 68.600 153.630 68.920 153.690 ;
        RECT 70.915 153.830 71.205 153.875 ;
        RECT 74.580 153.830 74.900 153.890 ;
        RECT 70.915 153.690 74.900 153.830 ;
        RECT 70.915 153.645 71.205 153.690 ;
        RECT 74.580 153.630 74.900 153.690 ;
        RECT 64.935 153.490 65.225 153.535 ;
        RECT 63.540 153.350 65.225 153.490 ;
        RECT 63.540 153.290 63.860 153.350 ;
        RECT 64.935 153.305 65.225 153.350 ;
        RECT 66.775 153.305 67.065 153.535 ;
        RECT 68.140 153.290 68.460 153.550 ;
        RECT 69.520 153.490 69.840 153.550 ;
        RECT 74.135 153.490 74.425 153.535 ;
        RECT 76.050 153.490 76.190 154.325 ;
        RECT 78.720 154.310 79.040 154.370 ;
        RECT 76.420 153.830 76.740 153.890 ;
        RECT 76.895 153.830 77.185 153.875 ;
        RECT 76.420 153.690 77.185 153.830 ;
        RECT 76.420 153.630 76.740 153.690 ;
        RECT 76.895 153.645 77.185 153.690 ;
        RECT 69.520 153.350 76.190 153.490 ;
        RECT 69.520 153.290 69.840 153.350 ;
        RECT 74.135 153.305 74.425 153.350 ;
        RECT 11.950 152.670 90.610 153.150 ;
        RECT 48.820 152.270 49.140 152.530 ;
        RECT 58.480 152.470 58.800 152.530 ;
        RECT 62.620 152.470 62.940 152.530 ;
        RECT 63.095 152.470 63.385 152.515 ;
        RECT 58.480 152.330 62.390 152.470 ;
        RECT 58.480 152.270 58.800 152.330 ;
        RECT 18.040 152.130 18.330 152.175 ;
        RECT 20.140 152.130 20.430 152.175 ;
        RECT 21.710 152.130 22.000 152.175 ;
        RECT 18.040 151.990 22.000 152.130 ;
        RECT 18.040 151.945 18.330 151.990 ;
        RECT 20.140 151.945 20.430 151.990 ;
        RECT 21.710 151.945 22.000 151.990 ;
        RECT 35.955 152.130 36.245 152.175 ;
        RECT 53.420 152.130 53.740 152.190 ;
        RECT 62.250 152.130 62.390 152.330 ;
        RECT 62.620 152.330 63.385 152.470 ;
        RECT 62.620 152.270 62.940 152.330 ;
        RECT 63.095 152.285 63.385 152.330 ;
        RECT 100.010 152.500 100.880 155.840 ;
        RECT 108.930 155.540 116.850 155.550 ;
        RECT 105.160 155.530 116.850 155.540 ;
        RECT 101.540 155.410 116.850 155.530 ;
        RECT 101.540 155.400 116.875 155.410 ;
        RECT 101.500 155.280 116.875 155.400 ;
        RECT 101.500 155.170 105.500 155.280 ;
        RECT 101.110 154.830 101.340 155.120 ;
        RECT 101.560 154.830 105.450 155.170 ;
        RECT 105.660 154.830 105.890 155.120 ;
        RECT 101.110 153.460 105.890 154.830 ;
        RECT 101.110 153.160 101.340 153.460 ;
        RECT 105.660 153.160 105.890 153.460 ;
        RECT 101.500 152.880 105.500 153.110 ;
        RECT 101.750 152.650 105.320 152.880 ;
        RECT 101.750 152.500 105.440 152.650 ;
        RECT 100.010 152.220 105.440 152.500 ;
        RECT 106.690 152.330 107.310 155.280 ;
        RECT 108.875 155.180 116.875 155.280 ;
        RECT 108.930 155.170 116.850 155.180 ;
        RECT 108.440 154.470 108.670 155.130 ;
        RECT 109.450 154.470 110.450 154.560 ;
        RECT 117.080 154.470 117.310 155.130 ;
        RECT 108.440 153.650 117.310 154.470 ;
        RECT 108.440 153.170 108.670 153.650 ;
        RECT 109.450 153.560 110.450 153.650 ;
        RECT 117.080 153.170 117.310 153.650 ;
        RECT 108.875 152.890 116.875 153.120 ;
        RECT 70.900 152.130 71.220 152.190 ;
        RECT 72.280 152.130 72.600 152.190 ;
        RECT 35.955 151.990 43.990 152.130 ;
        RECT 35.955 151.945 36.245 151.990 ;
        RECT 18.435 151.790 18.725 151.835 ;
        RECT 19.625 151.790 19.915 151.835 ;
        RECT 22.145 151.790 22.435 151.835 ;
        RECT 18.435 151.650 22.435 151.790 ;
        RECT 18.435 151.605 18.725 151.650 ;
        RECT 19.625 151.605 19.915 151.650 ;
        RECT 22.145 151.605 22.435 151.650 ;
        RECT 24.900 151.790 25.220 151.850 ;
        RECT 29.960 151.790 30.280 151.850 ;
        RECT 35.480 151.790 35.800 151.850 ;
        RECT 24.900 151.650 27.890 151.790 ;
        RECT 24.900 151.590 25.220 151.650 ;
        RECT 17.540 151.250 17.860 151.510 ;
        RECT 27.750 151.495 27.890 151.650 ;
        RECT 29.960 151.650 31.575 151.790 ;
        RECT 29.960 151.590 30.280 151.650 ;
        RECT 31.435 151.495 31.575 151.650 ;
        RECT 32.350 151.650 35.800 151.790 ;
        RECT 32.350 151.495 32.490 151.650 ;
        RECT 35.480 151.590 35.800 151.650 ;
        RECT 26.295 151.265 26.585 151.495 ;
        RECT 27.675 151.265 27.965 151.495 ;
        RECT 30.895 151.265 31.185 151.495 ;
        RECT 31.360 151.265 31.650 151.495 ;
        RECT 32.275 151.265 32.565 151.495 ;
        RECT 33.425 151.450 33.715 151.495 ;
        RECT 36.030 151.450 36.170 151.945 ;
        RECT 40.095 151.605 40.385 151.835 ;
        RECT 33.425 151.310 36.170 151.450 ;
        RECT 33.425 151.265 33.715 151.310 ;
        RECT 18.920 151.155 19.240 151.170 ;
        RECT 18.890 150.925 19.240 151.155 ;
        RECT 26.370 151.110 26.510 151.265 ;
        RECT 30.970 151.110 31.110 151.265 ;
        RECT 37.320 151.250 37.640 151.510 ;
        RECT 37.780 151.250 38.100 151.510 ;
        RECT 38.240 151.450 38.560 151.510 ;
        RECT 39.635 151.450 39.925 151.495 ;
        RECT 38.240 151.310 39.925 151.450 ;
        RECT 40.170 151.450 40.310 151.605 ;
        RECT 41.460 151.590 41.780 151.850 ;
        RECT 43.850 151.835 43.990 151.990 ;
        RECT 48.910 151.990 53.740 152.130 ;
        RECT 48.910 151.835 49.050 151.990 ;
        RECT 53.420 151.930 53.740 151.990 ;
        RECT 58.110 151.990 61.930 152.130 ;
        RECT 62.250 151.990 72.600 152.130 ;
        RECT 43.775 151.605 44.065 151.835 ;
        RECT 48.835 151.605 49.125 151.835 ;
        RECT 50.200 151.790 50.520 151.850 ;
        RECT 55.275 151.790 55.565 151.835 ;
        RECT 50.200 151.650 55.565 151.790 ;
        RECT 50.200 151.590 50.520 151.650 ;
        RECT 55.275 151.605 55.565 151.650 ;
        RECT 40.540 151.450 40.860 151.510 ;
        RECT 43.300 151.450 43.620 151.510 ;
        RECT 40.170 151.310 43.620 151.450 ;
        RECT 38.240 151.250 38.560 151.310 ;
        RECT 39.635 151.265 39.925 151.310 ;
        RECT 40.540 151.250 40.860 151.310 ;
        RECT 43.300 151.250 43.620 151.310 ;
        RECT 44.235 151.450 44.525 151.495 ;
        RECT 44.235 151.310 49.050 151.450 ;
        RECT 44.235 151.265 44.525 151.310 ;
        RECT 18.920 150.910 19.240 150.925 ;
        RECT 24.530 150.970 31.110 151.110 ;
        RECT 32.735 151.110 33.025 151.155 ;
        RECT 32.735 150.970 33.410 151.110 ;
        RECT 24.530 150.830 24.670 150.970 ;
        RECT 32.735 150.925 33.025 150.970 ;
        RECT 33.270 150.830 33.410 150.970 ;
        RECT 47.915 150.925 48.205 151.155 ;
        RECT 48.910 151.110 49.050 151.310 ;
        RECT 49.280 151.250 49.600 151.510 ;
        RECT 51.595 151.450 51.885 151.495 ;
        RECT 49.830 151.310 51.885 151.450 ;
        RECT 49.830 151.170 49.970 151.310 ;
        RECT 51.595 151.265 51.885 151.310 ;
        RECT 53.880 151.250 54.200 151.510 ;
        RECT 57.115 151.450 57.405 151.495 ;
        RECT 58.110 151.450 58.250 151.990 ;
        RECT 58.480 151.590 58.800 151.850 ;
        RECT 59.860 151.495 60.180 151.510 ;
        RECT 57.115 151.310 58.250 151.450 ;
        RECT 57.115 151.265 57.405 151.310 ;
        RECT 58.955 151.265 59.245 151.495 ;
        RECT 59.695 151.265 60.180 151.495 ;
        RECT 49.740 151.110 50.060 151.170 ;
        RECT 57.560 151.110 57.880 151.170 ;
        RECT 59.030 151.110 59.170 151.265 ;
        RECT 59.860 151.250 60.180 151.265 ;
        RECT 60.320 151.250 60.640 151.510 ;
        RECT 61.280 151.265 61.570 151.495 ;
        RECT 61.790 151.450 61.930 151.990 ;
        RECT 70.900 151.930 71.220 151.990 ;
        RECT 72.280 151.930 72.600 151.990 ;
        RECT 74.135 151.790 74.425 151.835 ;
        RECT 73.290 151.650 74.425 151.790 ;
        RECT 61.790 151.310 62.390 151.450 ;
        RECT 48.910 150.970 50.060 151.110 ;
        RECT 24.440 150.570 24.760 150.830 ;
        RECT 25.360 150.570 25.680 150.830 ;
        RECT 25.820 150.770 26.140 150.830 ;
        RECT 27.215 150.770 27.505 150.815 ;
        RECT 33.180 150.770 33.500 150.830 ;
        RECT 25.820 150.630 33.500 150.770 ;
        RECT 25.820 150.570 26.140 150.630 ;
        RECT 27.215 150.585 27.505 150.630 ;
        RECT 33.180 150.570 33.500 150.630 ;
        RECT 34.100 150.570 34.420 150.830 ;
        RECT 46.075 150.770 46.365 150.815 ;
        RECT 47.990 150.770 48.130 150.925 ;
        RECT 49.740 150.910 50.060 150.970 ;
        RECT 50.290 150.970 59.170 151.110 ;
        RECT 50.290 150.815 50.430 150.970 ;
        RECT 57.560 150.910 57.880 150.970 ;
        RECT 60.780 150.910 61.100 151.170 ;
        RECT 46.075 150.630 48.130 150.770 ;
        RECT 46.075 150.585 46.365 150.630 ;
        RECT 50.215 150.585 50.505 150.815 ;
        RECT 52.060 150.770 52.350 150.815 ;
        RECT 58.500 150.770 58.790 150.815 ;
        RECT 52.060 150.630 58.790 150.770 ;
        RECT 52.060 150.585 52.350 150.630 ;
        RECT 58.500 150.585 58.790 150.630 ;
        RECT 59.400 150.770 59.720 150.830 ;
        RECT 61.330 150.770 61.470 151.265 ;
        RECT 62.250 150.815 62.390 151.310 ;
        RECT 62.635 151.265 62.925 151.495 ;
        RECT 63.555 151.450 63.845 151.495 ;
        RECT 66.300 151.450 66.620 151.510 ;
        RECT 63.555 151.310 66.620 151.450 ;
        RECT 63.555 151.265 63.845 151.310 ;
        RECT 62.710 151.110 62.850 151.265 ;
        RECT 66.300 151.250 66.620 151.310 ;
        RECT 68.140 151.450 68.460 151.510 ;
        RECT 73.290 151.495 73.430 151.650 ;
        RECT 74.135 151.605 74.425 151.650 ;
        RECT 100.010 151.760 105.450 152.220 ;
        RECT 72.295 151.450 72.585 151.495 ;
        RECT 68.140 151.310 72.585 151.450 ;
        RECT 68.140 151.250 68.460 151.310 ;
        RECT 72.295 151.265 72.585 151.310 ;
        RECT 73.215 151.265 73.505 151.495 ;
        RECT 73.660 151.250 73.980 151.510 ;
        RECT 74.580 151.450 74.900 151.510 ;
        RECT 80.560 151.450 80.880 151.510 ;
        RECT 74.580 151.310 80.880 151.450 ;
        RECT 74.580 151.250 74.900 151.310 ;
        RECT 80.560 151.250 80.880 151.310 ;
        RECT 64.460 151.110 64.780 151.170 ;
        RECT 67.220 151.110 67.540 151.170 ;
        RECT 62.710 150.970 67.540 151.110 ;
        RECT 64.460 150.910 64.780 150.970 ;
        RECT 67.220 150.910 67.540 150.970 ;
        RECT 59.400 150.630 61.470 150.770 ;
        RECT 59.400 150.570 59.720 150.630 ;
        RECT 62.175 150.585 62.465 150.815 ;
        RECT 70.900 150.770 71.220 150.830 ;
        RECT 72.755 150.770 73.045 150.815 ;
        RECT 70.900 150.630 73.045 150.770 ;
        RECT 70.900 150.570 71.220 150.630 ;
        RECT 72.755 150.585 73.045 150.630 ;
        RECT 11.950 149.950 90.610 150.430 ;
        RECT 100.010 150.410 102.050 151.760 ;
        RECT 103.800 151.750 105.450 151.760 ;
        RECT 102.490 150.480 103.490 151.200 ;
        RECT 103.800 150.940 104.110 151.750 ;
        RECT 104.570 151.470 105.450 151.750 ;
        RECT 105.690 151.930 107.310 152.330 ;
        RECT 108.960 151.980 116.830 152.890 ;
        RECT 104.510 151.240 105.510 151.470 ;
        RECT 105.690 151.280 106.040 151.930 ;
        RECT 106.690 151.920 107.310 151.930 ;
        RECT 108.875 151.750 116.875 151.980 ;
        RECT 108.960 151.740 116.830 151.750 ;
        RECT 104.570 151.030 105.450 151.050 ;
        RECT 103.840 150.650 104.110 150.940 ;
        RECT 104.510 150.800 105.510 151.030 ;
        RECT 105.670 150.990 106.040 151.280 ;
        RECT 105.700 150.930 106.040 150.990 ;
        RECT 106.800 151.600 107.560 151.650 ;
        RECT 108.440 151.600 108.670 151.700 ;
        RECT 106.800 151.390 108.670 151.600 ;
        RECT 117.080 151.390 117.310 151.700 ;
        RECT 106.800 150.970 109.340 151.390 ;
        RECT 116.710 150.970 117.310 151.390 ;
        RECT 104.570 150.650 105.450 150.800 ;
        RECT 104.580 150.480 105.310 150.650 ;
        RECT 18.920 149.550 19.240 149.810 ;
        RECT 19.855 149.750 20.145 149.795 ;
        RECT 21.220 149.750 21.540 149.810 ;
        RECT 19.855 149.610 21.540 149.750 ;
        RECT 19.855 149.565 20.145 149.610 ;
        RECT 21.220 149.550 21.540 149.610 ;
        RECT 23.455 149.750 23.745 149.795 ;
        RECT 24.900 149.750 25.220 149.810 ;
        RECT 23.455 149.610 25.220 149.750 ;
        RECT 23.455 149.565 23.745 149.610 ;
        RECT 24.900 149.550 25.220 149.610 ;
        RECT 29.960 149.750 30.280 149.810 ;
        RECT 38.240 149.750 38.560 149.810 ;
        RECT 48.375 149.750 48.665 149.795 ;
        RECT 29.960 149.610 38.010 149.750 ;
        RECT 29.960 149.550 30.280 149.610 ;
        RECT 24.440 149.210 24.760 149.470 ;
        RECT 34.100 149.410 34.420 149.470 ;
        RECT 31.890 149.270 34.420 149.410 ;
        RECT 37.870 149.410 38.010 149.610 ;
        RECT 38.240 149.610 48.665 149.750 ;
        RECT 38.240 149.550 38.560 149.610 ;
        RECT 48.375 149.565 48.665 149.610 ;
        RECT 50.215 149.750 50.505 149.795 ;
        RECT 53.420 149.750 53.740 149.810 ;
        RECT 50.215 149.610 53.740 149.750 ;
        RECT 50.215 149.565 50.505 149.610 ;
        RECT 53.420 149.550 53.740 149.610 ;
        RECT 59.400 149.550 59.720 149.810 ;
        RECT 59.860 149.550 60.180 149.810 ;
        RECT 71.360 149.750 71.680 149.810 ;
        RECT 71.835 149.750 72.125 149.795 ;
        RECT 71.360 149.610 72.125 149.750 ;
        RECT 71.360 149.550 71.680 149.610 ;
        RECT 71.835 149.565 72.125 149.610 ;
        RECT 73.215 149.565 73.505 149.795 ;
        RECT 63.540 149.410 63.860 149.470 ;
        RECT 37.870 149.270 47.670 149.410 ;
        RECT 30.420 148.870 30.740 149.130 ;
        RECT 30.880 149.070 31.200 149.130 ;
        RECT 31.890 149.115 32.030 149.270 ;
        RECT 34.100 149.210 34.420 149.270 ;
        RECT 31.355 149.070 31.645 149.115 ;
        RECT 30.880 148.930 31.645 149.070 ;
        RECT 30.880 148.870 31.200 148.930 ;
        RECT 31.355 148.885 31.645 148.930 ;
        RECT 31.815 148.885 32.105 149.115 ;
        RECT 33.180 148.870 33.500 149.130 ;
        RECT 42.380 149.070 42.700 149.130 ;
        RECT 43.820 149.070 44.110 149.115 ;
        RECT 42.380 148.930 44.110 149.070 ;
        RECT 47.530 149.070 47.670 149.270 ;
        RECT 62.250 149.270 63.860 149.410 ;
        RECT 47.900 149.070 48.220 149.130 ;
        RECT 47.530 148.930 48.220 149.070 ;
        RECT 42.380 148.870 42.700 148.930 ;
        RECT 43.820 148.885 44.110 148.930 ;
        RECT 47.900 148.870 48.220 148.930 ;
        RECT 48.820 149.070 49.140 149.130 ;
        RECT 49.295 149.070 49.585 149.115 ;
        RECT 48.820 148.930 49.585 149.070 ;
        RECT 48.820 148.870 49.140 148.930 ;
        RECT 49.295 148.885 49.585 148.930 ;
        RECT 57.560 148.870 57.880 149.130 ;
        RECT 58.495 149.070 58.785 149.115 ;
        RECT 59.400 149.070 59.720 149.130 ;
        RECT 62.250 149.115 62.390 149.270 ;
        RECT 63.540 149.210 63.860 149.270 ;
        RECT 64.015 149.225 64.305 149.455 ;
        RECT 64.920 149.410 65.240 149.470 ;
        RECT 67.695 149.410 67.985 149.455 ;
        RECT 69.980 149.410 70.300 149.470 ;
        RECT 64.920 149.270 66.070 149.410 ;
        RECT 61.255 149.070 61.545 149.115 ;
        RECT 58.495 148.930 61.545 149.070 ;
        RECT 58.495 148.885 58.785 148.930 ;
        RECT 59.400 148.870 59.720 148.930 ;
        RECT 61.255 148.885 61.545 148.930 ;
        RECT 61.715 148.885 62.005 149.115 ;
        RECT 62.175 148.885 62.465 149.115 ;
        RECT 63.095 149.070 63.385 149.115 ;
        RECT 64.090 149.070 64.230 149.225 ;
        RECT 64.920 149.210 65.240 149.270 ;
        RECT 63.095 148.930 64.230 149.070 ;
        RECT 63.095 148.885 63.385 148.930 ;
        RECT 32.370 148.730 32.660 148.775 ;
        RECT 33.640 148.730 33.960 148.790 ;
        RECT 32.370 148.590 33.960 148.730 ;
        RECT 32.370 148.545 32.660 148.590 ;
        RECT 33.640 148.530 33.960 148.590 ;
        RECT 40.565 148.730 40.855 148.775 ;
        RECT 43.085 148.730 43.375 148.775 ;
        RECT 44.275 148.730 44.565 148.775 ;
        RECT 40.565 148.590 44.565 148.730 ;
        RECT 40.565 148.545 40.855 148.590 ;
        RECT 43.085 148.545 43.375 148.590 ;
        RECT 44.275 148.545 44.565 148.590 ;
        RECT 45.140 148.530 45.460 148.790 ;
        RECT 57.650 148.730 57.790 148.870 ;
        RECT 61.790 148.730 61.930 148.885 ;
        RECT 65.380 148.870 65.700 149.130 ;
        RECT 65.930 149.115 66.070 149.270 ;
        RECT 66.390 149.270 67.985 149.410 ;
        RECT 66.390 149.130 66.530 149.270 ;
        RECT 67.695 149.225 67.985 149.270 ;
        RECT 69.150 149.270 70.300 149.410 ;
        RECT 73.290 149.410 73.430 149.565 ;
        RECT 80.560 149.550 80.880 149.810 ;
        RECT 74.900 149.410 75.190 149.455 ;
        RECT 73.290 149.270 75.190 149.410 ;
        RECT 65.855 148.885 66.145 149.115 ;
        RECT 66.300 148.870 66.620 149.130 ;
        RECT 67.220 148.870 67.540 149.130 ;
        RECT 69.150 149.115 69.290 149.270 ;
        RECT 69.980 149.210 70.300 149.270 ;
        RECT 74.900 149.225 75.190 149.270 ;
        RECT 69.070 148.885 69.360 149.115 ;
        RECT 69.535 148.885 69.825 149.115 ;
        RECT 70.440 149.070 70.760 149.130 ;
        RECT 71.375 149.070 71.665 149.115 ;
        RECT 71.820 149.070 72.140 149.130 ;
        RECT 70.440 148.930 72.140 149.070 ;
        RECT 57.650 148.590 61.930 148.730 ;
        RECT 66.760 148.730 67.080 148.790 ;
        RECT 69.610 148.730 69.750 148.885 ;
        RECT 70.440 148.870 70.760 148.930 ;
        RECT 71.375 148.885 71.665 148.930 ;
        RECT 71.820 148.870 72.140 148.930 ;
        RECT 66.760 148.590 69.750 148.730 ;
        RECT 66.760 148.530 67.080 148.590 ;
        RECT 69.980 148.530 70.300 148.790 ;
        RECT 70.900 148.730 71.220 148.790 ;
        RECT 72.420 148.730 72.710 148.775 ;
        RECT 70.900 148.590 72.710 148.730 ;
        RECT 70.900 148.530 71.220 148.590 ;
        RECT 72.420 148.545 72.710 148.590 ;
        RECT 73.660 148.530 73.980 148.790 ;
        RECT 74.555 148.730 74.845 148.775 ;
        RECT 75.745 148.730 76.035 148.775 ;
        RECT 78.265 148.730 78.555 148.775 ;
        RECT 74.555 148.590 78.555 148.730 ;
        RECT 74.555 148.545 74.845 148.590 ;
        RECT 75.745 148.545 76.035 148.590 ;
        RECT 78.265 148.545 78.555 148.590 ;
        RECT 21.695 148.390 21.985 148.435 ;
        RECT 22.600 148.390 22.920 148.450 ;
        RECT 25.360 148.390 25.680 148.450 ;
        RECT 21.695 148.250 22.920 148.390 ;
        RECT 21.695 148.205 21.985 148.250 ;
        RECT 22.600 148.190 22.920 148.250 ;
        RECT 23.150 148.250 25.680 148.390 ;
        RECT 19.855 148.050 20.145 148.095 ;
        RECT 23.150 148.050 23.290 148.250 ;
        RECT 25.360 148.190 25.680 148.250 ;
        RECT 30.895 148.390 31.185 148.435 ;
        RECT 40.080 148.390 40.400 148.450 ;
        RECT 30.895 148.250 40.400 148.390 ;
        RECT 30.895 148.205 31.185 148.250 ;
        RECT 40.080 148.190 40.400 148.250 ;
        RECT 41.000 148.390 41.290 148.435 ;
        RECT 42.570 148.390 42.860 148.435 ;
        RECT 44.670 148.390 44.960 148.435 ;
        RECT 41.000 148.250 44.960 148.390 ;
        RECT 41.000 148.205 41.290 148.250 ;
        RECT 42.570 148.205 42.860 148.250 ;
        RECT 44.670 148.205 44.960 148.250 ;
        RECT 74.160 148.390 74.450 148.435 ;
        RECT 76.260 148.390 76.550 148.435 ;
        RECT 77.830 148.390 78.120 148.435 ;
        RECT 74.160 148.250 78.120 148.390 ;
        RECT 74.160 148.205 74.450 148.250 ;
        RECT 76.260 148.205 76.550 148.250 ;
        RECT 77.830 148.205 78.120 148.250 ;
        RECT 19.855 147.910 23.290 148.050 ;
        RECT 23.535 148.050 23.825 148.095 ;
        RECT 25.820 148.050 26.140 148.110 ;
        RECT 23.535 147.910 26.140 148.050 ;
        RECT 19.855 147.865 20.145 147.910 ;
        RECT 23.535 147.865 23.825 147.910 ;
        RECT 25.820 147.850 26.140 147.910 ;
        RECT 11.950 147.230 90.610 147.710 ;
        RECT 29.055 147.030 29.345 147.075 ;
        RECT 30.420 147.030 30.740 147.090 ;
        RECT 29.055 146.890 30.740 147.030 ;
        RECT 29.055 146.845 29.345 146.890 ;
        RECT 30.420 146.830 30.740 146.890 ;
        RECT 35.480 147.030 35.800 147.090 ;
        RECT 37.335 147.030 37.625 147.075 ;
        RECT 35.480 146.890 37.625 147.030 ;
        RECT 35.480 146.830 35.800 146.890 ;
        RECT 37.335 146.845 37.625 146.890 ;
        RECT 42.380 146.830 42.700 147.090 ;
        RECT 57.560 147.030 57.880 147.090 ;
        RECT 58.955 147.030 59.245 147.075 ;
        RECT 59.875 147.030 60.165 147.075 ;
        RECT 57.560 146.890 60.165 147.030 ;
        RECT 57.560 146.830 57.880 146.890 ;
        RECT 58.955 146.845 59.245 146.890 ;
        RECT 59.875 146.845 60.165 146.890 ;
        RECT 61.700 147.030 62.020 147.090 ;
        RECT 62.175 147.030 62.465 147.075 ;
        RECT 61.700 146.890 62.465 147.030 ;
        RECT 61.700 146.830 62.020 146.890 ;
        RECT 62.175 146.845 62.465 146.890 ;
        RECT 27.660 146.690 27.980 146.750 ;
        RECT 33.180 146.690 33.500 146.750 ;
        RECT 45.600 146.690 45.920 146.750 ;
        RECT 27.660 146.550 33.500 146.690 ;
        RECT 27.660 146.490 27.980 146.550 ;
        RECT 33.180 146.490 33.500 146.550 ;
        RECT 41.090 146.550 45.920 146.690 ;
        RECT 41.090 146.410 41.230 146.550 ;
        RECT 45.600 146.490 45.920 146.550 ;
        RECT 73.200 146.690 73.520 146.750 ;
        RECT 74.595 146.690 74.885 146.735 ;
        RECT 76.895 146.690 77.185 146.735 ;
        RECT 73.200 146.550 77.185 146.690 ;
        RECT 73.200 146.490 73.520 146.550 ;
        RECT 74.595 146.505 74.885 146.550 ;
        RECT 76.895 146.505 77.185 146.550 ;
        RECT 100.010 146.720 100.780 150.410 ;
        RECT 102.460 149.360 105.310 150.480 ;
        RECT 105.700 150.180 106.050 150.930 ;
        RECT 106.800 150.810 108.670 150.970 ;
        RECT 106.800 150.760 107.560 150.810 ;
        RECT 108.440 150.740 108.670 150.810 ;
        RECT 117.080 150.740 117.310 150.970 ;
        RECT 108.875 150.460 116.875 150.690 ;
        RECT 105.700 150.120 105.990 150.180 ;
        RECT 105.610 150.000 105.990 150.120 ;
        RECT 108.970 150.060 116.830 150.460 ;
        RECT 117.640 150.060 118.600 159.540 ;
        RECT 119.930 159.670 120.770 161.800 ;
        RECT 126.430 161.380 127.680 161.820 ;
        RECT 137.600 161.800 138.460 163.870 ;
        RECT 124.370 161.370 129.610 161.380 ;
        RECT 121.420 161.270 136.720 161.370 ;
        RECT 121.420 161.260 136.755 161.270 ;
        RECT 121.380 161.140 136.755 161.260 ;
        RECT 121.380 161.030 125.380 161.140 ;
        RECT 126.430 161.060 128.170 161.140 ;
        RECT 128.750 161.060 136.755 161.140 ;
        RECT 126.430 160.980 127.680 161.060 ;
        RECT 128.755 161.040 136.755 161.060 ;
        RECT 120.990 160.730 121.220 160.980 ;
        RECT 125.540 160.840 125.770 160.980 ;
        RECT 128.320 160.840 128.550 160.990 ;
        RECT 125.540 160.730 128.550 160.840 ;
        RECT 136.960 160.730 137.190 160.990 ;
        RECT 120.990 160.290 137.190 160.730 ;
        RECT 120.990 160.020 121.220 160.290 ;
        RECT 125.540 160.260 137.190 160.290 ;
        RECT 125.540 160.170 128.550 160.260 ;
        RECT 125.540 160.020 125.770 160.170 ;
        RECT 128.320 160.030 128.550 160.170 ;
        RECT 136.960 160.030 137.190 160.260 ;
        RECT 121.380 159.740 125.380 159.970 ;
        RECT 128.755 159.760 136.755 159.980 ;
        RECT 137.520 159.760 138.480 161.800 ;
        RECT 128.755 159.750 138.480 159.760 ;
        RECT 121.380 159.670 125.370 159.740 ;
        RECT 119.930 159.560 125.370 159.670 ;
        RECT 128.810 159.590 138.480 159.750 ;
        RECT 119.930 159.470 123.060 159.560 ;
        RECT 136.550 159.540 138.480 159.590 ;
        RECT 119.930 156.200 120.770 159.470 ;
        RECT 124.410 159.010 129.660 159.020 ;
        RECT 124.410 158.900 136.720 159.010 ;
        RECT 121.440 158.840 136.720 158.900 ;
        RECT 121.440 158.830 136.755 158.840 ;
        RECT 121.380 158.700 136.755 158.830 ;
        RECT 121.380 158.690 126.540 158.700 ;
        RECT 121.380 158.600 125.380 158.690 ;
        RECT 128.755 158.610 136.755 158.700 ;
        RECT 128.840 158.600 136.730 158.610 ;
        RECT 120.990 158.240 121.220 158.550 ;
        RECT 121.440 158.240 125.340 158.600 ;
        RECT 125.540 158.240 125.770 158.550 ;
        RECT 120.990 156.900 125.770 158.240 ;
        RECT 120.990 156.590 121.220 156.900 ;
        RECT 125.540 156.590 125.770 156.900 ;
        RECT 128.320 158.020 128.550 158.560 ;
        RECT 129.360 158.020 130.370 158.050 ;
        RECT 136.960 158.020 137.190 158.560 ;
        RECT 128.320 157.120 137.190 158.020 ;
        RECT 128.320 156.600 128.550 157.120 ;
        RECT 129.360 157.050 130.370 157.120 ;
        RECT 136.960 156.600 137.190 157.120 ;
        RECT 121.380 156.310 125.380 156.540 ;
        RECT 128.755 156.320 136.755 156.550 ;
        RECT 119.930 156.160 121.060 156.200 ;
        RECT 119.930 156.080 121.300 156.160 ;
        RECT 121.670 156.090 125.330 156.310 ;
        RECT 121.670 156.080 123.110 156.090 ;
        RECT 119.930 156.040 123.110 156.080 ;
        RECT 119.930 155.950 122.620 156.040 ;
        RECT 128.820 156.030 136.710 156.320 ;
        RECT 119.930 155.890 121.950 155.950 ;
        RECT 119.930 155.840 121.700 155.890 ;
        RECT 119.930 152.500 120.770 155.840 ;
        RECT 128.810 155.540 136.730 155.550 ;
        RECT 125.040 155.530 136.730 155.540 ;
        RECT 121.420 155.410 136.730 155.530 ;
        RECT 121.420 155.400 136.755 155.410 ;
        RECT 121.380 155.280 136.755 155.400 ;
        RECT 121.380 155.170 125.380 155.280 ;
        RECT 120.990 154.830 121.220 155.120 ;
        RECT 121.440 154.830 125.330 155.170 ;
        RECT 125.540 154.830 125.770 155.120 ;
        RECT 120.990 153.460 125.770 154.830 ;
        RECT 120.990 153.160 121.220 153.460 ;
        RECT 125.540 153.160 125.770 153.460 ;
        RECT 121.380 152.880 125.380 153.110 ;
        RECT 121.630 152.650 125.200 152.880 ;
        RECT 121.630 152.500 125.320 152.650 ;
        RECT 119.930 152.220 125.320 152.500 ;
        RECT 126.570 152.330 127.190 155.280 ;
        RECT 128.755 155.180 136.755 155.280 ;
        RECT 128.810 155.170 136.730 155.180 ;
        RECT 128.320 154.470 128.550 155.130 ;
        RECT 129.330 154.470 130.330 154.560 ;
        RECT 136.960 154.470 137.190 155.130 ;
        RECT 128.320 153.650 137.190 154.470 ;
        RECT 128.320 153.170 128.550 153.650 ;
        RECT 129.330 153.560 130.330 153.650 ;
        RECT 136.960 153.170 137.190 153.650 ;
        RECT 128.755 152.890 136.755 153.120 ;
        RECT 119.930 151.760 125.330 152.220 ;
        RECT 119.930 150.420 121.930 151.760 ;
        RECT 123.680 151.750 125.330 151.760 ;
        RECT 122.370 150.480 123.370 151.200 ;
        RECT 123.680 150.940 123.990 151.750 ;
        RECT 124.450 151.470 125.330 151.750 ;
        RECT 125.570 151.930 127.190 152.330 ;
        RECT 128.840 151.980 136.710 152.890 ;
        RECT 124.390 151.240 125.390 151.470 ;
        RECT 125.570 151.280 125.920 151.930 ;
        RECT 126.570 151.920 127.190 151.930 ;
        RECT 128.755 151.750 136.755 151.980 ;
        RECT 128.840 151.740 136.710 151.750 ;
        RECT 124.450 151.030 125.330 151.050 ;
        RECT 123.720 150.650 123.990 150.940 ;
        RECT 124.390 150.800 125.390 151.030 ;
        RECT 125.550 150.990 125.920 151.280 ;
        RECT 125.580 150.930 125.920 150.990 ;
        RECT 126.680 151.600 127.440 151.650 ;
        RECT 128.320 151.600 128.550 151.700 ;
        RECT 126.680 151.390 128.550 151.600 ;
        RECT 136.960 151.390 137.190 151.700 ;
        RECT 126.680 150.970 129.220 151.390 ;
        RECT 136.590 150.970 137.190 151.390 ;
        RECT 124.450 150.650 125.330 150.800 ;
        RECT 124.460 150.480 125.190 150.650 ;
        RECT 102.400 149.130 105.400 149.360 ;
        RECT 105.610 149.170 105.950 150.000 ;
        RECT 107.960 149.990 118.600 150.060 ;
        RECT 102.450 149.100 105.310 149.130 ;
        RECT 102.450 149.080 103.620 149.100 ;
        RECT 104.580 149.090 105.310 149.100 ;
        RECT 102.400 148.690 105.400 148.920 ;
        RECT 105.605 148.880 105.950 149.170 ;
        RECT 106.140 148.950 118.600 149.990 ;
        RECT 120.000 150.410 121.930 150.420 ;
        RECT 106.140 148.930 118.560 148.950 ;
        RECT 105.610 148.770 105.950 148.880 ;
        RECT 106.180 148.920 111.850 148.930 ;
        RECT 112.850 148.920 118.560 148.930 ;
        RECT 102.490 148.520 105.350 148.690 ;
        RECT 106.180 148.520 106.610 148.920 ;
        RECT 102.460 148.150 106.610 148.520 ;
        RECT 26.280 146.350 26.600 146.410 ;
        RECT 26.280 146.210 32.490 146.350 ;
        RECT 26.280 146.150 26.600 146.210 ;
        RECT 26.740 145.810 27.060 146.070 ;
        RECT 27.660 145.810 27.980 146.070 ;
        RECT 28.120 146.010 28.440 146.070 ;
        RECT 29.960 146.010 30.280 146.070 ;
        RECT 31.430 146.055 31.570 146.210 ;
        RECT 28.120 145.870 30.280 146.010 ;
        RECT 28.120 145.810 28.440 145.870 ;
        RECT 29.960 145.810 30.280 145.870 ;
        RECT 31.355 145.825 31.645 146.055 ;
        RECT 31.815 145.825 32.105 146.055 ;
        RECT 31.890 145.670 32.030 145.825 ;
        RECT 30.970 145.530 32.030 145.670 ;
        RECT 32.350 145.670 32.490 146.210 ;
        RECT 41.000 146.150 41.320 146.410 ;
        RECT 41.460 146.395 41.780 146.410 ;
        RECT 41.460 146.165 41.890 146.395 ;
        RECT 69.995 146.350 70.285 146.395 ;
        RECT 73.660 146.350 73.980 146.410 ;
        RECT 69.995 146.210 73.980 146.350 ;
        RECT 69.995 146.165 70.285 146.210 ;
        RECT 41.460 146.150 41.780 146.165 ;
        RECT 35.035 146.010 35.325 146.055 ;
        RECT 37.795 146.010 38.085 146.055 ;
        RECT 35.035 145.870 38.085 146.010 ;
        RECT 35.035 145.825 35.325 145.870 ;
        RECT 37.795 145.825 38.085 145.870 ;
        RECT 39.175 146.010 39.465 146.055 ;
        RECT 47.440 146.010 47.760 146.070 ;
        RECT 39.175 145.870 47.760 146.010 ;
        RECT 39.175 145.825 39.465 145.870 ;
        RECT 47.440 145.810 47.760 145.870 ;
        RECT 57.575 145.825 57.865 146.055 ;
        RECT 58.035 146.010 58.325 146.055 ;
        RECT 58.940 146.010 59.260 146.070 ;
        RECT 58.035 145.870 59.260 146.010 ;
        RECT 58.035 145.825 58.325 145.870 ;
        RECT 35.495 145.670 35.785 145.715 ;
        RECT 32.350 145.530 35.785 145.670 ;
        RECT 24.900 145.330 25.220 145.390 ;
        RECT 27.215 145.330 27.505 145.375 ;
        RECT 24.900 145.190 27.505 145.330 ;
        RECT 24.900 145.130 25.220 145.190 ;
        RECT 27.215 145.145 27.505 145.190 ;
        RECT 30.420 145.330 30.740 145.390 ;
        RECT 30.970 145.375 31.110 145.530 ;
        RECT 35.495 145.485 35.785 145.530 ;
        RECT 36.415 145.485 36.705 145.715 ;
        RECT 40.555 145.670 40.845 145.715 ;
        RECT 46.060 145.670 46.380 145.730 ;
        RECT 48.360 145.670 48.680 145.730 ;
        RECT 40.555 145.530 48.680 145.670 ;
        RECT 57.650 145.670 57.790 145.825 ;
        RECT 58.940 145.810 59.260 145.870 ;
        RECT 59.400 145.810 59.720 146.070 ;
        RECT 61.255 146.010 61.545 146.055 ;
        RECT 64.000 146.010 64.320 146.070 ;
        RECT 61.255 145.870 64.320 146.010 ;
        RECT 61.255 145.825 61.545 145.870 ;
        RECT 64.000 145.810 64.320 145.870 ;
        RECT 65.395 146.010 65.685 146.055 ;
        RECT 70.070 146.010 70.210 146.165 ;
        RECT 73.660 146.150 73.980 146.210 ;
        RECT 65.395 145.870 68.600 146.010 ;
        RECT 65.395 145.825 65.685 145.870 ;
        RECT 68.460 145.730 68.600 145.870 ;
        RECT 59.860 145.670 60.180 145.730 ;
        RECT 57.650 145.530 60.180 145.670 ;
        RECT 40.555 145.485 40.845 145.530 ;
        RECT 30.895 145.330 31.185 145.375 ;
        RECT 36.490 145.330 36.630 145.485 ;
        RECT 46.060 145.470 46.380 145.530 ;
        RECT 48.360 145.470 48.680 145.530 ;
        RECT 59.860 145.470 60.180 145.530 ;
        RECT 63.540 145.670 63.860 145.730 ;
        RECT 65.840 145.670 66.160 145.730 ;
        RECT 63.540 145.530 66.160 145.670 ;
        RECT 63.540 145.470 63.860 145.530 ;
        RECT 65.840 145.470 66.160 145.530 ;
        RECT 68.140 145.670 68.600 145.730 ;
        RECT 69.150 145.870 70.210 146.010 ;
        RECT 69.150 145.670 69.290 145.870 ;
        RECT 72.280 145.810 72.600 146.070 ;
        RECT 75.500 146.010 75.820 146.070 ;
        RECT 77.815 146.010 78.105 146.055 ;
        RECT 75.500 145.870 78.105 146.010 ;
        RECT 75.500 145.810 75.820 145.870 ;
        RECT 77.815 145.825 78.105 145.870 ;
        RECT 68.140 145.530 69.290 145.670 ;
        RECT 69.520 145.670 69.840 145.730 ;
        RECT 71.835 145.670 72.125 145.715 ;
        RECT 74.120 145.670 74.440 145.730 ;
        RECT 69.520 145.530 74.440 145.670 ;
        RECT 68.140 145.470 68.460 145.530 ;
        RECT 69.520 145.470 69.840 145.530 ;
        RECT 71.835 145.485 72.125 145.530 ;
        RECT 74.120 145.470 74.440 145.530 ;
        RECT 74.595 145.670 74.885 145.715 ;
        RECT 75.040 145.670 75.360 145.730 ;
        RECT 74.595 145.530 75.360 145.670 ;
        RECT 74.595 145.485 74.885 145.530 ;
        RECT 75.040 145.470 75.360 145.530 ;
        RECT 30.420 145.190 36.630 145.330 ;
        RECT 37.780 145.330 38.100 145.390 ;
        RECT 38.255 145.330 38.545 145.375 ;
        RECT 37.780 145.190 38.545 145.330 ;
        RECT 30.420 145.130 30.740 145.190 ;
        RECT 30.895 145.145 31.185 145.190 ;
        RECT 37.780 145.130 38.100 145.190 ;
        RECT 38.255 145.145 38.545 145.190 ;
        RECT 70.900 145.130 71.220 145.390 ;
        RECT 11.950 144.510 90.610 144.990 ;
        RECT 100.010 144.620 100.880 146.720 ;
        RECT 106.550 146.330 107.800 146.770 ;
        RECT 117.700 146.750 118.560 148.920 ;
        RECT 120.000 146.750 120.770 150.410 ;
        RECT 122.340 149.360 125.190 150.480 ;
        RECT 125.580 150.180 125.930 150.930 ;
        RECT 126.680 150.810 128.550 150.970 ;
        RECT 126.680 150.760 127.440 150.810 ;
        RECT 128.320 150.740 128.550 150.810 ;
        RECT 136.960 150.740 137.190 150.970 ;
        RECT 128.755 150.460 136.755 150.690 ;
        RECT 125.580 150.120 125.870 150.180 ;
        RECT 125.490 150.000 125.870 150.120 ;
        RECT 128.850 150.060 136.710 150.460 ;
        RECT 137.520 150.060 138.480 159.540 ;
        RECT 122.280 149.130 125.280 149.360 ;
        RECT 125.490 149.170 125.830 150.000 ;
        RECT 127.840 149.990 138.480 150.060 ;
        RECT 122.330 149.100 125.190 149.130 ;
        RECT 122.330 149.080 123.500 149.100 ;
        RECT 124.460 149.090 125.190 149.100 ;
        RECT 122.280 148.690 125.280 148.920 ;
        RECT 125.485 148.880 125.830 149.170 ;
        RECT 126.020 148.950 138.480 149.990 ;
        RECT 139.930 161.720 140.700 165.410 ;
        RECT 142.370 164.360 145.220 165.480 ;
        RECT 145.610 165.180 145.960 165.930 ;
        RECT 146.710 165.810 148.580 165.970 ;
        RECT 146.710 165.760 147.470 165.810 ;
        RECT 148.350 165.740 148.580 165.810 ;
        RECT 156.990 165.740 157.220 165.970 ;
        RECT 148.785 165.460 156.785 165.690 ;
        RECT 145.610 165.120 145.900 165.180 ;
        RECT 145.520 165.000 145.900 165.120 ;
        RECT 148.880 165.060 156.740 165.460 ;
        RECT 157.550 165.060 158.510 174.540 ;
        RECT 142.310 164.130 145.310 164.360 ;
        RECT 145.520 164.170 145.860 165.000 ;
        RECT 147.870 164.990 158.510 165.060 ;
        RECT 142.360 164.100 145.220 164.130 ;
        RECT 142.360 164.080 143.530 164.100 ;
        RECT 144.490 164.090 145.220 164.100 ;
        RECT 142.310 163.690 145.310 163.920 ;
        RECT 145.515 163.880 145.860 164.170 ;
        RECT 146.050 163.950 158.510 164.990 ;
        RECT 146.050 163.930 158.500 163.950 ;
        RECT 145.520 163.770 145.860 163.880 ;
        RECT 146.090 163.920 151.760 163.930 ;
        RECT 152.760 163.920 158.500 163.930 ;
        RECT 142.400 163.520 145.260 163.690 ;
        RECT 146.090 163.520 146.520 163.920 ;
        RECT 142.370 163.150 146.520 163.520 ;
        RECT 139.930 159.620 140.840 161.720 ;
        RECT 146.510 161.330 147.760 161.770 ;
        RECT 157.640 161.750 158.500 163.920 ;
        RECT 144.450 161.320 149.690 161.330 ;
        RECT 141.500 161.220 156.800 161.320 ;
        RECT 141.500 161.210 156.835 161.220 ;
        RECT 141.460 161.090 156.835 161.210 ;
        RECT 141.460 160.980 145.460 161.090 ;
        RECT 146.510 161.010 148.250 161.090 ;
        RECT 148.830 161.010 156.835 161.090 ;
        RECT 146.510 160.930 147.760 161.010 ;
        RECT 148.835 160.990 156.835 161.010 ;
        RECT 141.070 160.680 141.300 160.930 ;
        RECT 145.620 160.790 145.850 160.930 ;
        RECT 148.400 160.790 148.630 160.940 ;
        RECT 145.620 160.680 148.630 160.790 ;
        RECT 157.040 160.680 157.270 160.940 ;
        RECT 141.070 160.240 157.270 160.680 ;
        RECT 141.070 159.970 141.300 160.240 ;
        RECT 145.620 160.210 157.270 160.240 ;
        RECT 145.620 160.120 148.630 160.210 ;
        RECT 145.620 159.970 145.850 160.120 ;
        RECT 148.400 159.980 148.630 160.120 ;
        RECT 157.040 159.980 157.270 160.210 ;
        RECT 141.460 159.690 145.460 159.920 ;
        RECT 148.835 159.710 156.835 159.930 ;
        RECT 157.600 159.710 158.560 161.750 ;
        RECT 148.835 159.700 158.560 159.710 ;
        RECT 141.460 159.620 145.450 159.690 ;
        RECT 139.930 159.510 145.450 159.620 ;
        RECT 148.890 159.540 158.560 159.700 ;
        RECT 139.930 159.420 143.140 159.510 ;
        RECT 156.630 159.490 158.560 159.540 ;
        RECT 139.930 156.150 140.840 159.420 ;
        RECT 144.490 158.960 149.740 158.970 ;
        RECT 144.490 158.850 156.800 158.960 ;
        RECT 141.520 158.790 156.800 158.850 ;
        RECT 141.520 158.780 156.835 158.790 ;
        RECT 141.460 158.650 156.835 158.780 ;
        RECT 141.460 158.640 146.620 158.650 ;
        RECT 141.460 158.550 145.460 158.640 ;
        RECT 148.835 158.560 156.835 158.650 ;
        RECT 148.920 158.550 156.810 158.560 ;
        RECT 141.070 158.190 141.300 158.500 ;
        RECT 141.520 158.190 145.420 158.550 ;
        RECT 145.620 158.190 145.850 158.500 ;
        RECT 141.070 156.850 145.850 158.190 ;
        RECT 141.070 156.540 141.300 156.850 ;
        RECT 145.620 156.540 145.850 156.850 ;
        RECT 148.400 157.970 148.630 158.510 ;
        RECT 149.440 157.970 150.450 158.000 ;
        RECT 157.040 157.970 157.270 158.510 ;
        RECT 148.400 157.070 157.270 157.970 ;
        RECT 148.400 156.550 148.630 157.070 ;
        RECT 149.440 157.000 150.450 157.070 ;
        RECT 157.040 156.550 157.270 157.070 ;
        RECT 141.460 156.260 145.460 156.490 ;
        RECT 148.835 156.270 156.835 156.500 ;
        RECT 139.930 156.110 141.140 156.150 ;
        RECT 139.930 156.030 141.380 156.110 ;
        RECT 141.750 156.040 145.410 156.260 ;
        RECT 141.750 156.030 143.190 156.040 ;
        RECT 139.930 155.990 143.190 156.030 ;
        RECT 139.930 155.900 142.700 155.990 ;
        RECT 148.900 155.980 156.790 156.270 ;
        RECT 139.930 155.840 142.030 155.900 ;
        RECT 139.930 155.790 141.780 155.840 ;
        RECT 139.930 152.450 140.840 155.790 ;
        RECT 148.890 155.490 156.810 155.500 ;
        RECT 145.120 155.480 156.810 155.490 ;
        RECT 141.500 155.360 156.810 155.480 ;
        RECT 141.500 155.350 156.835 155.360 ;
        RECT 141.460 155.230 156.835 155.350 ;
        RECT 141.460 155.120 145.460 155.230 ;
        RECT 141.070 154.780 141.300 155.070 ;
        RECT 141.520 154.780 145.410 155.120 ;
        RECT 145.620 154.780 145.850 155.070 ;
        RECT 141.070 153.410 145.850 154.780 ;
        RECT 141.070 153.110 141.300 153.410 ;
        RECT 145.620 153.110 145.850 153.410 ;
        RECT 141.460 152.830 145.460 153.060 ;
        RECT 141.710 152.600 145.280 152.830 ;
        RECT 141.710 152.450 145.400 152.600 ;
        RECT 139.930 152.170 145.400 152.450 ;
        RECT 146.650 152.280 147.270 155.230 ;
        RECT 148.835 155.130 156.835 155.230 ;
        RECT 148.890 155.120 156.810 155.130 ;
        RECT 148.400 154.420 148.630 155.080 ;
        RECT 149.410 154.420 150.410 154.510 ;
        RECT 157.040 154.420 157.270 155.080 ;
        RECT 148.400 153.600 157.270 154.420 ;
        RECT 148.400 153.120 148.630 153.600 ;
        RECT 149.410 153.510 150.410 153.600 ;
        RECT 157.040 153.120 157.270 153.600 ;
        RECT 148.835 152.840 156.835 153.070 ;
        RECT 139.930 151.710 145.410 152.170 ;
        RECT 139.930 150.360 142.010 151.710 ;
        RECT 143.760 151.700 145.410 151.710 ;
        RECT 142.450 150.430 143.450 151.150 ;
        RECT 143.760 150.890 144.070 151.700 ;
        RECT 144.530 151.420 145.410 151.700 ;
        RECT 145.650 151.880 147.270 152.280 ;
        RECT 148.920 151.930 156.790 152.840 ;
        RECT 144.470 151.190 145.470 151.420 ;
        RECT 145.650 151.230 146.000 151.880 ;
        RECT 146.650 151.870 147.270 151.880 ;
        RECT 148.835 151.700 156.835 151.930 ;
        RECT 148.920 151.690 156.790 151.700 ;
        RECT 144.530 150.980 145.410 151.000 ;
        RECT 143.800 150.600 144.070 150.890 ;
        RECT 144.470 150.750 145.470 150.980 ;
        RECT 145.630 150.940 146.000 151.230 ;
        RECT 145.660 150.880 146.000 150.940 ;
        RECT 146.760 151.550 147.520 151.600 ;
        RECT 148.400 151.550 148.630 151.650 ;
        RECT 146.760 151.340 148.630 151.550 ;
        RECT 157.040 151.340 157.270 151.650 ;
        RECT 146.760 150.920 149.300 151.340 ;
        RECT 156.670 150.920 157.270 151.340 ;
        RECT 144.530 150.600 145.410 150.750 ;
        RECT 144.540 150.430 145.270 150.600 ;
        RECT 126.020 148.930 138.460 148.950 ;
        RECT 125.490 148.770 125.830 148.880 ;
        RECT 126.060 148.920 131.730 148.930 ;
        RECT 132.730 148.920 138.460 148.930 ;
        RECT 122.370 148.520 125.230 148.690 ;
        RECT 126.060 148.520 126.490 148.920 ;
        RECT 122.340 148.150 126.490 148.520 ;
        RECT 104.490 146.320 109.730 146.330 ;
        RECT 101.540 146.220 116.840 146.320 ;
        RECT 101.540 146.210 116.875 146.220 ;
        RECT 101.500 146.090 116.875 146.210 ;
        RECT 101.500 145.980 105.500 146.090 ;
        RECT 106.550 146.010 108.290 146.090 ;
        RECT 108.870 146.010 116.875 146.090 ;
        RECT 106.550 145.930 107.800 146.010 ;
        RECT 108.875 145.990 116.875 146.010 ;
        RECT 101.110 145.680 101.340 145.930 ;
        RECT 105.660 145.790 105.890 145.930 ;
        RECT 108.440 145.790 108.670 145.940 ;
        RECT 105.660 145.680 108.670 145.790 ;
        RECT 117.080 145.680 117.310 145.940 ;
        RECT 101.110 145.240 117.310 145.680 ;
        RECT 101.110 144.970 101.340 145.240 ;
        RECT 105.660 145.210 117.310 145.240 ;
        RECT 105.660 145.120 108.670 145.210 ;
        RECT 105.660 144.970 105.890 145.120 ;
        RECT 108.440 144.980 108.670 145.120 ;
        RECT 117.080 144.980 117.310 145.210 ;
        RECT 101.500 144.690 105.500 144.920 ;
        RECT 108.875 144.710 116.875 144.930 ;
        RECT 117.640 144.710 118.600 146.750 ;
        RECT 108.875 144.700 118.600 144.710 ;
        RECT 101.500 144.620 105.490 144.690 ;
        RECT 100.010 144.510 105.490 144.620 ;
        RECT 108.930 144.540 118.600 144.700 ;
        RECT 100.010 144.420 103.180 144.510 ;
        RECT 116.670 144.490 118.600 144.540 ;
        RECT 21.695 144.310 21.985 144.355 ;
        RECT 24.440 144.310 24.760 144.370 ;
        RECT 26.740 144.310 27.060 144.370 ;
        RECT 21.695 144.170 27.060 144.310 ;
        RECT 21.695 144.125 21.985 144.170 ;
        RECT 24.440 144.110 24.760 144.170 ;
        RECT 26.740 144.110 27.060 144.170 ;
        RECT 49.740 144.310 50.060 144.370 ;
        RECT 50.215 144.310 50.505 144.355 ;
        RECT 49.740 144.170 50.505 144.310 ;
        RECT 49.740 144.110 50.060 144.170 ;
        RECT 50.215 144.125 50.505 144.170 ;
        RECT 58.495 144.310 58.785 144.355 ;
        RECT 59.400 144.310 59.720 144.370 ;
        RECT 58.495 144.170 59.720 144.310 ;
        RECT 58.495 144.125 58.785 144.170 ;
        RECT 59.400 144.110 59.720 144.170 ;
        RECT 64.000 144.110 64.320 144.370 ;
        RECT 75.040 144.310 75.360 144.370 ;
        RECT 75.515 144.310 75.805 144.355 ;
        RECT 75.040 144.170 75.805 144.310 ;
        RECT 75.040 144.110 75.360 144.170 ;
        RECT 75.515 144.125 75.805 144.170 ;
        RECT 27.660 143.970 27.980 144.030 ;
        RECT 26.370 143.830 27.980 143.970 ;
        RECT 22.600 143.630 22.920 143.690 ;
        RECT 23.995 143.630 24.285 143.675 ;
        RECT 22.600 143.490 24.285 143.630 ;
        RECT 22.600 143.430 22.920 143.490 ;
        RECT 23.995 143.445 24.285 143.490 ;
        RECT 24.915 143.630 25.205 143.675 ;
        RECT 25.820 143.630 26.140 143.690 ;
        RECT 26.370 143.675 26.510 143.830 ;
        RECT 27.660 143.770 27.980 143.830 ;
        RECT 29.975 143.970 30.265 144.015 ;
        RECT 32.720 143.970 33.040 144.030 ;
        RECT 37.780 143.970 38.100 144.030 ;
        RECT 45.140 143.970 45.460 144.030 ;
        RECT 48.820 143.970 49.140 144.030 ;
        RECT 29.975 143.830 33.040 143.970 ;
        RECT 29.975 143.785 30.265 143.830 ;
        RECT 32.720 143.770 33.040 143.830 ;
        RECT 36.950 143.830 38.100 143.970 ;
        RECT 24.915 143.490 26.140 143.630 ;
        RECT 24.915 143.445 25.205 143.490 ;
        RECT 23.535 143.290 23.825 143.335 ;
        RECT 24.990 143.290 25.130 143.445 ;
        RECT 25.820 143.430 26.140 143.490 ;
        RECT 26.295 143.445 26.585 143.675 ;
        RECT 23.535 143.150 25.130 143.290 ;
        RECT 25.360 143.290 25.680 143.350 ;
        RECT 26.370 143.290 26.510 143.445 ;
        RECT 28.120 143.430 28.440 143.690 ;
        RECT 36.950 143.675 37.090 143.830 ;
        RECT 37.780 143.770 38.100 143.830 ;
        RECT 38.330 143.830 45.460 143.970 ;
        RECT 38.330 143.690 38.470 143.830 ;
        RECT 45.140 143.770 45.460 143.830 ;
        RECT 47.070 143.830 49.140 143.970 ;
        RECT 28.595 143.630 28.885 143.675 ;
        RECT 36.875 143.630 37.165 143.675 ;
        RECT 28.595 143.490 37.165 143.630 ;
        RECT 28.595 143.445 28.885 143.490 ;
        RECT 36.875 143.445 37.165 143.490 ;
        RECT 37.335 143.445 37.625 143.675 ;
        RECT 25.360 143.150 26.510 143.290 ;
        RECT 29.500 143.290 29.820 143.350 ;
        RECT 33.655 143.290 33.945 143.335 ;
        RECT 29.500 143.150 33.945 143.290 ;
        RECT 23.535 143.105 23.825 143.150 ;
        RECT 25.360 143.090 25.680 143.150 ;
        RECT 29.500 143.090 29.820 143.150 ;
        RECT 33.655 143.105 33.945 143.150 ;
        RECT 35.020 143.090 35.340 143.350 ;
        RECT 24.900 142.950 25.220 143.010 ;
        RECT 37.410 142.950 37.550 143.445 ;
        RECT 38.240 143.430 38.560 143.690 ;
        RECT 40.080 143.630 40.400 143.690 ;
        RECT 41.935 143.630 42.225 143.675 ;
        RECT 40.080 143.490 42.225 143.630 ;
        RECT 40.080 143.430 40.400 143.490 ;
        RECT 41.935 143.445 42.225 143.490 ;
        RECT 43.300 143.630 43.620 143.690 ;
        RECT 47.070 143.675 47.210 143.830 ;
        RECT 48.820 143.770 49.140 143.830 ;
        RECT 49.295 143.970 49.585 144.015 ;
        RECT 58.020 143.970 58.340 144.030 ;
        RECT 69.950 143.970 70.240 144.015 ;
        RECT 70.900 143.970 71.220 144.030 ;
        RECT 49.295 143.830 57.790 143.970 ;
        RECT 49.295 143.785 49.585 143.830 ;
        RECT 43.300 143.490 43.990 143.630 ;
        RECT 43.300 143.430 43.620 143.490 ;
        RECT 24.900 142.810 37.550 142.950 ;
        RECT 43.850 142.950 43.990 143.490 ;
        RECT 44.235 143.445 44.525 143.675 ;
        RECT 46.995 143.445 47.285 143.675 ;
        RECT 44.310 143.290 44.450 143.445 ;
        RECT 47.900 143.430 48.220 143.690 ;
        RECT 55.720 143.675 56.040 143.690 ;
        RECT 55.720 143.445 56.070 143.675 ;
        RECT 57.650 143.630 57.790 143.830 ;
        RECT 58.020 143.830 65.610 143.970 ;
        RECT 58.020 143.770 58.340 143.830 ;
        RECT 58.480 143.630 58.800 143.690 ;
        RECT 57.650 143.490 58.800 143.630 ;
        RECT 55.720 143.430 56.040 143.445 ;
        RECT 58.480 143.430 58.800 143.490 ;
        RECT 58.940 143.630 59.260 143.690 ;
        RECT 59.415 143.630 59.705 143.675 ;
        RECT 58.940 143.490 59.705 143.630 ;
        RECT 58.940 143.430 59.260 143.490 ;
        RECT 59.415 143.445 59.705 143.490 ;
        RECT 59.860 143.430 60.180 143.690 ;
        RECT 61.330 143.675 61.470 143.830 ;
        RECT 61.255 143.445 61.545 143.675 ;
        RECT 64.920 143.430 65.240 143.690 ;
        RECT 47.455 143.290 47.745 143.335 ;
        RECT 44.310 143.150 47.745 143.290 ;
        RECT 47.455 143.105 47.745 143.150 ;
        RECT 52.525 143.290 52.815 143.335 ;
        RECT 55.045 143.290 55.335 143.335 ;
        RECT 56.235 143.290 56.525 143.335 ;
        RECT 52.525 143.150 56.525 143.290 ;
        RECT 52.525 143.105 52.815 143.150 ;
        RECT 55.045 143.105 55.335 143.150 ;
        RECT 56.235 143.105 56.525 143.150 ;
        RECT 57.100 143.090 57.420 143.350 ;
        RECT 60.795 143.290 61.085 143.335 ;
        RECT 65.010 143.290 65.150 143.430 ;
        RECT 60.795 143.150 65.150 143.290 ;
        RECT 65.470 143.290 65.610 143.830 ;
        RECT 69.950 143.830 71.220 143.970 ;
        RECT 69.950 143.785 70.240 143.830 ;
        RECT 70.900 143.770 71.220 143.830 ;
        RECT 65.855 143.630 66.145 143.675 ;
        RECT 66.760 143.630 67.080 143.690 ;
        RECT 65.855 143.490 67.080 143.630 ;
        RECT 65.855 143.445 66.145 143.490 ;
        RECT 66.760 143.430 67.080 143.490 ;
        RECT 66.315 143.290 66.605 143.335 ;
        RECT 65.470 143.150 66.605 143.290 ;
        RECT 60.795 143.105 61.085 143.150 ;
        RECT 66.315 143.105 66.605 143.150 ;
        RECT 68.140 143.290 68.460 143.350 ;
        RECT 68.615 143.290 68.905 143.335 ;
        RECT 68.140 143.150 68.905 143.290 ;
        RECT 68.140 143.090 68.460 143.150 ;
        RECT 68.615 143.105 68.905 143.150 ;
        RECT 69.495 143.290 69.785 143.335 ;
        RECT 70.685 143.290 70.975 143.335 ;
        RECT 73.205 143.290 73.495 143.335 ;
        RECT 69.495 143.150 73.495 143.290 ;
        RECT 69.495 143.105 69.785 143.150 ;
        RECT 70.685 143.105 70.975 143.150 ;
        RECT 73.205 143.105 73.495 143.150 ;
        RECT 48.360 142.950 48.680 143.010 ;
        RECT 43.850 142.810 48.680 142.950 ;
        RECT 24.900 142.750 25.220 142.810 ;
        RECT 48.360 142.750 48.680 142.810 ;
        RECT 52.960 142.950 53.250 142.995 ;
        RECT 54.530 142.950 54.820 142.995 ;
        RECT 56.630 142.950 56.920 142.995 ;
        RECT 52.960 142.810 56.920 142.950 ;
        RECT 52.960 142.765 53.250 142.810 ;
        RECT 54.530 142.765 54.820 142.810 ;
        RECT 56.630 142.765 56.920 142.810 ;
        RECT 69.100 142.950 69.390 142.995 ;
        RECT 71.200 142.950 71.490 142.995 ;
        RECT 72.770 142.950 73.060 142.995 ;
        RECT 69.100 142.810 73.060 142.950 ;
        RECT 69.100 142.765 69.390 142.810 ;
        RECT 71.200 142.765 71.490 142.810 ;
        RECT 72.770 142.765 73.060 142.810 ;
        RECT 25.820 142.410 26.140 142.670 ;
        RECT 26.280 142.610 26.600 142.670 ;
        RECT 26.755 142.610 27.045 142.655 ;
        RECT 26.280 142.470 27.045 142.610 ;
        RECT 26.280 142.410 26.600 142.470 ;
        RECT 26.755 142.425 27.045 142.470 ;
        RECT 29.515 142.610 29.805 142.655 ;
        RECT 29.960 142.610 30.280 142.670 ;
        RECT 29.515 142.470 30.280 142.610 ;
        RECT 29.515 142.425 29.805 142.470 ;
        RECT 29.960 142.410 30.280 142.470 ;
        RECT 35.955 142.610 36.245 142.655 ;
        RECT 37.780 142.610 38.100 142.670 ;
        RECT 35.955 142.470 38.100 142.610 ;
        RECT 35.955 142.425 36.245 142.470 ;
        RECT 37.780 142.410 38.100 142.470 ;
        RECT 41.000 142.410 41.320 142.670 ;
        RECT 44.220 142.410 44.540 142.670 ;
        RECT 46.060 142.610 46.380 142.670 ;
        RECT 48.835 142.610 49.125 142.655 ;
        RECT 52.040 142.610 52.360 142.670 ;
        RECT 46.060 142.470 52.360 142.610 ;
        RECT 46.060 142.410 46.380 142.470 ;
        RECT 48.835 142.425 49.125 142.470 ;
        RECT 52.040 142.410 52.360 142.470 ;
        RECT 11.950 141.790 90.610 142.270 ;
        RECT 24.455 141.590 24.745 141.635 ;
        RECT 26.280 141.590 26.600 141.650 ;
        RECT 35.020 141.590 35.340 141.650 ;
        RECT 24.455 141.450 26.600 141.590 ;
        RECT 24.455 141.405 24.745 141.450 ;
        RECT 26.280 141.390 26.600 141.450 ;
        RECT 26.830 141.450 35.340 141.590 ;
        RECT 26.830 141.310 26.970 141.450 ;
        RECT 35.020 141.390 35.340 141.450 ;
        RECT 47.455 141.590 47.745 141.635 ;
        RECT 48.820 141.590 49.140 141.650 ;
        RECT 47.455 141.450 49.140 141.590 ;
        RECT 47.455 141.405 47.745 141.450 ;
        RECT 48.820 141.390 49.140 141.450 ;
        RECT 49.295 141.590 49.585 141.635 ;
        RECT 53.880 141.590 54.200 141.650 ;
        RECT 55.720 141.590 56.040 141.650 ;
        RECT 49.295 141.450 54.200 141.590 ;
        RECT 49.295 141.405 49.585 141.450 ;
        RECT 53.880 141.390 54.200 141.450 ;
        RECT 54.430 141.450 56.040 141.590 ;
        RECT 18.040 141.250 18.330 141.295 ;
        RECT 20.140 141.250 20.430 141.295 ;
        RECT 21.710 141.250 22.000 141.295 ;
        RECT 18.040 141.110 22.000 141.250 ;
        RECT 18.040 141.065 18.330 141.110 ;
        RECT 20.140 141.065 20.430 141.110 ;
        RECT 21.710 141.065 22.000 141.110 ;
        RECT 26.740 141.050 27.060 141.310 ;
        RECT 30.420 141.250 30.710 141.295 ;
        RECT 31.990 141.250 32.280 141.295 ;
        RECT 34.090 141.250 34.380 141.295 ;
        RECT 30.420 141.110 34.380 141.250 ;
        RECT 30.420 141.065 30.710 141.110 ;
        RECT 31.990 141.065 32.280 141.110 ;
        RECT 34.090 141.065 34.380 141.110 ;
        RECT 41.040 141.250 41.330 141.295 ;
        RECT 43.140 141.250 43.430 141.295 ;
        RECT 44.710 141.250 45.000 141.295 ;
        RECT 41.040 141.110 45.000 141.250 ;
        RECT 41.040 141.065 41.330 141.110 ;
        RECT 43.140 141.065 43.430 141.110 ;
        RECT 44.710 141.065 45.000 141.110 ;
        RECT 47.900 141.250 48.220 141.310 ;
        RECT 50.215 141.250 50.505 141.295 ;
        RECT 51.120 141.250 51.440 141.310 ;
        RECT 54.430 141.295 54.570 141.450 ;
        RECT 55.720 141.390 56.040 141.450 ;
        RECT 47.900 141.110 51.440 141.250 ;
        RECT 47.900 141.050 48.220 141.110 ;
        RECT 50.215 141.065 50.505 141.110 ;
        RECT 51.120 141.050 51.440 141.110 ;
        RECT 51.670 141.110 54.110 141.250 ;
        RECT 17.540 140.710 17.860 140.970 ;
        RECT 18.435 140.910 18.725 140.955 ;
        RECT 19.625 140.910 19.915 140.955 ;
        RECT 22.145 140.910 22.435 140.955 ;
        RECT 18.435 140.770 22.435 140.910 ;
        RECT 18.435 140.725 18.725 140.770 ;
        RECT 19.625 140.725 19.915 140.770 ;
        RECT 22.145 140.725 22.435 140.770 ;
        RECT 29.985 140.910 30.275 140.955 ;
        RECT 32.505 140.910 32.795 140.955 ;
        RECT 33.695 140.910 33.985 140.955 ;
        RECT 38.240 140.910 38.560 140.970 ;
        RECT 40.555 140.910 40.845 140.955 ;
        RECT 29.985 140.770 33.985 140.910 ;
        RECT 29.985 140.725 30.275 140.770 ;
        RECT 32.505 140.725 32.795 140.770 ;
        RECT 33.695 140.725 33.985 140.770 ;
        RECT 35.570 140.770 40.845 140.910 ;
        RECT 17.630 140.570 17.770 140.710 ;
        RECT 35.570 140.630 35.710 140.770 ;
        RECT 38.240 140.710 38.560 140.770 ;
        RECT 40.555 140.725 40.845 140.770 ;
        RECT 41.435 140.910 41.725 140.955 ;
        RECT 42.625 140.910 42.915 140.955 ;
        RECT 45.145 140.910 45.435 140.955 ;
        RECT 49.740 140.910 50.060 140.970 ;
        RECT 51.670 140.910 51.810 141.110 ;
        RECT 41.435 140.770 45.435 140.910 ;
        RECT 41.435 140.725 41.725 140.770 ;
        RECT 42.625 140.725 42.915 140.770 ;
        RECT 45.145 140.725 45.435 140.770 ;
        RECT 48.450 140.770 50.060 140.910 ;
        RECT 21.680 140.570 22.000 140.630 ;
        RECT 29.500 140.570 29.820 140.630 ;
        RECT 17.630 140.430 29.820 140.570 ;
        RECT 21.680 140.370 22.000 140.430 ;
        RECT 29.500 140.370 29.820 140.430 ;
        RECT 34.575 140.570 34.865 140.615 ;
        RECT 35.480 140.570 35.800 140.630 ;
        RECT 34.575 140.430 35.800 140.570 ;
        RECT 34.575 140.385 34.865 140.430 ;
        RECT 35.480 140.370 35.800 140.430 ;
        RECT 37.780 140.370 38.100 140.630 ;
        RECT 18.890 140.230 19.180 140.275 ;
        RECT 19.840 140.230 20.160 140.290 ;
        RECT 18.890 140.090 20.160 140.230 ;
        RECT 18.890 140.045 19.180 140.090 ;
        RECT 19.840 140.030 20.160 140.090 ;
        RECT 23.980 140.230 24.300 140.290 ;
        RECT 26.295 140.230 26.585 140.275 ;
        RECT 23.980 140.090 26.585 140.230 ;
        RECT 23.980 140.030 24.300 140.090 ;
        RECT 26.295 140.045 26.585 140.090 ;
        RECT 33.350 140.230 33.640 140.275 ;
        RECT 35.035 140.230 35.325 140.275 ;
        RECT 33.350 140.090 35.325 140.230 ;
        RECT 33.350 140.045 33.640 140.090 ;
        RECT 35.035 140.045 35.325 140.090 ;
        RECT 41.890 140.230 42.180 140.275 ;
        RECT 43.760 140.230 44.080 140.290 ;
        RECT 48.450 140.275 48.590 140.770 ;
        RECT 49.740 140.710 50.060 140.770 ;
        RECT 50.750 140.770 51.810 140.910 ;
        RECT 53.970 140.910 54.110 141.110 ;
        RECT 54.355 141.065 54.645 141.295 ;
        RECT 54.800 141.050 55.120 141.310 ;
        RECT 100.010 141.150 100.880 144.420 ;
        RECT 104.530 143.960 109.780 143.970 ;
        RECT 104.530 143.850 116.840 143.960 ;
        RECT 101.560 143.790 116.840 143.850 ;
        RECT 101.560 143.780 116.875 143.790 ;
        RECT 101.500 143.650 116.875 143.780 ;
        RECT 101.500 143.640 106.660 143.650 ;
        RECT 101.500 143.550 105.500 143.640 ;
        RECT 108.875 143.560 116.875 143.650 ;
        RECT 108.960 143.550 116.850 143.560 ;
        RECT 101.110 143.190 101.340 143.500 ;
        RECT 101.560 143.190 105.460 143.550 ;
        RECT 105.660 143.190 105.890 143.500 ;
        RECT 101.110 141.850 105.890 143.190 ;
        RECT 101.110 141.540 101.340 141.850 ;
        RECT 105.660 141.540 105.890 141.850 ;
        RECT 108.440 142.970 108.670 143.510 ;
        RECT 109.480 142.970 110.490 143.000 ;
        RECT 117.080 142.970 117.310 143.510 ;
        RECT 108.440 142.070 117.310 142.970 ;
        RECT 108.440 141.550 108.670 142.070 ;
        RECT 109.480 142.000 110.490 142.070 ;
        RECT 117.080 141.550 117.310 142.070 ;
        RECT 101.500 141.260 105.500 141.490 ;
        RECT 108.875 141.270 116.875 141.500 ;
        RECT 100.010 141.110 101.180 141.150 ;
        RECT 100.010 141.030 101.420 141.110 ;
        RECT 101.790 141.040 105.450 141.260 ;
        RECT 101.790 141.030 103.230 141.040 ;
        RECT 100.010 140.990 103.230 141.030 ;
        RECT 53.970 140.770 56.410 140.910 ;
        RECT 49.280 140.275 49.600 140.290 ;
        RECT 41.890 140.090 44.080 140.230 ;
        RECT 41.890 140.045 42.180 140.090 ;
        RECT 43.760 140.030 44.080 140.090 ;
        RECT 48.375 140.045 48.665 140.275 ;
        RECT 49.280 140.230 49.745 140.275 ;
        RECT 50.750 140.230 50.890 140.770 ;
        RECT 51.135 140.385 51.425 140.615 ;
        RECT 52.040 140.570 52.360 140.630 ;
        RECT 52.515 140.570 52.805 140.615 ;
        RECT 52.960 140.570 53.280 140.630 ;
        RECT 56.270 140.615 56.410 140.770 ;
        RECT 57.100 140.710 57.420 140.970 ;
        RECT 60.320 140.910 60.640 140.970 ;
        RECT 63.095 140.910 63.385 140.955 ;
        RECT 57.650 140.770 63.385 140.910 ;
        RECT 52.040 140.430 53.280 140.570 ;
        RECT 49.280 140.090 50.890 140.230 ;
        RECT 49.280 140.045 49.745 140.090 ;
        RECT 49.280 140.030 49.600 140.045 ;
        RECT 21.220 139.890 21.540 139.950 ;
        RECT 26.740 139.890 27.060 139.950 ;
        RECT 21.220 139.750 27.060 139.890 ;
        RECT 21.220 139.690 21.540 139.750 ;
        RECT 26.740 139.690 27.060 139.750 ;
        RECT 27.675 139.890 27.965 139.935 ;
        RECT 30.420 139.890 30.740 139.950 ;
        RECT 27.675 139.750 30.740 139.890 ;
        RECT 27.675 139.705 27.965 139.750 ;
        RECT 30.420 139.690 30.740 139.750 ;
        RECT 47.440 139.890 47.760 139.950 ;
        RECT 51.210 139.890 51.350 140.385 ;
        RECT 52.040 140.370 52.360 140.430 ;
        RECT 52.515 140.385 52.805 140.430 ;
        RECT 52.960 140.370 53.280 140.430 ;
        RECT 56.195 140.570 56.485 140.615 ;
        RECT 57.650 140.570 57.790 140.770 ;
        RECT 60.320 140.710 60.640 140.770 ;
        RECT 63.095 140.725 63.385 140.770 ;
        RECT 100.010 140.900 102.740 140.990 ;
        RECT 108.940 140.980 116.830 141.270 ;
        RECT 100.010 140.840 102.070 140.900 ;
        RECT 100.010 140.790 101.820 140.840 ;
        RECT 56.195 140.430 57.790 140.570 ;
        RECT 62.160 140.570 62.480 140.630 ;
        RECT 64.920 140.570 65.240 140.630 ;
        RECT 65.855 140.570 66.145 140.615 ;
        RECT 62.160 140.430 66.145 140.570 ;
        RECT 56.195 140.385 56.485 140.430 ;
        RECT 62.160 140.370 62.480 140.430 ;
        RECT 64.920 140.370 65.240 140.430 ;
        RECT 65.855 140.385 66.145 140.430 ;
        RECT 51.580 140.230 51.900 140.290 ;
        RECT 53.560 140.230 53.850 140.275 ;
        RECT 51.580 140.090 53.850 140.230 ;
        RECT 51.580 140.030 51.900 140.090 ;
        RECT 53.560 140.045 53.850 140.090 ;
        RECT 54.340 140.230 54.660 140.290 ;
        RECT 54.815 140.230 55.105 140.275 ;
        RECT 54.340 140.090 55.105 140.230 ;
        RECT 54.340 140.030 54.660 140.090 ;
        RECT 54.815 140.045 55.105 140.090 ;
        RECT 57.560 140.230 57.880 140.290 ;
        RECT 61.255 140.230 61.545 140.275 ;
        RECT 63.540 140.230 63.860 140.290 ;
        RECT 57.560 140.090 63.860 140.230 ;
        RECT 57.560 140.030 57.880 140.090 ;
        RECT 61.255 140.045 61.545 140.090 ;
        RECT 63.540 140.030 63.860 140.090 ;
        RECT 64.015 140.230 64.305 140.275 ;
        RECT 65.380 140.230 65.700 140.290 ;
        RECT 67.680 140.230 68.000 140.290 ;
        RECT 64.015 140.090 68.000 140.230 ;
        RECT 64.015 140.045 64.305 140.090 ;
        RECT 65.380 140.030 65.700 140.090 ;
        RECT 67.680 140.030 68.000 140.090 ;
        RECT 47.440 139.750 51.350 139.890 ;
        RECT 47.440 139.690 47.760 139.750 ;
        RECT 52.960 139.690 53.280 139.950 ;
        RECT 55.260 139.890 55.580 139.950 ;
        RECT 55.735 139.890 56.025 139.935 ;
        RECT 59.400 139.890 59.720 139.950 ;
        RECT 55.260 139.750 59.720 139.890 ;
        RECT 55.260 139.690 55.580 139.750 ;
        RECT 55.735 139.705 56.025 139.750 ;
        RECT 59.400 139.690 59.720 139.750 ;
        RECT 64.460 139.690 64.780 139.950 ;
        RECT 64.935 139.890 65.225 139.935 ;
        RECT 66.760 139.890 67.080 139.950 ;
        RECT 64.935 139.750 67.080 139.890 ;
        RECT 64.935 139.705 65.225 139.750 ;
        RECT 66.760 139.690 67.080 139.750 ;
        RECT 11.950 139.070 90.610 139.550 ;
        RECT 19.840 138.670 20.160 138.930 ;
        RECT 20.775 138.870 21.065 138.915 ;
        RECT 21.220 138.870 21.540 138.930 ;
        RECT 20.775 138.730 21.540 138.870 ;
        RECT 20.775 138.685 21.065 138.730 ;
        RECT 21.220 138.670 21.540 138.730 ;
        RECT 26.295 138.870 26.585 138.915 ;
        RECT 27.755 138.870 28.045 138.915 ;
        RECT 26.295 138.730 28.045 138.870 ;
        RECT 26.295 138.685 26.585 138.730 ;
        RECT 27.755 138.685 28.045 138.730 ;
        RECT 28.595 138.685 28.885 138.915 ;
        RECT 43.760 138.870 44.080 138.930 ;
        RECT 44.235 138.870 44.525 138.915 ;
        RECT 43.760 138.730 44.525 138.870 ;
        RECT 24.440 138.530 24.760 138.590 ;
        RECT 22.690 138.390 24.760 138.530 ;
        RECT 22.690 138.235 22.830 138.390 ;
        RECT 24.440 138.330 24.760 138.390 ;
        RECT 26.740 138.330 27.060 138.590 ;
        RECT 28.670 138.530 28.810 138.685 ;
        RECT 43.760 138.670 44.080 138.730 ;
        RECT 44.235 138.685 44.525 138.730 ;
        RECT 45.600 138.670 45.920 138.930 ;
        RECT 46.060 138.670 46.380 138.930 ;
        RECT 47.915 138.870 48.205 138.915 ;
        RECT 48.360 138.870 48.680 138.930 ;
        RECT 47.915 138.730 48.680 138.870 ;
        RECT 47.915 138.685 48.205 138.730 ;
        RECT 48.360 138.670 48.680 138.730 ;
        RECT 48.820 138.870 49.140 138.930 ;
        RECT 49.755 138.870 50.045 138.915 ;
        RECT 48.820 138.730 50.045 138.870 ;
        RECT 48.820 138.670 49.140 138.730 ;
        RECT 49.755 138.685 50.045 138.730 ;
        RECT 51.580 138.670 51.900 138.930 ;
        RECT 58.480 138.870 58.800 138.930 ;
        RECT 69.520 138.870 69.840 138.930 ;
        RECT 70.455 138.870 70.745 138.915 ;
        RECT 58.480 138.730 70.745 138.870 ;
        RECT 58.480 138.670 58.800 138.730 ;
        RECT 69.520 138.670 69.840 138.730 ;
        RECT 70.455 138.685 70.745 138.730 ;
        RECT 71.835 138.685 72.125 138.915 ;
        RECT 30.280 138.530 30.570 138.575 ;
        RECT 28.670 138.390 30.570 138.530 ;
        RECT 30.280 138.345 30.570 138.390 ;
        RECT 34.100 138.530 34.420 138.590 ;
        RECT 39.175 138.530 39.465 138.575 ;
        RECT 57.560 138.530 57.880 138.590 ;
        RECT 34.100 138.390 57.880 138.530 ;
        RECT 34.100 138.330 34.420 138.390 ;
        RECT 39.175 138.345 39.465 138.390 ;
        RECT 57.560 138.330 57.880 138.390 ;
        RECT 59.860 138.530 60.180 138.590 ;
        RECT 68.600 138.530 68.920 138.590 ;
        RECT 69.980 138.530 70.300 138.590 ;
        RECT 59.860 138.390 70.300 138.530 ;
        RECT 71.910 138.530 72.050 138.685 ;
        RECT 77.860 138.530 78.150 138.575 ;
        RECT 71.910 138.390 78.150 138.530 ;
        RECT 59.860 138.330 60.180 138.390 ;
        RECT 68.600 138.330 68.920 138.390 ;
        RECT 69.980 138.330 70.300 138.390 ;
        RECT 77.860 138.345 78.150 138.390 ;
        RECT 14.795 138.190 15.085 138.235 ;
        RECT 14.795 138.050 20.300 138.190 ;
        RECT 14.795 138.005 15.085 138.050 ;
        RECT 20.160 137.850 20.300 138.050 ;
        RECT 22.615 138.005 22.905 138.235 ;
        RECT 25.360 138.190 25.680 138.250 ;
        RECT 29.055 138.190 29.345 138.235 ;
        RECT 29.500 138.190 29.820 138.250 ;
        RECT 25.360 138.050 28.810 138.190 ;
        RECT 25.360 137.990 25.680 138.050 ;
        RECT 26.740 137.850 27.060 137.910 ;
        RECT 20.160 137.710 27.060 137.850 ;
        RECT 26.740 137.650 27.060 137.710 ;
        RECT 24.900 137.510 25.220 137.570 ;
        RECT 24.900 137.370 27.890 137.510 ;
        RECT 24.900 137.310 25.220 137.370 ;
        RECT 10.640 137.170 10.960 137.230 ;
        RECT 13.875 137.170 14.165 137.215 ;
        RECT 10.640 137.030 14.165 137.170 ;
        RECT 10.640 136.970 10.960 137.030 ;
        RECT 13.875 136.985 14.165 137.030 ;
        RECT 20.775 137.170 21.065 137.215 ;
        RECT 25.820 137.170 26.140 137.230 ;
        RECT 27.750 137.215 27.890 137.370 ;
        RECT 20.775 137.030 26.140 137.170 ;
        RECT 20.775 136.985 21.065 137.030 ;
        RECT 25.820 136.970 26.140 137.030 ;
        RECT 27.675 136.985 27.965 137.215 ;
        RECT 28.670 137.170 28.810 138.050 ;
        RECT 29.055 138.050 29.820 138.190 ;
        RECT 29.055 138.005 29.345 138.050 ;
        RECT 29.500 137.990 29.820 138.050 ;
        RECT 44.220 138.190 44.540 138.250 ;
        RECT 45.030 138.190 45.320 138.235 ;
        RECT 44.220 138.050 45.320 138.190 ;
        RECT 44.220 137.990 44.540 138.050 ;
        RECT 45.030 138.005 45.320 138.050 ;
        RECT 48.820 137.990 49.140 138.250 ;
        RECT 49.295 138.005 49.585 138.235 ;
        RECT 49.740 138.190 50.060 138.250 ;
        RECT 50.675 138.190 50.965 138.235 ;
        RECT 49.740 138.050 50.965 138.190 ;
        RECT 29.935 137.850 30.225 137.895 ;
        RECT 31.125 137.850 31.415 137.895 ;
        RECT 33.645 137.850 33.935 137.895 ;
        RECT 29.935 137.710 33.935 137.850 ;
        RECT 29.935 137.665 30.225 137.710 ;
        RECT 31.125 137.665 31.415 137.710 ;
        RECT 33.645 137.665 33.935 137.710 ;
        RECT 35.480 137.850 35.800 137.910 ;
        RECT 42.855 137.850 43.145 137.895 ;
        RECT 35.480 137.710 43.145 137.850 ;
        RECT 35.480 137.650 35.800 137.710 ;
        RECT 42.855 137.665 43.145 137.710 ;
        RECT 47.440 137.650 47.760 137.910 ;
        RECT 49.370 137.850 49.510 138.005 ;
        RECT 49.740 137.990 50.060 138.050 ;
        RECT 50.675 138.005 50.965 138.050 ;
        RECT 50.750 137.850 50.890 138.005 ;
        RECT 51.120 137.990 51.440 138.250 ;
        RECT 52.055 138.190 52.345 138.235 ;
        RECT 54.800 138.190 55.120 138.250 ;
        RECT 52.055 138.050 55.120 138.190 ;
        RECT 52.055 138.005 52.345 138.050 ;
        RECT 54.800 137.990 55.120 138.050 ;
        RECT 57.100 137.990 57.420 138.250 ;
        RECT 64.460 138.190 64.780 138.250 ;
        RECT 65.855 138.190 66.145 138.235 ;
        RECT 64.460 138.050 66.145 138.190 ;
        RECT 64.460 137.990 64.780 138.050 ;
        RECT 65.855 138.005 66.145 138.050 ;
        RECT 66.760 137.990 67.080 138.250 ;
        RECT 75.500 138.190 75.820 138.250 ;
        RECT 67.310 138.050 75.820 138.190 ;
        RECT 54.340 137.850 54.660 137.910 ;
        RECT 67.310 137.850 67.450 138.050 ;
        RECT 75.500 137.990 75.820 138.050 ;
        RECT 75.960 138.190 76.280 138.250 ;
        RECT 79.195 138.190 79.485 138.235 ;
        RECT 75.960 138.050 79.485 138.190 ;
        RECT 75.960 137.990 76.280 138.050 ;
        RECT 79.195 138.005 79.485 138.050 ;
        RECT 49.370 137.710 49.970 137.850 ;
        RECT 50.750 137.710 54.660 137.850 ;
        RECT 29.540 137.510 29.830 137.555 ;
        RECT 31.640 137.510 31.930 137.555 ;
        RECT 33.210 137.510 33.500 137.555 ;
        RECT 29.540 137.370 33.500 137.510 ;
        RECT 29.540 137.325 29.830 137.370 ;
        RECT 31.640 137.325 31.930 137.370 ;
        RECT 33.210 137.325 33.500 137.370 ;
        RECT 35.955 137.170 36.245 137.215 ;
        RECT 28.670 137.030 36.245 137.170 ;
        RECT 35.955 136.985 36.245 137.030 ;
        RECT 48.360 137.170 48.680 137.230 ;
        RECT 49.830 137.170 49.970 137.710 ;
        RECT 54.340 137.650 54.660 137.710 ;
        RECT 54.890 137.710 67.450 137.850 ;
        RECT 52.040 137.510 52.360 137.570 ;
        RECT 54.890 137.510 55.030 137.710 ;
        RECT 68.600 137.650 68.920 137.910 ;
        RECT 69.980 137.650 70.300 137.910 ;
        RECT 71.040 137.850 71.330 137.895 ;
        RECT 71.820 137.850 72.140 137.910 ;
        RECT 71.040 137.710 72.140 137.850 ;
        RECT 71.040 137.665 71.330 137.710 ;
        RECT 71.820 137.650 72.140 137.710 ;
        RECT 74.605 137.850 74.895 137.895 ;
        RECT 77.125 137.850 77.415 137.895 ;
        RECT 78.315 137.850 78.605 137.895 ;
        RECT 74.605 137.710 78.605 137.850 ;
        RECT 74.605 137.665 74.895 137.710 ;
        RECT 77.125 137.665 77.415 137.710 ;
        RECT 78.315 137.665 78.605 137.710 ;
        RECT 52.040 137.370 55.030 137.510 ;
        RECT 64.920 137.510 65.240 137.570 ;
        RECT 72.295 137.510 72.585 137.555 ;
        RECT 64.920 137.370 72.585 137.510 ;
        RECT 52.040 137.310 52.360 137.370 ;
        RECT 64.920 137.310 65.240 137.370 ;
        RECT 72.295 137.325 72.585 137.370 ;
        RECT 75.040 137.510 75.330 137.555 ;
        RECT 76.610 137.510 76.900 137.555 ;
        RECT 78.710 137.510 79.000 137.555 ;
        RECT 75.040 137.370 79.000 137.510 ;
        RECT 75.040 137.325 75.330 137.370 ;
        RECT 76.610 137.325 76.900 137.370 ;
        RECT 78.710 137.325 79.000 137.370 ;
        RECT 100.010 137.450 100.880 140.790 ;
        RECT 108.930 140.490 116.850 140.500 ;
        RECT 105.160 140.480 116.850 140.490 ;
        RECT 101.540 140.360 116.850 140.480 ;
        RECT 101.540 140.350 116.875 140.360 ;
        RECT 101.500 140.230 116.875 140.350 ;
        RECT 101.500 140.120 105.500 140.230 ;
        RECT 101.110 139.780 101.340 140.070 ;
        RECT 101.560 139.780 105.450 140.120 ;
        RECT 105.660 139.780 105.890 140.070 ;
        RECT 101.110 138.410 105.890 139.780 ;
        RECT 101.110 138.110 101.340 138.410 ;
        RECT 105.660 138.110 105.890 138.410 ;
        RECT 101.500 137.830 105.500 138.060 ;
        RECT 101.750 137.600 105.320 137.830 ;
        RECT 101.750 137.450 105.440 137.600 ;
        RECT 55.260 137.170 55.580 137.230 ;
        RECT 48.360 137.030 55.580 137.170 ;
        RECT 48.360 136.970 48.680 137.030 ;
        RECT 55.260 136.970 55.580 137.030 ;
        RECT 66.775 137.170 67.065 137.215 ;
        RECT 67.220 137.170 67.540 137.230 ;
        RECT 66.775 137.030 67.540 137.170 ;
        RECT 66.775 136.985 67.065 137.030 ;
        RECT 67.220 136.970 67.540 137.030 ;
        RECT 100.010 137.170 105.440 137.450 ;
        RECT 106.690 137.280 107.310 140.230 ;
        RECT 108.875 140.130 116.875 140.230 ;
        RECT 108.930 140.120 116.850 140.130 ;
        RECT 108.440 139.420 108.670 140.080 ;
        RECT 109.450 139.420 110.450 139.510 ;
        RECT 117.080 139.420 117.310 140.080 ;
        RECT 108.440 138.600 117.310 139.420 ;
        RECT 108.440 138.120 108.670 138.600 ;
        RECT 109.450 138.510 110.450 138.600 ;
        RECT 117.080 138.120 117.310 138.600 ;
        RECT 108.875 137.840 116.875 138.070 ;
        RECT 11.950 136.350 90.610 136.830 ;
        RECT 100.010 136.710 105.450 137.170 ;
        RECT 41.460 136.150 41.780 136.210 ;
        RECT 45.600 136.150 45.920 136.210 ;
        RECT 52.960 136.150 53.280 136.210 ;
        RECT 41.460 136.010 53.280 136.150 ;
        RECT 41.460 135.950 41.780 136.010 ;
        RECT 45.600 135.950 45.920 136.010 ;
        RECT 52.960 135.950 53.280 136.010 ;
        RECT 64.460 135.950 64.780 136.210 ;
        RECT 64.920 136.150 65.240 136.210 ;
        RECT 65.395 136.150 65.685 136.195 ;
        RECT 64.920 136.010 65.685 136.150 ;
        RECT 64.920 135.950 65.240 136.010 ;
        RECT 65.395 135.965 65.685 136.010 ;
        RECT 32.720 135.610 33.040 135.870 ;
        RECT 37.360 135.810 37.650 135.855 ;
        RECT 39.460 135.810 39.750 135.855 ;
        RECT 41.030 135.810 41.320 135.855 ;
        RECT 63.540 135.810 63.860 135.870 ;
        RECT 37.360 135.670 41.320 135.810 ;
        RECT 37.360 135.625 37.650 135.670 ;
        RECT 39.460 135.625 39.750 135.670 ;
        RECT 41.030 135.625 41.320 135.670 ;
        RECT 58.110 135.670 63.860 135.810 ;
        RECT 58.110 135.530 58.250 135.670 ;
        RECT 63.540 135.610 63.860 135.670 ;
        RECT 37.755 135.470 38.045 135.515 ;
        RECT 38.945 135.470 39.235 135.515 ;
        RECT 41.465 135.470 41.755 135.515 ;
        RECT 37.755 135.330 41.755 135.470 ;
        RECT 37.755 135.285 38.045 135.330 ;
        RECT 38.945 135.285 39.235 135.330 ;
        RECT 41.465 135.285 41.755 135.330 ;
        RECT 47.440 135.470 47.760 135.530 ;
        RECT 51.135 135.470 51.425 135.515 ;
        RECT 47.440 135.330 56.870 135.470 ;
        RECT 47.440 135.270 47.760 135.330 ;
        RECT 51.135 135.285 51.425 135.330 ;
        RECT 29.500 135.130 29.820 135.190 ;
        RECT 29.975 135.130 30.265 135.175 ;
        RECT 29.500 134.990 30.265 135.130 ;
        RECT 29.500 134.930 29.820 134.990 ;
        RECT 29.975 134.945 30.265 134.990 ;
        RECT 30.420 135.130 30.740 135.190 ;
        RECT 34.115 135.130 34.405 135.175 ;
        RECT 30.420 134.990 34.405 135.130 ;
        RECT 30.420 134.930 30.740 134.990 ;
        RECT 34.115 134.945 34.405 134.990 ;
        RECT 35.480 135.130 35.800 135.190 ;
        RECT 36.875 135.130 37.165 135.175 ;
        RECT 41.000 135.130 41.320 135.190 ;
        RECT 35.480 134.990 37.165 135.130 ;
        RECT 35.480 134.930 35.800 134.990 ;
        RECT 36.875 134.945 37.165 134.990 ;
        RECT 37.410 134.990 41.320 135.130 ;
        RECT 32.735 134.790 33.025 134.835 ;
        RECT 33.180 134.790 33.500 134.850 ;
        RECT 32.735 134.650 33.500 134.790 ;
        RECT 32.735 134.605 33.025 134.650 ;
        RECT 33.180 134.590 33.500 134.650 ;
        RECT 33.655 134.790 33.945 134.835 ;
        RECT 37.410 134.790 37.550 134.990 ;
        RECT 41.000 134.930 41.320 134.990 ;
        RECT 52.040 134.930 52.360 135.190 ;
        RECT 56.730 135.175 56.870 135.330 ;
        RECT 58.020 135.270 58.340 135.530 ;
        RECT 58.480 135.270 58.800 135.530 ;
        RECT 56.655 135.130 56.945 135.175 ;
        RECT 59.860 135.130 60.180 135.190 ;
        RECT 56.655 134.990 60.180 135.130 ;
        RECT 56.655 134.945 56.945 134.990 ;
        RECT 59.860 134.930 60.180 134.990 ;
        RECT 60.320 134.930 60.640 135.190 ;
        RECT 61.255 134.945 61.545 135.175 ;
        RECT 38.240 134.835 38.560 134.850 ;
        RECT 33.655 134.650 37.550 134.790 ;
        RECT 33.655 134.605 33.945 134.650 ;
        RECT 38.210 134.605 38.560 134.835 ;
        RECT 59.080 134.790 59.370 134.835 ;
        RECT 60.795 134.790 61.085 134.835 ;
        RECT 59.080 134.650 61.085 134.790 ;
        RECT 61.330 134.790 61.470 134.945 ;
        RECT 62.160 134.930 62.480 135.190 ;
        RECT 63.095 135.130 63.385 135.175 ;
        RECT 64.550 135.130 64.690 135.950 ;
        RECT 65.470 135.470 65.610 135.965 ;
        RECT 66.760 135.950 67.080 136.210 ;
        RECT 67.680 136.150 68.000 136.210 ;
        RECT 71.820 136.150 72.140 136.210 ;
        RECT 72.295 136.150 72.585 136.195 ;
        RECT 67.680 136.010 68.600 136.150 ;
        RECT 67.680 135.950 68.000 136.010 ;
        RECT 68.460 135.470 68.600 136.010 ;
        RECT 71.820 136.010 72.585 136.150 ;
        RECT 71.820 135.950 72.140 136.010 ;
        RECT 72.295 135.965 72.585 136.010 ;
        RECT 69.995 135.470 70.285 135.515 ;
        RECT 65.470 135.330 67.450 135.470 ;
        RECT 63.095 134.990 64.690 135.130 ;
        RECT 67.310 135.130 67.450 135.330 ;
        RECT 68.230 135.330 70.285 135.470 ;
        RECT 68.230 135.175 68.370 135.330 ;
        RECT 69.995 135.285 70.285 135.330 ;
        RECT 100.010 135.360 102.050 136.710 ;
        RECT 103.800 136.700 105.450 136.710 ;
        RECT 102.490 135.430 103.490 136.150 ;
        RECT 103.800 135.890 104.110 136.700 ;
        RECT 104.570 136.420 105.450 136.700 ;
        RECT 105.690 136.880 107.310 137.280 ;
        RECT 108.960 136.930 116.830 137.840 ;
        RECT 104.510 136.190 105.510 136.420 ;
        RECT 105.690 136.230 106.040 136.880 ;
        RECT 106.690 136.870 107.310 136.880 ;
        RECT 108.875 136.700 116.875 136.930 ;
        RECT 108.960 136.690 116.830 136.700 ;
        RECT 104.570 135.980 105.450 136.000 ;
        RECT 103.840 135.600 104.110 135.890 ;
        RECT 104.510 135.750 105.510 135.980 ;
        RECT 105.670 135.940 106.040 136.230 ;
        RECT 105.700 135.880 106.040 135.940 ;
        RECT 106.800 136.550 107.560 136.600 ;
        RECT 108.440 136.550 108.670 136.650 ;
        RECT 106.800 136.340 108.670 136.550 ;
        RECT 117.080 136.340 117.310 136.650 ;
        RECT 106.800 135.920 109.340 136.340 ;
        RECT 116.710 135.920 117.310 136.340 ;
        RECT 104.570 135.600 105.450 135.750 ;
        RECT 104.580 135.430 105.310 135.600 ;
        RECT 67.695 135.130 67.985 135.175 ;
        RECT 67.310 134.990 67.985 135.130 ;
        RECT 63.095 134.945 63.385 134.990 ;
        RECT 67.695 134.945 67.985 134.990 ;
        RECT 68.155 134.945 68.445 135.175 ;
        RECT 70.455 134.945 70.745 135.175 ;
        RECT 65.380 134.835 65.700 134.850 ;
        RECT 62.635 134.790 62.925 134.835 ;
        RECT 61.330 134.650 62.925 134.790 ;
        RECT 59.080 134.605 59.370 134.650 ;
        RECT 60.795 134.605 61.085 134.650 ;
        RECT 62.635 134.605 62.925 134.650 ;
        RECT 65.315 134.605 65.700 134.835 ;
        RECT 27.660 134.450 27.980 134.510 ;
        RECT 33.730 134.450 33.870 134.605 ;
        RECT 38.240 134.590 38.560 134.605 ;
        RECT 65.380 134.590 65.700 134.605 ;
        RECT 66.300 134.790 66.620 134.850 ;
        RECT 66.775 134.790 67.065 134.835 ;
        RECT 66.300 134.650 67.065 134.790 ;
        RECT 67.770 134.790 67.910 134.945 ;
        RECT 70.530 134.790 70.670 134.945 ;
        RECT 67.770 134.650 70.670 134.790 ;
        RECT 66.300 134.590 66.620 134.650 ;
        RECT 66.775 134.605 67.065 134.650 ;
        RECT 27.660 134.310 33.870 134.450 ;
        RECT 43.775 134.450 44.065 134.495 ;
        RECT 46.060 134.450 46.380 134.510 ;
        RECT 43.775 134.310 46.380 134.450 ;
        RECT 27.660 134.250 27.980 134.310 ;
        RECT 43.775 134.265 44.065 134.310 ;
        RECT 46.060 134.250 46.380 134.310 ;
        RECT 59.860 134.250 60.180 134.510 ;
        RECT 11.950 133.630 90.610 134.110 ;
        RECT 23.980 133.430 24.300 133.490 ;
        RECT 25.835 133.430 26.125 133.475 ;
        RECT 23.980 133.290 26.125 133.430 ;
        RECT 23.980 133.230 24.300 133.290 ;
        RECT 25.835 133.245 26.125 133.290 ;
        RECT 26.755 133.430 27.045 133.475 ;
        RECT 29.960 133.430 30.280 133.490 ;
        RECT 26.755 133.290 30.280 133.430 ;
        RECT 26.755 133.245 27.045 133.290 ;
        RECT 29.960 133.230 30.280 133.290 ;
        RECT 39.175 133.430 39.465 133.475 ;
        RECT 52.515 133.430 52.805 133.475 ;
        RECT 52.960 133.430 53.280 133.490 ;
        RECT 39.175 133.290 48.590 133.430 ;
        RECT 39.175 133.245 39.465 133.290 ;
        RECT 38.255 133.090 38.545 133.135 ;
        RECT 47.440 133.090 47.760 133.150 ;
        RECT 38.255 132.950 47.760 133.090 ;
        RECT 48.450 133.090 48.590 133.290 ;
        RECT 52.515 133.290 53.280 133.430 ;
        RECT 52.515 133.245 52.805 133.290 ;
        RECT 52.960 133.230 53.280 133.290 ;
        RECT 62.160 133.430 62.480 133.490 ;
        RECT 63.095 133.430 63.385 133.475 ;
        RECT 62.160 133.290 63.385 133.430 ;
        RECT 62.160 133.230 62.480 133.290 ;
        RECT 63.095 133.245 63.385 133.290 ;
        RECT 66.300 133.430 66.620 133.490 ;
        RECT 71.835 133.430 72.125 133.475 ;
        RECT 66.300 133.290 72.125 133.430 ;
        RECT 66.300 133.230 66.620 133.290 ;
        RECT 71.835 133.245 72.125 133.290 ;
        RECT 51.580 133.090 51.900 133.150 ;
        RECT 52.055 133.090 52.345 133.135 ;
        RECT 48.450 132.950 52.345 133.090 ;
        RECT 38.255 132.905 38.545 132.950 ;
        RECT 47.440 132.890 47.760 132.950 ;
        RECT 51.580 132.890 51.900 132.950 ;
        RECT 52.055 132.905 52.345 132.950 ;
        RECT 57.530 133.090 57.820 133.135 ;
        RECT 59.860 133.090 60.180 133.150 ;
        RECT 68.140 133.090 68.460 133.150 ;
        RECT 72.740 133.090 73.060 133.150 ;
        RECT 75.040 133.090 75.360 133.150 ;
        RECT 57.530 132.950 60.180 133.090 ;
        RECT 57.530 132.905 57.820 132.950 ;
        RECT 59.860 132.890 60.180 132.950 ;
        RECT 65.010 132.950 75.360 133.090 ;
        RECT 39.635 132.750 39.925 132.795 ;
        RECT 41.460 132.750 41.780 132.810 ;
        RECT 39.635 132.610 41.780 132.750 ;
        RECT 39.635 132.565 39.925 132.610 ;
        RECT 41.460 132.550 41.780 132.610 ;
        RECT 45.155 132.750 45.445 132.795 ;
        RECT 45.600 132.750 45.920 132.810 ;
        RECT 45.155 132.610 45.920 132.750 ;
        RECT 45.155 132.565 45.445 132.610 ;
        RECT 45.600 132.550 45.920 132.610 ;
        RECT 46.060 132.550 46.380 132.810 ;
        RECT 48.360 132.550 48.680 132.810 ;
        RECT 53.100 132.750 53.390 132.795 ;
        RECT 50.290 132.610 53.390 132.750 ;
        RECT 28.595 132.410 28.885 132.455 ;
        RECT 29.500 132.410 29.820 132.470 ;
        RECT 28.595 132.270 29.820 132.410 ;
        RECT 28.595 132.225 28.885 132.270 ;
        RECT 29.500 132.210 29.820 132.270 ;
        RECT 34.560 132.210 34.880 132.470 ;
        RECT 44.695 132.410 44.985 132.455 ;
        RECT 46.150 132.410 46.290 132.550 ;
        RECT 44.695 132.270 46.290 132.410 ;
        RECT 44.695 132.225 44.985 132.270 ;
        RECT 48.820 132.210 49.140 132.470 ;
        RECT 50.290 132.455 50.430 132.610 ;
        RECT 53.100 132.565 53.390 132.610 ;
        RECT 56.195 132.750 56.485 132.795 ;
        RECT 56.640 132.750 56.960 132.810 ;
        RECT 65.010 132.795 65.150 132.950 ;
        RECT 68.140 132.890 68.460 132.950 ;
        RECT 72.740 132.890 73.060 132.950 ;
        RECT 75.040 132.890 75.360 132.950 ;
        RECT 66.300 132.795 66.620 132.810 ;
        RECT 56.195 132.610 56.960 132.750 ;
        RECT 56.195 132.565 56.485 132.610 ;
        RECT 56.640 132.550 56.960 132.610 ;
        RECT 64.935 132.565 65.225 132.795 ;
        RECT 66.270 132.565 66.620 132.795 ;
        RECT 66.300 132.550 66.620 132.565 ;
        RECT 50.215 132.225 50.505 132.455 ;
        RECT 50.675 132.225 50.965 132.455 ;
        RECT 57.075 132.410 57.365 132.455 ;
        RECT 58.265 132.410 58.555 132.455 ;
        RECT 60.785 132.410 61.075 132.455 ;
        RECT 57.075 132.270 61.075 132.410 ;
        RECT 57.075 132.225 57.365 132.270 ;
        RECT 58.265 132.225 58.555 132.270 ;
        RECT 60.785 132.225 61.075 132.270 ;
        RECT 65.815 132.410 66.105 132.455 ;
        RECT 67.005 132.410 67.295 132.455 ;
        RECT 69.525 132.410 69.815 132.455 ;
        RECT 65.815 132.270 69.815 132.410 ;
        RECT 65.815 132.225 66.105 132.270 ;
        RECT 67.005 132.225 67.295 132.270 ;
        RECT 69.525 132.225 69.815 132.270 ;
        RECT 38.240 131.870 38.560 132.130 ;
        RECT 47.440 132.070 47.760 132.130 ;
        RECT 50.750 132.070 50.890 132.225 ;
        RECT 47.440 131.930 50.890 132.070 ;
        RECT 56.680 132.070 56.970 132.115 ;
        RECT 58.780 132.070 59.070 132.115 ;
        RECT 60.350 132.070 60.640 132.115 ;
        RECT 56.680 131.930 60.640 132.070 ;
        RECT 47.440 131.870 47.760 131.930 ;
        RECT 56.680 131.885 56.970 131.930 ;
        RECT 58.780 131.885 59.070 131.930 ;
        RECT 60.350 131.885 60.640 131.930 ;
        RECT 65.420 132.070 65.710 132.115 ;
        RECT 67.520 132.070 67.810 132.115 ;
        RECT 69.090 132.070 69.380 132.115 ;
        RECT 65.420 131.930 69.380 132.070 ;
        RECT 65.420 131.885 65.710 131.930 ;
        RECT 67.520 131.885 67.810 131.930 ;
        RECT 69.090 131.885 69.380 131.930 ;
        RECT 26.755 131.730 27.045 131.775 ;
        RECT 27.660 131.730 27.980 131.790 ;
        RECT 26.755 131.590 27.980 131.730 ;
        RECT 26.755 131.545 27.045 131.590 ;
        RECT 27.660 131.530 27.980 131.590 ;
        RECT 29.960 131.730 30.280 131.790 ;
        RECT 32.735 131.730 33.025 131.775 ;
        RECT 33.180 131.730 33.500 131.790 ;
        RECT 29.960 131.590 33.500 131.730 ;
        RECT 29.960 131.530 30.280 131.590 ;
        RECT 32.735 131.545 33.025 131.590 ;
        RECT 33.180 131.530 33.500 131.590 ;
        RECT 36.400 131.730 36.720 131.790 ;
        RECT 37.335 131.730 37.625 131.775 ;
        RECT 36.400 131.590 37.625 131.730 ;
        RECT 36.400 131.530 36.720 131.590 ;
        RECT 37.335 131.545 37.625 131.590 ;
        RECT 41.460 131.530 41.780 131.790 ;
        RECT 44.220 131.730 44.540 131.790 ;
        RECT 45.615 131.730 45.905 131.775 ;
        RECT 44.220 131.590 45.905 131.730 ;
        RECT 44.220 131.530 44.540 131.590 ;
        RECT 45.615 131.545 45.905 131.590 ;
        RECT 53.880 131.530 54.200 131.790 ;
        RECT 100.010 131.720 100.780 135.360 ;
        RECT 102.460 134.310 105.310 135.430 ;
        RECT 105.700 135.130 106.050 135.880 ;
        RECT 106.800 135.760 108.670 135.920 ;
        RECT 106.800 135.710 107.560 135.760 ;
        RECT 108.440 135.690 108.670 135.760 ;
        RECT 117.080 135.690 117.310 135.920 ;
        RECT 108.875 135.410 116.875 135.640 ;
        RECT 105.700 135.070 105.990 135.130 ;
        RECT 105.610 134.950 105.990 135.070 ;
        RECT 108.970 135.010 116.830 135.410 ;
        RECT 117.640 135.010 118.600 144.490 ;
        RECT 119.930 144.620 120.770 146.750 ;
        RECT 126.430 146.330 127.680 146.770 ;
        RECT 137.600 146.750 138.460 148.920 ;
        RECT 124.370 146.320 129.610 146.330 ;
        RECT 121.420 146.220 136.720 146.320 ;
        RECT 121.420 146.210 136.755 146.220 ;
        RECT 121.380 146.090 136.755 146.210 ;
        RECT 121.380 145.980 125.380 146.090 ;
        RECT 126.430 146.010 128.170 146.090 ;
        RECT 128.750 146.010 136.755 146.090 ;
        RECT 126.430 145.930 127.680 146.010 ;
        RECT 128.755 145.990 136.755 146.010 ;
        RECT 120.990 145.680 121.220 145.930 ;
        RECT 125.540 145.790 125.770 145.930 ;
        RECT 128.320 145.790 128.550 145.940 ;
        RECT 125.540 145.680 128.550 145.790 ;
        RECT 136.960 145.680 137.190 145.940 ;
        RECT 120.990 145.240 137.190 145.680 ;
        RECT 120.990 144.970 121.220 145.240 ;
        RECT 125.540 145.210 137.190 145.240 ;
        RECT 125.540 145.120 128.550 145.210 ;
        RECT 125.540 144.970 125.770 145.120 ;
        RECT 128.320 144.980 128.550 145.120 ;
        RECT 136.960 144.980 137.190 145.210 ;
        RECT 121.380 144.690 125.380 144.920 ;
        RECT 128.755 144.710 136.755 144.930 ;
        RECT 137.520 144.710 138.480 146.750 ;
        RECT 128.755 144.700 138.480 144.710 ;
        RECT 121.380 144.620 125.370 144.690 ;
        RECT 119.930 144.510 125.370 144.620 ;
        RECT 128.810 144.540 138.480 144.700 ;
        RECT 119.930 144.420 123.060 144.510 ;
        RECT 136.550 144.490 138.480 144.540 ;
        RECT 119.930 141.150 120.770 144.420 ;
        RECT 124.410 143.960 129.660 143.970 ;
        RECT 124.410 143.850 136.720 143.960 ;
        RECT 121.440 143.790 136.720 143.850 ;
        RECT 121.440 143.780 136.755 143.790 ;
        RECT 121.380 143.650 136.755 143.780 ;
        RECT 121.380 143.640 126.540 143.650 ;
        RECT 121.380 143.550 125.380 143.640 ;
        RECT 128.755 143.560 136.755 143.650 ;
        RECT 128.840 143.550 136.730 143.560 ;
        RECT 120.990 143.190 121.220 143.500 ;
        RECT 121.440 143.190 125.340 143.550 ;
        RECT 125.540 143.190 125.770 143.500 ;
        RECT 120.990 141.850 125.770 143.190 ;
        RECT 120.990 141.540 121.220 141.850 ;
        RECT 125.540 141.540 125.770 141.850 ;
        RECT 128.320 142.970 128.550 143.510 ;
        RECT 129.360 142.970 130.370 143.000 ;
        RECT 136.960 142.970 137.190 143.510 ;
        RECT 128.320 142.070 137.190 142.970 ;
        RECT 128.320 141.550 128.550 142.070 ;
        RECT 129.360 142.000 130.370 142.070 ;
        RECT 136.960 141.550 137.190 142.070 ;
        RECT 121.380 141.260 125.380 141.490 ;
        RECT 128.755 141.270 136.755 141.500 ;
        RECT 119.930 141.110 121.060 141.150 ;
        RECT 119.930 141.030 121.300 141.110 ;
        RECT 121.670 141.040 125.330 141.260 ;
        RECT 121.670 141.030 123.110 141.040 ;
        RECT 119.930 140.990 123.110 141.030 ;
        RECT 119.930 140.900 122.620 140.990 ;
        RECT 128.820 140.980 136.710 141.270 ;
        RECT 119.930 140.840 121.950 140.900 ;
        RECT 119.930 140.790 121.700 140.840 ;
        RECT 119.930 137.450 120.770 140.790 ;
        RECT 128.810 140.490 136.730 140.500 ;
        RECT 125.040 140.480 136.730 140.490 ;
        RECT 121.420 140.360 136.730 140.480 ;
        RECT 121.420 140.350 136.755 140.360 ;
        RECT 121.380 140.230 136.755 140.350 ;
        RECT 121.380 140.120 125.380 140.230 ;
        RECT 120.990 139.780 121.220 140.070 ;
        RECT 121.440 139.780 125.330 140.120 ;
        RECT 125.540 139.780 125.770 140.070 ;
        RECT 120.990 138.410 125.770 139.780 ;
        RECT 120.990 138.110 121.220 138.410 ;
        RECT 125.540 138.110 125.770 138.410 ;
        RECT 121.380 137.830 125.380 138.060 ;
        RECT 121.630 137.600 125.200 137.830 ;
        RECT 121.630 137.450 125.320 137.600 ;
        RECT 119.930 137.170 125.320 137.450 ;
        RECT 126.570 137.280 127.190 140.230 ;
        RECT 128.755 140.130 136.755 140.230 ;
        RECT 128.810 140.120 136.730 140.130 ;
        RECT 128.320 139.420 128.550 140.080 ;
        RECT 129.330 139.420 130.330 139.510 ;
        RECT 136.960 139.420 137.190 140.080 ;
        RECT 128.320 138.600 137.190 139.420 ;
        RECT 128.320 138.120 128.550 138.600 ;
        RECT 129.330 138.510 130.330 138.600 ;
        RECT 136.960 138.120 137.190 138.600 ;
        RECT 128.755 137.840 136.755 138.070 ;
        RECT 119.930 136.710 125.330 137.170 ;
        RECT 119.930 135.370 121.930 136.710 ;
        RECT 123.680 136.700 125.330 136.710 ;
        RECT 122.370 135.430 123.370 136.150 ;
        RECT 123.680 135.890 123.990 136.700 ;
        RECT 124.450 136.420 125.330 136.700 ;
        RECT 125.570 136.880 127.190 137.280 ;
        RECT 128.840 136.930 136.710 137.840 ;
        RECT 124.390 136.190 125.390 136.420 ;
        RECT 125.570 136.230 125.920 136.880 ;
        RECT 126.570 136.870 127.190 136.880 ;
        RECT 128.755 136.700 136.755 136.930 ;
        RECT 128.840 136.690 136.710 136.700 ;
        RECT 124.450 135.980 125.330 136.000 ;
        RECT 123.720 135.600 123.990 135.890 ;
        RECT 124.390 135.750 125.390 135.980 ;
        RECT 125.550 135.940 125.920 136.230 ;
        RECT 125.580 135.880 125.920 135.940 ;
        RECT 126.680 136.550 127.440 136.600 ;
        RECT 128.320 136.550 128.550 136.650 ;
        RECT 126.680 136.340 128.550 136.550 ;
        RECT 136.960 136.340 137.190 136.650 ;
        RECT 126.680 135.920 129.220 136.340 ;
        RECT 136.590 135.920 137.190 136.340 ;
        RECT 124.450 135.600 125.330 135.750 ;
        RECT 124.460 135.430 125.190 135.600 ;
        RECT 102.400 134.080 105.400 134.310 ;
        RECT 105.610 134.120 105.950 134.950 ;
        RECT 107.960 134.940 118.600 135.010 ;
        RECT 102.450 134.050 105.310 134.080 ;
        RECT 102.450 134.030 103.620 134.050 ;
        RECT 104.580 134.040 105.310 134.050 ;
        RECT 102.400 133.640 105.400 133.870 ;
        RECT 105.605 133.830 105.950 134.120 ;
        RECT 106.140 133.900 118.600 134.940 ;
        RECT 120.000 135.360 121.930 135.370 ;
        RECT 106.140 133.880 118.560 133.900 ;
        RECT 105.610 133.720 105.950 133.830 ;
        RECT 106.180 133.870 111.850 133.880 ;
        RECT 112.850 133.870 118.560 133.880 ;
        RECT 102.490 133.470 105.350 133.640 ;
        RECT 106.180 133.470 106.610 133.870 ;
        RECT 102.460 133.100 106.610 133.470 ;
        RECT 11.950 130.910 90.610 131.390 ;
        RECT 59.400 130.510 59.720 130.770 ;
        RECT 66.300 130.710 66.620 130.770 ;
        RECT 67.235 130.710 67.525 130.755 ;
        RECT 66.300 130.570 67.525 130.710 ;
        RECT 66.300 130.510 66.620 130.570 ;
        RECT 67.235 130.525 67.525 130.570 ;
        RECT 28.120 130.370 28.410 130.415 ;
        RECT 29.690 130.370 29.980 130.415 ;
        RECT 31.790 130.370 32.080 130.415 ;
        RECT 28.120 130.230 32.080 130.370 ;
        RECT 28.120 130.185 28.410 130.230 ;
        RECT 29.690 130.185 29.980 130.230 ;
        RECT 31.790 130.185 32.080 130.230 ;
        RECT 35.520 130.370 35.810 130.415 ;
        RECT 37.620 130.370 37.910 130.415 ;
        RECT 39.190 130.370 39.480 130.415 ;
        RECT 35.520 130.230 39.480 130.370 ;
        RECT 35.520 130.185 35.810 130.230 ;
        RECT 37.620 130.185 37.910 130.230 ;
        RECT 39.190 130.185 39.480 130.230 ;
        RECT 41.000 130.370 41.320 130.430 ;
        RECT 45.615 130.370 45.905 130.415 ;
        RECT 41.000 130.230 45.905 130.370 ;
        RECT 41.000 130.170 41.320 130.230 ;
        RECT 45.615 130.185 45.905 130.230 ;
        RECT 53.000 130.370 53.290 130.415 ;
        RECT 55.100 130.370 55.390 130.415 ;
        RECT 56.670 130.370 56.960 130.415 ;
        RECT 68.600 130.370 68.920 130.430 ;
        RECT 53.000 130.230 56.960 130.370 ;
        RECT 53.000 130.185 53.290 130.230 ;
        RECT 55.100 130.185 55.390 130.230 ;
        RECT 56.670 130.185 56.960 130.230 ;
        RECT 64.090 130.230 68.920 130.370 ;
        RECT 27.685 130.030 27.975 130.075 ;
        RECT 30.205 130.030 30.495 130.075 ;
        RECT 31.395 130.030 31.685 130.075 ;
        RECT 32.720 130.030 33.040 130.090 ;
        RECT 27.685 129.890 31.685 130.030 ;
        RECT 27.685 129.845 27.975 129.890 ;
        RECT 30.205 129.845 30.495 129.890 ;
        RECT 31.395 129.845 31.685 129.890 ;
        RECT 31.890 129.890 33.040 130.030 ;
        RECT 30.995 129.690 31.285 129.735 ;
        RECT 31.890 129.690 32.030 129.890 ;
        RECT 32.720 129.830 33.040 129.890 ;
        RECT 35.915 130.030 36.205 130.075 ;
        RECT 37.105 130.030 37.395 130.075 ;
        RECT 39.625 130.030 39.915 130.075 ;
        RECT 44.695 130.030 44.985 130.075 ;
        RECT 35.915 129.890 39.915 130.030 ;
        RECT 35.915 129.845 36.205 129.890 ;
        RECT 37.105 129.845 37.395 129.890 ;
        RECT 39.625 129.845 39.915 129.890 ;
        RECT 43.390 129.890 44.985 130.030 ;
        RECT 30.995 129.550 32.030 129.690 ;
        RECT 32.275 129.690 32.565 129.735 ;
        RECT 35.035 129.690 35.325 129.735 ;
        RECT 35.480 129.690 35.800 129.750 ;
        RECT 36.400 129.735 36.720 129.750 ;
        RECT 36.370 129.690 36.720 129.735 ;
        RECT 39.160 129.690 39.480 129.750 ;
        RECT 32.275 129.550 35.800 129.690 ;
        RECT 36.205 129.550 36.720 129.690 ;
        RECT 30.995 129.505 31.285 129.550 ;
        RECT 32.275 129.505 32.565 129.550 ;
        RECT 35.035 129.505 35.325 129.550 ;
        RECT 35.480 129.490 35.800 129.550 ;
        RECT 36.370 129.505 36.720 129.550 ;
        RECT 36.400 129.490 36.720 129.505 ;
        RECT 37.410 129.550 39.480 129.690 ;
        RECT 27.200 129.350 27.520 129.410 ;
        RECT 33.655 129.350 33.945 129.395 ;
        RECT 27.200 129.210 33.945 129.350 ;
        RECT 27.200 129.150 27.520 129.210 ;
        RECT 33.655 129.165 33.945 129.210 ;
        RECT 34.575 129.350 34.865 129.395 ;
        RECT 37.410 129.350 37.550 129.550 ;
        RECT 39.160 129.490 39.480 129.550 ;
        RECT 41.920 129.690 42.240 129.750 ;
        RECT 42.855 129.690 43.145 129.735 ;
        RECT 41.920 129.550 43.145 129.690 ;
        RECT 41.920 129.490 42.240 129.550 ;
        RECT 42.855 129.505 43.145 129.550 ;
        RECT 42.395 129.350 42.685 129.395 ;
        RECT 34.575 129.210 37.550 129.350 ;
        RECT 37.870 129.210 42.685 129.350 ;
        RECT 34.575 129.165 34.865 129.210 ;
        RECT 25.360 128.810 25.680 129.070 ;
        RECT 32.735 129.010 33.025 129.055 ;
        RECT 37.870 129.010 38.010 129.210 ;
        RECT 42.395 129.165 42.685 129.210 ;
        RECT 32.735 128.870 38.010 129.010 ;
        RECT 39.160 129.010 39.480 129.070 ;
        RECT 41.935 129.010 42.225 129.055 ;
        RECT 43.390 129.010 43.530 129.890 ;
        RECT 44.695 129.845 44.985 129.890 ;
        RECT 46.060 130.030 46.380 130.090 ;
        RECT 64.090 130.075 64.230 130.230 ;
        RECT 68.600 130.170 68.920 130.230 ;
        RECT 53.395 130.030 53.685 130.075 ;
        RECT 54.585 130.030 54.875 130.075 ;
        RECT 57.105 130.030 57.395 130.075 ;
        RECT 46.060 129.890 52.270 130.030 ;
        RECT 44.220 129.490 44.540 129.750 ;
        RECT 44.770 129.690 44.910 129.845 ;
        RECT 46.060 129.830 46.380 129.890 ;
        RECT 47.900 129.690 48.220 129.750 ;
        RECT 52.130 129.735 52.270 129.890 ;
        RECT 53.395 129.890 57.395 130.030 ;
        RECT 53.395 129.845 53.685 129.890 ;
        RECT 54.585 129.845 54.875 129.890 ;
        RECT 57.105 129.845 57.395 129.890 ;
        RECT 64.015 129.845 64.305 130.075 ;
        RECT 66.440 130.030 66.730 130.075 ;
        RECT 67.220 130.030 67.540 130.090 ;
        RECT 66.440 129.890 67.540 130.030 ;
        RECT 66.440 129.845 66.730 129.890 ;
        RECT 67.220 129.830 67.540 129.890 ;
        RECT 48.835 129.690 49.125 129.735 ;
        RECT 51.135 129.690 51.425 129.735 ;
        RECT 44.770 129.550 51.425 129.690 ;
        RECT 47.900 129.490 48.220 129.550 ;
        RECT 48.835 129.505 49.125 129.550 ;
        RECT 51.135 129.505 51.425 129.550 ;
        RECT 52.055 129.505 52.345 129.735 ;
        RECT 52.515 129.690 52.805 129.735 ;
        RECT 56.640 129.690 56.960 129.750 ;
        RECT 52.515 129.550 56.960 129.690 ;
        RECT 52.515 129.505 52.805 129.550 ;
        RECT 56.640 129.490 56.960 129.550 ;
        RECT 63.540 129.690 63.860 129.750 ;
        RECT 65.395 129.690 65.685 129.735 ;
        RECT 63.540 129.550 65.685 129.690 ;
        RECT 63.540 129.490 63.860 129.550 ;
        RECT 65.395 129.505 65.685 129.550 ;
        RECT 100.010 129.620 100.880 131.720 ;
        RECT 106.550 131.330 107.800 131.770 ;
        RECT 117.700 131.750 118.560 133.870 ;
        RECT 120.000 131.810 120.770 135.360 ;
        RECT 122.340 134.310 125.190 135.430 ;
        RECT 125.580 135.130 125.930 135.880 ;
        RECT 126.680 135.760 128.550 135.920 ;
        RECT 126.680 135.710 127.440 135.760 ;
        RECT 128.320 135.690 128.550 135.760 ;
        RECT 136.960 135.690 137.190 135.920 ;
        RECT 128.755 135.410 136.755 135.640 ;
        RECT 125.580 135.070 125.870 135.130 ;
        RECT 125.490 134.950 125.870 135.070 ;
        RECT 128.850 135.010 136.710 135.410 ;
        RECT 137.520 135.010 138.480 144.490 ;
        RECT 122.280 134.080 125.280 134.310 ;
        RECT 125.490 134.120 125.830 134.950 ;
        RECT 127.840 134.940 138.480 135.010 ;
        RECT 122.330 134.050 125.190 134.080 ;
        RECT 122.330 134.030 123.500 134.050 ;
        RECT 124.460 134.040 125.190 134.050 ;
        RECT 122.280 133.640 125.280 133.870 ;
        RECT 125.485 133.830 125.830 134.120 ;
        RECT 126.020 133.900 138.480 134.940 ;
        RECT 139.930 146.720 140.700 150.360 ;
        RECT 142.420 149.310 145.270 150.430 ;
        RECT 145.660 150.130 146.010 150.880 ;
        RECT 146.760 150.760 148.630 150.920 ;
        RECT 146.760 150.710 147.520 150.760 ;
        RECT 148.400 150.690 148.630 150.760 ;
        RECT 157.040 150.690 157.270 150.920 ;
        RECT 148.835 150.410 156.835 150.640 ;
        RECT 145.660 150.070 145.950 150.130 ;
        RECT 145.570 149.950 145.950 150.070 ;
        RECT 148.930 150.010 156.790 150.410 ;
        RECT 157.600 150.010 158.560 159.490 ;
        RECT 142.360 149.080 145.360 149.310 ;
        RECT 145.570 149.120 145.910 149.950 ;
        RECT 147.920 149.940 158.560 150.010 ;
        RECT 142.410 149.050 145.270 149.080 ;
        RECT 142.410 149.030 143.580 149.050 ;
        RECT 144.540 149.040 145.270 149.050 ;
        RECT 142.360 148.640 145.360 148.870 ;
        RECT 145.565 148.830 145.910 149.120 ;
        RECT 146.100 148.900 158.560 149.940 ;
        RECT 146.100 148.880 158.500 148.900 ;
        RECT 145.570 148.720 145.910 148.830 ;
        RECT 146.140 148.870 151.810 148.880 ;
        RECT 152.810 148.870 158.500 148.880 ;
        RECT 142.450 148.470 145.310 148.640 ;
        RECT 146.140 148.470 146.570 148.870 ;
        RECT 142.420 148.100 146.570 148.470 ;
        RECT 139.930 144.620 140.790 146.720 ;
        RECT 146.460 146.330 147.710 146.770 ;
        RECT 157.640 146.750 158.500 148.870 ;
        RECT 144.400 146.320 149.640 146.330 ;
        RECT 141.450 146.220 156.750 146.320 ;
        RECT 141.450 146.210 156.785 146.220 ;
        RECT 141.410 146.090 156.785 146.210 ;
        RECT 141.410 145.980 145.410 146.090 ;
        RECT 146.460 146.010 148.200 146.090 ;
        RECT 148.780 146.010 156.785 146.090 ;
        RECT 146.460 145.930 147.710 146.010 ;
        RECT 148.785 145.990 156.785 146.010 ;
        RECT 141.020 145.680 141.250 145.930 ;
        RECT 145.570 145.790 145.800 145.930 ;
        RECT 148.350 145.790 148.580 145.940 ;
        RECT 145.570 145.680 148.580 145.790 ;
        RECT 156.990 145.680 157.220 145.940 ;
        RECT 141.020 145.240 157.220 145.680 ;
        RECT 141.020 144.970 141.250 145.240 ;
        RECT 145.570 145.210 157.220 145.240 ;
        RECT 145.570 145.120 148.580 145.210 ;
        RECT 145.570 144.970 145.800 145.120 ;
        RECT 148.350 144.980 148.580 145.120 ;
        RECT 156.990 144.980 157.220 145.210 ;
        RECT 141.410 144.690 145.410 144.920 ;
        RECT 148.785 144.710 156.785 144.930 ;
        RECT 157.550 144.710 158.510 146.750 ;
        RECT 148.785 144.700 158.510 144.710 ;
        RECT 141.410 144.620 145.400 144.690 ;
        RECT 139.930 144.510 145.400 144.620 ;
        RECT 148.840 144.540 158.510 144.700 ;
        RECT 139.930 144.420 143.090 144.510 ;
        RECT 156.580 144.490 158.510 144.540 ;
        RECT 139.930 141.150 140.790 144.420 ;
        RECT 144.440 143.960 149.690 143.970 ;
        RECT 144.440 143.850 156.750 143.960 ;
        RECT 141.470 143.790 156.750 143.850 ;
        RECT 141.470 143.780 156.785 143.790 ;
        RECT 141.410 143.650 156.785 143.780 ;
        RECT 141.410 143.640 146.570 143.650 ;
        RECT 141.410 143.550 145.410 143.640 ;
        RECT 148.785 143.560 156.785 143.650 ;
        RECT 148.870 143.550 156.760 143.560 ;
        RECT 141.020 143.190 141.250 143.500 ;
        RECT 141.470 143.190 145.370 143.550 ;
        RECT 145.570 143.190 145.800 143.500 ;
        RECT 141.020 141.850 145.800 143.190 ;
        RECT 141.020 141.540 141.250 141.850 ;
        RECT 145.570 141.540 145.800 141.850 ;
        RECT 148.350 142.970 148.580 143.510 ;
        RECT 149.390 142.970 150.400 143.000 ;
        RECT 156.990 142.970 157.220 143.510 ;
        RECT 148.350 142.070 157.220 142.970 ;
        RECT 148.350 141.550 148.580 142.070 ;
        RECT 149.390 142.000 150.400 142.070 ;
        RECT 156.990 141.550 157.220 142.070 ;
        RECT 141.410 141.260 145.410 141.490 ;
        RECT 148.785 141.270 156.785 141.500 ;
        RECT 139.930 141.110 141.090 141.150 ;
        RECT 139.930 141.030 141.330 141.110 ;
        RECT 141.700 141.040 145.360 141.260 ;
        RECT 141.700 141.030 143.140 141.040 ;
        RECT 139.930 140.990 143.140 141.030 ;
        RECT 139.930 140.900 142.650 140.990 ;
        RECT 148.850 140.980 156.740 141.270 ;
        RECT 139.930 140.840 141.980 140.900 ;
        RECT 139.930 140.790 141.730 140.840 ;
        RECT 139.930 137.450 140.790 140.790 ;
        RECT 148.840 140.490 156.760 140.500 ;
        RECT 145.070 140.480 156.760 140.490 ;
        RECT 141.450 140.360 156.760 140.480 ;
        RECT 141.450 140.350 156.785 140.360 ;
        RECT 141.410 140.230 156.785 140.350 ;
        RECT 141.410 140.120 145.410 140.230 ;
        RECT 141.020 139.780 141.250 140.070 ;
        RECT 141.470 139.780 145.360 140.120 ;
        RECT 145.570 139.780 145.800 140.070 ;
        RECT 141.020 138.410 145.800 139.780 ;
        RECT 141.020 138.110 141.250 138.410 ;
        RECT 145.570 138.110 145.800 138.410 ;
        RECT 141.410 137.830 145.410 138.060 ;
        RECT 141.660 137.600 145.230 137.830 ;
        RECT 141.660 137.450 145.350 137.600 ;
        RECT 139.930 137.170 145.350 137.450 ;
        RECT 146.600 137.280 147.220 140.230 ;
        RECT 148.785 140.130 156.785 140.230 ;
        RECT 148.840 140.120 156.760 140.130 ;
        RECT 148.350 139.420 148.580 140.080 ;
        RECT 149.360 139.420 150.360 139.510 ;
        RECT 156.990 139.420 157.220 140.080 ;
        RECT 148.350 138.600 157.220 139.420 ;
        RECT 148.350 138.120 148.580 138.600 ;
        RECT 149.360 138.510 150.360 138.600 ;
        RECT 156.990 138.120 157.220 138.600 ;
        RECT 148.785 137.840 156.785 138.070 ;
        RECT 139.930 136.710 145.360 137.170 ;
        RECT 139.930 135.360 141.960 136.710 ;
        RECT 143.710 136.700 145.360 136.710 ;
        RECT 142.400 135.430 143.400 136.150 ;
        RECT 143.710 135.890 144.020 136.700 ;
        RECT 144.480 136.420 145.360 136.700 ;
        RECT 145.600 136.880 147.220 137.280 ;
        RECT 148.870 136.930 156.740 137.840 ;
        RECT 144.420 136.190 145.420 136.420 ;
        RECT 145.600 136.230 145.950 136.880 ;
        RECT 146.600 136.870 147.220 136.880 ;
        RECT 148.785 136.700 156.785 136.930 ;
        RECT 148.870 136.690 156.740 136.700 ;
        RECT 144.480 135.980 145.360 136.000 ;
        RECT 143.750 135.600 144.020 135.890 ;
        RECT 144.420 135.750 145.420 135.980 ;
        RECT 145.580 135.940 145.950 136.230 ;
        RECT 145.610 135.880 145.950 135.940 ;
        RECT 146.710 136.550 147.470 136.600 ;
        RECT 148.350 136.550 148.580 136.650 ;
        RECT 146.710 136.340 148.580 136.550 ;
        RECT 156.990 136.340 157.220 136.650 ;
        RECT 146.710 135.920 149.250 136.340 ;
        RECT 156.620 135.920 157.220 136.340 ;
        RECT 144.480 135.600 145.360 135.750 ;
        RECT 144.490 135.430 145.220 135.600 ;
        RECT 126.020 133.880 138.460 133.900 ;
        RECT 125.490 133.720 125.830 133.830 ;
        RECT 126.060 133.870 131.730 133.880 ;
        RECT 132.730 133.870 138.460 133.880 ;
        RECT 122.370 133.470 125.230 133.640 ;
        RECT 126.060 133.470 126.490 133.870 ;
        RECT 122.340 133.100 126.490 133.470 ;
        RECT 104.490 131.320 109.730 131.330 ;
        RECT 101.540 131.220 116.840 131.320 ;
        RECT 101.540 131.210 116.875 131.220 ;
        RECT 101.500 131.090 116.875 131.210 ;
        RECT 101.500 130.980 105.500 131.090 ;
        RECT 106.550 131.010 108.290 131.090 ;
        RECT 108.870 131.010 116.875 131.090 ;
        RECT 106.550 130.930 107.800 131.010 ;
        RECT 108.875 130.990 116.875 131.010 ;
        RECT 101.110 130.680 101.340 130.930 ;
        RECT 105.660 130.790 105.890 130.930 ;
        RECT 108.440 130.790 108.670 130.940 ;
        RECT 105.660 130.680 108.670 130.790 ;
        RECT 117.080 130.680 117.310 130.940 ;
        RECT 101.110 130.240 117.310 130.680 ;
        RECT 101.110 129.970 101.340 130.240 ;
        RECT 105.660 130.210 117.310 130.240 ;
        RECT 105.660 130.120 108.670 130.210 ;
        RECT 105.660 129.970 105.890 130.120 ;
        RECT 108.440 129.980 108.670 130.120 ;
        RECT 117.080 129.980 117.310 130.210 ;
        RECT 101.500 129.690 105.500 129.920 ;
        RECT 108.875 129.710 116.875 129.930 ;
        RECT 117.640 129.710 118.600 131.750 ;
        RECT 108.875 129.700 118.600 129.710 ;
        RECT 101.500 129.620 105.490 129.690 ;
        RECT 100.010 129.510 105.490 129.620 ;
        RECT 108.930 129.540 118.600 129.700 ;
        RECT 100.010 129.420 103.180 129.510 ;
        RECT 116.670 129.490 118.600 129.540 ;
        RECT 43.760 129.350 44.080 129.410 ;
        RECT 53.880 129.395 54.200 129.410 ;
        RECT 46.075 129.350 46.365 129.395 ;
        RECT 53.850 129.350 54.200 129.395 ;
        RECT 43.760 129.210 46.365 129.350 ;
        RECT 53.685 129.210 54.200 129.350 ;
        RECT 43.760 129.150 44.080 129.210 ;
        RECT 46.075 129.165 46.365 129.210 ;
        RECT 53.850 129.165 54.200 129.210 ;
        RECT 53.880 129.150 54.200 129.165 ;
        RECT 39.160 128.870 43.530 129.010 ;
        RECT 44.680 129.010 45.000 129.070 ;
        RECT 48.360 129.010 48.680 129.070 ;
        RECT 51.135 129.010 51.425 129.055 ;
        RECT 44.680 128.870 51.425 129.010 ;
        RECT 32.735 128.825 33.025 128.870 ;
        RECT 39.160 128.810 39.480 128.870 ;
        RECT 41.935 128.825 42.225 128.870 ;
        RECT 44.680 128.810 45.000 128.870 ;
        RECT 48.360 128.810 48.680 128.870 ;
        RECT 51.135 128.825 51.425 128.870 ;
        RECT 52.960 129.010 53.280 129.070 ;
        RECT 65.855 129.010 66.145 129.055 ;
        RECT 52.960 128.870 66.145 129.010 ;
        RECT 52.960 128.810 53.280 128.870 ;
        RECT 65.855 128.825 66.145 128.870 ;
        RECT 11.950 128.190 90.610 128.670 ;
        RECT 27.200 127.790 27.520 128.050 ;
        RECT 34.560 127.790 34.880 128.050 ;
        RECT 46.075 127.805 46.365 128.035 ;
        RECT 44.220 127.650 44.540 127.710 ;
        RECT 36.030 127.510 44.540 127.650 ;
        RECT 32.835 127.310 33.125 127.355 ;
        RECT 33.640 127.310 33.960 127.370 ;
        RECT 32.835 127.170 33.960 127.310 ;
        RECT 32.835 127.125 33.125 127.170 ;
        RECT 33.640 127.110 33.960 127.170 ;
        RECT 36.030 127.030 36.170 127.510 ;
        RECT 44.220 127.450 44.540 127.510 ;
        RECT 36.415 127.310 36.705 127.355 ;
        RECT 43.760 127.310 44.080 127.370 ;
        RECT 36.415 127.170 44.080 127.310 ;
        RECT 36.415 127.125 36.705 127.170 ;
        RECT 43.760 127.110 44.080 127.170 ;
        RECT 44.680 127.110 45.000 127.370 ;
        RECT 46.150 127.310 46.290 127.805 ;
        RECT 47.815 127.310 48.105 127.355 ;
        RECT 46.150 127.170 48.105 127.310 ;
        RECT 47.815 127.125 48.105 127.170 ;
        RECT 29.525 126.970 29.815 127.015 ;
        RECT 32.045 126.970 32.335 127.015 ;
        RECT 33.235 126.970 33.525 127.015 ;
        RECT 29.525 126.830 33.525 126.970 ;
        RECT 29.525 126.785 29.815 126.830 ;
        RECT 32.045 126.785 32.335 126.830 ;
        RECT 33.235 126.785 33.525 126.830 ;
        RECT 34.115 126.785 34.405 127.015 ;
        RECT 29.960 126.630 30.250 126.675 ;
        RECT 31.530 126.630 31.820 126.675 ;
        RECT 33.630 126.630 33.920 126.675 ;
        RECT 29.960 126.490 33.920 126.630 ;
        RECT 34.190 126.630 34.330 126.785 ;
        RECT 35.940 126.770 36.260 127.030 ;
        RECT 38.700 126.970 39.020 127.030 ;
        RECT 39.175 126.970 39.465 127.015 ;
        RECT 38.700 126.830 39.465 126.970 ;
        RECT 38.700 126.770 39.020 126.830 ;
        RECT 39.175 126.785 39.465 126.830 ;
        RECT 40.540 126.970 40.860 127.030 ;
        RECT 42.840 126.970 43.160 127.030 ;
        RECT 40.540 126.830 43.160 126.970 ;
        RECT 40.540 126.770 40.860 126.830 ;
        RECT 42.840 126.770 43.160 126.830 ;
        RECT 43.315 126.970 43.605 127.015 ;
        RECT 44.220 126.970 44.540 127.030 ;
        RECT 43.315 126.830 44.540 126.970 ;
        RECT 43.315 126.785 43.605 126.830 ;
        RECT 44.220 126.770 44.540 126.830 ;
        RECT 45.140 126.770 45.460 127.030 ;
        RECT 46.535 126.785 46.825 127.015 ;
        RECT 47.415 126.970 47.705 127.015 ;
        RECT 48.605 126.970 48.895 127.015 ;
        RECT 51.125 126.970 51.415 127.015 ;
        RECT 47.415 126.830 51.415 126.970 ;
        RECT 47.415 126.785 47.705 126.830 ;
        RECT 48.605 126.785 48.895 126.830 ;
        RECT 51.125 126.785 51.415 126.830 ;
        RECT 35.480 126.630 35.800 126.690 ;
        RECT 46.610 126.630 46.750 126.785 ;
        RECT 34.190 126.490 46.750 126.630 ;
        RECT 47.020 126.630 47.310 126.675 ;
        RECT 49.120 126.630 49.410 126.675 ;
        RECT 50.690 126.630 50.980 126.675 ;
        RECT 47.020 126.490 50.980 126.630 ;
        RECT 29.960 126.445 30.250 126.490 ;
        RECT 31.530 126.445 31.820 126.490 ;
        RECT 33.630 126.445 33.920 126.490 ;
        RECT 35.480 126.430 35.800 126.490 ;
        RECT 43.390 126.350 43.530 126.490 ;
        RECT 47.020 126.445 47.310 126.490 ;
        RECT 49.120 126.445 49.410 126.490 ;
        RECT 50.690 126.445 50.980 126.490 ;
        RECT 52.040 126.630 52.360 126.690 ;
        RECT 53.435 126.630 53.725 126.675 ;
        RECT 52.040 126.490 53.725 126.630 ;
        RECT 52.040 126.430 52.360 126.490 ;
        RECT 53.435 126.445 53.725 126.490 ;
        RECT 38.240 126.290 38.560 126.350 ;
        RECT 40.540 126.290 40.860 126.350 ;
        RECT 38.240 126.150 40.860 126.290 ;
        RECT 38.240 126.090 38.560 126.150 ;
        RECT 40.540 126.090 40.860 126.150 ;
        RECT 42.380 126.090 42.700 126.350 ;
        RECT 43.300 126.090 43.620 126.350 ;
        RECT 44.220 126.290 44.540 126.350 ;
        RECT 47.440 126.290 47.760 126.350 ;
        RECT 44.220 126.150 47.760 126.290 ;
        RECT 44.220 126.090 44.540 126.150 ;
        RECT 47.440 126.090 47.760 126.150 ;
        RECT 100.010 126.150 100.880 129.420 ;
        RECT 104.530 128.960 109.780 128.970 ;
        RECT 104.530 128.850 116.840 128.960 ;
        RECT 101.560 128.790 116.840 128.850 ;
        RECT 101.560 128.780 116.875 128.790 ;
        RECT 101.500 128.650 116.875 128.780 ;
        RECT 101.500 128.640 106.660 128.650 ;
        RECT 101.500 128.550 105.500 128.640 ;
        RECT 108.875 128.560 116.875 128.650 ;
        RECT 108.960 128.550 116.850 128.560 ;
        RECT 101.110 128.190 101.340 128.500 ;
        RECT 101.560 128.190 105.460 128.550 ;
        RECT 105.660 128.190 105.890 128.500 ;
        RECT 101.110 126.850 105.890 128.190 ;
        RECT 101.110 126.540 101.340 126.850 ;
        RECT 105.660 126.540 105.890 126.850 ;
        RECT 108.440 127.970 108.670 128.510 ;
        RECT 109.480 127.970 110.490 128.000 ;
        RECT 117.080 127.970 117.310 128.510 ;
        RECT 108.440 127.070 117.310 127.970 ;
        RECT 108.440 126.550 108.670 127.070 ;
        RECT 109.480 127.000 110.490 127.070 ;
        RECT 117.080 126.550 117.310 127.070 ;
        RECT 101.500 126.260 105.500 126.490 ;
        RECT 108.875 126.270 116.875 126.500 ;
        RECT 100.010 126.110 101.180 126.150 ;
        RECT 100.010 126.030 101.420 126.110 ;
        RECT 101.790 126.040 105.450 126.260 ;
        RECT 101.790 126.030 103.230 126.040 ;
        RECT 100.010 125.990 103.230 126.030 ;
        RECT 11.950 125.470 90.610 125.950 ;
        RECT 100.010 125.900 102.740 125.990 ;
        RECT 108.940 125.980 116.830 126.270 ;
        RECT 100.010 125.840 102.070 125.900 ;
        RECT 100.010 125.790 101.820 125.840 ;
        RECT 33.640 125.070 33.960 125.330 ;
        RECT 38.700 125.070 39.020 125.330 ;
        RECT 39.175 125.270 39.465 125.315 ;
        RECT 41.460 125.270 41.780 125.330 ;
        RECT 39.175 125.130 41.780 125.270 ;
        RECT 39.175 125.085 39.465 125.130 ;
        RECT 41.460 125.070 41.780 125.130 ;
        RECT 43.760 125.270 44.080 125.330 ;
        RECT 45.600 125.270 45.920 125.330 ;
        RECT 46.980 125.270 47.300 125.330 ;
        RECT 47.455 125.270 47.745 125.315 ;
        RECT 43.760 125.130 44.865 125.270 ;
        RECT 43.760 125.070 44.080 125.130 ;
        RECT 35.035 124.930 35.325 124.975 ;
        RECT 35.940 124.930 36.260 124.990 ;
        RECT 35.035 124.790 36.260 124.930 ;
        RECT 35.035 124.745 35.325 124.790 ;
        RECT 35.940 124.730 36.260 124.790 ;
        RECT 40.080 124.730 40.400 124.990 ;
        RECT 40.580 124.930 40.870 124.975 ;
        RECT 42.680 124.930 42.970 124.975 ;
        RECT 44.250 124.930 44.540 124.975 ;
        RECT 40.580 124.790 44.540 124.930 ;
        RECT 44.725 124.930 44.865 125.130 ;
        RECT 45.600 125.130 47.745 125.270 ;
        RECT 45.600 125.070 45.920 125.130 ;
        RECT 46.980 125.070 47.300 125.130 ;
        RECT 47.455 125.085 47.745 125.130 ;
        RECT 52.515 124.930 52.805 124.975 ;
        RECT 44.725 124.790 52.805 124.930 ;
        RECT 40.580 124.745 40.870 124.790 ;
        RECT 42.680 124.745 42.970 124.790 ;
        RECT 44.250 124.745 44.540 124.790 ;
        RECT 52.515 124.745 52.805 124.790 ;
        RECT 25.360 124.590 25.680 124.650 ;
        RECT 26.755 124.590 27.045 124.635 ;
        RECT 25.360 124.450 27.045 124.590 ;
        RECT 25.360 124.390 25.680 124.450 ;
        RECT 26.755 124.405 27.045 124.450 ;
        RECT 35.480 124.390 35.800 124.650 ;
        RECT 40.170 124.590 40.310 124.730 ;
        RECT 36.950 124.450 40.310 124.590 ;
        RECT 40.975 124.590 41.265 124.635 ;
        RECT 42.165 124.590 42.455 124.635 ;
        RECT 44.685 124.590 44.975 124.635 ;
        RECT 40.975 124.450 44.975 124.590 ;
        RECT 34.575 124.065 34.865 124.295 ;
        RECT 35.955 124.250 36.245 124.295 ;
        RECT 36.400 124.250 36.720 124.310 ;
        RECT 36.950 124.295 37.090 124.450 ;
        RECT 40.975 124.405 41.265 124.450 ;
        RECT 42.165 124.405 42.455 124.450 ;
        RECT 44.685 124.405 44.975 124.450 ;
        RECT 47.900 124.390 48.220 124.650 ;
        RECT 64.475 124.590 64.765 124.635 ;
        RECT 64.935 124.590 65.225 124.635 ;
        RECT 64.475 124.450 65.225 124.590 ;
        RECT 64.475 124.405 64.765 124.450 ;
        RECT 64.935 124.405 65.225 124.450 ;
        RECT 35.955 124.110 36.720 124.250 ;
        RECT 35.955 124.065 36.245 124.110 ;
        RECT 34.650 123.910 34.790 124.065 ;
        RECT 36.400 124.050 36.720 124.110 ;
        RECT 36.875 124.065 37.165 124.295 ;
        RECT 37.780 124.050 38.100 124.310 ;
        RECT 38.240 124.050 38.560 124.310 ;
        RECT 39.635 124.065 39.925 124.295 ;
        RECT 40.095 124.250 40.385 124.295 ;
        RECT 43.300 124.250 43.620 124.310 ;
        RECT 40.095 124.110 43.620 124.250 ;
        RECT 40.095 124.065 40.385 124.110 ;
        RECT 39.160 123.910 39.480 123.970 ;
        RECT 34.650 123.770 39.480 123.910 ;
        RECT 39.160 123.710 39.480 123.770 ;
        RECT 29.975 123.570 30.265 123.615 ;
        RECT 30.420 123.570 30.740 123.630 ;
        RECT 29.975 123.430 30.740 123.570 ;
        RECT 39.710 123.570 39.850 124.065 ;
        RECT 43.300 124.050 43.620 124.110 ;
        RECT 47.440 124.050 47.760 124.310 ;
        RECT 58.480 124.050 58.800 124.310 ;
        RECT 66.300 124.050 66.620 124.310 ;
        RECT 66.760 124.050 67.080 124.310 ;
        RECT 67.235 124.065 67.525 124.295 ;
        RECT 67.680 124.250 68.000 124.310 ;
        RECT 68.155 124.250 68.445 124.295 ;
        RECT 67.680 124.110 68.445 124.250 ;
        RECT 41.430 123.910 41.720 123.955 ;
        RECT 42.380 123.910 42.700 123.970 ;
        RECT 41.430 123.770 42.700 123.910 ;
        RECT 41.430 123.725 41.720 123.770 ;
        RECT 42.380 123.710 42.700 123.770 ;
        RECT 51.595 123.725 51.885 123.955 ;
        RECT 64.460 123.910 64.780 123.970 ;
        RECT 67.310 123.910 67.450 124.065 ;
        RECT 67.680 124.050 68.000 124.110 ;
        RECT 68.155 124.065 68.445 124.110 ;
        RECT 64.460 123.770 67.450 123.910 ;
        RECT 45.140 123.570 45.460 123.630 ;
        RECT 39.710 123.430 45.460 123.570 ;
        RECT 29.975 123.385 30.265 123.430 ;
        RECT 30.420 123.370 30.740 123.430 ;
        RECT 45.140 123.370 45.460 123.430 ;
        RECT 49.295 123.570 49.585 123.615 ;
        RECT 49.740 123.570 50.060 123.630 ;
        RECT 51.670 123.570 51.810 123.725 ;
        RECT 64.460 123.710 64.780 123.770 ;
        RECT 49.295 123.430 51.810 123.570 ;
        RECT 55.260 123.570 55.580 123.630 ;
        RECT 55.735 123.570 56.025 123.615 ;
        RECT 55.260 123.430 56.025 123.570 ;
        RECT 49.295 123.385 49.585 123.430 ;
        RECT 49.740 123.370 50.060 123.430 ;
        RECT 55.260 123.370 55.580 123.430 ;
        RECT 55.735 123.385 56.025 123.430 ;
        RECT 60.320 123.570 60.640 123.630 ;
        RECT 61.255 123.570 61.545 123.615 ;
        RECT 60.320 123.430 61.545 123.570 ;
        RECT 60.320 123.370 60.640 123.430 ;
        RECT 61.255 123.385 61.545 123.430 ;
        RECT 11.950 122.750 90.610 123.230 ;
        RECT 28.595 122.550 28.885 122.595 ;
        RECT 29.500 122.550 29.820 122.610 ;
        RECT 28.595 122.410 29.820 122.550 ;
        RECT 28.595 122.365 28.885 122.410 ;
        RECT 29.500 122.350 29.820 122.410 ;
        RECT 45.140 122.550 45.460 122.610 ;
        RECT 46.535 122.550 46.825 122.595 ;
        RECT 45.140 122.410 46.825 122.550 ;
        RECT 45.140 122.350 45.460 122.410 ;
        RECT 46.535 122.365 46.825 122.410 ;
        RECT 47.440 122.550 47.760 122.610 ;
        RECT 61.715 122.550 62.005 122.595 ;
        RECT 47.440 122.410 62.005 122.550 ;
        RECT 47.440 122.350 47.760 122.410 ;
        RECT 61.715 122.365 62.005 122.410 ;
        RECT 100.010 122.450 100.880 125.790 ;
        RECT 108.930 125.490 116.850 125.500 ;
        RECT 105.160 125.480 116.850 125.490 ;
        RECT 101.540 125.360 116.850 125.480 ;
        RECT 101.540 125.350 116.875 125.360 ;
        RECT 101.500 125.230 116.875 125.350 ;
        RECT 101.500 125.120 105.500 125.230 ;
        RECT 101.110 124.780 101.340 125.070 ;
        RECT 101.560 124.780 105.450 125.120 ;
        RECT 105.660 124.780 105.890 125.070 ;
        RECT 101.110 123.410 105.890 124.780 ;
        RECT 101.110 123.110 101.340 123.410 ;
        RECT 105.660 123.110 105.890 123.410 ;
        RECT 101.500 122.830 105.500 123.060 ;
        RECT 101.750 122.600 105.320 122.830 ;
        RECT 101.750 122.450 105.440 122.600 ;
        RECT 44.695 122.210 44.985 122.255 ;
        RECT 56.640 122.210 56.960 122.270 ;
        RECT 44.695 122.070 47.210 122.210 ;
        RECT 44.695 122.025 44.985 122.070 ;
        RECT 47.070 121.930 47.210 122.070 ;
        RECT 53.970 122.070 56.960 122.210 ;
        RECT 21.680 121.670 22.000 121.930 ;
        RECT 22.140 121.870 22.460 121.930 ;
        RECT 22.975 121.870 23.265 121.915 ;
        RECT 22.140 121.730 23.265 121.870 ;
        RECT 22.140 121.670 22.460 121.730 ;
        RECT 22.975 121.685 23.265 121.730 ;
        RECT 45.615 121.685 45.905 121.915 ;
        RECT 46.980 121.870 47.300 121.930 ;
        RECT 47.455 121.870 47.745 121.915 ;
        RECT 46.980 121.730 47.745 121.870 ;
        RECT 22.575 121.530 22.865 121.575 ;
        RECT 23.765 121.530 24.055 121.575 ;
        RECT 26.285 121.530 26.575 121.575 ;
        RECT 22.575 121.390 26.575 121.530 ;
        RECT 45.690 121.530 45.830 121.685 ;
        RECT 46.980 121.670 47.300 121.730 ;
        RECT 47.455 121.685 47.745 121.730 ;
        RECT 48.360 121.670 48.680 121.930 ;
        RECT 53.970 121.915 54.110 122.070 ;
        RECT 56.640 122.010 56.960 122.070 ;
        RECT 100.010 122.170 105.440 122.450 ;
        RECT 106.690 122.280 107.310 125.230 ;
        RECT 108.875 125.130 116.875 125.230 ;
        RECT 108.930 125.120 116.850 125.130 ;
        RECT 108.440 124.420 108.670 125.080 ;
        RECT 109.450 124.420 110.450 124.510 ;
        RECT 117.080 124.420 117.310 125.080 ;
        RECT 108.440 123.600 117.310 124.420 ;
        RECT 108.440 123.120 108.670 123.600 ;
        RECT 109.450 123.510 110.450 123.600 ;
        RECT 117.080 123.120 117.310 123.600 ;
        RECT 108.875 122.840 116.875 123.070 ;
        RECT 55.260 121.915 55.580 121.930 ;
        RECT 53.895 121.685 54.185 121.915 ;
        RECT 55.230 121.870 55.580 121.915 ;
        RECT 61.255 121.870 61.545 121.915 ;
        RECT 55.065 121.730 55.580 121.870 ;
        RECT 55.230 121.685 55.580 121.730 ;
        RECT 55.260 121.670 55.580 121.685 ;
        RECT 60.870 121.730 61.545 121.870 ;
        RECT 48.450 121.530 48.590 121.670 ;
        RECT 45.690 121.390 48.590 121.530 ;
        RECT 54.775 121.530 55.065 121.575 ;
        RECT 55.965 121.530 56.255 121.575 ;
        RECT 58.485 121.530 58.775 121.575 ;
        RECT 54.775 121.390 58.775 121.530 ;
        RECT 22.575 121.345 22.865 121.390 ;
        RECT 23.765 121.345 24.055 121.390 ;
        RECT 26.285 121.345 26.575 121.390 ;
        RECT 54.775 121.345 55.065 121.390 ;
        RECT 55.965 121.345 56.255 121.390 ;
        RECT 58.485 121.345 58.775 121.390 ;
        RECT 22.180 121.190 22.470 121.235 ;
        RECT 24.280 121.190 24.570 121.235 ;
        RECT 25.850 121.190 26.140 121.235 ;
        RECT 22.180 121.050 26.140 121.190 ;
        RECT 22.180 121.005 22.470 121.050 ;
        RECT 24.280 121.005 24.570 121.050 ;
        RECT 25.850 121.005 26.140 121.050 ;
        RECT 39.620 121.190 39.940 121.250 ;
        RECT 60.870 121.235 61.010 121.730 ;
        RECT 61.255 121.685 61.545 121.730 ;
        RECT 62.175 121.870 62.465 121.915 ;
        RECT 65.840 121.870 66.160 121.930 ;
        RECT 62.175 121.730 66.160 121.870 ;
        RECT 62.175 121.685 62.465 121.730 ;
        RECT 65.840 121.670 66.160 121.730 ;
        RECT 71.475 121.870 71.765 121.915 ;
        RECT 72.280 121.870 72.600 121.930 ;
        RECT 71.475 121.730 72.600 121.870 ;
        RECT 71.475 121.685 71.765 121.730 ;
        RECT 72.280 121.670 72.600 121.730 ;
        RECT 72.740 121.870 73.060 121.930 ;
        RECT 75.500 121.870 75.820 121.930 ;
        RECT 72.740 121.730 75.820 121.870 ;
        RECT 72.740 121.670 73.060 121.730 ;
        RECT 75.500 121.670 75.820 121.730 ;
        RECT 100.010 121.710 105.450 122.170 ;
        RECT 68.165 121.530 68.455 121.575 ;
        RECT 70.685 121.530 70.975 121.575 ;
        RECT 71.875 121.530 72.165 121.575 ;
        RECT 68.165 121.390 72.165 121.530 ;
        RECT 68.165 121.345 68.455 121.390 ;
        RECT 70.685 121.345 70.975 121.390 ;
        RECT 71.875 121.345 72.165 121.390 ;
        RECT 48.375 121.190 48.665 121.235 ;
        RECT 39.620 121.050 48.665 121.190 ;
        RECT 39.620 120.990 39.940 121.050 ;
        RECT 48.375 121.005 48.665 121.050 ;
        RECT 54.380 121.190 54.670 121.235 ;
        RECT 56.480 121.190 56.770 121.235 ;
        RECT 58.050 121.190 58.340 121.235 ;
        RECT 54.380 121.050 58.340 121.190 ;
        RECT 54.380 121.005 54.670 121.050 ;
        RECT 56.480 121.005 56.770 121.050 ;
        RECT 58.050 121.005 58.340 121.050 ;
        RECT 60.795 121.005 61.085 121.235 ;
        RECT 68.600 121.190 68.890 121.235 ;
        RECT 70.170 121.190 70.460 121.235 ;
        RECT 72.270 121.190 72.560 121.235 ;
        RECT 68.600 121.050 72.560 121.190 ;
        RECT 68.600 121.005 68.890 121.050 ;
        RECT 70.170 121.005 70.460 121.050 ;
        RECT 72.270 121.005 72.560 121.050 ;
        RECT 43.760 120.650 44.080 120.910 ;
        RECT 65.855 120.850 66.145 120.895 ;
        RECT 67.220 120.850 67.540 120.910 ;
        RECT 65.855 120.710 67.540 120.850 ;
        RECT 65.855 120.665 66.145 120.710 ;
        RECT 67.220 120.650 67.540 120.710 ;
        RECT 11.950 120.030 90.610 120.510 ;
        RECT 100.010 120.360 102.050 121.710 ;
        RECT 103.800 121.700 105.450 121.710 ;
        RECT 102.490 120.430 103.490 121.150 ;
        RECT 103.800 120.890 104.110 121.700 ;
        RECT 104.570 121.420 105.450 121.700 ;
        RECT 105.690 121.880 107.310 122.280 ;
        RECT 108.960 121.930 116.830 122.840 ;
        RECT 104.510 121.190 105.510 121.420 ;
        RECT 105.690 121.230 106.040 121.880 ;
        RECT 106.690 121.870 107.310 121.880 ;
        RECT 108.875 121.700 116.875 121.930 ;
        RECT 108.960 121.690 116.830 121.700 ;
        RECT 104.570 120.980 105.450 121.000 ;
        RECT 103.840 120.600 104.110 120.890 ;
        RECT 104.510 120.750 105.510 120.980 ;
        RECT 105.670 120.940 106.040 121.230 ;
        RECT 105.700 120.880 106.040 120.940 ;
        RECT 106.800 121.550 107.560 121.600 ;
        RECT 108.440 121.550 108.670 121.650 ;
        RECT 106.800 121.340 108.670 121.550 ;
        RECT 117.080 121.340 117.310 121.650 ;
        RECT 106.800 120.920 109.340 121.340 ;
        RECT 116.710 120.920 117.310 121.340 ;
        RECT 104.570 120.600 105.450 120.750 ;
        RECT 104.580 120.430 105.310 120.600 ;
        RECT 22.140 119.630 22.460 119.890 ;
        RECT 23.060 119.830 23.380 119.890 ;
        RECT 29.960 119.830 30.280 119.890 ;
        RECT 23.060 119.690 30.280 119.830 ;
        RECT 23.060 119.630 23.380 119.690 ;
        RECT 29.960 119.630 30.280 119.690 ;
        RECT 65.840 119.630 66.160 119.890 ;
        RECT 66.300 119.630 66.620 119.890 ;
        RECT 72.280 119.830 72.600 119.890 ;
        RECT 72.755 119.830 73.045 119.875 ;
        RECT 72.280 119.690 73.045 119.830 ;
        RECT 72.280 119.630 72.600 119.690 ;
        RECT 72.755 119.645 73.045 119.690 ;
        RECT 17.540 119.490 17.830 119.535 ;
        RECT 19.110 119.490 19.400 119.535 ;
        RECT 21.210 119.490 21.500 119.535 ;
        RECT 25.860 119.490 26.150 119.535 ;
        RECT 27.960 119.490 28.250 119.535 ;
        RECT 29.530 119.490 29.820 119.535 ;
        RECT 17.540 119.350 21.500 119.490 ;
        RECT 17.540 119.305 17.830 119.350 ;
        RECT 19.110 119.305 19.400 119.350 ;
        RECT 21.210 119.305 21.500 119.350 ;
        RECT 21.770 119.350 25.590 119.490 ;
        RECT 21.770 119.210 21.910 119.350 ;
        RECT 17.105 119.150 17.395 119.195 ;
        RECT 19.625 119.150 19.915 119.195 ;
        RECT 20.815 119.150 21.105 119.195 ;
        RECT 17.105 119.010 21.105 119.150 ;
        RECT 17.105 118.965 17.395 119.010 ;
        RECT 19.625 118.965 19.915 119.010 ;
        RECT 20.815 118.965 21.105 119.010 ;
        RECT 21.680 118.950 22.000 119.210 ;
        RECT 25.450 119.195 25.590 119.350 ;
        RECT 25.860 119.350 29.820 119.490 ;
        RECT 25.860 119.305 26.150 119.350 ;
        RECT 27.960 119.305 28.250 119.350 ;
        RECT 29.530 119.305 29.820 119.350 ;
        RECT 51.620 119.490 51.910 119.535 ;
        RECT 53.720 119.490 54.010 119.535 ;
        RECT 55.290 119.490 55.580 119.535 ;
        RECT 51.620 119.350 55.580 119.490 ;
        RECT 51.620 119.305 51.910 119.350 ;
        RECT 53.720 119.305 54.010 119.350 ;
        RECT 55.290 119.305 55.580 119.350 ;
        RECT 59.440 119.490 59.730 119.535 ;
        RECT 61.540 119.490 61.830 119.535 ;
        RECT 63.110 119.490 63.400 119.535 ;
        RECT 59.440 119.350 63.400 119.490 ;
        RECT 59.440 119.305 59.730 119.350 ;
        RECT 61.540 119.305 61.830 119.350 ;
        RECT 63.110 119.305 63.400 119.350 ;
        RECT 25.375 118.965 25.665 119.195 ;
        RECT 26.255 119.150 26.545 119.195 ;
        RECT 27.445 119.150 27.735 119.195 ;
        RECT 29.965 119.150 30.255 119.195 ;
        RECT 26.255 119.010 30.255 119.150 ;
        RECT 26.255 118.965 26.545 119.010 ;
        RECT 27.445 118.965 27.735 119.010 ;
        RECT 29.965 118.965 30.255 119.010 ;
        RECT 52.015 119.150 52.305 119.195 ;
        RECT 53.205 119.150 53.495 119.195 ;
        RECT 55.725 119.150 56.015 119.195 ;
        RECT 52.015 119.010 56.015 119.150 ;
        RECT 52.015 118.965 52.305 119.010 ;
        RECT 53.205 118.965 53.495 119.010 ;
        RECT 55.725 118.965 56.015 119.010 ;
        RECT 59.835 119.150 60.125 119.195 ;
        RECT 61.025 119.150 61.315 119.195 ;
        RECT 63.545 119.150 63.835 119.195 ;
        RECT 59.835 119.010 63.835 119.150 ;
        RECT 65.930 119.150 66.070 119.630 ;
        RECT 69.075 119.150 69.365 119.195 ;
        RECT 65.930 119.010 69.365 119.150 ;
        RECT 59.835 118.965 60.125 119.010 ;
        RECT 61.025 118.965 61.315 119.010 ;
        RECT 63.545 118.965 63.835 119.010 ;
        RECT 69.075 118.965 69.365 119.010 ;
        RECT 23.060 118.610 23.380 118.870 ;
        RECT 23.520 118.810 23.840 118.870 ;
        RECT 23.995 118.810 24.285 118.855 ;
        RECT 23.520 118.670 24.285 118.810 ;
        RECT 23.520 118.610 23.840 118.670 ;
        RECT 23.995 118.625 24.285 118.670 ;
        RECT 24.455 118.625 24.745 118.855 ;
        RECT 35.495 118.810 35.785 118.855 ;
        RECT 32.350 118.670 35.785 118.810 ;
        RECT 20.470 118.470 20.760 118.515 ;
        RECT 22.600 118.470 22.920 118.530 ;
        RECT 20.470 118.330 22.920 118.470 ;
        RECT 20.470 118.285 20.760 118.330 ;
        RECT 22.600 118.270 22.920 118.330 ;
        RECT 14.795 118.130 15.085 118.175 ;
        RECT 16.620 118.130 16.940 118.190 ;
        RECT 14.795 117.990 16.940 118.130 ;
        RECT 14.795 117.945 15.085 117.990 ;
        RECT 16.620 117.930 16.940 117.990 ;
        RECT 23.060 118.130 23.380 118.190 ;
        RECT 24.530 118.130 24.670 118.625 ;
        RECT 24.900 118.470 25.220 118.530 ;
        RECT 26.600 118.470 26.890 118.515 ;
        RECT 24.900 118.330 26.890 118.470 ;
        RECT 24.900 118.270 25.220 118.330 ;
        RECT 26.600 118.285 26.890 118.330 ;
        RECT 23.060 117.990 24.670 118.130 ;
        RECT 29.500 118.130 29.820 118.190 ;
        RECT 32.350 118.175 32.490 118.670 ;
        RECT 35.495 118.625 35.785 118.670 ;
        RECT 39.620 118.610 39.940 118.870 ;
        RECT 48.820 118.810 49.140 118.870 ;
        RECT 51.135 118.810 51.425 118.855 ;
        RECT 56.640 118.810 56.960 118.870 ;
        RECT 60.320 118.855 60.640 118.870 ;
        RECT 58.955 118.810 59.245 118.855 ;
        RECT 60.290 118.810 60.640 118.855 ;
        RECT 48.820 118.670 59.245 118.810 ;
        RECT 60.125 118.670 60.640 118.810 ;
        RECT 48.820 118.610 49.140 118.670 ;
        RECT 51.135 118.625 51.425 118.670 ;
        RECT 56.640 118.610 56.960 118.670 ;
        RECT 58.955 118.625 59.245 118.670 ;
        RECT 60.290 118.625 60.640 118.670 ;
        RECT 60.320 118.610 60.640 118.625 ;
        RECT 67.220 118.810 67.540 118.870 ;
        RECT 69.995 118.810 70.285 118.855 ;
        RECT 70.440 118.810 70.760 118.870 ;
        RECT 67.220 118.670 70.760 118.810 ;
        RECT 67.220 118.610 67.540 118.670 ;
        RECT 69.995 118.625 70.285 118.670 ;
        RECT 70.440 118.610 70.760 118.670 ;
        RECT 71.820 118.610 72.140 118.870 ;
        RECT 52.500 118.515 52.820 118.530 ;
        RECT 52.470 118.285 52.820 118.515 ;
        RECT 52.500 118.270 52.820 118.285 ;
        RECT 64.920 118.470 65.240 118.530 ;
        RECT 70.915 118.470 71.205 118.515 ;
        RECT 64.920 118.330 71.205 118.470 ;
        RECT 64.920 118.270 65.240 118.330 ;
        RECT 70.915 118.285 71.205 118.330 ;
        RECT 71.360 118.270 71.680 118.530 ;
        RECT 32.275 118.130 32.565 118.175 ;
        RECT 29.500 117.990 32.565 118.130 ;
        RECT 23.060 117.930 23.380 117.990 ;
        RECT 29.500 117.930 29.820 117.990 ;
        RECT 32.275 117.945 32.565 117.990 ;
        RECT 32.720 117.930 33.040 118.190 ;
        RECT 36.400 118.130 36.720 118.190 ;
        RECT 36.875 118.130 37.165 118.175 ;
        RECT 36.400 117.990 37.165 118.130 ;
        RECT 36.400 117.930 36.720 117.990 ;
        RECT 36.875 117.945 37.165 117.990 ;
        RECT 55.720 118.130 56.040 118.190 ;
        RECT 58.035 118.130 58.325 118.175 ;
        RECT 55.720 117.990 58.325 118.130 ;
        RECT 55.720 117.930 56.040 117.990 ;
        RECT 58.035 117.945 58.325 117.990 ;
        RECT 11.950 117.310 90.610 117.790 ;
        RECT 24.455 116.925 24.745 117.155 ;
        RECT 37.780 117.110 38.100 117.170 ;
        RECT 38.715 117.110 39.005 117.155 ;
        RECT 37.780 116.970 39.005 117.110 ;
        RECT 22.600 116.770 22.920 116.830 ;
        RECT 24.530 116.770 24.670 116.925 ;
        RECT 37.780 116.910 38.100 116.970 ;
        RECT 38.715 116.925 39.005 116.970 ;
        RECT 55.735 117.110 56.025 117.155 ;
        RECT 58.480 117.110 58.800 117.170 ;
        RECT 55.735 116.970 58.800 117.110 ;
        RECT 55.735 116.925 56.025 116.970 ;
        RECT 58.480 116.910 58.800 116.970 ;
        RECT 64.920 116.910 65.240 117.170 ;
        RECT 66.760 117.110 67.080 117.170 ;
        RECT 67.695 117.110 67.985 117.155 ;
        RECT 66.760 116.970 67.985 117.110 ;
        RECT 66.760 116.910 67.080 116.970 ;
        RECT 67.695 116.925 67.985 116.970 ;
        RECT 22.600 116.630 24.670 116.770 ;
        RECT 25.295 116.770 25.585 116.815 ;
        RECT 25.820 116.770 26.140 116.830 ;
        RECT 25.295 116.630 26.140 116.770 ;
        RECT 22.600 116.570 22.920 116.630 ;
        RECT 25.295 116.585 25.585 116.630 ;
        RECT 25.820 116.570 26.140 116.630 ;
        RECT 26.295 116.770 26.585 116.815 ;
        RECT 32.720 116.770 33.040 116.830 ;
        RECT 37.870 116.770 38.010 116.910 ;
        RECT 26.295 116.630 33.040 116.770 ;
        RECT 26.295 116.585 26.585 116.630 ;
        RECT 32.720 116.570 33.040 116.630 ;
        RECT 36.030 116.630 38.010 116.770 ;
        RECT 10.640 116.430 10.960 116.490 ;
        RECT 13.875 116.430 14.165 116.475 ;
        RECT 10.640 116.290 14.165 116.430 ;
        RECT 10.640 116.230 10.960 116.290 ;
        RECT 13.875 116.245 14.165 116.290 ;
        RECT 23.520 116.230 23.840 116.490 ;
        RECT 23.995 116.430 24.285 116.475 ;
        RECT 26.755 116.430 27.045 116.475 ;
        RECT 23.995 116.290 27.045 116.430 ;
        RECT 23.995 116.245 24.285 116.290 ;
        RECT 26.755 116.245 27.045 116.290 ;
        RECT 30.420 116.230 30.740 116.490 ;
        RECT 36.030 116.475 36.170 116.630 ;
        RECT 31.355 116.245 31.645 116.475 ;
        RECT 35.955 116.245 36.245 116.475 ;
        RECT 23.610 116.090 23.750 116.230 ;
        RECT 25.820 116.090 26.140 116.150 ;
        RECT 23.610 115.950 26.140 116.090 ;
        RECT 25.820 115.890 26.140 115.950 ;
        RECT 29.975 116.090 30.265 116.135 ;
        RECT 30.895 116.090 31.185 116.135 ;
        RECT 29.975 115.950 31.185 116.090 ;
        RECT 29.975 115.905 30.265 115.950 ;
        RECT 30.895 115.905 31.185 115.950 ;
        RECT 14.795 115.750 15.085 115.795 ;
        RECT 15.240 115.750 15.560 115.810 ;
        RECT 14.795 115.610 15.560 115.750 ;
        RECT 14.795 115.565 15.085 115.610 ;
        RECT 15.240 115.550 15.560 115.610 ;
        RECT 22.615 115.750 22.905 115.795 ;
        RECT 24.900 115.750 25.220 115.810 ;
        RECT 22.615 115.610 25.220 115.750 ;
        RECT 22.615 115.565 22.905 115.610 ;
        RECT 24.900 115.550 25.220 115.610 ;
        RECT 29.500 115.750 29.820 115.810 ;
        RECT 31.430 115.750 31.570 116.245 ;
        RECT 35.480 115.890 35.800 116.150 ;
        RECT 29.500 115.610 31.570 115.750 ;
        RECT 29.500 115.550 29.820 115.610 ;
        RECT 36.030 115.470 36.170 116.245 ;
        RECT 36.400 116.230 36.720 116.490 ;
        RECT 38.715 116.245 39.005 116.475 ;
        RECT 39.160 116.430 39.480 116.490 ;
        RECT 39.635 116.430 39.925 116.475 ;
        RECT 40.540 116.430 40.860 116.490 ;
        RECT 39.160 116.290 40.860 116.430 ;
        RECT 36.875 115.905 37.165 116.135 ;
        RECT 38.790 116.090 38.930 116.245 ;
        RECT 39.160 116.230 39.480 116.290 ;
        RECT 39.635 116.245 39.925 116.290 ;
        RECT 40.540 116.230 40.860 116.290 ;
        RECT 42.840 116.430 43.160 116.490 ;
        RECT 43.760 116.430 44.080 116.490 ;
        RECT 42.840 116.290 44.080 116.430 ;
        RECT 42.840 116.230 43.160 116.290 ;
        RECT 43.760 116.230 44.080 116.290 ;
        RECT 44.695 116.245 44.985 116.475 ;
        RECT 40.080 116.090 40.400 116.150 ;
        RECT 38.790 115.950 40.400 116.090 ;
        RECT 36.950 115.750 37.090 115.905 ;
        RECT 40.080 115.890 40.400 115.950 ;
        RECT 41.460 115.750 41.780 115.810 ;
        RECT 36.950 115.610 41.780 115.750 ;
        RECT 41.460 115.550 41.780 115.610 ;
        RECT 43.760 115.750 44.080 115.810 ;
        RECT 44.770 115.750 44.910 116.245 ;
        RECT 48.820 116.230 49.140 116.490 ;
        RECT 50.200 116.475 50.520 116.490 ;
        RECT 50.170 116.245 50.520 116.475 ;
        RECT 50.200 116.230 50.520 116.245 ;
        RECT 64.460 116.230 64.780 116.490 ;
        RECT 65.395 116.430 65.685 116.475 ;
        RECT 66.850 116.430 66.990 116.910 ;
        RECT 100.010 116.810 100.780 120.360 ;
        RECT 102.460 119.310 105.310 120.430 ;
        RECT 105.700 120.130 106.050 120.880 ;
        RECT 106.800 120.760 108.670 120.920 ;
        RECT 106.800 120.710 107.560 120.760 ;
        RECT 108.440 120.690 108.670 120.760 ;
        RECT 117.080 120.690 117.310 120.920 ;
        RECT 108.875 120.410 116.875 120.640 ;
        RECT 105.700 120.070 105.990 120.130 ;
        RECT 105.610 119.950 105.990 120.070 ;
        RECT 108.970 120.010 116.830 120.410 ;
        RECT 117.640 120.010 118.600 129.490 ;
        RECT 119.930 129.680 120.770 131.810 ;
        RECT 126.430 131.390 127.680 131.830 ;
        RECT 137.600 131.810 138.460 133.870 ;
        RECT 124.370 131.380 129.610 131.390 ;
        RECT 121.420 131.280 136.720 131.380 ;
        RECT 121.420 131.270 136.755 131.280 ;
        RECT 121.380 131.150 136.755 131.270 ;
        RECT 121.380 131.040 125.380 131.150 ;
        RECT 126.430 131.070 128.170 131.150 ;
        RECT 128.750 131.070 136.755 131.150 ;
        RECT 126.430 130.990 127.680 131.070 ;
        RECT 128.755 131.050 136.755 131.070 ;
        RECT 120.990 130.740 121.220 130.990 ;
        RECT 125.540 130.850 125.770 130.990 ;
        RECT 128.320 130.850 128.550 131.000 ;
        RECT 125.540 130.740 128.550 130.850 ;
        RECT 136.960 130.740 137.190 131.000 ;
        RECT 120.990 130.300 137.190 130.740 ;
        RECT 120.990 130.030 121.220 130.300 ;
        RECT 125.540 130.270 137.190 130.300 ;
        RECT 125.540 130.180 128.550 130.270 ;
        RECT 125.540 130.030 125.770 130.180 ;
        RECT 128.320 130.040 128.550 130.180 ;
        RECT 136.960 130.040 137.190 130.270 ;
        RECT 121.380 129.750 125.380 129.980 ;
        RECT 128.755 129.770 136.755 129.990 ;
        RECT 137.520 129.770 138.480 131.810 ;
        RECT 128.755 129.760 138.480 129.770 ;
        RECT 121.380 129.680 125.370 129.750 ;
        RECT 119.930 129.570 125.370 129.680 ;
        RECT 128.810 129.600 138.480 129.760 ;
        RECT 119.930 129.480 123.060 129.570 ;
        RECT 136.550 129.550 138.480 129.600 ;
        RECT 119.930 126.210 120.770 129.480 ;
        RECT 124.410 129.020 129.660 129.030 ;
        RECT 124.410 128.910 136.720 129.020 ;
        RECT 121.440 128.850 136.720 128.910 ;
        RECT 121.440 128.840 136.755 128.850 ;
        RECT 121.380 128.710 136.755 128.840 ;
        RECT 121.380 128.700 126.540 128.710 ;
        RECT 121.380 128.610 125.380 128.700 ;
        RECT 128.755 128.620 136.755 128.710 ;
        RECT 128.840 128.610 136.730 128.620 ;
        RECT 120.990 128.250 121.220 128.560 ;
        RECT 121.440 128.250 125.340 128.610 ;
        RECT 125.540 128.250 125.770 128.560 ;
        RECT 120.990 126.910 125.770 128.250 ;
        RECT 120.990 126.600 121.220 126.910 ;
        RECT 125.540 126.600 125.770 126.910 ;
        RECT 128.320 128.030 128.550 128.570 ;
        RECT 129.360 128.030 130.370 128.060 ;
        RECT 136.960 128.030 137.190 128.570 ;
        RECT 128.320 127.130 137.190 128.030 ;
        RECT 128.320 126.610 128.550 127.130 ;
        RECT 129.360 127.060 130.370 127.130 ;
        RECT 136.960 126.610 137.190 127.130 ;
        RECT 121.380 126.320 125.380 126.550 ;
        RECT 128.755 126.330 136.755 126.560 ;
        RECT 119.930 126.170 121.060 126.210 ;
        RECT 119.930 126.090 121.300 126.170 ;
        RECT 121.670 126.100 125.330 126.320 ;
        RECT 121.670 126.090 123.110 126.100 ;
        RECT 119.930 126.050 123.110 126.090 ;
        RECT 119.930 125.960 122.620 126.050 ;
        RECT 128.820 126.040 136.710 126.330 ;
        RECT 119.930 125.900 121.950 125.960 ;
        RECT 119.930 125.850 121.700 125.900 ;
        RECT 119.930 122.510 120.770 125.850 ;
        RECT 128.810 125.550 136.730 125.560 ;
        RECT 125.040 125.540 136.730 125.550 ;
        RECT 121.420 125.420 136.730 125.540 ;
        RECT 121.420 125.410 136.755 125.420 ;
        RECT 121.380 125.290 136.755 125.410 ;
        RECT 121.380 125.180 125.380 125.290 ;
        RECT 120.990 124.840 121.220 125.130 ;
        RECT 121.440 124.840 125.330 125.180 ;
        RECT 125.540 124.840 125.770 125.130 ;
        RECT 120.990 123.470 125.770 124.840 ;
        RECT 120.990 123.170 121.220 123.470 ;
        RECT 125.540 123.170 125.770 123.470 ;
        RECT 121.380 122.890 125.380 123.120 ;
        RECT 121.630 122.660 125.200 122.890 ;
        RECT 121.630 122.510 125.320 122.660 ;
        RECT 119.930 122.230 125.320 122.510 ;
        RECT 126.570 122.340 127.190 125.290 ;
        RECT 128.755 125.190 136.755 125.290 ;
        RECT 128.810 125.180 136.730 125.190 ;
        RECT 128.320 124.480 128.550 125.140 ;
        RECT 129.330 124.480 130.330 124.570 ;
        RECT 136.960 124.480 137.190 125.140 ;
        RECT 128.320 123.660 137.190 124.480 ;
        RECT 128.320 123.180 128.550 123.660 ;
        RECT 129.330 123.570 130.330 123.660 ;
        RECT 136.960 123.180 137.190 123.660 ;
        RECT 128.755 122.900 136.755 123.130 ;
        RECT 119.930 121.770 125.330 122.230 ;
        RECT 119.930 120.430 121.930 121.770 ;
        RECT 123.680 121.760 125.330 121.770 ;
        RECT 122.370 120.490 123.370 121.210 ;
        RECT 123.680 120.950 123.990 121.760 ;
        RECT 124.450 121.480 125.330 121.760 ;
        RECT 125.570 121.940 127.190 122.340 ;
        RECT 128.840 121.990 136.710 122.900 ;
        RECT 124.390 121.250 125.390 121.480 ;
        RECT 125.570 121.290 125.920 121.940 ;
        RECT 126.570 121.930 127.190 121.940 ;
        RECT 128.755 121.760 136.755 121.990 ;
        RECT 128.840 121.750 136.710 121.760 ;
        RECT 124.450 121.040 125.330 121.060 ;
        RECT 123.720 120.660 123.990 120.950 ;
        RECT 124.390 120.810 125.390 121.040 ;
        RECT 125.550 121.000 125.920 121.290 ;
        RECT 125.580 120.940 125.920 121.000 ;
        RECT 126.680 121.610 127.440 121.660 ;
        RECT 128.320 121.610 128.550 121.710 ;
        RECT 126.680 121.400 128.550 121.610 ;
        RECT 136.960 121.400 137.190 121.710 ;
        RECT 126.680 120.980 129.220 121.400 ;
        RECT 136.590 120.980 137.190 121.400 ;
        RECT 124.450 120.660 125.330 120.810 ;
        RECT 124.460 120.490 125.190 120.660 ;
        RECT 102.400 119.080 105.400 119.310 ;
        RECT 105.610 119.120 105.950 119.950 ;
        RECT 107.960 119.940 118.600 120.010 ;
        RECT 102.450 119.050 105.310 119.080 ;
        RECT 102.450 119.030 103.620 119.050 ;
        RECT 104.580 119.040 105.310 119.050 ;
        RECT 102.400 118.640 105.400 118.870 ;
        RECT 105.605 118.830 105.950 119.120 ;
        RECT 106.140 118.900 118.600 119.940 ;
        RECT 120.000 120.420 121.930 120.430 ;
        RECT 106.140 118.880 118.560 118.900 ;
        RECT 105.610 118.720 105.950 118.830 ;
        RECT 106.180 118.870 111.850 118.880 ;
        RECT 112.850 118.870 118.560 118.880 ;
        RECT 102.490 118.470 105.350 118.640 ;
        RECT 106.180 118.470 106.610 118.870 ;
        RECT 102.460 118.100 106.610 118.470 ;
        RECT 100.000 116.780 100.780 116.810 ;
        RECT 65.395 116.290 66.990 116.430 ;
        RECT 65.395 116.245 65.685 116.290 ;
        RECT 48.360 115.890 48.680 116.150 ;
        RECT 49.715 116.090 50.005 116.135 ;
        RECT 50.905 116.090 51.195 116.135 ;
        RECT 53.425 116.090 53.715 116.135 ;
        RECT 49.715 115.950 53.715 116.090 ;
        RECT 49.715 115.905 50.005 115.950 ;
        RECT 50.905 115.905 51.195 115.950 ;
        RECT 53.425 115.905 53.715 115.950 ;
        RECT 45.155 115.750 45.445 115.795 ;
        RECT 43.760 115.610 45.445 115.750 ;
        RECT 43.760 115.550 44.080 115.610 ;
        RECT 45.155 115.565 45.445 115.610 ;
        RECT 49.320 115.750 49.610 115.795 ;
        RECT 51.420 115.750 51.710 115.795 ;
        RECT 52.990 115.750 53.280 115.795 ;
        RECT 49.320 115.610 53.280 115.750 ;
        RECT 66.850 115.750 66.990 116.290 ;
        RECT 67.220 116.230 67.540 116.490 ;
        RECT 68.155 116.430 68.445 116.475 ;
        RECT 68.600 116.430 68.920 116.490 ;
        RECT 68.155 116.290 68.920 116.430 ;
        RECT 68.155 116.245 68.445 116.290 ;
        RECT 68.600 116.230 68.920 116.290 ;
        RECT 87.000 116.430 87.320 116.490 ;
        RECT 87.475 116.430 87.765 116.475 ;
        RECT 87.000 116.290 87.765 116.430 ;
        RECT 87.000 116.230 87.320 116.290 ;
        RECT 87.475 116.245 87.765 116.290 ;
        RECT 70.440 116.090 70.760 116.150 ;
        RECT 70.915 116.090 71.205 116.135 ;
        RECT 70.440 115.950 71.205 116.090 ;
        RECT 70.440 115.890 70.760 115.950 ;
        RECT 70.915 115.905 71.205 115.950 ;
        RECT 72.295 115.750 72.585 115.795 ;
        RECT 66.850 115.610 72.585 115.750 ;
        RECT 49.320 115.565 49.610 115.610 ;
        RECT 51.420 115.565 51.710 115.610 ;
        RECT 52.990 115.565 53.280 115.610 ;
        RECT 72.295 115.565 72.585 115.610 ;
        RECT 88.380 115.550 88.700 115.810 ;
        RECT 25.375 115.410 25.665 115.455 ;
        RECT 30.420 115.410 30.740 115.470 ;
        RECT 25.375 115.270 30.740 115.410 ;
        RECT 25.375 115.225 25.665 115.270 ;
        RECT 30.420 115.210 30.740 115.270 ;
        RECT 34.560 115.210 34.880 115.470 ;
        RECT 35.940 115.210 36.260 115.470 ;
        RECT 42.380 115.410 42.700 115.470 ;
        RECT 43.315 115.410 43.605 115.455 ;
        RECT 42.380 115.270 43.605 115.410 ;
        RECT 42.380 115.210 42.700 115.270 ;
        RECT 43.315 115.225 43.605 115.270 ;
        RECT 44.220 115.210 44.540 115.470 ;
        RECT 73.215 115.410 73.505 115.455 ;
        RECT 77.800 115.410 78.120 115.470 ;
        RECT 73.215 115.270 78.120 115.410 ;
        RECT 73.215 115.225 73.505 115.270 ;
        RECT 77.800 115.210 78.120 115.270 ;
        RECT 11.950 114.590 90.610 115.070 ;
        RECT 100.000 114.680 100.830 116.780 ;
        RECT 106.500 116.390 107.750 116.830 ;
        RECT 117.700 116.810 118.560 118.870 ;
        RECT 120.000 116.810 120.770 120.420 ;
        RECT 122.340 119.370 125.190 120.490 ;
        RECT 125.580 120.190 125.930 120.940 ;
        RECT 126.680 120.820 128.550 120.980 ;
        RECT 126.680 120.770 127.440 120.820 ;
        RECT 128.320 120.750 128.550 120.820 ;
        RECT 136.960 120.750 137.190 120.980 ;
        RECT 128.755 120.470 136.755 120.700 ;
        RECT 125.580 120.130 125.870 120.190 ;
        RECT 125.490 120.010 125.870 120.130 ;
        RECT 128.850 120.070 136.710 120.470 ;
        RECT 137.520 120.070 138.480 129.550 ;
        RECT 122.280 119.140 125.280 119.370 ;
        RECT 125.490 119.180 125.830 120.010 ;
        RECT 127.840 120.000 138.480 120.070 ;
        RECT 122.330 119.110 125.190 119.140 ;
        RECT 122.330 119.090 123.500 119.110 ;
        RECT 124.460 119.100 125.190 119.110 ;
        RECT 122.280 118.700 125.280 118.930 ;
        RECT 125.485 118.890 125.830 119.180 ;
        RECT 126.020 118.960 138.480 120.000 ;
        RECT 139.930 131.780 140.700 135.360 ;
        RECT 142.370 134.310 145.220 135.430 ;
        RECT 145.610 135.130 145.960 135.880 ;
        RECT 146.710 135.760 148.580 135.920 ;
        RECT 146.710 135.710 147.470 135.760 ;
        RECT 148.350 135.690 148.580 135.760 ;
        RECT 156.990 135.690 157.220 135.920 ;
        RECT 148.785 135.410 156.785 135.640 ;
        RECT 145.610 135.070 145.900 135.130 ;
        RECT 145.520 134.950 145.900 135.070 ;
        RECT 148.880 135.010 156.740 135.410 ;
        RECT 157.550 135.010 158.510 144.490 ;
        RECT 142.310 134.080 145.310 134.310 ;
        RECT 145.520 134.120 145.860 134.950 ;
        RECT 147.870 134.940 158.510 135.010 ;
        RECT 142.360 134.050 145.220 134.080 ;
        RECT 142.360 134.030 143.530 134.050 ;
        RECT 144.490 134.040 145.220 134.050 ;
        RECT 142.310 133.640 145.310 133.870 ;
        RECT 145.515 133.830 145.860 134.120 ;
        RECT 146.050 133.900 158.510 134.940 ;
        RECT 146.050 133.880 158.500 133.900 ;
        RECT 145.520 133.720 145.860 133.830 ;
        RECT 146.090 133.870 151.760 133.880 ;
        RECT 152.760 133.870 158.500 133.880 ;
        RECT 142.400 133.470 145.260 133.640 ;
        RECT 146.090 133.470 146.520 133.870 ;
        RECT 142.370 133.100 146.520 133.470 ;
        RECT 139.930 129.680 140.790 131.780 ;
        RECT 146.460 131.390 147.710 131.830 ;
        RECT 157.640 131.810 158.500 133.870 ;
        RECT 144.400 131.380 149.640 131.390 ;
        RECT 141.450 131.280 156.750 131.380 ;
        RECT 141.450 131.270 156.785 131.280 ;
        RECT 141.410 131.150 156.785 131.270 ;
        RECT 141.410 131.040 145.410 131.150 ;
        RECT 146.460 131.070 148.200 131.150 ;
        RECT 148.780 131.070 156.785 131.150 ;
        RECT 146.460 130.990 147.710 131.070 ;
        RECT 148.785 131.050 156.785 131.070 ;
        RECT 141.020 130.740 141.250 130.990 ;
        RECT 145.570 130.850 145.800 130.990 ;
        RECT 148.350 130.850 148.580 131.000 ;
        RECT 145.570 130.740 148.580 130.850 ;
        RECT 156.990 130.740 157.220 131.000 ;
        RECT 141.020 130.300 157.220 130.740 ;
        RECT 141.020 130.030 141.250 130.300 ;
        RECT 145.570 130.270 157.220 130.300 ;
        RECT 145.570 130.180 148.580 130.270 ;
        RECT 145.570 130.030 145.800 130.180 ;
        RECT 148.350 130.040 148.580 130.180 ;
        RECT 156.990 130.040 157.220 130.270 ;
        RECT 141.410 129.750 145.410 129.980 ;
        RECT 148.785 129.770 156.785 129.990 ;
        RECT 157.550 129.770 158.510 131.810 ;
        RECT 148.785 129.760 158.510 129.770 ;
        RECT 141.410 129.680 145.400 129.750 ;
        RECT 139.930 129.570 145.400 129.680 ;
        RECT 148.840 129.600 158.510 129.760 ;
        RECT 139.930 129.480 143.090 129.570 ;
        RECT 156.580 129.550 158.510 129.600 ;
        RECT 139.930 126.210 140.790 129.480 ;
        RECT 144.440 129.020 149.690 129.030 ;
        RECT 144.440 128.910 156.750 129.020 ;
        RECT 141.470 128.850 156.750 128.910 ;
        RECT 141.470 128.840 156.785 128.850 ;
        RECT 141.410 128.710 156.785 128.840 ;
        RECT 141.410 128.700 146.570 128.710 ;
        RECT 141.410 128.610 145.410 128.700 ;
        RECT 148.785 128.620 156.785 128.710 ;
        RECT 148.870 128.610 156.760 128.620 ;
        RECT 141.020 128.250 141.250 128.560 ;
        RECT 141.470 128.250 145.370 128.610 ;
        RECT 145.570 128.250 145.800 128.560 ;
        RECT 141.020 126.910 145.800 128.250 ;
        RECT 141.020 126.600 141.250 126.910 ;
        RECT 145.570 126.600 145.800 126.910 ;
        RECT 148.350 128.030 148.580 128.570 ;
        RECT 149.390 128.030 150.400 128.060 ;
        RECT 156.990 128.030 157.220 128.570 ;
        RECT 148.350 127.130 157.220 128.030 ;
        RECT 148.350 126.610 148.580 127.130 ;
        RECT 149.390 127.060 150.400 127.130 ;
        RECT 156.990 126.610 157.220 127.130 ;
        RECT 141.410 126.320 145.410 126.550 ;
        RECT 148.785 126.330 156.785 126.560 ;
        RECT 139.930 126.170 141.090 126.210 ;
        RECT 139.930 126.090 141.330 126.170 ;
        RECT 141.700 126.100 145.360 126.320 ;
        RECT 141.700 126.090 143.140 126.100 ;
        RECT 139.930 126.050 143.140 126.090 ;
        RECT 139.930 125.960 142.650 126.050 ;
        RECT 148.850 126.040 156.740 126.330 ;
        RECT 139.930 125.900 141.980 125.960 ;
        RECT 139.930 125.850 141.730 125.900 ;
        RECT 139.930 122.510 140.790 125.850 ;
        RECT 148.840 125.550 156.760 125.560 ;
        RECT 145.070 125.540 156.760 125.550 ;
        RECT 141.450 125.420 156.760 125.540 ;
        RECT 141.450 125.410 156.785 125.420 ;
        RECT 141.410 125.290 156.785 125.410 ;
        RECT 141.410 125.180 145.410 125.290 ;
        RECT 141.020 124.840 141.250 125.130 ;
        RECT 141.470 124.840 145.360 125.180 ;
        RECT 145.570 124.840 145.800 125.130 ;
        RECT 141.020 123.470 145.800 124.840 ;
        RECT 141.020 123.170 141.250 123.470 ;
        RECT 145.570 123.170 145.800 123.470 ;
        RECT 141.410 122.890 145.410 123.120 ;
        RECT 141.660 122.660 145.230 122.890 ;
        RECT 141.660 122.510 145.350 122.660 ;
        RECT 139.930 122.230 145.350 122.510 ;
        RECT 146.600 122.340 147.220 125.290 ;
        RECT 148.785 125.190 156.785 125.290 ;
        RECT 148.840 125.180 156.760 125.190 ;
        RECT 148.350 124.480 148.580 125.140 ;
        RECT 149.360 124.480 150.360 124.570 ;
        RECT 156.990 124.480 157.220 125.140 ;
        RECT 148.350 123.660 157.220 124.480 ;
        RECT 148.350 123.180 148.580 123.660 ;
        RECT 149.360 123.570 150.360 123.660 ;
        RECT 156.990 123.180 157.220 123.660 ;
        RECT 148.785 122.900 156.785 123.130 ;
        RECT 139.930 121.770 145.360 122.230 ;
        RECT 139.930 120.420 141.960 121.770 ;
        RECT 143.710 121.760 145.360 121.770 ;
        RECT 142.400 120.490 143.400 121.210 ;
        RECT 143.710 120.950 144.020 121.760 ;
        RECT 144.480 121.480 145.360 121.760 ;
        RECT 145.600 121.940 147.220 122.340 ;
        RECT 148.870 121.990 156.740 122.900 ;
        RECT 144.420 121.250 145.420 121.480 ;
        RECT 145.600 121.290 145.950 121.940 ;
        RECT 146.600 121.930 147.220 121.940 ;
        RECT 148.785 121.760 156.785 121.990 ;
        RECT 148.870 121.750 156.740 121.760 ;
        RECT 144.480 121.040 145.360 121.060 ;
        RECT 143.750 120.660 144.020 120.950 ;
        RECT 144.420 120.810 145.420 121.040 ;
        RECT 145.580 121.000 145.950 121.290 ;
        RECT 145.610 120.940 145.950 121.000 ;
        RECT 146.710 121.610 147.470 121.660 ;
        RECT 148.350 121.610 148.580 121.710 ;
        RECT 146.710 121.400 148.580 121.610 ;
        RECT 156.990 121.400 157.220 121.710 ;
        RECT 146.710 120.980 149.250 121.400 ;
        RECT 156.620 120.980 157.220 121.400 ;
        RECT 144.480 120.660 145.360 120.810 ;
        RECT 144.490 120.490 145.220 120.660 ;
        RECT 126.020 118.940 138.460 118.960 ;
        RECT 125.490 118.780 125.830 118.890 ;
        RECT 126.060 118.930 131.730 118.940 ;
        RECT 132.730 118.930 138.460 118.940 ;
        RECT 122.370 118.530 125.230 118.700 ;
        RECT 126.060 118.530 126.490 118.930 ;
        RECT 122.340 118.160 126.490 118.530 ;
        RECT 104.440 116.380 109.680 116.390 ;
        RECT 101.490 116.280 116.790 116.380 ;
        RECT 101.490 116.270 116.825 116.280 ;
        RECT 101.450 116.150 116.825 116.270 ;
        RECT 101.450 116.040 105.450 116.150 ;
        RECT 106.500 116.070 108.240 116.150 ;
        RECT 108.820 116.070 116.825 116.150 ;
        RECT 106.500 115.990 107.750 116.070 ;
        RECT 108.825 116.050 116.825 116.070 ;
        RECT 101.060 115.740 101.290 115.990 ;
        RECT 105.610 115.850 105.840 115.990 ;
        RECT 108.390 115.850 108.620 116.000 ;
        RECT 105.610 115.740 108.620 115.850 ;
        RECT 117.030 115.740 117.260 116.000 ;
        RECT 101.060 115.300 117.260 115.740 ;
        RECT 101.060 115.030 101.290 115.300 ;
        RECT 105.610 115.270 117.260 115.300 ;
        RECT 105.610 115.180 108.620 115.270 ;
        RECT 105.610 115.030 105.840 115.180 ;
        RECT 108.390 115.040 108.620 115.180 ;
        RECT 117.030 115.040 117.260 115.270 ;
        RECT 101.450 114.750 105.450 114.980 ;
        RECT 108.825 114.770 116.825 114.990 ;
        RECT 117.590 114.770 118.560 116.810 ;
        RECT 108.825 114.760 118.560 114.770 ;
        RECT 101.450 114.680 105.440 114.750 ;
        RECT 100.000 114.570 105.440 114.680 ;
        RECT 108.880 114.600 118.560 114.760 ;
        RECT 100.000 114.480 103.130 114.570 ;
        RECT 116.620 114.550 118.560 114.600 ;
        RECT 55.735 114.390 56.025 114.435 ;
        RECT 56.180 114.390 56.500 114.450 ;
        RECT 55.735 114.250 56.500 114.390 ;
        RECT 55.735 114.205 56.025 114.250 ;
        RECT 56.180 114.190 56.500 114.250 ;
        RECT 87.000 114.190 87.320 114.450 ;
        RECT 33.680 114.050 33.970 114.095 ;
        RECT 35.780 114.050 36.070 114.095 ;
        RECT 37.350 114.050 37.640 114.095 ;
        RECT 33.680 113.910 37.640 114.050 ;
        RECT 33.680 113.865 33.970 113.910 ;
        RECT 35.780 113.865 36.070 113.910 ;
        RECT 37.350 113.865 37.640 113.910 ;
        RECT 43.800 114.050 44.090 114.095 ;
        RECT 45.900 114.050 46.190 114.095 ;
        RECT 47.470 114.050 47.760 114.095 ;
        RECT 43.800 113.910 47.760 114.050 ;
        RECT 43.800 113.865 44.090 113.910 ;
        RECT 45.900 113.865 46.190 113.910 ;
        RECT 47.470 113.865 47.760 113.910 ;
        RECT 48.360 114.050 48.680 114.110 ;
        RECT 50.215 114.050 50.505 114.095 ;
        RECT 48.360 113.910 50.505 114.050 ;
        RECT 48.360 113.850 48.680 113.910 ;
        RECT 50.215 113.865 50.505 113.910 ;
        RECT 57.600 114.050 57.890 114.095 ;
        RECT 59.700 114.050 59.990 114.095 ;
        RECT 61.270 114.050 61.560 114.095 ;
        RECT 57.600 113.910 61.560 114.050 ;
        RECT 57.600 113.865 57.890 113.910 ;
        RECT 59.700 113.865 59.990 113.910 ;
        RECT 61.270 113.865 61.560 113.910 ;
        RECT 68.600 113.850 68.920 114.110 ;
        RECT 71.360 114.050 71.650 114.095 ;
        RECT 72.930 114.050 73.220 114.095 ;
        RECT 75.030 114.050 75.320 114.095 ;
        RECT 71.360 113.910 75.320 114.050 ;
        RECT 71.360 113.865 71.650 113.910 ;
        RECT 72.930 113.865 73.220 113.910 ;
        RECT 75.030 113.865 75.320 113.910 ;
        RECT 34.075 113.710 34.365 113.755 ;
        RECT 35.265 113.710 35.555 113.755 ;
        RECT 37.785 113.710 38.075 113.755 ;
        RECT 34.075 113.570 38.075 113.710 ;
        RECT 34.075 113.525 34.365 113.570 ;
        RECT 35.265 113.525 35.555 113.570 ;
        RECT 37.785 113.525 38.075 113.570 ;
        RECT 43.300 113.510 43.620 113.770 ;
        RECT 44.195 113.710 44.485 113.755 ;
        RECT 45.385 113.710 45.675 113.755 ;
        RECT 47.905 113.710 48.195 113.755 ;
        RECT 44.195 113.570 48.195 113.710 ;
        RECT 44.195 113.525 44.485 113.570 ;
        RECT 45.385 113.525 45.675 113.570 ;
        RECT 47.905 113.525 48.195 113.570 ;
        RECT 10.640 113.370 10.960 113.430 ;
        RECT 13.415 113.370 13.705 113.415 ;
        RECT 10.640 113.230 13.705 113.370 ;
        RECT 10.640 113.170 10.960 113.230 ;
        RECT 13.415 113.185 13.705 113.230 ;
        RECT 14.795 113.370 15.085 113.415 ;
        RECT 15.700 113.370 16.020 113.430 ;
        RECT 20.300 113.370 20.620 113.430 ;
        RECT 20.775 113.370 21.065 113.415 ;
        RECT 14.795 113.230 19.150 113.370 ;
        RECT 14.795 113.185 15.085 113.230 ;
        RECT 15.700 113.170 16.020 113.230 ;
        RECT 6.960 113.030 7.280 113.090 ;
        RECT 19.010 113.030 19.150 113.230 ;
        RECT 20.300 113.230 21.065 113.370 ;
        RECT 20.300 113.170 20.620 113.230 ;
        RECT 20.775 113.185 21.065 113.230 ;
        RECT 21.680 113.370 22.000 113.430 ;
        RECT 29.960 113.370 30.280 113.430 ;
        RECT 33.195 113.370 33.485 113.415 ;
        RECT 21.680 113.230 33.485 113.370 ;
        RECT 21.680 113.170 22.000 113.230 ;
        RECT 29.960 113.170 30.280 113.230 ;
        RECT 33.195 113.185 33.485 113.230 ;
        RECT 34.190 113.230 41.230 113.370 ;
        RECT 25.360 113.030 25.680 113.090 ;
        RECT 34.190 113.030 34.330 113.230 ;
        RECT 6.960 112.890 18.690 113.030 ;
        RECT 19.010 112.890 34.330 113.030 ;
        RECT 34.530 113.030 34.820 113.075 ;
        RECT 40.555 113.030 40.845 113.075 ;
        RECT 34.530 112.890 40.845 113.030 ;
        RECT 6.960 112.830 7.280 112.890 ;
        RECT 18.000 112.490 18.320 112.750 ;
        RECT 18.550 112.690 18.690 112.890 ;
        RECT 25.360 112.830 25.680 112.890 ;
        RECT 34.530 112.845 34.820 112.890 ;
        RECT 40.555 112.845 40.845 112.890 ;
        RECT 35.480 112.690 35.800 112.750 ;
        RECT 18.550 112.550 35.800 112.690 ;
        RECT 35.480 112.490 35.800 112.550 ;
        RECT 39.160 112.690 39.480 112.750 ;
        RECT 40.080 112.690 40.400 112.750 ;
        RECT 39.160 112.550 40.400 112.690 ;
        RECT 41.090 112.690 41.230 113.230 ;
        RECT 41.460 113.170 41.780 113.430 ;
        RECT 42.380 113.170 42.700 113.430 ;
        RECT 42.840 113.370 43.160 113.430 ;
        RECT 48.450 113.370 48.590 113.850 ;
        RECT 56.640 113.710 56.960 113.770 ;
        RECT 57.115 113.710 57.405 113.755 ;
        RECT 56.640 113.570 57.405 113.710 ;
        RECT 56.640 113.510 56.960 113.570 ;
        RECT 57.115 113.525 57.405 113.570 ;
        RECT 57.995 113.710 58.285 113.755 ;
        RECT 59.185 113.710 59.475 113.755 ;
        RECT 61.705 113.710 61.995 113.755 ;
        RECT 57.995 113.570 61.995 113.710 ;
        RECT 57.995 113.525 58.285 113.570 ;
        RECT 59.185 113.525 59.475 113.570 ;
        RECT 61.705 113.525 61.995 113.570 ;
        RECT 70.925 113.710 71.215 113.755 ;
        RECT 73.445 113.710 73.735 113.755 ;
        RECT 74.635 113.710 74.925 113.755 ;
        RECT 70.925 113.570 74.925 113.710 ;
        RECT 70.925 113.525 71.215 113.570 ;
        RECT 73.445 113.525 73.735 113.570 ;
        RECT 74.635 113.525 74.925 113.570 ;
        RECT 42.840 113.230 43.340 113.370 ;
        RECT 44.310 113.230 48.590 113.370 ;
        RECT 42.840 113.170 43.160 113.230 ;
        RECT 43.300 113.030 43.620 113.090 ;
        RECT 44.310 113.030 44.450 113.230 ;
        RECT 53.895 113.185 54.185 113.415 ;
        RECT 63.080 113.370 63.400 113.430 ;
        RECT 64.475 113.370 64.765 113.415 ;
        RECT 63.080 113.230 64.765 113.370 ;
        RECT 44.680 113.075 45.000 113.090 ;
        RECT 43.300 112.890 44.450 113.030 ;
        RECT 43.300 112.830 43.620 112.890 ;
        RECT 44.650 112.845 45.000 113.075 ;
        RECT 44.680 112.830 45.000 112.845 ;
        RECT 53.970 112.690 54.110 113.185 ;
        RECT 63.080 113.170 63.400 113.230 ;
        RECT 64.475 113.185 64.765 113.230 ;
        RECT 65.395 113.185 65.685 113.415 ;
        RECT 68.155 113.370 68.445 113.415 ;
        RECT 69.060 113.370 69.380 113.430 ;
        RECT 71.360 113.370 71.680 113.430 ;
        RECT 68.155 113.230 71.680 113.370 ;
        RECT 68.155 113.185 68.445 113.230 ;
        RECT 55.720 112.830 56.040 113.090 ;
        RECT 58.450 113.030 58.740 113.075 ;
        RECT 64.935 113.030 65.225 113.075 ;
        RECT 58.450 112.890 65.225 113.030 ;
        RECT 65.470 113.030 65.610 113.185 ;
        RECT 69.060 113.170 69.380 113.230 ;
        RECT 71.360 113.170 71.680 113.230 ;
        RECT 75.500 113.370 75.820 113.430 ;
        RECT 78.260 113.370 78.580 113.430 ;
        RECT 75.500 113.230 78.580 113.370 ;
        RECT 75.500 113.170 75.820 113.230 ;
        RECT 78.260 113.170 78.580 113.230 ;
        RECT 86.080 113.170 86.400 113.430 ;
        RECT 87.000 113.370 87.320 113.430 ;
        RECT 87.475 113.370 87.765 113.415 ;
        RECT 87.000 113.230 87.765 113.370 ;
        RECT 87.000 113.170 87.320 113.230 ;
        RECT 87.475 113.185 87.765 113.230 ;
        RECT 69.520 113.030 69.840 113.090 ;
        RECT 65.470 112.890 69.840 113.030 ;
        RECT 58.450 112.845 58.740 112.890 ;
        RECT 64.935 112.845 65.225 112.890 ;
        RECT 69.520 112.830 69.840 112.890 ;
        RECT 73.200 113.030 73.520 113.090 ;
        RECT 74.180 113.030 74.470 113.075 ;
        RECT 73.200 112.890 74.470 113.030 ;
        RECT 73.200 112.830 73.520 112.890 ;
        RECT 74.180 112.845 74.470 112.890 ;
        RECT 54.800 112.690 55.120 112.750 ;
        RECT 41.090 112.550 55.120 112.690 ;
        RECT 39.160 112.490 39.480 112.550 ;
        RECT 40.080 112.490 40.400 112.550 ;
        RECT 54.800 112.490 55.120 112.550 ;
        RECT 56.655 112.690 56.945 112.735 ;
        RECT 63.540 112.690 63.860 112.750 ;
        RECT 56.655 112.550 63.860 112.690 ;
        RECT 56.655 112.505 56.945 112.550 ;
        RECT 63.540 112.490 63.860 112.550 ;
        RECT 64.015 112.690 64.305 112.735 ;
        RECT 65.380 112.690 65.700 112.750 ;
        RECT 67.220 112.690 67.540 112.750 ;
        RECT 64.015 112.550 67.540 112.690 ;
        RECT 64.015 112.505 64.305 112.550 ;
        RECT 65.380 112.490 65.700 112.550 ;
        RECT 67.220 112.490 67.540 112.550 ;
        RECT 67.680 112.690 68.000 112.750 ;
        RECT 72.740 112.690 73.060 112.750 ;
        RECT 67.680 112.550 73.060 112.690 ;
        RECT 67.680 112.490 68.000 112.550 ;
        RECT 72.740 112.490 73.060 112.550 ;
        RECT 88.380 112.490 88.700 112.750 ;
        RECT 11.950 111.870 90.610 112.350 ;
        RECT 19.855 111.670 20.145 111.715 ;
        RECT 20.760 111.670 21.080 111.730 ;
        RECT 19.855 111.530 21.080 111.670 ;
        RECT 19.855 111.485 20.145 111.530 ;
        RECT 20.760 111.470 21.080 111.530 ;
        RECT 21.680 111.470 22.000 111.730 ;
        RECT 36.875 111.670 37.165 111.715 ;
        RECT 41.460 111.670 41.780 111.730 ;
        RECT 36.875 111.530 39.390 111.670 ;
        RECT 36.875 111.485 37.165 111.530 ;
        RECT 21.770 111.330 21.910 111.470 ;
        RECT 20.390 111.190 21.910 111.330 ;
        RECT 31.310 111.330 31.600 111.375 ;
        RECT 34.560 111.330 34.880 111.390 ;
        RECT 31.310 111.190 34.880 111.330 ;
        RECT 20.390 111.050 20.530 111.190 ;
        RECT 31.310 111.145 31.600 111.190 ;
        RECT 34.560 111.130 34.880 111.190 ;
        RECT 14.795 110.990 15.085 111.035 ;
        RECT 15.240 110.990 15.560 111.050 ;
        RECT 14.795 110.850 15.560 110.990 ;
        RECT 14.795 110.805 15.085 110.850 ;
        RECT 15.240 110.790 15.560 110.850 ;
        RECT 16.620 110.790 16.940 111.050 ;
        RECT 20.300 110.790 20.620 111.050 ;
        RECT 21.680 111.035 22.000 111.050 ;
        RECT 21.650 110.805 22.000 111.035 ;
        RECT 21.680 110.790 22.000 110.805 ;
        RECT 25.820 110.990 26.140 111.050 ;
        RECT 27.675 110.990 27.965 111.035 ;
        RECT 25.820 110.850 27.965 110.990 ;
        RECT 25.820 110.790 26.140 110.850 ;
        RECT 27.675 110.805 27.965 110.850 ;
        RECT 28.595 110.990 28.885 111.035 ;
        RECT 29.500 110.990 29.820 111.050 ;
        RECT 28.595 110.850 29.820 110.990 ;
        RECT 28.595 110.805 28.885 110.850 ;
        RECT 29.500 110.790 29.820 110.850 ;
        RECT 29.960 110.790 30.280 111.050 ;
        RECT 35.020 110.990 35.340 111.050 ;
        RECT 39.250 111.035 39.390 111.530 ;
        RECT 41.460 111.530 42.610 111.670 ;
        RECT 41.460 111.470 41.780 111.530 ;
        RECT 40.080 111.330 40.400 111.390 ;
        RECT 41.935 111.330 42.225 111.375 ;
        RECT 40.080 111.190 42.225 111.330 ;
        RECT 42.470 111.330 42.610 111.530 ;
        RECT 44.680 111.470 45.000 111.730 ;
        RECT 63.080 111.470 63.400 111.730 ;
        RECT 63.540 111.670 63.860 111.730 ;
        RECT 65.855 111.670 66.145 111.715 ;
        RECT 63.540 111.530 66.145 111.670 ;
        RECT 63.540 111.470 63.860 111.530 ;
        RECT 65.855 111.485 66.145 111.530 ;
        RECT 67.235 111.485 67.525 111.715 ;
        RECT 68.615 111.670 68.905 111.715 ;
        RECT 69.060 111.670 69.380 111.730 ;
        RECT 68.615 111.530 69.380 111.670 ;
        RECT 68.615 111.485 68.905 111.530 ;
        RECT 45.615 111.330 45.905 111.375 ;
        RECT 42.470 111.190 45.905 111.330 ;
        RECT 40.080 111.130 40.400 111.190 ;
        RECT 41.935 111.145 42.225 111.190 ;
        RECT 45.615 111.145 45.905 111.190 ;
        RECT 38.255 110.990 38.545 111.035 ;
        RECT 35.020 110.850 38.545 110.990 ;
        RECT 35.020 110.790 35.340 110.850 ;
        RECT 38.255 110.805 38.545 110.850 ;
        RECT 39.175 110.990 39.465 111.035 ;
        RECT 39.620 110.990 39.940 111.050 ;
        RECT 39.175 110.850 39.940 110.990 ;
        RECT 39.175 110.805 39.465 110.850 ;
        RECT 39.620 110.790 39.940 110.850 ;
        RECT 41.000 110.990 41.320 111.050 ;
        RECT 42.840 110.990 43.160 111.050 ;
        RECT 41.000 110.850 43.160 110.990 ;
        RECT 41.000 110.790 41.320 110.850 ;
        RECT 42.840 110.790 43.160 110.850 ;
        RECT 43.315 110.990 43.605 111.035 ;
        RECT 43.760 110.990 44.080 111.050 ;
        RECT 43.315 110.850 44.080 110.990 ;
        RECT 43.315 110.805 43.605 110.850 ;
        RECT 43.760 110.790 44.080 110.850 ;
        RECT 45.155 110.805 45.445 111.035 ;
        RECT 16.160 110.450 16.480 110.710 ;
        RECT 21.195 110.650 21.485 110.695 ;
        RECT 22.385 110.650 22.675 110.695 ;
        RECT 24.905 110.650 25.195 110.695 ;
        RECT 21.195 110.510 25.195 110.650 ;
        RECT 21.195 110.465 21.485 110.510 ;
        RECT 22.385 110.465 22.675 110.510 ;
        RECT 24.905 110.465 25.195 110.510 ;
        RECT 30.855 110.650 31.145 110.695 ;
        RECT 32.045 110.650 32.335 110.695 ;
        RECT 34.565 110.650 34.855 110.695 ;
        RECT 30.855 110.510 34.855 110.650 ;
        RECT 30.855 110.465 31.145 110.510 ;
        RECT 32.045 110.465 32.335 110.510 ;
        RECT 34.565 110.465 34.855 110.510 ;
        RECT 44.220 110.650 44.540 110.710 ;
        RECT 44.695 110.650 44.985 110.695 ;
        RECT 44.220 110.510 44.985 110.650 ;
        RECT 44.220 110.450 44.540 110.510 ;
        RECT 44.695 110.465 44.985 110.510 ;
        RECT 15.255 110.310 15.545 110.355 ;
        RECT 20.800 110.310 21.090 110.355 ;
        RECT 22.900 110.310 23.190 110.355 ;
        RECT 24.470 110.310 24.760 110.355 ;
        RECT 15.255 110.170 20.300 110.310 ;
        RECT 15.255 110.125 15.545 110.170 ;
        RECT 15.715 109.970 16.005 110.015 ;
        RECT 17.080 109.970 17.400 110.030 ;
        RECT 15.715 109.830 17.400 109.970 ;
        RECT 20.160 109.970 20.300 110.170 ;
        RECT 20.800 110.170 24.760 110.310 ;
        RECT 20.800 110.125 21.090 110.170 ;
        RECT 22.900 110.125 23.190 110.170 ;
        RECT 24.470 110.125 24.760 110.170 ;
        RECT 30.460 110.310 30.750 110.355 ;
        RECT 32.560 110.310 32.850 110.355 ;
        RECT 34.130 110.310 34.420 110.355 ;
        RECT 30.460 110.170 34.420 110.310 ;
        RECT 30.460 110.125 30.750 110.170 ;
        RECT 32.560 110.125 32.850 110.170 ;
        RECT 34.130 110.125 34.420 110.170 ;
        RECT 40.095 110.310 40.385 110.355 ;
        RECT 45.230 110.310 45.370 110.805 ;
        RECT 54.800 110.790 55.120 111.050 ;
        RECT 55.720 110.790 56.040 111.050 ;
        RECT 56.180 110.790 56.500 111.050 ;
        RECT 62.160 110.790 62.480 111.050 ;
        RECT 65.930 110.990 66.070 111.485 ;
        RECT 67.310 111.330 67.450 111.485 ;
        RECT 69.060 111.470 69.380 111.530 ;
        RECT 69.520 111.330 69.840 111.390 ;
        RECT 71.820 111.330 72.140 111.390 ;
        RECT 72.295 111.330 72.585 111.375 ;
        RECT 67.310 111.190 72.585 111.330 ;
        RECT 69.520 111.130 69.840 111.190 ;
        RECT 71.820 111.130 72.140 111.190 ;
        RECT 72.295 111.145 72.585 111.190 ;
        RECT 100.000 111.210 100.830 114.480 ;
        RECT 104.480 114.020 109.730 114.030 ;
        RECT 104.480 113.910 116.790 114.020 ;
        RECT 101.510 113.850 116.790 113.910 ;
        RECT 101.510 113.840 116.825 113.850 ;
        RECT 101.450 113.710 116.825 113.840 ;
        RECT 101.450 113.700 106.610 113.710 ;
        RECT 101.450 113.610 105.450 113.700 ;
        RECT 108.825 113.620 116.825 113.710 ;
        RECT 108.910 113.610 116.800 113.620 ;
        RECT 101.060 113.250 101.290 113.560 ;
        RECT 101.510 113.250 105.410 113.610 ;
        RECT 105.610 113.250 105.840 113.560 ;
        RECT 101.060 111.910 105.840 113.250 ;
        RECT 101.060 111.600 101.290 111.910 ;
        RECT 105.610 111.600 105.840 111.910 ;
        RECT 108.390 113.030 108.620 113.570 ;
        RECT 109.430 113.030 110.440 113.060 ;
        RECT 117.030 113.030 117.260 113.570 ;
        RECT 108.390 112.130 117.260 113.030 ;
        RECT 108.390 111.610 108.620 112.130 ;
        RECT 109.430 112.060 110.440 112.130 ;
        RECT 117.030 111.610 117.260 112.130 ;
        RECT 101.450 111.320 105.450 111.550 ;
        RECT 108.825 111.330 116.825 111.560 ;
        RECT 100.000 111.170 101.130 111.210 ;
        RECT 100.000 111.090 101.370 111.170 ;
        RECT 101.740 111.100 105.400 111.320 ;
        RECT 101.740 111.090 103.180 111.100 ;
        RECT 100.000 111.050 103.180 111.090 ;
        RECT 68.140 110.990 68.460 111.050 ;
        RECT 65.930 110.850 68.460 110.990 ;
        RECT 68.140 110.790 68.460 110.850 ;
        RECT 73.660 110.990 73.980 111.050 ;
        RECT 74.135 110.990 74.425 111.035 ;
        RECT 73.660 110.850 74.425 110.990 ;
        RECT 73.660 110.790 73.980 110.850 ;
        RECT 74.135 110.805 74.425 110.850 ;
        RECT 78.260 110.790 78.580 111.050 ;
        RECT 79.640 111.035 79.960 111.050 ;
        RECT 79.610 110.805 79.960 111.035 ;
        RECT 79.640 110.790 79.960 110.805 ;
        RECT 100.000 110.960 102.690 111.050 ;
        RECT 108.890 111.040 116.780 111.330 ;
        RECT 100.000 110.900 102.020 110.960 ;
        RECT 100.000 110.850 101.770 110.900 ;
        RECT 55.260 110.650 55.580 110.710 ;
        RECT 56.270 110.650 56.410 110.790 ;
        RECT 55.260 110.510 56.410 110.650 ;
        RECT 60.795 110.650 61.085 110.695 ;
        RECT 64.015 110.650 64.305 110.695 ;
        RECT 60.795 110.510 64.305 110.650 ;
        RECT 55.260 110.450 55.580 110.510 ;
        RECT 60.795 110.465 61.085 110.510 ;
        RECT 64.015 110.465 64.305 110.510 ;
        RECT 40.095 110.170 45.370 110.310 ;
        RECT 58.035 110.310 58.325 110.355 ;
        RECT 61.255 110.310 61.545 110.355 ;
        RECT 62.620 110.310 62.940 110.370 ;
        RECT 58.035 110.170 62.940 110.310 ;
        RECT 64.090 110.310 64.230 110.465 ;
        RECT 65.380 110.450 65.700 110.710 ;
        RECT 66.300 110.695 66.620 110.710 ;
        RECT 66.300 110.465 66.730 110.695 ;
        RECT 71.375 110.465 71.665 110.695 ;
        RECT 72.740 110.650 73.060 110.710 ;
        RECT 73.215 110.650 73.505 110.695 ;
        RECT 72.740 110.510 73.505 110.650 ;
        RECT 66.300 110.450 66.620 110.465 ;
        RECT 67.220 110.310 67.540 110.370 ;
        RECT 64.090 110.170 67.540 110.310 ;
        RECT 40.095 110.125 40.385 110.170 ;
        RECT 58.035 110.125 58.325 110.170 ;
        RECT 61.255 110.125 61.545 110.170 ;
        RECT 62.620 110.110 62.940 110.170 ;
        RECT 67.220 110.110 67.540 110.170 ;
        RECT 69.060 110.310 69.380 110.370 ;
        RECT 70.900 110.310 71.220 110.370 ;
        RECT 71.450 110.310 71.590 110.465 ;
        RECT 72.740 110.450 73.060 110.510 ;
        RECT 73.215 110.465 73.505 110.510 ;
        RECT 79.155 110.650 79.445 110.695 ;
        RECT 80.345 110.650 80.635 110.695 ;
        RECT 82.865 110.650 83.155 110.695 ;
        RECT 86.080 110.650 86.400 110.710 ;
        RECT 88.395 110.650 88.685 110.695 ;
        RECT 79.155 110.510 83.155 110.650 ;
        RECT 79.155 110.465 79.445 110.510 ;
        RECT 80.345 110.465 80.635 110.510 ;
        RECT 82.865 110.465 83.155 110.510 ;
        RECT 85.250 110.510 88.685 110.650 ;
        RECT 73.675 110.310 73.965 110.355 ;
        RECT 77.340 110.310 77.660 110.370 ;
        RECT 85.250 110.355 85.390 110.510 ;
        RECT 86.080 110.450 86.400 110.510 ;
        RECT 88.395 110.465 88.685 110.510 ;
        RECT 69.060 110.170 71.590 110.310 ;
        RECT 72.830 110.170 77.660 110.310 ;
        RECT 69.060 110.110 69.380 110.170 ;
        RECT 70.900 110.110 71.220 110.170 ;
        RECT 26.280 109.970 26.600 110.030 ;
        RECT 20.160 109.830 26.600 109.970 ;
        RECT 15.715 109.785 16.005 109.830 ;
        RECT 17.080 109.770 17.400 109.830 ;
        RECT 26.280 109.770 26.600 109.830 ;
        RECT 26.740 109.970 27.060 110.030 ;
        RECT 27.215 109.970 27.505 110.015 ;
        RECT 26.740 109.830 27.505 109.970 ;
        RECT 26.740 109.770 27.060 109.830 ;
        RECT 27.215 109.785 27.505 109.830 ;
        RECT 27.675 109.970 27.965 110.015 ;
        RECT 38.700 109.970 39.020 110.030 ;
        RECT 27.675 109.830 39.020 109.970 ;
        RECT 27.675 109.785 27.965 109.830 ;
        RECT 38.700 109.770 39.020 109.830 ;
        RECT 39.160 109.770 39.480 110.030 ;
        RECT 42.855 109.970 43.145 110.015 ;
        RECT 43.300 109.970 43.620 110.030 ;
        RECT 43.775 109.970 44.065 110.015 ;
        RECT 42.855 109.830 44.065 109.970 ;
        RECT 42.855 109.785 43.145 109.830 ;
        RECT 43.300 109.770 43.620 109.830 ;
        RECT 43.775 109.785 44.065 109.830 ;
        RECT 64.460 109.970 64.780 110.030 ;
        RECT 72.830 109.970 72.970 110.170 ;
        RECT 73.675 110.125 73.965 110.170 ;
        RECT 77.340 110.110 77.660 110.170 ;
        RECT 78.760 110.310 79.050 110.355 ;
        RECT 80.860 110.310 81.150 110.355 ;
        RECT 82.430 110.310 82.720 110.355 ;
        RECT 78.760 110.170 82.720 110.310 ;
        RECT 78.760 110.125 79.050 110.170 ;
        RECT 80.860 110.125 81.150 110.170 ;
        RECT 82.430 110.125 82.720 110.170 ;
        RECT 85.175 110.125 85.465 110.355 ;
        RECT 64.460 109.830 72.970 109.970 ;
        RECT 64.460 109.770 64.780 109.830 ;
        RECT 73.200 109.770 73.520 110.030 ;
        RECT 85.620 109.770 85.940 110.030 ;
        RECT 11.950 109.150 90.610 109.630 ;
        RECT 19.840 108.950 20.160 109.010 ;
        RECT 20.315 108.950 20.605 108.995 ;
        RECT 19.840 108.810 20.605 108.950 ;
        RECT 19.840 108.750 20.160 108.810 ;
        RECT 20.315 108.765 20.605 108.810 ;
        RECT 21.680 108.750 22.000 109.010 ;
        RECT 22.615 108.950 22.905 108.995 ;
        RECT 25.820 108.950 26.140 109.010 ;
        RECT 22.615 108.810 26.140 108.950 ;
        RECT 22.615 108.765 22.905 108.810 ;
        RECT 13.900 108.610 14.190 108.655 ;
        RECT 16.000 108.610 16.290 108.655 ;
        RECT 17.570 108.610 17.860 108.655 ;
        RECT 13.900 108.470 17.860 108.610 ;
        RECT 13.900 108.425 14.190 108.470 ;
        RECT 16.000 108.425 16.290 108.470 ;
        RECT 17.570 108.425 17.860 108.470 ;
        RECT 21.235 108.610 21.525 108.655 ;
        RECT 22.690 108.610 22.830 108.765 ;
        RECT 25.820 108.750 26.140 108.810 ;
        RECT 26.280 108.950 26.600 109.010 ;
        RECT 29.515 108.950 29.805 108.995 ;
        RECT 26.280 108.810 29.805 108.950 ;
        RECT 26.280 108.750 26.600 108.810 ;
        RECT 29.515 108.765 29.805 108.810 ;
        RECT 30.435 108.765 30.725 108.995 ;
        RECT 35.020 108.950 35.340 109.010 ;
        RECT 35.495 108.950 35.785 108.995 ;
        RECT 35.020 108.810 35.785 108.950 ;
        RECT 24.900 108.610 25.220 108.670 ;
        RECT 26.740 108.610 27.060 108.670 ;
        RECT 30.510 108.610 30.650 108.765 ;
        RECT 35.020 108.750 35.340 108.810 ;
        RECT 35.495 108.765 35.785 108.810 ;
        RECT 37.795 108.950 38.085 108.995 ;
        RECT 41.000 108.950 41.320 109.010 ;
        RECT 37.795 108.810 41.320 108.950 ;
        RECT 37.795 108.765 38.085 108.810 ;
        RECT 41.000 108.750 41.320 108.810 ;
        RECT 49.295 108.765 49.585 108.995 ;
        RECT 21.235 108.470 22.830 108.610 ;
        RECT 24.070 108.470 30.650 108.610 ;
        RECT 21.235 108.425 21.525 108.470 ;
        RECT 14.295 108.270 14.585 108.315 ;
        RECT 15.485 108.270 15.775 108.315 ;
        RECT 18.005 108.270 18.295 108.315 ;
        RECT 14.295 108.130 18.295 108.270 ;
        RECT 14.295 108.085 14.585 108.130 ;
        RECT 15.485 108.085 15.775 108.130 ;
        RECT 18.005 108.085 18.295 108.130 ;
        RECT 22.140 108.070 22.460 108.330 ;
        RECT 13.415 107.930 13.705 107.975 ;
        RECT 20.300 107.930 20.620 107.990 ;
        RECT 13.415 107.790 20.620 107.930 ;
        RECT 13.415 107.745 13.705 107.790 ;
        RECT 20.300 107.730 20.620 107.790 ;
        RECT 20.775 107.930 21.065 107.975 ;
        RECT 21.220 107.930 21.540 107.990 ;
        RECT 23.060 107.930 23.380 107.990 ;
        RECT 20.775 107.790 23.380 107.930 ;
        RECT 20.775 107.745 21.065 107.790 ;
        RECT 21.220 107.730 21.540 107.790 ;
        RECT 23.060 107.730 23.380 107.790 ;
        RECT 23.535 107.940 23.825 107.975 ;
        RECT 24.070 107.940 24.210 108.470 ;
        RECT 24.900 108.410 25.220 108.470 ;
        RECT 26.740 108.410 27.060 108.470 ;
        RECT 35.110 108.270 35.250 108.750 ;
        RECT 38.240 108.610 38.560 108.670 ;
        RECT 38.715 108.610 39.005 108.655 ;
        RECT 38.240 108.470 39.005 108.610 ;
        RECT 38.240 108.410 38.560 108.470 ;
        RECT 38.715 108.425 39.005 108.470 ;
        RECT 39.160 108.610 39.480 108.670 ;
        RECT 49.370 108.610 49.510 108.765 ;
        RECT 57.560 108.750 57.880 109.010 ;
        RECT 62.160 108.950 62.480 109.010 ;
        RECT 64.000 108.950 64.320 109.010 ;
        RECT 65.395 108.950 65.685 108.995 ;
        RECT 62.160 108.810 65.685 108.950 ;
        RECT 62.160 108.750 62.480 108.810 ;
        RECT 64.000 108.750 64.320 108.810 ;
        RECT 65.395 108.765 65.685 108.810 ;
        RECT 67.680 108.950 68.000 109.010 ;
        RECT 68.615 108.950 68.905 108.995 ;
        RECT 67.680 108.810 68.905 108.950 ;
        RECT 55.720 108.610 56.040 108.670 ;
        RECT 39.160 108.470 56.040 108.610 ;
        RECT 39.160 108.410 39.480 108.470 ;
        RECT 55.720 108.410 56.040 108.470 ;
        RECT 24.530 108.130 31.570 108.270 ;
        RECT 24.530 107.990 24.670 108.130 ;
        RECT 23.535 107.800 24.210 107.940 ;
        RECT 23.535 107.745 23.825 107.800 ;
        RECT 24.440 107.730 24.760 107.990 ;
        RECT 27.215 107.930 27.505 107.975 ;
        RECT 29.055 107.930 29.345 107.975 ;
        RECT 24.990 107.790 27.505 107.930 ;
        RECT 13.860 107.590 14.180 107.650 ;
        RECT 14.640 107.590 14.930 107.635 ;
        RECT 13.860 107.450 14.930 107.590 ;
        RECT 13.860 107.390 14.180 107.450 ;
        RECT 14.640 107.405 14.930 107.450 ;
        RECT 15.240 107.590 15.560 107.650 ;
        RECT 24.990 107.590 25.130 107.790 ;
        RECT 27.215 107.745 27.505 107.790 ;
        RECT 27.750 107.790 29.345 107.930 ;
        RECT 15.240 107.450 25.130 107.590 ;
        RECT 15.240 107.390 15.560 107.450 ;
        RECT 24.990 107.250 25.130 107.450 ;
        RECT 25.360 107.590 25.680 107.650 ;
        RECT 27.750 107.590 27.890 107.790 ;
        RECT 29.055 107.745 29.345 107.790 ;
        RECT 29.500 107.930 29.820 107.990 ;
        RECT 31.430 107.975 31.570 108.130 ;
        RECT 34.190 108.130 35.250 108.270 ;
        RECT 35.480 108.270 35.800 108.330 ;
        RECT 65.470 108.270 65.610 108.765 ;
        RECT 67.680 108.750 68.000 108.810 ;
        RECT 68.615 108.765 68.905 108.810 ;
        RECT 70.900 108.750 71.220 109.010 ;
        RECT 71.820 108.950 72.140 109.010 ;
        RECT 73.660 108.950 73.980 109.010 ;
        RECT 71.820 108.810 73.980 108.950 ;
        RECT 71.820 108.750 72.140 108.810 ;
        RECT 73.660 108.750 73.980 108.810 ;
        RECT 79.640 108.950 79.960 109.010 ;
        RECT 80.575 108.950 80.865 108.995 ;
        RECT 79.640 108.810 80.865 108.950 ;
        RECT 79.640 108.750 79.960 108.810 ;
        RECT 80.575 108.765 80.865 108.810 ;
        RECT 87.000 108.750 87.320 109.010 ;
        RECT 67.220 108.610 67.540 108.670 ;
        RECT 70.440 108.610 70.760 108.670 ;
        RECT 72.755 108.610 73.045 108.655 ;
        RECT 74.120 108.610 74.440 108.670 ;
        RECT 67.220 108.470 71.590 108.610 ;
        RECT 67.220 108.410 67.540 108.470 ;
        RECT 70.440 108.410 70.760 108.470 ;
        RECT 71.450 108.315 71.590 108.470 ;
        RECT 72.755 108.470 77.110 108.610 ;
        RECT 72.755 108.425 73.045 108.470 ;
        RECT 74.120 108.410 74.440 108.470 ;
        RECT 35.480 108.130 51.350 108.270 ;
        RECT 65.470 108.130 71.130 108.270 ;
        RECT 34.190 107.975 34.330 108.130 ;
        RECT 35.480 108.070 35.800 108.130 ;
        RECT 30.435 107.930 30.725 107.975 ;
        RECT 29.500 107.790 30.725 107.930 ;
        RECT 29.500 107.730 29.820 107.790 ;
        RECT 30.435 107.745 30.725 107.790 ;
        RECT 31.355 107.745 31.645 107.975 ;
        RECT 34.115 107.745 34.405 107.975 ;
        RECT 35.035 107.930 35.325 107.975 ;
        RECT 35.940 107.930 36.260 107.990 ;
        RECT 35.035 107.790 36.260 107.930 ;
        RECT 35.035 107.745 35.325 107.790 ;
        RECT 35.940 107.730 36.260 107.790 ;
        RECT 36.875 107.745 37.165 107.975 ;
        RECT 38.255 107.930 38.545 107.975 ;
        RECT 40.540 107.930 40.860 107.990 ;
        RECT 38.255 107.790 40.860 107.930 ;
        RECT 38.255 107.745 38.545 107.790 ;
        RECT 25.360 107.450 27.890 107.590 ;
        RECT 28.265 107.590 28.555 107.635 ;
        RECT 29.960 107.590 30.280 107.650 ;
        RECT 36.950 107.590 37.090 107.745 ;
        RECT 40.540 107.730 40.860 107.790 ;
        RECT 41.475 107.745 41.765 107.975 ;
        RECT 37.320 107.590 37.640 107.650 ;
        RECT 41.550 107.590 41.690 107.745 ;
        RECT 42.840 107.730 43.160 107.990 ;
        RECT 43.315 107.930 43.605 107.975 ;
        RECT 43.760 107.930 44.080 107.990 ;
        RECT 43.315 107.790 44.080 107.930 ;
        RECT 43.315 107.745 43.605 107.790 ;
        RECT 43.760 107.730 44.080 107.790 ;
        RECT 44.220 107.730 44.540 107.990 ;
        RECT 51.210 107.975 51.350 108.130 ;
        RECT 51.135 107.745 51.425 107.975 ;
        RECT 64.935 107.930 65.225 107.975 ;
        RECT 65.380 107.930 65.700 107.990 ;
        RECT 67.220 107.930 67.540 107.990 ;
        RECT 70.990 107.975 71.130 108.130 ;
        RECT 71.375 108.085 71.665 108.315 ;
        RECT 71.910 108.130 74.350 108.270 ;
        RECT 64.935 107.790 70.670 107.930 ;
        RECT 64.935 107.745 65.225 107.790 ;
        RECT 65.380 107.730 65.700 107.790 ;
        RECT 67.220 107.730 67.540 107.790 ;
        RECT 45.600 107.590 45.920 107.650 ;
        RECT 28.265 107.450 30.280 107.590 ;
        RECT 25.360 107.390 25.680 107.450 ;
        RECT 28.265 107.405 28.555 107.450 ;
        RECT 29.960 107.390 30.280 107.450 ;
        RECT 34.650 107.450 36.630 107.590 ;
        RECT 36.950 107.450 45.920 107.590 ;
        RECT 34.650 107.250 34.790 107.450 ;
        RECT 24.990 107.110 34.790 107.250 ;
        RECT 35.020 107.050 35.340 107.310 ;
        RECT 36.490 107.250 36.630 107.450 ;
        RECT 37.320 107.390 37.640 107.450 ;
        RECT 45.600 107.390 45.920 107.450 ;
        RECT 48.360 107.390 48.680 107.650 ;
        RECT 55.260 107.590 55.580 107.650 ;
        RECT 70.530 107.590 70.670 107.790 ;
        RECT 70.915 107.745 71.205 107.975 ;
        RECT 71.910 107.930 72.050 108.130 ;
        RECT 74.210 107.975 74.350 108.130 ;
        RECT 76.970 107.975 77.110 108.470 ;
        RECT 83.320 108.070 83.640 108.330 ;
        RECT 73.215 107.930 73.505 107.975 ;
        RECT 71.450 107.790 72.050 107.930 ;
        RECT 72.370 107.790 73.505 107.930 ;
        RECT 71.450 107.590 71.590 107.790 ;
        RECT 48.910 107.450 55.580 107.590 ;
        RECT 48.910 107.250 49.050 107.450 ;
        RECT 55.260 107.390 55.580 107.450 ;
        RECT 67.770 107.450 70.210 107.590 ;
        RECT 70.530 107.450 71.590 107.590 ;
        RECT 67.770 107.310 67.910 107.450 ;
        RECT 36.490 107.110 49.050 107.250 ;
        RECT 49.280 107.295 49.600 107.310 ;
        RECT 49.280 107.065 49.665 107.295 ;
        RECT 49.280 107.050 49.600 107.065 ;
        RECT 50.200 107.050 50.520 107.310 ;
        RECT 67.680 107.050 68.000 107.310 ;
        RECT 68.600 107.050 68.920 107.310 ;
        RECT 70.070 107.250 70.210 107.450 ;
        RECT 72.370 107.250 72.510 107.790 ;
        RECT 73.215 107.745 73.505 107.790 ;
        RECT 74.135 107.745 74.425 107.975 ;
        RECT 76.895 107.745 77.185 107.975 ;
        RECT 77.340 107.930 77.660 107.990 ;
        RECT 82.415 107.930 82.705 107.975 ;
        RECT 85.620 107.930 85.940 107.990 ;
        RECT 77.340 107.790 77.855 107.930 ;
        RECT 82.415 107.790 85.940 107.930 ;
        RECT 77.340 107.730 77.660 107.790 ;
        RECT 82.415 107.745 82.705 107.790 ;
        RECT 85.620 107.730 85.940 107.790 ;
        RECT 86.080 107.730 86.400 107.990 ;
        RECT 100.000 107.510 100.830 110.850 ;
        RECT 108.880 110.550 116.800 110.560 ;
        RECT 105.110 110.540 116.800 110.550 ;
        RECT 101.490 110.420 116.800 110.540 ;
        RECT 101.490 110.410 116.825 110.420 ;
        RECT 101.450 110.290 116.825 110.410 ;
        RECT 101.450 110.180 105.450 110.290 ;
        RECT 101.060 109.840 101.290 110.130 ;
        RECT 101.510 109.840 105.400 110.180 ;
        RECT 105.610 109.840 105.840 110.130 ;
        RECT 101.060 108.470 105.840 109.840 ;
        RECT 101.060 108.170 101.290 108.470 ;
        RECT 105.610 108.170 105.840 108.470 ;
        RECT 101.450 107.890 105.450 108.120 ;
        RECT 101.700 107.660 105.270 107.890 ;
        RECT 101.700 107.510 105.390 107.660 ;
        RECT 70.070 107.110 72.510 107.250 ;
        RECT 75.500 107.250 75.820 107.310 ;
        RECT 78.735 107.250 79.025 107.295 ;
        RECT 75.500 107.110 79.025 107.250 ;
        RECT 75.500 107.050 75.820 107.110 ;
        RECT 78.735 107.065 79.025 107.110 ;
        RECT 81.480 107.250 81.800 107.310 ;
        RECT 82.875 107.250 83.165 107.295 ;
        RECT 81.480 107.110 83.165 107.250 ;
        RECT 81.480 107.050 81.800 107.110 ;
        RECT 82.875 107.065 83.165 107.110 ;
        RECT 100.000 107.230 105.390 107.510 ;
        RECT 106.640 107.340 107.260 110.290 ;
        RECT 108.825 110.190 116.825 110.290 ;
        RECT 108.880 110.180 116.800 110.190 ;
        RECT 108.390 109.480 108.620 110.140 ;
        RECT 109.400 109.480 110.400 109.570 ;
        RECT 117.030 109.480 117.260 110.140 ;
        RECT 108.390 108.660 117.260 109.480 ;
        RECT 108.390 108.180 108.620 108.660 ;
        RECT 109.400 108.570 110.400 108.660 ;
        RECT 117.030 108.180 117.260 108.660 ;
        RECT 108.825 107.900 116.825 108.130 ;
        RECT 11.950 106.430 90.610 106.910 ;
        RECT 100.000 106.770 105.400 107.230 ;
        RECT 13.860 106.030 14.180 106.290 ;
        RECT 22.140 106.230 22.460 106.290 ;
        RECT 23.535 106.230 23.825 106.275 ;
        RECT 22.140 106.090 23.825 106.230 ;
        RECT 22.140 106.030 22.460 106.090 ;
        RECT 23.535 106.045 23.825 106.090 ;
        RECT 37.320 106.030 37.640 106.290 ;
        RECT 38.240 106.230 38.560 106.290 ;
        RECT 38.715 106.230 39.005 106.275 ;
        RECT 38.240 106.090 39.005 106.230 ;
        RECT 38.240 106.030 38.560 106.090 ;
        RECT 38.715 106.045 39.005 106.090 ;
        RECT 40.540 106.230 40.860 106.290 ;
        RECT 41.475 106.230 41.765 106.275 ;
        RECT 43.760 106.230 44.080 106.290 ;
        RECT 55.720 106.275 56.040 106.290 ;
        RECT 49.295 106.230 49.585 106.275 ;
        RECT 40.540 106.090 41.765 106.230 ;
        RECT 40.540 106.030 40.860 106.090 ;
        RECT 41.475 106.045 41.765 106.090 ;
        RECT 42.010 106.090 49.585 106.230 ;
        RECT 15.240 105.690 15.560 105.950 ;
        RECT 15.700 105.690 16.020 105.950 ;
        RECT 16.405 105.890 16.695 105.935 ;
        RECT 18.000 105.890 18.320 105.950 ;
        RECT 20.760 105.890 21.080 105.950 ;
        RECT 23.980 105.890 24.300 105.950 ;
        RECT 35.020 105.890 35.340 105.950 ;
        RECT 16.405 105.750 18.320 105.890 ;
        RECT 16.405 105.705 16.695 105.750 ;
        RECT 18.000 105.690 18.320 105.750 ;
        RECT 20.390 105.750 21.080 105.890 ;
        RECT 14.795 105.365 15.085 105.595 ;
        RECT 14.870 105.210 15.010 105.365 ;
        RECT 17.080 105.350 17.400 105.610 ;
        RECT 18.935 105.550 19.225 105.595 ;
        RECT 19.840 105.550 20.160 105.610 ;
        RECT 20.390 105.595 20.530 105.750 ;
        RECT 20.760 105.690 21.080 105.750 ;
        RECT 21.310 105.750 25.130 105.890 ;
        RECT 21.310 105.595 21.450 105.750 ;
        RECT 23.980 105.690 24.300 105.750 ;
        RECT 24.990 105.610 25.130 105.750 ;
        RECT 35.020 105.750 39.850 105.890 ;
        RECT 35.020 105.690 35.340 105.750 ;
        RECT 18.935 105.410 20.160 105.550 ;
        RECT 18.935 105.365 19.225 105.410 ;
        RECT 19.840 105.350 20.160 105.410 ;
        RECT 20.315 105.365 20.605 105.595 ;
        RECT 21.235 105.365 21.525 105.595 ;
        RECT 21.680 105.350 22.000 105.610 ;
        RECT 24.900 105.350 25.220 105.610 ;
        RECT 25.360 105.550 25.680 105.610 ;
        RECT 30.435 105.550 30.725 105.595 ;
        RECT 25.360 105.410 30.725 105.550 ;
        RECT 25.360 105.350 25.680 105.410 ;
        RECT 30.435 105.365 30.725 105.410 ;
        RECT 31.770 105.550 32.060 105.595 ;
        RECT 31.770 105.410 36.170 105.550 ;
        RECT 31.770 105.365 32.060 105.410 ;
        RECT 16.160 105.210 16.480 105.270 ;
        RECT 20.775 105.210 21.065 105.255 ;
        RECT 22.140 105.210 22.460 105.270 ;
        RECT 23.535 105.210 23.825 105.255 ;
        RECT 14.870 105.070 18.690 105.210 ;
        RECT 16.160 105.010 16.480 105.070 ;
        RECT 12.940 104.870 13.260 104.930 ;
        RECT 18.015 104.870 18.305 104.915 ;
        RECT 12.940 104.730 18.305 104.870 ;
        RECT 18.550 104.870 18.690 105.070 ;
        RECT 20.775 105.070 23.825 105.210 ;
        RECT 20.775 105.025 21.065 105.070 ;
        RECT 22.140 105.010 22.460 105.070 ;
        RECT 23.535 105.025 23.825 105.070 ;
        RECT 24.440 105.210 24.760 105.270 ;
        RECT 29.515 105.210 29.805 105.255 ;
        RECT 24.440 105.070 29.805 105.210 ;
        RECT 24.440 105.010 24.760 105.070 ;
        RECT 29.515 105.025 29.805 105.070 ;
        RECT 31.315 105.210 31.605 105.255 ;
        RECT 32.505 105.210 32.795 105.255 ;
        RECT 35.025 105.210 35.315 105.255 ;
        RECT 31.315 105.070 35.315 105.210 ;
        RECT 36.030 105.210 36.170 105.410 ;
        RECT 38.240 105.350 38.560 105.610 ;
        RECT 39.710 105.595 39.850 105.750 ;
        RECT 39.635 105.365 39.925 105.595 ;
        RECT 41.015 105.550 41.305 105.595 ;
        RECT 41.460 105.550 41.780 105.610 ;
        RECT 42.010 105.595 42.150 106.090 ;
        RECT 43.760 106.030 44.080 106.090 ;
        RECT 49.295 106.045 49.585 106.090 ;
        RECT 55.720 106.045 56.105 106.275 ;
        RECT 62.620 106.230 62.940 106.290 ;
        RECT 65.840 106.230 66.160 106.290 ;
        RECT 74.580 106.230 74.900 106.290 ;
        RECT 77.355 106.230 77.645 106.275 ;
        RECT 83.320 106.230 83.640 106.290 ;
        RECT 62.620 106.090 76.190 106.230 ;
        RECT 55.720 106.030 56.040 106.045 ;
        RECT 62.620 106.030 62.940 106.090 ;
        RECT 65.840 106.030 66.160 106.090 ;
        RECT 74.580 106.030 74.900 106.090 ;
        RECT 54.800 105.690 55.120 105.950 ;
        RECT 65.380 105.890 65.700 105.950 ;
        RECT 66.300 105.890 66.620 105.950 ;
        RECT 65.380 105.750 75.730 105.890 ;
        RECT 65.380 105.690 65.700 105.750 ;
        RECT 66.300 105.690 66.620 105.750 ;
        RECT 75.590 105.610 75.730 105.750 ;
        RECT 41.015 105.410 41.780 105.550 ;
        RECT 41.015 105.365 41.305 105.410 ;
        RECT 41.460 105.350 41.780 105.410 ;
        RECT 41.935 105.365 42.225 105.595 ;
        RECT 43.730 105.550 44.020 105.595 ;
        RECT 45.140 105.550 45.460 105.610 ;
        RECT 43.730 105.410 45.460 105.550 ;
        RECT 43.730 105.365 44.020 105.410 ;
        RECT 45.140 105.350 45.460 105.410 ;
        RECT 64.000 105.350 64.320 105.610 ;
        RECT 67.680 105.550 68.000 105.610 ;
        RECT 71.835 105.550 72.125 105.595 ;
        RECT 67.680 105.410 72.125 105.550 ;
        RECT 67.680 105.350 68.000 105.410 ;
        RECT 71.835 105.365 72.125 105.410 ;
        RECT 72.755 105.550 73.045 105.595 ;
        RECT 73.660 105.550 73.980 105.610 ;
        RECT 72.755 105.410 73.980 105.550 ;
        RECT 72.755 105.365 73.045 105.410 ;
        RECT 73.660 105.350 73.980 105.410 ;
        RECT 74.135 105.365 74.425 105.595 ;
        RECT 40.555 105.210 40.845 105.255 ;
        RECT 36.030 105.070 40.845 105.210 ;
        RECT 31.315 105.025 31.605 105.070 ;
        RECT 32.505 105.025 32.795 105.070 ;
        RECT 35.025 105.025 35.315 105.070 ;
        RECT 40.555 105.025 40.845 105.070 ;
        RECT 42.380 105.010 42.700 105.270 ;
        RECT 43.275 105.210 43.565 105.255 ;
        RECT 44.465 105.210 44.755 105.255 ;
        RECT 46.985 105.210 47.275 105.255 ;
        RECT 43.275 105.070 47.275 105.210 ;
        RECT 43.275 105.025 43.565 105.070 ;
        RECT 44.465 105.025 44.755 105.070 ;
        RECT 46.985 105.025 47.275 105.070 ;
        RECT 52.500 105.210 52.820 105.270 ;
        RECT 53.435 105.210 53.725 105.255 ;
        RECT 52.500 105.070 53.725 105.210 ;
        RECT 52.500 105.010 52.820 105.070 ;
        RECT 53.435 105.025 53.725 105.070 ;
        RECT 53.880 105.210 54.200 105.270 ;
        RECT 57.115 105.210 57.405 105.255 ;
        RECT 53.880 105.070 57.405 105.210 ;
        RECT 53.880 105.010 54.200 105.070 ;
        RECT 57.115 105.025 57.405 105.070 ;
        RECT 65.395 105.210 65.685 105.255 ;
        RECT 67.770 105.210 67.910 105.350 ;
        RECT 65.395 105.070 67.910 105.210 ;
        RECT 72.280 105.210 72.600 105.270 ;
        RECT 74.210 105.210 74.350 105.365 ;
        RECT 75.040 105.350 75.360 105.610 ;
        RECT 75.500 105.350 75.820 105.610 ;
        RECT 76.050 105.595 76.190 106.090 ;
        RECT 77.355 106.090 83.640 106.230 ;
        RECT 77.355 106.045 77.645 106.090 ;
        RECT 83.320 106.030 83.640 106.090 ;
        RECT 75.975 105.365 76.265 105.595 ;
        RECT 79.195 105.365 79.485 105.595 ;
        RECT 100.000 105.430 102.000 106.770 ;
        RECT 103.750 106.760 105.400 106.770 ;
        RECT 102.440 105.490 103.440 106.210 ;
        RECT 103.750 105.950 104.060 106.760 ;
        RECT 104.520 106.480 105.400 106.760 ;
        RECT 105.640 106.940 107.260 107.340 ;
        RECT 108.910 106.990 116.780 107.900 ;
        RECT 104.460 106.250 105.460 106.480 ;
        RECT 105.640 106.290 105.990 106.940 ;
        RECT 106.640 106.930 107.260 106.940 ;
        RECT 108.825 106.760 116.825 106.990 ;
        RECT 108.910 106.750 116.780 106.760 ;
        RECT 104.520 106.040 105.400 106.060 ;
        RECT 103.790 105.660 104.060 105.950 ;
        RECT 104.460 105.810 105.460 106.040 ;
        RECT 105.620 106.000 105.990 106.290 ;
        RECT 105.650 105.940 105.990 106.000 ;
        RECT 106.750 106.610 107.510 106.660 ;
        RECT 108.390 106.610 108.620 106.710 ;
        RECT 106.750 106.400 108.620 106.610 ;
        RECT 117.030 106.400 117.260 106.710 ;
        RECT 106.750 105.980 109.290 106.400 ;
        RECT 116.660 105.980 117.260 106.400 ;
        RECT 104.520 105.660 105.400 105.810 ;
        RECT 104.530 105.490 105.260 105.660 ;
        RECT 100.080 105.420 102.000 105.430 ;
        RECT 72.280 105.070 74.350 105.210 ;
        RECT 65.395 105.025 65.685 105.070 ;
        RECT 72.280 105.010 72.600 105.070 ;
        RECT 22.615 104.870 22.905 104.915 ;
        RECT 23.060 104.870 23.380 104.930 ;
        RECT 30.920 104.870 31.210 104.915 ;
        RECT 33.020 104.870 33.310 104.915 ;
        RECT 34.590 104.870 34.880 104.915 ;
        RECT 18.550 104.730 27.430 104.870 ;
        RECT 12.940 104.670 13.260 104.730 ;
        RECT 18.015 104.685 18.305 104.730 ;
        RECT 22.615 104.685 22.905 104.730 ;
        RECT 23.060 104.670 23.380 104.730 ;
        RECT 24.440 104.330 24.760 104.590 ;
        RECT 24.900 104.530 25.220 104.590 ;
        RECT 26.755 104.530 27.045 104.575 ;
        RECT 24.900 104.390 27.045 104.530 ;
        RECT 27.290 104.530 27.430 104.730 ;
        RECT 30.920 104.730 34.880 104.870 ;
        RECT 30.920 104.685 31.210 104.730 ;
        RECT 33.020 104.685 33.310 104.730 ;
        RECT 34.590 104.685 34.880 104.730 ;
        RECT 42.880 104.870 43.170 104.915 ;
        RECT 44.980 104.870 45.270 104.915 ;
        RECT 46.550 104.870 46.840 104.915 ;
        RECT 42.880 104.730 46.840 104.870 ;
        RECT 42.880 104.685 43.170 104.730 ;
        RECT 44.980 104.685 45.270 104.730 ;
        RECT 46.550 104.685 46.840 104.730 ;
        RECT 56.655 104.870 56.945 104.915 ;
        RECT 78.720 104.870 79.040 104.930 ;
        RECT 79.270 104.870 79.410 105.365 ;
        RECT 86.080 105.210 86.400 105.270 ;
        RECT 87.475 105.210 87.765 105.255 ;
        RECT 86.080 105.070 87.765 105.210 ;
        RECT 86.080 105.010 86.400 105.070 ;
        RECT 87.475 105.025 87.765 105.070 ;
        RECT 56.655 104.730 79.410 104.870 ;
        RECT 56.655 104.685 56.945 104.730 ;
        RECT 78.720 104.670 79.040 104.730 ;
        RECT 48.360 104.530 48.680 104.590 ;
        RECT 27.290 104.390 48.680 104.530 ;
        RECT 24.900 104.330 25.220 104.390 ;
        RECT 26.755 104.345 27.045 104.390 ;
        RECT 48.360 104.330 48.680 104.390 ;
        RECT 50.660 104.330 50.980 104.590 ;
        RECT 55.260 104.530 55.580 104.590 ;
        RECT 55.735 104.530 56.025 104.575 ;
        RECT 55.260 104.390 56.025 104.530 ;
        RECT 55.260 104.330 55.580 104.390 ;
        RECT 55.735 104.345 56.025 104.390 ;
        RECT 60.320 104.330 60.640 104.590 ;
        RECT 64.000 104.530 64.320 104.590 ;
        RECT 64.475 104.530 64.765 104.575 ;
        RECT 64.000 104.390 64.765 104.530 ;
        RECT 64.000 104.330 64.320 104.390 ;
        RECT 64.475 104.345 64.765 104.390 ;
        RECT 64.935 104.530 65.225 104.575 ;
        RECT 66.300 104.530 66.620 104.590 ;
        RECT 64.935 104.390 66.620 104.530 ;
        RECT 64.935 104.345 65.225 104.390 ;
        RECT 66.300 104.330 66.620 104.390 ;
        RECT 72.280 104.530 72.600 104.590 ;
        RECT 73.215 104.530 73.505 104.575 ;
        RECT 72.280 104.390 73.505 104.530 ;
        RECT 72.280 104.330 72.600 104.390 ;
        RECT 73.215 104.345 73.505 104.390 ;
        RECT 73.660 104.530 73.980 104.590 ;
        RECT 75.500 104.530 75.820 104.590 ;
        RECT 78.275 104.530 78.565 104.575 ;
        RECT 73.660 104.390 78.565 104.530 ;
        RECT 73.660 104.330 73.980 104.390 ;
        RECT 75.500 104.330 75.820 104.390 ;
        RECT 78.275 104.345 78.565 104.390 ;
        RECT 82.860 104.530 83.180 104.590 ;
        RECT 84.715 104.530 85.005 104.575 ;
        RECT 82.860 104.390 85.005 104.530 ;
        RECT 82.860 104.330 83.180 104.390 ;
        RECT 84.715 104.345 85.005 104.390 ;
        RECT 102.410 104.370 105.260 105.490 ;
        RECT 105.650 105.190 106.000 105.940 ;
        RECT 106.750 105.820 108.620 105.980 ;
        RECT 106.750 105.770 107.510 105.820 ;
        RECT 108.390 105.750 108.620 105.820 ;
        RECT 117.030 105.750 117.260 105.980 ;
        RECT 108.825 105.470 116.825 105.700 ;
        RECT 105.650 105.130 105.940 105.190 ;
        RECT 105.560 105.010 105.940 105.130 ;
        RECT 108.920 105.070 116.780 105.470 ;
        RECT 117.590 105.070 118.560 114.550 ;
        RECT 119.930 114.680 120.770 116.810 ;
        RECT 126.430 116.390 127.680 116.830 ;
        RECT 137.600 116.810 138.460 118.930 ;
        RECT 124.370 116.380 129.610 116.390 ;
        RECT 121.420 116.280 136.720 116.380 ;
        RECT 121.420 116.270 136.755 116.280 ;
        RECT 121.380 116.150 136.755 116.270 ;
        RECT 121.380 116.040 125.380 116.150 ;
        RECT 126.430 116.070 128.170 116.150 ;
        RECT 128.750 116.070 136.755 116.150 ;
        RECT 126.430 115.990 127.680 116.070 ;
        RECT 128.755 116.050 136.755 116.070 ;
        RECT 120.990 115.740 121.220 115.990 ;
        RECT 125.540 115.850 125.770 115.990 ;
        RECT 128.320 115.850 128.550 116.000 ;
        RECT 125.540 115.740 128.550 115.850 ;
        RECT 136.960 115.740 137.190 116.000 ;
        RECT 120.990 115.300 137.190 115.740 ;
        RECT 120.990 115.030 121.220 115.300 ;
        RECT 125.540 115.270 137.190 115.300 ;
        RECT 125.540 115.180 128.550 115.270 ;
        RECT 125.540 115.030 125.770 115.180 ;
        RECT 128.320 115.040 128.550 115.180 ;
        RECT 136.960 115.040 137.190 115.270 ;
        RECT 121.380 114.750 125.380 114.980 ;
        RECT 128.755 114.770 136.755 114.990 ;
        RECT 137.520 114.770 138.480 116.810 ;
        RECT 128.755 114.760 138.480 114.770 ;
        RECT 121.380 114.680 125.370 114.750 ;
        RECT 119.930 114.570 125.370 114.680 ;
        RECT 128.810 114.600 138.480 114.760 ;
        RECT 119.930 114.480 123.060 114.570 ;
        RECT 136.550 114.550 138.480 114.600 ;
        RECT 119.930 111.210 120.770 114.480 ;
        RECT 124.410 114.020 129.660 114.030 ;
        RECT 124.410 113.910 136.720 114.020 ;
        RECT 121.440 113.850 136.720 113.910 ;
        RECT 121.440 113.840 136.755 113.850 ;
        RECT 121.380 113.710 136.755 113.840 ;
        RECT 121.380 113.700 126.540 113.710 ;
        RECT 121.380 113.610 125.380 113.700 ;
        RECT 128.755 113.620 136.755 113.710 ;
        RECT 128.840 113.610 136.730 113.620 ;
        RECT 120.990 113.250 121.220 113.560 ;
        RECT 121.440 113.250 125.340 113.610 ;
        RECT 125.540 113.250 125.770 113.560 ;
        RECT 120.990 111.910 125.770 113.250 ;
        RECT 120.990 111.600 121.220 111.910 ;
        RECT 125.540 111.600 125.770 111.910 ;
        RECT 128.320 113.030 128.550 113.570 ;
        RECT 129.360 113.030 130.370 113.060 ;
        RECT 136.960 113.030 137.190 113.570 ;
        RECT 128.320 112.130 137.190 113.030 ;
        RECT 128.320 111.610 128.550 112.130 ;
        RECT 129.360 112.060 130.370 112.130 ;
        RECT 136.960 111.610 137.190 112.130 ;
        RECT 121.380 111.320 125.380 111.550 ;
        RECT 128.755 111.330 136.755 111.560 ;
        RECT 119.930 111.170 121.060 111.210 ;
        RECT 119.930 111.090 121.300 111.170 ;
        RECT 121.670 111.100 125.330 111.320 ;
        RECT 121.670 111.090 123.110 111.100 ;
        RECT 119.930 111.050 123.110 111.090 ;
        RECT 119.930 110.960 122.620 111.050 ;
        RECT 128.820 111.040 136.710 111.330 ;
        RECT 119.930 110.900 121.950 110.960 ;
        RECT 119.930 110.850 121.700 110.900 ;
        RECT 119.930 107.510 120.770 110.850 ;
        RECT 128.810 110.550 136.730 110.560 ;
        RECT 125.040 110.540 136.730 110.550 ;
        RECT 121.420 110.420 136.730 110.540 ;
        RECT 121.420 110.410 136.755 110.420 ;
        RECT 121.380 110.290 136.755 110.410 ;
        RECT 121.380 110.180 125.380 110.290 ;
        RECT 120.990 109.840 121.220 110.130 ;
        RECT 121.440 109.840 125.330 110.180 ;
        RECT 125.540 109.840 125.770 110.130 ;
        RECT 120.990 108.470 125.770 109.840 ;
        RECT 120.990 108.170 121.220 108.470 ;
        RECT 125.540 108.170 125.770 108.470 ;
        RECT 121.380 107.890 125.380 108.120 ;
        RECT 121.630 107.660 125.200 107.890 ;
        RECT 121.630 107.510 125.320 107.660 ;
        RECT 119.930 107.230 125.320 107.510 ;
        RECT 126.570 107.340 127.190 110.290 ;
        RECT 128.755 110.190 136.755 110.290 ;
        RECT 128.810 110.180 136.730 110.190 ;
        RECT 128.320 109.480 128.550 110.140 ;
        RECT 129.330 109.480 130.330 109.570 ;
        RECT 136.960 109.480 137.190 110.140 ;
        RECT 128.320 108.660 137.190 109.480 ;
        RECT 128.320 108.180 128.550 108.660 ;
        RECT 129.330 108.570 130.330 108.660 ;
        RECT 136.960 108.180 137.190 108.660 ;
        RECT 128.755 107.900 136.755 108.130 ;
        RECT 119.930 106.770 125.330 107.230 ;
        RECT 119.930 105.880 121.930 106.770 ;
        RECT 123.680 106.760 125.330 106.770 ;
        RECT 11.950 103.710 90.610 104.190 ;
        RECT 102.350 104.140 105.350 104.370 ;
        RECT 105.560 104.180 105.900 105.010 ;
        RECT 107.910 105.000 118.560 105.070 ;
        RECT 102.400 104.110 105.260 104.140 ;
        RECT 102.400 104.090 103.570 104.110 ;
        RECT 104.530 104.100 105.260 104.110 ;
        RECT 102.350 103.700 105.350 103.930 ;
        RECT 105.555 103.890 105.900 104.180 ;
        RECT 106.090 104.040 118.560 105.000 ;
        RECT 119.900 105.420 121.930 105.880 ;
        RECT 122.370 105.490 123.370 106.210 ;
        RECT 123.680 105.950 123.990 106.760 ;
        RECT 124.450 106.480 125.330 106.760 ;
        RECT 125.570 106.940 127.190 107.340 ;
        RECT 128.840 106.990 136.710 107.900 ;
        RECT 124.390 106.250 125.390 106.480 ;
        RECT 125.570 106.290 125.920 106.940 ;
        RECT 126.570 106.930 127.190 106.940 ;
        RECT 128.755 106.760 136.755 106.990 ;
        RECT 128.840 106.750 136.710 106.760 ;
        RECT 124.450 106.040 125.330 106.060 ;
        RECT 123.720 105.660 123.990 105.950 ;
        RECT 124.390 105.810 125.390 106.040 ;
        RECT 125.550 106.000 125.920 106.290 ;
        RECT 125.580 105.940 125.920 106.000 ;
        RECT 126.680 106.610 127.440 106.660 ;
        RECT 128.320 106.610 128.550 106.710 ;
        RECT 126.680 106.400 128.550 106.610 ;
        RECT 136.960 106.400 137.190 106.710 ;
        RECT 126.680 105.980 129.220 106.400 ;
        RECT 136.590 105.980 137.190 106.400 ;
        RECT 124.450 105.660 125.330 105.810 ;
        RECT 124.460 105.490 125.190 105.660 ;
        RECT 106.090 103.960 118.550 104.040 ;
        RECT 106.090 103.940 118.420 103.960 ;
        RECT 105.560 103.780 105.900 103.890 ;
        RECT 106.130 103.930 111.800 103.940 ;
        RECT 112.800 103.930 118.420 103.940 ;
        RECT 14.335 103.510 14.625 103.555 ;
        RECT 20.300 103.510 20.620 103.570 ;
        RECT 21.220 103.510 21.540 103.570 ;
        RECT 32.275 103.510 32.565 103.555 ;
        RECT 14.335 103.370 21.540 103.510 ;
        RECT 14.335 103.325 14.625 103.370 ;
        RECT 20.300 103.310 20.620 103.370 ;
        RECT 21.220 103.310 21.540 103.370 ;
        RECT 22.690 103.370 32.565 103.510 ;
        RECT 22.690 103.230 22.830 103.370 ;
        RECT 32.275 103.325 32.565 103.370 ;
        RECT 37.335 103.510 37.625 103.555 ;
        RECT 38.240 103.510 38.560 103.570 ;
        RECT 37.335 103.370 38.560 103.510 ;
        RECT 37.335 103.325 37.625 103.370 ;
        RECT 38.240 103.310 38.560 103.370 ;
        RECT 38.715 103.510 39.005 103.555 ;
        RECT 41.920 103.510 42.240 103.570 ;
        RECT 38.715 103.370 42.240 103.510 ;
        RECT 38.715 103.325 39.005 103.370 ;
        RECT 41.920 103.310 42.240 103.370 ;
        RECT 45.140 103.310 45.460 103.570 ;
        RECT 49.280 103.510 49.600 103.570 ;
        RECT 49.755 103.510 50.045 103.555 ;
        RECT 49.280 103.370 50.045 103.510 ;
        RECT 49.280 103.310 49.600 103.370 ;
        RECT 49.755 103.325 50.045 103.370 ;
        RECT 52.055 103.510 52.345 103.555 ;
        RECT 53.880 103.510 54.200 103.570 ;
        RECT 52.055 103.370 54.200 103.510 ;
        RECT 52.055 103.325 52.345 103.370 ;
        RECT 53.880 103.310 54.200 103.370 ;
        RECT 86.080 103.310 86.400 103.570 ;
        RECT 102.440 103.530 105.300 103.700 ;
        RECT 106.130 103.530 107.465 103.930 ;
        RECT 22.600 103.170 22.920 103.230 ;
        RECT 17.170 103.030 22.920 103.170 ;
        RECT 10.640 102.490 10.960 102.550 ;
        RECT 13.875 102.490 14.165 102.535 ;
        RECT 10.640 102.350 14.165 102.490 ;
        RECT 10.640 102.290 10.960 102.350 ;
        RECT 13.875 102.305 14.165 102.350 ;
        RECT 16.175 102.490 16.465 102.535 ;
        RECT 16.620 102.490 16.940 102.550 ;
        RECT 17.170 102.535 17.310 103.030 ;
        RECT 22.600 102.970 22.920 103.030 ;
        RECT 25.860 103.170 26.150 103.215 ;
        RECT 27.960 103.170 28.250 103.215 ;
        RECT 29.530 103.170 29.820 103.215 ;
        RECT 43.775 103.170 44.065 103.215 ;
        RECT 25.860 103.030 29.820 103.170 ;
        RECT 25.860 102.985 26.150 103.030 ;
        RECT 27.960 102.985 28.250 103.030 ;
        RECT 29.530 102.985 29.820 103.030 ;
        RECT 40.170 103.030 44.065 103.170 ;
        RECT 22.140 102.630 22.460 102.890 ;
        RECT 25.360 102.630 25.680 102.890 ;
        RECT 26.255 102.830 26.545 102.875 ;
        RECT 27.445 102.830 27.735 102.875 ;
        RECT 29.965 102.830 30.255 102.875 ;
        RECT 40.170 102.830 40.310 103.030 ;
        RECT 43.775 102.985 44.065 103.030 ;
        RECT 54.800 103.170 55.090 103.215 ;
        RECT 56.370 103.170 56.660 103.215 ;
        RECT 58.470 103.170 58.760 103.215 ;
        RECT 54.800 103.030 58.760 103.170 ;
        RECT 54.800 102.985 55.090 103.030 ;
        RECT 56.370 102.985 56.660 103.030 ;
        RECT 58.470 102.985 58.760 103.030 ;
        RECT 64.475 103.170 64.765 103.215 ;
        RECT 66.760 103.170 67.080 103.230 ;
        RECT 75.960 103.170 76.280 103.230 ;
        RECT 64.475 103.030 67.080 103.170 ;
        RECT 64.475 102.985 64.765 103.030 ;
        RECT 66.760 102.970 67.080 103.030 ;
        RECT 72.830 103.030 76.280 103.170 ;
        RECT 43.300 102.830 43.620 102.890 ;
        RECT 26.255 102.690 30.255 102.830 ;
        RECT 26.255 102.645 26.545 102.690 ;
        RECT 27.445 102.645 27.735 102.690 ;
        RECT 29.965 102.645 30.255 102.690 ;
        RECT 37.870 102.690 40.310 102.830 ;
        RECT 16.175 102.350 16.940 102.490 ;
        RECT 16.175 102.305 16.465 102.350 ;
        RECT 16.620 102.290 16.940 102.350 ;
        RECT 17.095 102.305 17.385 102.535 ;
        RECT 18.000 102.290 18.320 102.550 ;
        RECT 22.615 102.490 22.905 102.535 ;
        RECT 24.900 102.490 25.220 102.550 ;
        RECT 37.870 102.535 38.010 102.690 ;
        RECT 22.615 102.350 25.220 102.490 ;
        RECT 22.615 102.305 22.905 102.350 ;
        RECT 24.900 102.290 25.220 102.350 ;
        RECT 36.875 102.305 37.165 102.535 ;
        RECT 37.795 102.305 38.085 102.535 ;
        RECT 16.710 102.150 16.850 102.290 ;
        RECT 22.140 102.150 22.460 102.210 ;
        RECT 26.600 102.150 26.890 102.195 ;
        RECT 16.710 102.010 22.460 102.150 ;
        RECT 22.140 101.950 22.460 102.010 ;
        RECT 24.530 102.010 26.890 102.150 ;
        RECT 36.950 102.150 37.090 102.305 ;
        RECT 39.620 102.290 39.940 102.550 ;
        RECT 40.170 102.535 40.310 102.690 ;
        RECT 41.090 102.690 43.620 102.830 ;
        RECT 40.095 102.490 40.385 102.535 ;
        RECT 40.540 102.490 40.860 102.550 ;
        RECT 41.090 102.535 41.230 102.690 ;
        RECT 43.300 102.630 43.620 102.690 ;
        RECT 54.365 102.830 54.655 102.875 ;
        RECT 56.885 102.830 57.175 102.875 ;
        RECT 58.075 102.830 58.365 102.875 ;
        RECT 54.365 102.690 58.365 102.830 ;
        RECT 54.365 102.645 54.655 102.690 ;
        RECT 56.885 102.645 57.175 102.690 ;
        RECT 58.075 102.645 58.365 102.690 ;
        RECT 60.320 102.830 60.640 102.890 ;
        RECT 61.715 102.830 62.005 102.875 ;
        RECT 60.320 102.690 62.005 102.830 ;
        RECT 60.320 102.630 60.640 102.690 ;
        RECT 61.715 102.645 62.005 102.690 ;
        RECT 62.635 102.830 62.925 102.875 ;
        RECT 71.835 102.830 72.125 102.875 ;
        RECT 62.635 102.690 72.125 102.830 ;
        RECT 62.635 102.645 62.925 102.690 ;
        RECT 71.835 102.645 72.125 102.690 ;
        RECT 40.095 102.350 40.860 102.490 ;
        RECT 40.095 102.305 40.385 102.350 ;
        RECT 40.540 102.290 40.860 102.350 ;
        RECT 41.015 102.305 41.305 102.535 ;
        RECT 41.460 102.290 41.780 102.550 ;
        RECT 41.935 102.305 42.225 102.535 ;
        RECT 42.855 102.490 43.145 102.535 ;
        RECT 43.760 102.490 44.080 102.550 ;
        RECT 42.855 102.350 44.080 102.490 ;
        RECT 42.855 102.305 43.145 102.350 ;
        RECT 42.010 102.150 42.150 102.305 ;
        RECT 43.760 102.290 44.080 102.350 ;
        RECT 44.220 102.290 44.540 102.550 ;
        RECT 50.215 102.490 50.505 102.535 ;
        RECT 55.720 102.490 56.040 102.550 ;
        RECT 58.955 102.490 59.245 102.535 ;
        RECT 50.215 102.350 54.570 102.490 ;
        RECT 50.215 102.305 50.505 102.350 ;
        RECT 54.430 102.210 54.570 102.350 ;
        RECT 55.720 102.350 59.245 102.490 ;
        RECT 55.720 102.290 56.040 102.350 ;
        RECT 58.955 102.305 59.245 102.350 ;
        RECT 63.540 102.290 63.860 102.550 ;
        RECT 65.380 102.290 65.700 102.550 ;
        RECT 65.840 102.490 66.160 102.550 ;
        RECT 72.830 102.535 72.970 103.030 ;
        RECT 75.960 102.970 76.280 103.030 ;
        RECT 79.680 103.170 79.970 103.215 ;
        RECT 81.780 103.170 82.070 103.215 ;
        RECT 83.350 103.170 83.640 103.215 ;
        RECT 79.680 103.030 83.640 103.170 ;
        RECT 102.410 103.160 107.465 103.530 ;
        RECT 79.680 102.985 79.970 103.030 ;
        RECT 81.780 102.985 82.070 103.030 ;
        RECT 83.350 102.985 83.640 103.030 ;
        RECT 106.195 102.975 107.465 103.160 ;
        RECT 73.215 102.830 73.505 102.875 ;
        RECT 73.660 102.830 73.980 102.890 ;
        RECT 75.500 102.830 75.820 102.890 ;
        RECT 73.215 102.690 73.980 102.830 ;
        RECT 73.215 102.645 73.505 102.690 ;
        RECT 73.660 102.630 73.980 102.690 ;
        RECT 74.210 102.690 75.820 102.830 ;
        RECT 74.210 102.535 74.350 102.690 ;
        RECT 75.500 102.630 75.820 102.690 ;
        RECT 80.075 102.830 80.365 102.875 ;
        RECT 81.265 102.830 81.555 102.875 ;
        RECT 83.785 102.830 84.075 102.875 ;
        RECT 80.075 102.690 84.075 102.830 ;
        RECT 80.075 102.645 80.365 102.690 ;
        RECT 81.265 102.645 81.555 102.690 ;
        RECT 83.785 102.645 84.075 102.690 ;
        RECT 66.315 102.490 66.605 102.535 ;
        RECT 65.840 102.350 66.605 102.490 ;
        RECT 65.840 102.290 66.160 102.350 ;
        RECT 66.315 102.305 66.605 102.350 ;
        RECT 71.375 102.305 71.665 102.535 ;
        RECT 72.295 102.305 72.585 102.535 ;
        RECT 72.755 102.305 73.045 102.535 ;
        RECT 74.135 102.305 74.425 102.535 ;
        RECT 74.595 102.305 74.885 102.535 ;
        RECT 36.950 102.010 42.150 102.150 ;
        RECT 17.080 101.610 17.400 101.870 ;
        RECT 20.760 101.610 21.080 101.870 ;
        RECT 24.530 101.855 24.670 102.010 ;
        RECT 26.600 101.965 26.890 102.010 ;
        RECT 40.170 101.870 40.310 102.010 ;
        RECT 54.340 101.950 54.660 102.210 ;
        RECT 57.730 102.150 58.020 102.195 ;
        RECT 61.255 102.150 61.545 102.195 ;
        RECT 65.470 102.150 65.610 102.290 ;
        RECT 57.730 102.010 59.630 102.150 ;
        RECT 57.730 101.965 58.020 102.010 ;
        RECT 24.455 101.625 24.745 101.855 ;
        RECT 40.080 101.610 40.400 101.870 ;
        RECT 59.490 101.855 59.630 102.010 ;
        RECT 61.255 102.010 65.610 102.150 ;
        RECT 61.255 101.965 61.545 102.010 ;
        RECT 59.415 101.625 59.705 101.855 ;
        RECT 64.920 101.810 65.240 101.870 ;
        RECT 65.855 101.810 66.145 101.855 ;
        RECT 64.920 101.670 66.145 101.810 ;
        RECT 71.450 101.810 71.590 102.305 ;
        RECT 72.370 102.150 72.510 102.305 ;
        RECT 73.200 102.150 73.520 102.210 ;
        RECT 74.670 102.150 74.810 102.305 ;
        RECT 79.180 102.290 79.500 102.550 ;
        RECT 72.370 102.010 74.810 102.150 ;
        RECT 80.530 102.150 80.820 102.195 ;
        RECT 81.020 102.150 81.340 102.210 ;
        RECT 80.530 102.010 81.340 102.150 ;
        RECT 73.200 101.950 73.520 102.010 ;
        RECT 80.530 101.965 80.820 102.010 ;
        RECT 81.020 101.950 81.340 102.010 ;
        RECT 73.660 101.810 73.980 101.870 ;
        RECT 71.450 101.670 73.980 101.810 ;
        RECT 64.920 101.610 65.240 101.670 ;
        RECT 65.855 101.625 66.145 101.670 ;
        RECT 73.660 101.610 73.980 101.670 ;
        RECT 75.515 101.810 75.805 101.855 ;
        RECT 83.780 101.810 84.100 101.870 ;
        RECT 75.515 101.670 84.100 101.810 ;
        RECT 75.515 101.625 75.805 101.670 ;
        RECT 83.780 101.610 84.100 101.670 ;
        RECT 11.950 100.990 90.610 101.470 ;
        RECT 106.195 101.085 107.455 102.975 ;
        RECT 119.900 102.760 120.990 105.420 ;
        RECT 122.340 104.370 125.190 105.490 ;
        RECT 125.580 105.190 125.930 105.940 ;
        RECT 126.680 105.820 128.550 105.980 ;
        RECT 126.680 105.770 127.440 105.820 ;
        RECT 128.320 105.750 128.550 105.820 ;
        RECT 136.960 105.750 137.190 105.980 ;
        RECT 128.755 105.470 136.755 105.700 ;
        RECT 125.580 105.130 125.870 105.190 ;
        RECT 125.490 105.010 125.870 105.130 ;
        RECT 128.850 105.070 136.710 105.470 ;
        RECT 137.520 105.070 138.480 114.550 ;
        RECT 139.930 116.780 140.700 120.420 ;
        RECT 142.370 119.370 145.220 120.490 ;
        RECT 145.610 120.190 145.960 120.940 ;
        RECT 146.710 120.820 148.580 120.980 ;
        RECT 146.710 120.770 147.470 120.820 ;
        RECT 148.350 120.750 148.580 120.820 ;
        RECT 156.990 120.750 157.220 120.980 ;
        RECT 148.785 120.470 156.785 120.700 ;
        RECT 145.610 120.130 145.900 120.190 ;
        RECT 145.520 120.010 145.900 120.130 ;
        RECT 148.880 120.070 156.740 120.470 ;
        RECT 157.550 120.070 158.510 129.550 ;
        RECT 142.310 119.140 145.310 119.370 ;
        RECT 145.520 119.180 145.860 120.010 ;
        RECT 147.870 120.000 158.510 120.070 ;
        RECT 142.360 119.110 145.220 119.140 ;
        RECT 142.360 119.090 143.530 119.110 ;
        RECT 144.490 119.100 145.220 119.110 ;
        RECT 142.310 118.700 145.310 118.930 ;
        RECT 145.515 118.890 145.860 119.180 ;
        RECT 146.050 118.960 158.510 120.000 ;
        RECT 146.050 118.940 158.500 118.960 ;
        RECT 145.520 118.780 145.860 118.890 ;
        RECT 146.090 118.930 151.760 118.940 ;
        RECT 152.760 118.930 158.500 118.940 ;
        RECT 142.400 118.530 145.260 118.700 ;
        RECT 146.090 118.530 146.520 118.930 ;
        RECT 142.370 118.160 146.520 118.530 ;
        RECT 139.930 114.680 140.790 116.780 ;
        RECT 146.460 116.390 147.710 116.830 ;
        RECT 157.640 116.810 158.500 118.930 ;
        RECT 144.400 116.380 149.640 116.390 ;
        RECT 141.450 116.280 156.750 116.380 ;
        RECT 141.450 116.270 156.785 116.280 ;
        RECT 141.410 116.150 156.785 116.270 ;
        RECT 141.410 116.040 145.410 116.150 ;
        RECT 146.460 116.070 148.200 116.150 ;
        RECT 148.780 116.070 156.785 116.150 ;
        RECT 146.460 115.990 147.710 116.070 ;
        RECT 148.785 116.050 156.785 116.070 ;
        RECT 141.020 115.740 141.250 115.990 ;
        RECT 145.570 115.850 145.800 115.990 ;
        RECT 148.350 115.850 148.580 116.000 ;
        RECT 145.570 115.740 148.580 115.850 ;
        RECT 156.990 115.740 157.220 116.000 ;
        RECT 141.020 115.300 157.220 115.740 ;
        RECT 141.020 115.030 141.250 115.300 ;
        RECT 145.570 115.270 157.220 115.300 ;
        RECT 145.570 115.180 148.580 115.270 ;
        RECT 145.570 115.030 145.800 115.180 ;
        RECT 148.350 115.040 148.580 115.180 ;
        RECT 156.990 115.040 157.220 115.270 ;
        RECT 141.410 114.750 145.410 114.980 ;
        RECT 148.785 114.770 156.785 114.990 ;
        RECT 157.550 114.770 158.510 116.810 ;
        RECT 148.785 114.760 158.510 114.770 ;
        RECT 141.410 114.680 145.400 114.750 ;
        RECT 139.930 114.570 145.400 114.680 ;
        RECT 148.840 114.600 158.510 114.760 ;
        RECT 139.930 114.480 143.090 114.570 ;
        RECT 156.580 114.550 158.510 114.600 ;
        RECT 139.930 111.210 140.790 114.480 ;
        RECT 144.440 114.020 149.690 114.030 ;
        RECT 144.440 113.910 156.750 114.020 ;
        RECT 141.470 113.850 156.750 113.910 ;
        RECT 141.470 113.840 156.785 113.850 ;
        RECT 141.410 113.710 156.785 113.840 ;
        RECT 141.410 113.700 146.570 113.710 ;
        RECT 141.410 113.610 145.410 113.700 ;
        RECT 148.785 113.620 156.785 113.710 ;
        RECT 148.870 113.610 156.760 113.620 ;
        RECT 141.020 113.250 141.250 113.560 ;
        RECT 141.470 113.250 145.370 113.610 ;
        RECT 145.570 113.250 145.800 113.560 ;
        RECT 141.020 111.910 145.800 113.250 ;
        RECT 141.020 111.600 141.250 111.910 ;
        RECT 145.570 111.600 145.800 111.910 ;
        RECT 148.350 113.030 148.580 113.570 ;
        RECT 149.390 113.030 150.400 113.060 ;
        RECT 156.990 113.030 157.220 113.570 ;
        RECT 148.350 112.130 157.220 113.030 ;
        RECT 148.350 111.610 148.580 112.130 ;
        RECT 149.390 112.060 150.400 112.130 ;
        RECT 156.990 111.610 157.220 112.130 ;
        RECT 141.410 111.320 145.410 111.550 ;
        RECT 148.785 111.330 156.785 111.560 ;
        RECT 139.930 111.170 141.090 111.210 ;
        RECT 139.930 111.090 141.330 111.170 ;
        RECT 141.700 111.100 145.360 111.320 ;
        RECT 141.700 111.090 143.140 111.100 ;
        RECT 139.930 111.050 143.140 111.090 ;
        RECT 139.930 110.960 142.650 111.050 ;
        RECT 148.850 111.040 156.740 111.330 ;
        RECT 139.930 110.900 141.980 110.960 ;
        RECT 139.930 110.850 141.730 110.900 ;
        RECT 139.930 107.510 140.790 110.850 ;
        RECT 148.840 110.550 156.760 110.560 ;
        RECT 145.070 110.540 156.760 110.550 ;
        RECT 141.450 110.420 156.760 110.540 ;
        RECT 141.450 110.410 156.785 110.420 ;
        RECT 141.410 110.290 156.785 110.410 ;
        RECT 141.410 110.180 145.410 110.290 ;
        RECT 141.020 109.840 141.250 110.130 ;
        RECT 141.470 109.840 145.360 110.180 ;
        RECT 145.570 109.840 145.800 110.130 ;
        RECT 141.020 108.470 145.800 109.840 ;
        RECT 141.020 108.170 141.250 108.470 ;
        RECT 145.570 108.170 145.800 108.470 ;
        RECT 141.410 107.890 145.410 108.120 ;
        RECT 141.660 107.660 145.230 107.890 ;
        RECT 141.660 107.510 145.350 107.660 ;
        RECT 139.930 107.230 145.350 107.510 ;
        RECT 146.600 107.340 147.220 110.290 ;
        RECT 148.785 110.190 156.785 110.290 ;
        RECT 148.840 110.180 156.760 110.190 ;
        RECT 148.350 109.480 148.580 110.140 ;
        RECT 149.360 109.480 150.360 109.570 ;
        RECT 156.990 109.480 157.220 110.140 ;
        RECT 148.350 108.660 157.220 109.480 ;
        RECT 148.350 108.180 148.580 108.660 ;
        RECT 149.360 108.570 150.360 108.660 ;
        RECT 156.990 108.180 157.220 108.660 ;
        RECT 148.785 107.900 156.785 108.130 ;
        RECT 139.930 106.770 145.360 107.230 ;
        RECT 139.930 106.630 141.960 106.770 ;
        RECT 139.960 105.430 141.960 106.630 ;
        RECT 143.710 106.760 145.360 106.770 ;
        RECT 142.400 105.490 143.400 106.210 ;
        RECT 143.710 105.950 144.020 106.760 ;
        RECT 144.480 106.480 145.360 106.760 ;
        RECT 145.600 106.940 147.220 107.340 ;
        RECT 148.870 106.990 156.740 107.900 ;
        RECT 144.420 106.250 145.420 106.480 ;
        RECT 145.600 106.290 145.950 106.940 ;
        RECT 146.600 106.930 147.220 106.940 ;
        RECT 148.785 106.760 156.785 106.990 ;
        RECT 148.870 106.750 156.740 106.760 ;
        RECT 144.480 106.040 145.360 106.060 ;
        RECT 143.750 105.660 144.020 105.950 ;
        RECT 144.420 105.810 145.420 106.040 ;
        RECT 145.580 106.000 145.950 106.290 ;
        RECT 145.610 105.940 145.950 106.000 ;
        RECT 146.710 106.610 147.470 106.660 ;
        RECT 148.350 106.610 148.580 106.710 ;
        RECT 146.710 106.400 148.580 106.610 ;
        RECT 156.990 106.400 157.220 106.710 ;
        RECT 146.710 105.980 149.250 106.400 ;
        RECT 156.620 105.980 157.220 106.400 ;
        RECT 144.480 105.660 145.360 105.810 ;
        RECT 144.490 105.490 145.220 105.660 ;
        RECT 140.040 105.420 141.960 105.430 ;
        RECT 122.280 104.140 125.280 104.370 ;
        RECT 125.490 104.180 125.830 105.010 ;
        RECT 127.840 105.000 138.480 105.070 ;
        RECT 122.330 104.110 125.190 104.140 ;
        RECT 122.330 104.090 123.500 104.110 ;
        RECT 124.460 104.100 125.190 104.110 ;
        RECT 122.280 103.700 125.280 103.930 ;
        RECT 125.485 103.890 125.830 104.180 ;
        RECT 126.020 103.960 138.480 105.000 ;
        RECT 142.370 104.370 145.220 105.490 ;
        RECT 145.610 105.190 145.960 105.940 ;
        RECT 146.710 105.820 148.580 105.980 ;
        RECT 146.710 105.770 147.470 105.820 ;
        RECT 148.350 105.750 148.580 105.820 ;
        RECT 156.990 105.750 157.220 105.980 ;
        RECT 148.785 105.470 156.785 105.700 ;
        RECT 145.610 105.130 145.900 105.190 ;
        RECT 145.520 105.010 145.900 105.130 ;
        RECT 148.880 105.070 156.740 105.470 ;
        RECT 157.550 105.070 158.510 114.550 ;
        RECT 142.310 104.140 145.310 104.370 ;
        RECT 145.520 104.180 145.860 105.010 ;
        RECT 147.870 105.000 158.510 105.070 ;
        RECT 142.360 104.110 145.220 104.140 ;
        RECT 142.360 104.090 143.530 104.110 ;
        RECT 144.490 104.100 145.220 104.110 ;
        RECT 126.020 103.940 138.350 103.960 ;
        RECT 125.490 103.780 125.830 103.890 ;
        RECT 126.060 103.930 131.730 103.940 ;
        RECT 132.730 103.930 138.350 103.940 ;
        RECT 122.370 103.530 125.230 103.700 ;
        RECT 126.060 103.530 126.490 103.930 ;
        RECT 142.310 103.700 145.310 103.930 ;
        RECT 145.515 103.890 145.860 104.180 ;
        RECT 146.050 103.960 158.510 105.000 ;
        RECT 146.050 103.940 158.460 103.960 ;
        RECT 145.520 103.780 145.860 103.890 ;
        RECT 146.090 103.930 151.760 103.940 ;
        RECT 152.760 103.930 158.460 103.940 ;
        RECT 142.400 103.530 145.260 103.700 ;
        RECT 146.090 103.530 146.520 103.930 ;
        RECT 122.340 103.160 126.490 103.530 ;
        RECT 142.370 103.160 146.520 103.530 ;
        RECT 113.040 102.695 116.730 102.710 ;
        RECT 119.900 102.695 135.450 102.760 ;
        RECT 113.040 101.710 135.450 102.695 ;
        RECT 113.040 101.690 132.370 101.710 ;
        RECT 113.040 101.675 123.360 101.690 ;
        RECT 113.040 101.660 116.730 101.675 ;
        RECT 99.990 101.065 112.800 101.085 ;
        RECT 22.140 100.590 22.460 100.850 ;
        RECT 22.600 100.590 22.920 100.850 ;
        RECT 39.620 100.790 39.940 100.850 ;
        RECT 41.475 100.790 41.765 100.835 ;
        RECT 39.620 100.650 41.765 100.790 ;
        RECT 39.620 100.590 39.940 100.650 ;
        RECT 41.475 100.605 41.765 100.650 ;
        RECT 43.315 100.790 43.605 100.835 ;
        RECT 52.500 100.790 52.820 100.850 ;
        RECT 43.315 100.650 52.820 100.790 ;
        RECT 43.315 100.605 43.605 100.650 ;
        RECT 52.500 100.590 52.820 100.650 ;
        RECT 63.095 100.790 63.385 100.835 ;
        RECT 63.540 100.790 63.860 100.850 ;
        RECT 63.095 100.650 63.860 100.790 ;
        RECT 63.095 100.605 63.385 100.650 ;
        RECT 63.540 100.590 63.860 100.650 ;
        RECT 64.015 100.605 64.305 100.835 ;
        RECT 64.460 100.790 64.780 100.850 ;
        RECT 66.300 100.790 66.620 100.850 ;
        RECT 64.460 100.650 66.620 100.790 ;
        RECT 14.750 100.450 15.040 100.495 ;
        RECT 24.915 100.450 25.205 100.495 ;
        RECT 14.750 100.310 25.205 100.450 ;
        RECT 14.750 100.265 15.040 100.310 ;
        RECT 24.915 100.265 25.205 100.310 ;
        RECT 42.380 100.450 42.700 100.510 ;
        RECT 47.440 100.450 47.760 100.510 ;
        RECT 42.380 100.310 47.760 100.450 ;
        RECT 42.380 100.250 42.700 100.310 ;
        RECT 13.400 99.910 13.720 100.170 ;
        RECT 20.760 100.110 21.080 100.170 ;
        RECT 24.455 100.110 24.745 100.155 ;
        RECT 20.760 99.970 24.745 100.110 ;
        RECT 20.760 99.910 21.080 99.970 ;
        RECT 24.455 99.925 24.745 99.970 ;
        RECT 25.375 99.925 25.665 100.155 ;
        RECT 43.775 100.110 44.065 100.155 ;
        RECT 44.680 100.110 45.000 100.170 ;
        RECT 45.690 100.155 45.830 100.310 ;
        RECT 47.440 100.250 47.760 100.310 ;
        RECT 55.260 100.450 55.580 100.510 ;
        RECT 55.735 100.450 56.025 100.495 ;
        RECT 55.260 100.310 56.025 100.450 ;
        RECT 55.260 100.250 55.580 100.310 ;
        RECT 55.735 100.265 56.025 100.310 ;
        RECT 57.530 100.450 57.820 100.495 ;
        RECT 64.090 100.450 64.230 100.605 ;
        RECT 64.460 100.590 64.780 100.650 ;
        RECT 66.300 100.590 66.620 100.650 ;
        RECT 73.200 100.590 73.520 100.850 ;
        RECT 75.040 100.790 75.360 100.850 ;
        RECT 75.975 100.790 76.265 100.835 ;
        RECT 75.040 100.650 76.265 100.790 ;
        RECT 75.040 100.590 75.360 100.650 ;
        RECT 75.975 100.605 76.265 100.650 ;
        RECT 81.020 100.590 81.340 100.850 ;
        RECT 82.860 100.590 83.180 100.850 ;
        RECT 79.195 100.450 79.485 100.495 ;
        RECT 57.530 100.310 64.230 100.450 ;
        RECT 75.130 100.310 79.485 100.450 ;
        RECT 57.530 100.265 57.820 100.310 ;
        RECT 46.980 100.155 47.300 100.170 ;
        RECT 43.775 99.970 45.000 100.110 ;
        RECT 43.775 99.925 44.065 99.970 ;
        RECT 14.295 99.770 14.585 99.815 ;
        RECT 15.485 99.770 15.775 99.815 ;
        RECT 18.005 99.770 18.295 99.815 ;
        RECT 21.570 99.770 21.860 99.815 ;
        RECT 14.295 99.630 18.295 99.770 ;
        RECT 14.295 99.585 14.585 99.630 ;
        RECT 15.485 99.585 15.775 99.630 ;
        RECT 18.005 99.585 18.295 99.630 ;
        RECT 20.390 99.630 21.860 99.770 ;
        RECT 13.900 99.430 14.190 99.475 ;
        RECT 16.000 99.430 16.290 99.475 ;
        RECT 17.570 99.430 17.860 99.475 ;
        RECT 13.900 99.290 17.860 99.430 ;
        RECT 13.900 99.245 14.190 99.290 ;
        RECT 16.000 99.245 16.290 99.290 ;
        RECT 17.570 99.245 17.860 99.290 ;
        RECT 20.390 99.150 20.530 99.630 ;
        RECT 21.570 99.585 21.860 99.630 ;
        RECT 23.980 99.570 24.300 99.830 ;
        RECT 24.900 99.770 25.220 99.830 ;
        RECT 25.450 99.770 25.590 99.925 ;
        RECT 44.680 99.910 45.000 99.970 ;
        RECT 45.615 99.925 45.905 100.155 ;
        RECT 46.950 99.925 47.300 100.155 ;
        RECT 46.980 99.910 47.300 99.925 ;
        RECT 54.800 99.910 55.120 100.170 ;
        RECT 64.920 100.110 65.240 100.170 ;
        RECT 65.855 100.110 66.145 100.155 ;
        RECT 64.920 99.970 66.145 100.110 ;
        RECT 64.920 99.910 65.240 99.970 ;
        RECT 65.855 99.925 66.145 99.970 ;
        RECT 67.680 100.110 68.000 100.170 ;
        RECT 70.915 100.110 71.205 100.155 ;
        RECT 67.680 99.970 71.205 100.110 ;
        RECT 67.680 99.910 68.000 99.970 ;
        RECT 70.915 99.925 71.205 99.970 ;
        RECT 72.295 100.110 72.585 100.155 ;
        RECT 72.740 100.110 73.060 100.170 ;
        RECT 72.295 99.970 73.060 100.110 ;
        RECT 72.295 99.925 72.585 99.970 ;
        RECT 72.740 99.910 73.060 99.970 ;
        RECT 74.120 99.910 74.440 100.170 ;
        RECT 74.580 100.110 74.900 100.170 ;
        RECT 75.130 100.155 75.270 100.310 ;
        RECT 79.195 100.265 79.485 100.310 ;
        RECT 99.970 100.255 112.810 101.065 ;
        RECT 99.990 100.195 112.800 100.255 ;
        RECT 75.055 100.110 75.345 100.155 ;
        RECT 77.815 100.110 78.105 100.155 ;
        RECT 74.580 99.970 75.345 100.110 ;
        RECT 74.580 99.910 74.900 99.970 ;
        RECT 75.055 99.925 75.345 99.970 ;
        RECT 75.590 99.970 78.105 100.110 ;
        RECT 24.900 99.630 25.590 99.770 ;
        RECT 24.900 99.570 25.220 99.630 ;
        RECT 44.235 99.585 44.525 99.815 ;
        RECT 46.495 99.770 46.785 99.815 ;
        RECT 47.685 99.770 47.975 99.815 ;
        RECT 50.205 99.770 50.495 99.815 ;
        RECT 56.195 99.770 56.485 99.815 ;
        RECT 46.495 99.630 50.495 99.770 ;
        RECT 46.495 99.585 46.785 99.630 ;
        RECT 47.685 99.585 47.975 99.630 ;
        RECT 50.205 99.585 50.495 99.630 ;
        RECT 55.810 99.630 56.485 99.770 ;
        RECT 44.310 99.430 44.450 99.585 ;
        RECT 55.810 99.490 55.950 99.630 ;
        RECT 56.195 99.585 56.485 99.630 ;
        RECT 57.075 99.770 57.365 99.815 ;
        RECT 58.265 99.770 58.555 99.815 ;
        RECT 60.785 99.770 61.075 99.815 ;
        RECT 57.075 99.630 61.075 99.770 ;
        RECT 57.075 99.585 57.365 99.630 ;
        RECT 58.265 99.585 58.555 99.630 ;
        RECT 60.785 99.585 61.075 99.630 ;
        RECT 66.760 99.770 67.080 99.830 ;
        RECT 69.060 99.770 69.380 99.830 ;
        RECT 66.760 99.630 69.380 99.770 ;
        RECT 66.760 99.570 67.080 99.630 ;
        RECT 69.060 99.570 69.380 99.630 ;
        RECT 71.835 99.770 72.125 99.815 ;
        RECT 73.200 99.770 73.520 99.830 ;
        RECT 74.210 99.770 74.350 99.910 ;
        RECT 71.835 99.630 74.350 99.770 ;
        RECT 71.835 99.585 72.125 99.630 ;
        RECT 73.200 99.570 73.520 99.630 ;
        RECT 45.600 99.430 45.920 99.490 ;
        RECT 44.310 99.290 45.920 99.430 ;
        RECT 45.600 99.230 45.920 99.290 ;
        RECT 46.100 99.430 46.390 99.475 ;
        RECT 48.200 99.430 48.490 99.475 ;
        RECT 49.770 99.430 50.060 99.475 ;
        RECT 46.100 99.290 50.060 99.430 ;
        RECT 46.100 99.245 46.390 99.290 ;
        RECT 48.200 99.245 48.490 99.290 ;
        RECT 49.770 99.245 50.060 99.290 ;
        RECT 50.290 99.290 55.030 99.430 ;
        RECT 20.300 98.890 20.620 99.150 ;
        RECT 20.760 98.890 21.080 99.150 ;
        RECT 32.720 99.090 33.040 99.150 ;
        RECT 50.290 99.090 50.430 99.290 ;
        RECT 32.720 98.950 50.430 99.090 ;
        RECT 32.720 98.890 33.040 98.950 ;
        RECT 54.340 98.890 54.660 99.150 ;
        RECT 54.890 99.090 55.030 99.290 ;
        RECT 55.720 99.230 56.040 99.490 ;
        RECT 56.680 99.430 56.970 99.475 ;
        RECT 58.780 99.430 59.070 99.475 ;
        RECT 60.350 99.430 60.640 99.475 ;
        RECT 56.680 99.290 60.640 99.430 ;
        RECT 56.680 99.245 56.970 99.290 ;
        RECT 58.780 99.245 59.070 99.290 ;
        RECT 60.350 99.245 60.640 99.290 ;
        RECT 71.360 99.230 71.680 99.490 ;
        RECT 74.120 99.230 74.440 99.490 ;
        RECT 75.040 99.430 75.360 99.490 ;
        RECT 75.590 99.430 75.730 99.970 ;
        RECT 77.815 99.925 78.105 99.970 ;
        RECT 78.260 99.910 78.580 100.170 ;
        RECT 100.990 99.835 101.430 100.195 ;
        RECT 102.570 100.085 103.730 100.195 ;
        RECT 102.570 99.835 103.010 100.085 ;
        RECT 104.160 99.835 104.600 100.195 ;
        RECT 105.750 99.835 106.190 100.195 ;
        RECT 76.880 99.770 77.200 99.830 ;
        RECT 77.355 99.770 77.645 99.815 ;
        RECT 76.880 99.630 77.645 99.770 ;
        RECT 76.880 99.570 77.200 99.630 ;
        RECT 77.355 99.585 77.645 99.630 ;
        RECT 83.320 99.570 83.640 99.830 ;
        RECT 83.780 99.570 84.100 99.830 ;
        RECT 100.130 99.785 100.360 99.815 ;
        RECT 100.520 99.785 100.750 99.835 ;
        RECT 75.040 99.290 75.730 99.430 ;
        RECT 75.960 99.430 76.280 99.490 ;
        RECT 80.100 99.430 80.420 99.490 ;
        RECT 75.960 99.290 80.420 99.430 ;
        RECT 75.040 99.230 75.360 99.290 ;
        RECT 75.960 99.230 76.280 99.290 ;
        RECT 80.100 99.230 80.420 99.290 ;
        RECT 76.420 99.090 76.740 99.150 ;
        RECT 54.890 98.950 76.740 99.090 ;
        RECT 76.420 98.890 76.740 98.950 ;
        RECT 77.800 98.890 78.120 99.150 ;
        RECT 11.950 98.270 90.610 98.750 ;
        RECT 17.080 98.070 17.400 98.130 ;
        RECT 17.555 98.070 17.845 98.115 ;
        RECT 17.080 97.930 17.845 98.070 ;
        RECT 17.080 97.870 17.400 97.930 ;
        RECT 17.555 97.885 17.845 97.930 ;
        RECT 18.000 97.870 18.320 98.130 ;
        RECT 36.400 98.070 36.720 98.130 ;
        RECT 40.095 98.070 40.385 98.115 ;
        RECT 36.400 97.930 40.385 98.070 ;
        RECT 36.400 97.870 36.720 97.930 ;
        RECT 40.095 97.885 40.385 97.930 ;
        RECT 46.535 98.070 46.825 98.115 ;
        RECT 46.980 98.070 47.300 98.130 ;
        RECT 46.535 97.930 47.300 98.070 ;
        RECT 46.535 97.885 46.825 97.930 ;
        RECT 46.980 97.870 47.300 97.930 ;
        RECT 66.775 98.070 67.065 98.115 ;
        RECT 67.680 98.070 68.000 98.130 ;
        RECT 66.775 97.930 68.000 98.070 ;
        RECT 66.775 97.885 67.065 97.930 ;
        RECT 67.680 97.870 68.000 97.930 ;
        RECT 73.200 97.870 73.520 98.130 ;
        RECT 73.660 98.070 73.980 98.130 ;
        RECT 74.595 98.070 74.885 98.115 ;
        RECT 76.880 98.070 77.200 98.130 ;
        RECT 73.660 97.930 74.885 98.070 ;
        RECT 73.660 97.870 73.980 97.930 ;
        RECT 74.595 97.885 74.885 97.930 ;
        RECT 76.050 97.930 77.200 98.070 ;
        RECT 33.220 97.730 33.510 97.775 ;
        RECT 35.320 97.730 35.610 97.775 ;
        RECT 36.890 97.730 37.180 97.775 ;
        RECT 33.220 97.590 37.180 97.730 ;
        RECT 33.220 97.545 33.510 97.590 ;
        RECT 35.320 97.545 35.610 97.590 ;
        RECT 36.890 97.545 37.180 97.590 ;
        RECT 39.635 97.730 39.925 97.775 ;
        RECT 49.280 97.730 49.600 97.790 ;
        RECT 72.740 97.730 73.060 97.790 ;
        RECT 76.050 97.730 76.190 97.930 ;
        RECT 76.880 97.870 77.200 97.930 ;
        RECT 81.495 98.070 81.785 98.115 ;
        RECT 83.320 98.070 83.640 98.130 ;
        RECT 81.495 97.930 83.640 98.070 ;
        RECT 81.495 97.885 81.785 97.930 ;
        RECT 83.320 97.870 83.640 97.930 ;
        RECT 39.635 97.590 43.070 97.730 ;
        RECT 39.635 97.545 39.925 97.590 ;
        RECT 18.475 97.390 18.765 97.435 ;
        RECT 18.935 97.390 19.225 97.435 ;
        RECT 18.475 97.250 19.225 97.390 ;
        RECT 18.475 97.205 18.765 97.250 ;
        RECT 18.935 97.205 19.225 97.250 ;
        RECT 25.360 97.390 25.680 97.450 ;
        RECT 42.930 97.435 43.070 97.590 ;
        RECT 49.280 97.590 53.190 97.730 ;
        RECT 49.280 97.530 49.600 97.590 ;
        RECT 32.735 97.390 33.025 97.435 ;
        RECT 25.360 97.250 33.025 97.390 ;
        RECT 25.360 97.190 25.680 97.250 ;
        RECT 32.735 97.205 33.025 97.250 ;
        RECT 33.615 97.390 33.905 97.435 ;
        RECT 34.805 97.390 35.095 97.435 ;
        RECT 37.325 97.390 37.615 97.435 ;
        RECT 33.615 97.250 37.615 97.390 ;
        RECT 33.615 97.205 33.905 97.250 ;
        RECT 34.805 97.205 35.095 97.250 ;
        RECT 37.325 97.205 37.615 97.250 ;
        RECT 42.855 97.390 43.145 97.435 ;
        RECT 43.760 97.390 44.080 97.450 ;
        RECT 42.855 97.250 44.080 97.390 ;
        RECT 42.855 97.205 43.145 97.250 ;
        RECT 43.760 97.190 44.080 97.250 ;
        RECT 49.740 97.190 50.060 97.450 ;
        RECT 17.095 96.865 17.385 97.095 ;
        RECT 20.300 97.050 20.620 97.110 ;
        RECT 21.695 97.050 21.985 97.095 ;
        RECT 20.300 96.910 21.985 97.050 ;
        RECT 17.170 96.710 17.310 96.865 ;
        RECT 20.300 96.850 20.620 96.910 ;
        RECT 21.695 96.865 21.985 96.910 ;
        RECT 48.835 97.050 49.125 97.095 ;
        RECT 50.660 97.050 50.980 97.110 ;
        RECT 53.050 97.095 53.190 97.590 ;
        RECT 72.740 97.590 76.190 97.730 ;
        RECT 76.420 97.730 76.740 97.790 ;
        RECT 76.420 97.590 79.410 97.730 ;
        RECT 72.740 97.530 73.060 97.590 ;
        RECT 76.420 97.530 76.740 97.590 ;
        RECT 54.340 97.390 54.660 97.450 ;
        RECT 57.100 97.390 57.420 97.450 ;
        RECT 54.340 97.250 57.420 97.390 ;
        RECT 54.340 97.190 54.660 97.250 ;
        RECT 57.100 97.190 57.420 97.250 ;
        RECT 64.000 97.390 64.320 97.450 ;
        RECT 64.000 97.250 68.370 97.390 ;
        RECT 64.000 97.190 64.320 97.250 ;
        RECT 68.230 97.110 68.370 97.250 ;
        RECT 78.720 97.190 79.040 97.450 ;
        RECT 79.270 97.435 79.410 97.590 ;
        RECT 79.195 97.205 79.485 97.435 ;
        RECT 48.835 96.910 50.980 97.050 ;
        RECT 48.835 96.865 49.125 96.910 ;
        RECT 50.660 96.850 50.980 96.910 ;
        RECT 52.975 96.865 53.265 97.095 ;
        RECT 60.320 96.850 60.640 97.110 ;
        RECT 63.555 97.050 63.845 97.095 ;
        RECT 66.760 97.050 67.080 97.110 ;
        RECT 63.555 96.910 67.080 97.050 ;
        RECT 63.555 96.865 63.845 96.910 ;
        RECT 66.760 96.850 67.080 96.910 ;
        RECT 68.140 96.850 68.460 97.110 ;
        RECT 69.060 96.850 69.380 97.110 ;
        RECT 71.360 97.050 71.680 97.110 ;
        RECT 72.755 97.050 73.045 97.095 ;
        RECT 71.360 96.910 73.045 97.050 ;
        RECT 71.360 96.850 71.680 96.910 ;
        RECT 72.755 96.865 73.045 96.910 ;
        RECT 73.200 96.850 73.520 97.110 ;
        RECT 21.220 96.710 21.540 96.770 ;
        RECT 23.980 96.710 24.300 96.770 ;
        RECT 34.100 96.755 34.420 96.770 ;
        RECT 17.170 96.570 24.300 96.710 ;
        RECT 21.220 96.510 21.540 96.570 ;
        RECT 23.980 96.510 24.300 96.570 ;
        RECT 34.070 96.525 34.420 96.755 ;
        RECT 48.375 96.710 48.665 96.755 ;
        RECT 53.435 96.710 53.725 96.755 ;
        RECT 53.880 96.710 54.200 96.770 ;
        RECT 48.375 96.570 51.350 96.710 ;
        RECT 48.375 96.525 48.665 96.570 ;
        RECT 34.100 96.510 34.420 96.525 ;
        RECT 51.210 96.415 51.350 96.570 ;
        RECT 53.435 96.570 54.200 96.710 ;
        RECT 53.435 96.525 53.725 96.570 ;
        RECT 53.880 96.510 54.200 96.570 ;
        RECT 67.220 96.710 67.540 96.770 ;
        RECT 67.695 96.710 67.985 96.755 ;
        RECT 70.900 96.710 71.220 96.770 ;
        RECT 67.220 96.570 67.985 96.710 ;
        RECT 67.220 96.510 67.540 96.570 ;
        RECT 67.695 96.525 67.985 96.570 ;
        RECT 68.230 96.570 71.220 96.710 ;
        RECT 51.135 96.185 51.425 96.415 ;
        RECT 65.840 96.170 66.160 96.430 ;
        RECT 66.695 96.370 66.985 96.415 ;
        RECT 68.230 96.370 68.370 96.570 ;
        RECT 70.900 96.510 71.220 96.570 ;
        RECT 66.695 96.230 68.370 96.370 ;
        RECT 68.600 96.370 68.920 96.430 ;
        RECT 75.040 96.370 75.360 96.430 ;
        RECT 68.600 96.230 75.360 96.370 ;
        RECT 66.695 96.185 66.985 96.230 ;
        RECT 68.600 96.170 68.920 96.230 ;
        RECT 75.040 96.170 75.360 96.230 ;
        RECT 79.640 96.170 79.960 96.430 ;
        RECT 11.950 95.550 90.610 96.030 ;
        RECT 21.235 95.350 21.525 95.395 ;
        RECT 21.680 95.350 22.000 95.410 ;
        RECT 24.900 95.350 25.220 95.410 ;
        RECT 21.235 95.210 25.220 95.350 ;
        RECT 21.235 95.165 21.525 95.210 ;
        RECT 21.680 95.150 22.000 95.210 ;
        RECT 24.900 95.150 25.220 95.210 ;
        RECT 31.815 95.350 32.105 95.395 ;
        RECT 32.720 95.350 33.040 95.410 ;
        RECT 31.815 95.210 33.040 95.350 ;
        RECT 31.815 95.165 32.105 95.210 ;
        RECT 32.720 95.150 33.040 95.210 ;
        RECT 33.655 95.350 33.945 95.395 ;
        RECT 34.100 95.350 34.420 95.410 ;
        RECT 43.760 95.395 44.080 95.410 ;
        RECT 33.655 95.210 34.420 95.350 ;
        RECT 33.655 95.165 33.945 95.210 ;
        RECT 34.100 95.150 34.420 95.210 ;
        RECT 35.495 95.350 35.785 95.395 ;
        RECT 38.715 95.350 39.005 95.395 ;
        RECT 35.495 95.210 39.005 95.350 ;
        RECT 35.495 95.165 35.785 95.210 ;
        RECT 38.715 95.165 39.005 95.210 ;
        RECT 43.760 95.165 44.145 95.395 ;
        RECT 53.895 95.350 54.185 95.395 ;
        RECT 60.320 95.350 60.640 95.410 ;
        RECT 53.895 95.210 60.640 95.350 ;
        RECT 53.895 95.165 54.185 95.210 ;
        RECT 43.760 95.150 44.080 95.165 ;
        RECT 17.080 95.010 17.400 95.070 ;
        RECT 35.955 95.010 36.245 95.055 ;
        RECT 36.400 95.010 36.720 95.070 ;
        RECT 17.080 94.870 19.610 95.010 ;
        RECT 17.080 94.810 17.400 94.870 ;
        RECT 19.470 94.715 19.610 94.870 ;
        RECT 35.955 94.870 36.720 95.010 ;
        RECT 35.955 94.825 36.245 94.870 ;
        RECT 36.400 94.810 36.720 94.870 ;
        RECT 42.840 94.810 43.160 95.070 ;
        RECT 16.635 94.670 16.925 94.715 ;
        RECT 16.635 94.530 19.150 94.670 ;
        RECT 16.635 94.485 16.925 94.530 ;
        RECT 17.095 94.145 17.385 94.375 ;
        RECT 17.170 93.990 17.310 94.145 ;
        RECT 17.540 94.130 17.860 94.390 ;
        RECT 19.010 94.330 19.150 94.530 ;
        RECT 19.395 94.485 19.685 94.715 ;
        RECT 20.315 94.670 20.605 94.715 ;
        RECT 21.220 94.670 21.540 94.730 ;
        RECT 20.315 94.530 21.540 94.670 ;
        RECT 20.315 94.485 20.605 94.530 ;
        RECT 21.220 94.470 21.540 94.530 ;
        RECT 24.915 94.670 25.205 94.715 ;
        RECT 25.360 94.670 25.680 94.730 ;
        RECT 26.280 94.715 26.600 94.730 ;
        RECT 24.915 94.530 25.680 94.670 ;
        RECT 24.915 94.485 25.205 94.530 ;
        RECT 25.360 94.470 25.680 94.530 ;
        RECT 26.250 94.485 26.600 94.715 ;
        RECT 26.280 94.470 26.600 94.485 ;
        RECT 40.540 94.470 40.860 94.730 ;
        RECT 41.015 94.670 41.305 94.715 ;
        RECT 53.970 94.670 54.110 95.165 ;
        RECT 60.320 95.150 60.640 95.210 ;
        RECT 64.015 95.165 64.305 95.395 ;
        RECT 74.595 95.350 74.885 95.395 ;
        RECT 79.640 95.350 79.960 95.410 ;
        RECT 74.595 95.210 79.960 95.350 ;
        RECT 74.595 95.165 74.885 95.210 ;
        RECT 59.570 95.010 59.860 95.055 ;
        RECT 64.090 95.010 64.230 95.165 ;
        RECT 79.640 95.150 79.960 95.210 ;
        RECT 81.035 95.350 81.325 95.395 ;
        RECT 81.480 95.350 81.800 95.410 ;
        RECT 81.035 95.210 81.800 95.350 ;
        RECT 81.035 95.165 81.325 95.210 ;
        RECT 81.480 95.150 81.800 95.210 ;
        RECT 59.570 94.870 64.230 95.010 ;
        RECT 59.570 94.825 59.860 94.870 ;
        RECT 65.380 94.810 65.700 95.070 ;
        RECT 65.855 95.010 66.145 95.055 ;
        RECT 67.695 95.010 67.985 95.055 ;
        RECT 65.855 94.870 67.985 95.010 ;
        RECT 65.855 94.825 66.145 94.870 ;
        RECT 67.695 94.825 67.985 94.870 ;
        RECT 69.610 94.870 79.870 95.010 ;
        RECT 41.015 94.530 54.110 94.670 ;
        RECT 54.890 94.530 61.470 94.670 ;
        RECT 41.015 94.485 41.305 94.530 ;
        RECT 19.840 94.330 20.160 94.390 ;
        RECT 23.980 94.330 24.300 94.390 ;
        RECT 19.010 94.190 24.300 94.330 ;
        RECT 19.840 94.130 20.160 94.190 ;
        RECT 23.980 94.130 24.300 94.190 ;
        RECT 25.795 94.330 26.085 94.375 ;
        RECT 26.985 94.330 27.275 94.375 ;
        RECT 29.505 94.330 29.795 94.375 ;
        RECT 25.795 94.190 29.795 94.330 ;
        RECT 25.795 94.145 26.085 94.190 ;
        RECT 26.985 94.145 27.275 94.190 ;
        RECT 29.505 94.145 29.795 94.190 ;
        RECT 36.860 94.130 37.180 94.390 ;
        RECT 41.935 94.330 42.225 94.375 ;
        RECT 54.340 94.330 54.660 94.390 ;
        RECT 41.935 94.190 54.660 94.330 ;
        RECT 41.935 94.145 42.225 94.190 ;
        RECT 54.340 94.130 54.660 94.190 ;
        RECT 21.220 93.990 21.540 94.050 ;
        RECT 23.520 93.990 23.840 94.050 ;
        RECT 25.400 93.990 25.690 94.035 ;
        RECT 27.500 93.990 27.790 94.035 ;
        RECT 29.070 93.990 29.360 94.035 ;
        RECT 54.890 93.990 55.030 94.530 ;
        RECT 56.205 94.330 56.495 94.375 ;
        RECT 58.725 94.330 59.015 94.375 ;
        RECT 59.915 94.330 60.205 94.375 ;
        RECT 56.205 94.190 60.205 94.330 ;
        RECT 56.205 94.145 56.495 94.190 ;
        RECT 58.725 94.145 59.015 94.190 ;
        RECT 59.915 94.145 60.205 94.190 ;
        RECT 60.795 94.145 61.085 94.375 ;
        RECT 17.170 93.850 25.130 93.990 ;
        RECT 21.220 93.790 21.540 93.850 ;
        RECT 23.520 93.790 23.840 93.850 ;
        RECT 14.780 93.450 15.100 93.710 ;
        RECT 20.300 93.450 20.620 93.710 ;
        RECT 24.990 93.650 25.130 93.850 ;
        RECT 25.400 93.850 29.360 93.990 ;
        RECT 25.400 93.805 25.690 93.850 ;
        RECT 27.500 93.805 27.790 93.850 ;
        RECT 29.070 93.805 29.360 93.850 ;
        RECT 30.050 93.850 55.030 93.990 ;
        RECT 56.640 93.990 56.930 94.035 ;
        RECT 58.210 93.990 58.500 94.035 ;
        RECT 60.310 93.990 60.600 94.035 ;
        RECT 56.640 93.850 60.600 93.990 ;
        RECT 30.050 93.650 30.190 93.850 ;
        RECT 56.640 93.805 56.930 93.850 ;
        RECT 58.210 93.805 58.500 93.850 ;
        RECT 60.310 93.805 60.600 93.850 ;
        RECT 24.990 93.510 30.190 93.650 ;
        RECT 43.760 93.450 44.080 93.710 ;
        RECT 44.695 93.650 44.985 93.695 ;
        RECT 46.980 93.650 47.300 93.710 ;
        RECT 44.695 93.510 47.300 93.650 ;
        RECT 44.695 93.465 44.985 93.510 ;
        RECT 46.980 93.450 47.300 93.510 ;
        RECT 55.720 93.650 56.040 93.710 ;
        RECT 60.870 93.650 61.010 94.145 ;
        RECT 61.330 93.990 61.470 94.530 ;
        RECT 64.935 94.485 65.225 94.715 ;
        RECT 65.010 94.330 65.150 94.485 ;
        RECT 66.760 94.470 67.080 94.730 ;
        RECT 68.600 94.470 68.920 94.730 ;
        RECT 69.060 94.470 69.380 94.730 ;
        RECT 67.680 94.330 68.000 94.390 ;
        RECT 65.010 94.190 68.000 94.330 ;
        RECT 67.680 94.130 68.000 94.190 ;
        RECT 69.610 93.990 69.750 94.870 ;
        RECT 69.995 94.485 70.285 94.715 ;
        RECT 70.070 94.330 70.210 94.485 ;
        RECT 70.440 94.470 70.760 94.730 ;
        RECT 71.360 94.670 71.680 94.730 ;
        RECT 72.755 94.670 73.045 94.715 ;
        RECT 71.360 94.530 73.045 94.670 ;
        RECT 71.360 94.470 71.680 94.530 ;
        RECT 72.755 94.485 73.045 94.530 ;
        RECT 75.040 94.470 75.360 94.730 ;
        RECT 75.975 94.670 76.265 94.715 ;
        RECT 76.420 94.670 76.740 94.730 ;
        RECT 75.975 94.530 76.740 94.670 ;
        RECT 75.975 94.485 76.265 94.530 ;
        RECT 76.420 94.470 76.740 94.530 ;
        RECT 76.895 94.670 77.185 94.715 ;
        RECT 78.275 94.670 78.565 94.715 ;
        RECT 76.895 94.530 78.565 94.670 ;
        RECT 76.895 94.485 77.185 94.530 ;
        RECT 78.275 94.485 78.565 94.530 ;
        RECT 78.720 94.670 79.040 94.730 ;
        RECT 79.730 94.715 79.870 94.870 ;
        RECT 79.195 94.670 79.485 94.715 ;
        RECT 78.720 94.530 79.485 94.670 ;
        RECT 78.720 94.470 79.040 94.530 ;
        RECT 79.195 94.485 79.485 94.530 ;
        RECT 79.655 94.485 79.945 94.715 ;
        RECT 80.115 94.485 80.405 94.715 ;
        RECT 71.820 94.330 72.140 94.390 ;
        RECT 70.070 94.190 72.140 94.330 ;
        RECT 71.820 94.130 72.140 94.190 ;
        RECT 73.215 94.145 73.505 94.375 ;
        RECT 75.500 94.330 75.820 94.390 ;
        RECT 77.800 94.330 78.120 94.390 ;
        RECT 80.190 94.330 80.330 94.485 ;
        RECT 75.500 94.190 80.330 94.330 ;
        RECT 61.330 93.850 69.750 93.990 ;
        RECT 73.290 93.990 73.430 94.145 ;
        RECT 75.500 94.130 75.820 94.190 ;
        RECT 77.800 94.130 78.120 94.190 ;
        RECT 76.420 93.990 76.740 94.050 ;
        RECT 73.290 93.850 76.740 93.990 ;
        RECT 76.420 93.790 76.740 93.850 ;
        RECT 100.130 93.895 100.750 99.785 ;
        RECT 55.720 93.510 61.010 93.650 ;
        RECT 65.840 93.650 66.160 93.710 ;
        RECT 68.140 93.650 68.460 93.710 ;
        RECT 70.440 93.650 70.760 93.710 ;
        RECT 65.840 93.510 70.760 93.650 ;
        RECT 55.720 93.450 56.040 93.510 ;
        RECT 65.840 93.450 66.160 93.510 ;
        RECT 68.140 93.450 68.460 93.510 ;
        RECT 70.440 93.450 70.760 93.510 ;
        RECT 73.675 93.650 73.965 93.695 ;
        RECT 77.340 93.650 77.660 93.710 ;
        RECT 73.675 93.510 77.660 93.650 ;
        RECT 73.675 93.465 73.965 93.510 ;
        RECT 77.340 93.450 77.660 93.510 ;
        RECT 100.130 93.615 100.370 93.895 ;
        RECT 100.520 93.835 100.750 93.895 ;
        RECT 100.960 93.895 101.430 99.835 ;
        RECT 102.100 99.765 102.330 99.835 ;
        RECT 101.800 93.915 102.330 99.765 ;
        RECT 101.800 93.895 101.960 93.915 ;
        RECT 100.960 93.835 101.190 93.895 ;
        RECT 101.810 93.655 101.960 93.895 ;
        RECT 102.100 93.835 102.330 93.915 ;
        RECT 102.540 93.915 103.010 99.835 ;
        RECT 103.680 99.765 103.910 99.835 ;
        RECT 103.310 95.175 103.920 99.765 ;
        RECT 102.540 93.835 102.770 93.915 ;
        RECT 103.290 93.885 103.920 95.175 ;
        RECT 104.120 93.925 104.600 99.835 ;
        RECT 105.260 99.785 105.490 99.835 ;
        RECT 11.950 92.830 90.610 93.310 ;
        RECT 20.315 92.630 20.605 92.675 ;
        RECT 21.220 92.630 21.540 92.690 ;
        RECT 20.315 92.490 21.540 92.630 ;
        RECT 20.315 92.445 20.605 92.490 ;
        RECT 21.220 92.430 21.540 92.490 ;
        RECT 23.060 92.430 23.380 92.690 ;
        RECT 23.995 92.630 24.285 92.675 ;
        RECT 24.440 92.630 24.760 92.690 ;
        RECT 23.995 92.490 24.760 92.630 ;
        RECT 23.995 92.445 24.285 92.490 ;
        RECT 24.440 92.430 24.760 92.490 ;
        RECT 25.835 92.630 26.125 92.675 ;
        RECT 26.280 92.630 26.600 92.690 ;
        RECT 25.835 92.490 26.600 92.630 ;
        RECT 25.835 92.445 26.125 92.490 ;
        RECT 26.280 92.430 26.600 92.490 ;
        RECT 47.455 92.630 47.745 92.675 ;
        RECT 47.900 92.630 48.220 92.690 ;
        RECT 47.455 92.490 48.220 92.630 ;
        RECT 47.455 92.445 47.745 92.490 ;
        RECT 47.900 92.430 48.220 92.490 ;
        RECT 70.915 92.445 71.205 92.675 ;
        RECT 71.360 92.630 71.680 92.690 ;
        RECT 71.835 92.630 72.125 92.675 ;
        RECT 71.360 92.490 72.125 92.630 ;
        RECT 13.900 92.290 14.190 92.335 ;
        RECT 16.000 92.290 16.290 92.335 ;
        RECT 17.570 92.290 17.860 92.335 ;
        RECT 13.900 92.150 17.860 92.290 ;
        RECT 13.900 92.105 14.190 92.150 ;
        RECT 16.000 92.105 16.290 92.150 ;
        RECT 17.570 92.105 17.860 92.150 ;
        RECT 13.400 91.750 13.720 92.010 ;
        RECT 14.295 91.950 14.585 91.995 ;
        RECT 15.485 91.950 15.775 91.995 ;
        RECT 18.005 91.950 18.295 91.995 ;
        RECT 21.680 91.950 22.000 92.010 ;
        RECT 14.295 91.810 18.295 91.950 ;
        RECT 14.295 91.765 14.585 91.810 ;
        RECT 15.485 91.765 15.775 91.810 ;
        RECT 18.005 91.765 18.295 91.810 ;
        RECT 20.850 91.810 22.000 91.950 ;
        RECT 24.530 91.950 24.670 92.430 ;
        RECT 28.595 91.950 28.885 91.995 ;
        RECT 24.530 91.810 28.885 91.950 ;
        RECT 13.490 91.610 13.630 91.750 ;
        RECT 20.300 91.610 20.620 91.670 ;
        RECT 13.490 91.470 20.620 91.610 ;
        RECT 20.300 91.410 20.620 91.470 ;
        RECT 14.780 91.315 15.100 91.330 ;
        RECT 14.750 91.270 15.100 91.315 ;
        RECT 14.585 91.130 15.100 91.270 ;
        RECT 14.750 91.085 15.100 91.130 ;
        RECT 14.780 91.070 15.100 91.085 ;
        RECT 17.540 91.270 17.860 91.330 ;
        RECT 20.850 91.270 20.990 91.810 ;
        RECT 21.680 91.750 22.000 91.810 ;
        RECT 28.595 91.765 28.885 91.810 ;
        RECT 37.320 91.950 37.640 92.010 ;
        RECT 39.635 91.950 39.925 91.995 ;
        RECT 40.540 91.950 40.860 92.010 ;
        RECT 67.220 91.950 67.540 92.010 ;
        RECT 70.990 91.950 71.130 92.445 ;
        RECT 71.360 92.430 71.680 92.490 ;
        RECT 71.835 92.445 72.125 92.490 ;
        RECT 37.320 91.810 40.860 91.950 ;
        RECT 37.320 91.750 37.640 91.810 ;
        RECT 39.635 91.765 39.925 91.810 ;
        RECT 40.540 91.750 40.860 91.810 ;
        RECT 66.850 91.810 71.130 91.950 ;
        RECT 23.980 91.610 24.300 91.670 ;
        RECT 26.280 91.610 26.600 91.670 ;
        RECT 28.135 91.610 28.425 91.655 ;
        RECT 23.980 91.470 28.425 91.610 ;
        RECT 23.980 91.410 24.300 91.470 ;
        RECT 26.280 91.410 26.600 91.470 ;
        RECT 28.135 91.425 28.425 91.470 ;
        RECT 46.535 91.425 46.825 91.655 ;
        RECT 46.980 91.610 47.300 91.670 ;
        RECT 66.850 91.655 66.990 91.810 ;
        RECT 67.220 91.750 67.540 91.810 ;
        RECT 78.720 91.750 79.040 92.010 ;
        RECT 47.455 91.610 47.745 91.655 ;
        RECT 46.980 91.470 47.745 91.610 ;
        RECT 17.540 91.130 20.990 91.270 ;
        RECT 21.680 91.270 22.000 91.330 ;
        RECT 22.155 91.270 22.445 91.315 ;
        RECT 21.680 91.130 22.445 91.270 ;
        RECT 17.540 91.070 17.860 91.130 ;
        RECT 21.680 91.070 22.000 91.130 ;
        RECT 22.155 91.085 22.445 91.130 ;
        RECT 27.675 91.270 27.965 91.315 ;
        RECT 32.720 91.270 33.040 91.330 ;
        RECT 27.675 91.130 33.040 91.270 ;
        RECT 27.675 91.085 27.965 91.130 ;
        RECT 32.720 91.070 33.040 91.130 ;
        RECT 45.155 91.270 45.445 91.315 ;
        RECT 45.600 91.270 45.920 91.330 ;
        RECT 45.155 91.130 45.920 91.270 ;
        RECT 46.610 91.270 46.750 91.425 ;
        RECT 46.980 91.410 47.300 91.470 ;
        RECT 47.455 91.425 47.745 91.470 ;
        RECT 66.775 91.425 67.065 91.655 ;
        RECT 67.695 91.610 67.985 91.655 ;
        RECT 71.360 91.610 71.680 91.670 ;
        RECT 67.695 91.470 71.680 91.610 ;
        RECT 67.695 91.425 67.985 91.470 ;
        RECT 71.070 91.410 71.680 91.470 ;
        RECT 77.340 91.410 77.660 91.670 ;
        RECT 77.800 91.410 78.120 91.670 ;
        RECT 80.115 91.610 80.405 91.655 ;
        RECT 80.560 91.610 80.880 91.670 ;
        RECT 80.115 91.470 80.880 91.610 ;
        RECT 80.115 91.425 80.405 91.470 ;
        RECT 80.560 91.410 80.880 91.470 ;
        RECT 88.380 91.410 88.700 91.670 ;
        RECT 51.120 91.270 51.440 91.330 ;
        RECT 46.610 91.130 51.440 91.270 ;
        RECT 45.155 91.085 45.445 91.130 ;
        RECT 45.600 91.070 45.920 91.130 ;
        RECT 51.120 91.070 51.440 91.130 ;
        RECT 65.840 91.070 66.160 91.330 ;
        RECT 69.060 91.270 69.380 91.330 ;
        RECT 69.995 91.270 70.285 91.315 ;
        RECT 71.070 91.300 71.435 91.410 ;
        RECT 69.060 91.130 70.285 91.270 ;
        RECT 71.145 91.255 71.435 91.300 ;
        RECT 69.060 91.070 69.380 91.130 ;
        RECT 69.995 91.085 70.285 91.130 ;
        RECT 100.130 91.185 100.510 93.615 ;
        RECT 100.710 93.605 101.000 93.630 ;
        RECT 100.700 92.905 101.020 93.605 ;
        RECT 100.650 91.875 101.650 92.905 ;
        RECT 100.700 91.185 101.020 91.875 ;
        RECT 20.760 90.930 21.080 90.990 ;
        RECT 23.155 90.930 23.445 90.975 ;
        RECT 20.760 90.790 23.445 90.930 ;
        RECT 20.760 90.730 21.080 90.790 ;
        RECT 23.155 90.745 23.445 90.790 ;
        RECT 40.080 90.930 40.400 90.990 ;
        RECT 42.395 90.930 42.685 90.975 ;
        RECT 40.080 90.790 42.685 90.930 ;
        RECT 40.080 90.730 40.400 90.790 ;
        RECT 42.395 90.745 42.685 90.790 ;
        RECT 48.360 90.730 48.680 90.990 ;
        RECT 68.600 90.930 68.920 90.990 ;
        RECT 76.420 90.930 76.740 90.990 ;
        RECT 79.655 90.930 79.945 90.975 ;
        RECT 68.600 90.790 79.945 90.930 ;
        RECT 68.600 90.730 68.920 90.790 ;
        RECT 76.420 90.730 76.740 90.790 ;
        RECT 79.655 90.745 79.945 90.790 ;
        RECT 85.620 90.730 85.940 90.990 ;
        RECT 100.130 90.875 100.370 91.185 ;
        RECT 100.720 91.145 101.020 91.185 ;
        RECT 100.720 91.135 101.010 91.145 ;
        RECT 101.810 91.125 102.010 93.655 ;
        RECT 102.290 93.625 102.580 93.630 ;
        RECT 102.280 92.955 102.620 93.625 ;
        RECT 102.150 91.925 103.150 92.955 ;
        RECT 102.280 91.155 102.620 91.925 ;
        RECT 102.300 91.135 102.590 91.155 ;
        RECT 100.530 90.875 100.760 90.975 ;
        RECT 100.130 90.865 100.760 90.875 ;
        RECT 11.950 90.110 90.610 90.590 ;
        RECT 15.715 89.910 16.005 89.955 ;
        RECT 17.080 89.910 17.400 89.970 ;
        RECT 23.060 89.910 23.380 89.970 ;
        RECT 15.715 89.770 17.400 89.910 ;
        RECT 15.715 89.725 16.005 89.770 ;
        RECT 17.080 89.710 17.400 89.770 ;
        RECT 17.630 89.770 23.380 89.910 ;
        RECT 17.630 89.570 17.770 89.770 ;
        RECT 23.060 89.710 23.380 89.770 ;
        RECT 24.900 89.910 25.220 89.970 ;
        RECT 24.900 89.770 25.590 89.910 ;
        RECT 24.900 89.710 25.220 89.770 ;
        RECT 20.300 89.570 20.620 89.630 ;
        RECT 25.450 89.615 25.590 89.770 ;
        RECT 37.320 89.710 37.640 89.970 ;
        RECT 38.255 89.725 38.545 89.955 ;
        RECT 16.710 89.430 17.770 89.570 ;
        RECT 18.090 89.430 25.130 89.570 ;
        RECT 16.710 88.255 16.850 89.430 ;
        RECT 17.540 89.030 17.860 89.290 ;
        RECT 18.090 89.275 18.230 89.430 ;
        RECT 20.300 89.370 20.620 89.430 ;
        RECT 18.015 89.045 18.305 89.275 ;
        RECT 19.350 89.230 19.640 89.275 ;
        RECT 20.760 89.230 21.080 89.290 ;
        RECT 19.350 89.090 21.080 89.230 ;
        RECT 24.990 89.230 25.130 89.430 ;
        RECT 25.375 89.385 25.665 89.615 ;
        RECT 25.820 89.570 26.140 89.630 ;
        RECT 26.375 89.570 26.665 89.615 ;
        RECT 25.820 89.430 26.665 89.570 ;
        RECT 25.820 89.370 26.140 89.430 ;
        RECT 26.375 89.385 26.665 89.430 ;
        RECT 31.770 89.570 32.060 89.615 ;
        RECT 38.330 89.570 38.470 89.725 ;
        RECT 40.080 89.710 40.400 89.970 ;
        RECT 41.460 89.910 41.780 89.970 ;
        RECT 44.235 89.910 44.525 89.955 ;
        RECT 41.460 89.770 44.525 89.910 ;
        RECT 41.460 89.710 41.780 89.770 ;
        RECT 44.235 89.725 44.525 89.770 ;
        RECT 47.900 89.710 48.220 89.970 ;
        RECT 50.660 89.910 50.980 89.970 ;
        RECT 48.450 89.770 50.980 89.910 ;
        RECT 48.450 89.570 48.590 89.770 ;
        RECT 50.660 89.710 50.980 89.770 ;
        RECT 51.120 89.710 51.440 89.970 ;
        RECT 62.635 89.910 62.925 89.955 ;
        RECT 67.220 89.910 67.540 89.970 ;
        RECT 62.635 89.770 67.540 89.910 ;
        RECT 62.635 89.725 62.925 89.770 ;
        RECT 67.220 89.710 67.540 89.770 ;
        RECT 70.900 89.710 71.220 89.970 ;
        RECT 72.755 89.910 73.045 89.955 ;
        RECT 73.200 89.910 73.520 89.970 ;
        RECT 72.755 89.770 73.520 89.910 ;
        RECT 72.755 89.725 73.045 89.770 ;
        RECT 73.200 89.710 73.520 89.770 ;
        RECT 86.080 89.910 86.400 89.970 ;
        RECT 87.015 89.910 87.305 89.955 ;
        RECT 88.380 89.910 88.700 89.970 ;
        RECT 86.080 89.770 88.700 89.910 ;
        RECT 86.080 89.710 86.400 89.770 ;
        RECT 87.015 89.725 87.305 89.770 ;
        RECT 88.380 89.710 88.700 89.770 ;
        RECT 31.770 89.430 38.470 89.570 ;
        RECT 45.690 89.430 48.590 89.570 ;
        RECT 48.835 89.570 49.125 89.615 ;
        RECT 55.260 89.570 55.580 89.630 ;
        RECT 48.835 89.430 55.580 89.570 ;
        RECT 31.770 89.385 32.060 89.430 ;
        RECT 42.840 89.230 43.160 89.290 ;
        RECT 45.690 89.275 45.830 89.430 ;
        RECT 48.835 89.385 49.125 89.430 ;
        RECT 55.260 89.370 55.580 89.430 ;
        RECT 65.855 89.570 66.145 89.615 ;
        RECT 68.140 89.570 68.460 89.630 ;
        RECT 65.855 89.430 72.050 89.570 ;
        RECT 65.855 89.385 66.145 89.430 ;
        RECT 68.140 89.370 68.460 89.430 ;
        RECT 45.615 89.230 45.905 89.275 ;
        RECT 24.990 89.090 25.590 89.230 ;
        RECT 19.350 89.045 19.640 89.090 ;
        RECT 20.760 89.030 21.080 89.090 ;
        RECT 25.450 88.950 25.590 89.090 ;
        RECT 42.840 89.090 45.905 89.230 ;
        RECT 42.840 89.030 43.160 89.090 ;
        RECT 45.615 89.045 45.905 89.090 ;
        RECT 46.075 89.045 46.365 89.275 ;
        RECT 17.095 88.705 17.385 88.935 ;
        RECT 18.895 88.890 19.185 88.935 ;
        RECT 20.085 88.890 20.375 88.935 ;
        RECT 22.605 88.890 22.895 88.935 ;
        RECT 18.895 88.750 22.895 88.890 ;
        RECT 18.895 88.705 19.185 88.750 ;
        RECT 20.085 88.705 20.375 88.750 ;
        RECT 22.605 88.705 22.895 88.750 ;
        RECT 25.360 88.890 25.680 88.950 ;
        RECT 30.435 88.890 30.725 88.935 ;
        RECT 25.360 88.750 30.725 88.890 ;
        RECT 16.635 88.025 16.925 88.255 ;
        RECT 17.170 88.210 17.310 88.705 ;
        RECT 25.360 88.690 25.680 88.750 ;
        RECT 30.435 88.705 30.725 88.750 ;
        RECT 31.315 88.890 31.605 88.935 ;
        RECT 32.505 88.890 32.795 88.935 ;
        RECT 35.025 88.890 35.315 88.935 ;
        RECT 31.315 88.750 35.315 88.890 ;
        RECT 31.315 88.705 31.605 88.750 ;
        RECT 32.505 88.705 32.795 88.750 ;
        RECT 35.025 88.705 35.315 88.750 ;
        RECT 35.480 88.890 35.800 88.950 ;
        RECT 40.555 88.890 40.845 88.935 ;
        RECT 35.480 88.750 40.845 88.890 ;
        RECT 35.480 88.690 35.800 88.750 ;
        RECT 40.555 88.705 40.845 88.750 ;
        RECT 41.475 88.705 41.765 88.935 ;
        RECT 46.150 88.890 46.290 89.045 ;
        RECT 46.520 89.030 46.840 89.290 ;
        RECT 47.455 89.230 47.745 89.275 ;
        RECT 48.360 89.230 48.680 89.290 ;
        RECT 47.455 89.090 48.680 89.230 ;
        RECT 47.455 89.045 47.745 89.090 ;
        RECT 48.360 89.030 48.680 89.090 ;
        RECT 50.660 89.030 50.980 89.290 ;
        RECT 57.070 89.230 57.360 89.275 ;
        RECT 64.015 89.230 64.305 89.275 ;
        RECT 57.070 89.090 64.305 89.230 ;
        RECT 57.070 89.045 57.360 89.090 ;
        RECT 64.015 89.045 64.305 89.090 ;
        RECT 64.920 89.030 65.240 89.290 ;
        RECT 65.380 89.030 65.700 89.290 ;
        RECT 66.445 89.230 66.735 89.275 ;
        RECT 65.930 89.090 66.735 89.230 ;
        RECT 53.435 88.890 53.725 88.935 ;
        RECT 46.150 88.750 53.725 88.890 ;
        RECT 18.500 88.550 18.790 88.595 ;
        RECT 20.600 88.550 20.890 88.595 ;
        RECT 22.170 88.550 22.460 88.595 ;
        RECT 18.500 88.410 22.460 88.550 ;
        RECT 18.500 88.365 18.790 88.410 ;
        RECT 20.600 88.365 20.890 88.410 ;
        RECT 22.170 88.365 22.460 88.410 ;
        RECT 23.060 88.550 23.380 88.610 ;
        RECT 30.920 88.550 31.210 88.595 ;
        RECT 33.020 88.550 33.310 88.595 ;
        RECT 34.590 88.550 34.880 88.595 ;
        RECT 23.060 88.410 26.510 88.550 ;
        RECT 23.060 88.350 23.380 88.410 ;
        RECT 21.680 88.210 22.000 88.270 ;
        RECT 24.900 88.210 25.220 88.270 ;
        RECT 26.370 88.255 26.510 88.410 ;
        RECT 30.920 88.410 34.880 88.550 ;
        RECT 41.550 88.550 41.690 88.705 ;
        RECT 47.900 88.550 48.220 88.610 ;
        RECT 41.550 88.410 48.220 88.550 ;
        RECT 30.920 88.365 31.210 88.410 ;
        RECT 33.020 88.365 33.310 88.410 ;
        RECT 34.590 88.365 34.880 88.410 ;
        RECT 47.900 88.350 48.220 88.410 ;
        RECT 48.910 88.270 49.050 88.750 ;
        RECT 53.435 88.705 53.725 88.750 ;
        RECT 55.720 88.690 56.040 88.950 ;
        RECT 56.615 88.890 56.905 88.935 ;
        RECT 57.805 88.890 58.095 88.935 ;
        RECT 60.325 88.890 60.615 88.935 ;
        RECT 56.615 88.750 60.615 88.890 ;
        RECT 56.615 88.705 56.905 88.750 ;
        RECT 57.805 88.705 58.095 88.750 ;
        RECT 60.325 88.705 60.615 88.750 ;
        RECT 64.460 88.890 64.780 88.950 ;
        RECT 65.930 88.890 66.070 89.090 ;
        RECT 66.445 89.045 66.735 89.090 ;
        RECT 67.220 89.230 67.540 89.290 ;
        RECT 68.615 89.230 68.905 89.275 ;
        RECT 69.060 89.230 69.380 89.290 ;
        RECT 67.220 89.090 69.380 89.230 ;
        RECT 67.220 89.030 67.540 89.090 ;
        RECT 68.615 89.045 68.905 89.090 ;
        RECT 69.060 89.030 69.380 89.090 ;
        RECT 71.360 89.030 71.680 89.290 ;
        RECT 71.910 89.275 72.050 89.430 ;
        RECT 71.835 89.045 72.125 89.275 ;
        RECT 73.290 89.230 73.430 89.710 ;
        RECT 77.340 89.570 77.660 89.630 ;
        RECT 78.720 89.570 79.040 89.630 ;
        RECT 77.340 89.430 79.040 89.570 ;
        RECT 77.340 89.370 77.660 89.430 ;
        RECT 78.720 89.370 79.040 89.430 ;
        RECT 76.435 89.230 76.725 89.275 ;
        RECT 73.290 89.090 76.725 89.230 ;
        RECT 76.435 89.045 76.725 89.090 ;
        RECT 77.800 89.030 78.120 89.290 ;
        RECT 78.260 89.030 78.580 89.290 ;
        RECT 79.180 89.230 79.500 89.290 ;
        RECT 81.480 89.275 81.800 89.290 ;
        RECT 80.115 89.230 80.405 89.275 ;
        RECT 79.180 89.090 80.405 89.230 ;
        RECT 79.180 89.030 79.500 89.090 ;
        RECT 80.115 89.045 80.405 89.090 ;
        RECT 81.450 89.045 81.800 89.275 ;
        RECT 81.480 89.030 81.800 89.045 ;
        RECT 87.460 89.030 87.780 89.290 ;
        RECT 100.100 89.065 100.760 90.865 ;
        RECT 100.130 89.045 100.360 89.065 ;
        RECT 64.460 88.750 66.070 88.890 ;
        RECT 64.460 88.690 64.780 88.750 ;
        RECT 52.040 88.350 52.360 88.610 ;
        RECT 56.220 88.550 56.510 88.595 ;
        RECT 58.320 88.550 58.610 88.595 ;
        RECT 59.890 88.550 60.180 88.595 ;
        RECT 56.220 88.410 60.180 88.550 ;
        RECT 56.220 88.365 56.510 88.410 ;
        RECT 58.320 88.365 58.610 88.410 ;
        RECT 59.890 88.365 60.180 88.410 ;
        RECT 70.455 88.550 70.745 88.595 ;
        RECT 71.450 88.550 71.590 89.030 ;
        RECT 100.530 88.975 100.760 89.065 ;
        RECT 100.970 90.905 101.200 90.975 ;
        RECT 100.970 89.095 101.530 90.905 ;
        RECT 101.810 90.865 101.960 91.125 ;
        RECT 102.110 90.865 102.340 90.975 ;
        RECT 101.810 90.855 102.340 90.865 ;
        RECT 100.970 88.975 101.200 89.095 ;
        RECT 72.740 88.890 73.060 88.950 ;
        RECT 73.660 88.890 73.980 88.950 ;
        RECT 72.740 88.750 73.980 88.890 ;
        RECT 72.740 88.690 73.060 88.750 ;
        RECT 73.660 88.690 73.980 88.750 ;
        RECT 80.995 88.890 81.285 88.935 ;
        RECT 82.185 88.890 82.475 88.935 ;
        RECT 84.705 88.890 84.995 88.935 ;
        RECT 80.995 88.750 84.995 88.890 ;
        RECT 101.360 88.775 101.530 89.095 ;
        RECT 101.770 89.055 102.340 90.855 ;
        RECT 101.820 89.045 102.340 89.055 ;
        RECT 102.110 88.975 102.340 89.045 ;
        RECT 102.550 90.925 102.780 90.975 ;
        RECT 102.550 90.895 103.060 90.925 ;
        RECT 102.550 89.085 103.090 90.895 ;
        RECT 103.290 90.875 103.480 93.885 ;
        RECT 103.680 93.835 103.910 93.885 ;
        RECT 104.120 93.835 104.350 93.925 ;
        RECT 104.870 93.885 105.490 99.785 ;
        RECT 103.840 92.955 104.200 93.635 ;
        RECT 103.660 91.925 104.660 92.955 ;
        RECT 103.840 91.135 104.200 91.925 ;
        RECT 103.690 90.875 103.920 90.975 ;
        RECT 103.290 90.205 103.920 90.875 ;
        RECT 102.550 88.975 102.780 89.085 ;
        RECT 102.920 88.855 103.090 89.085 ;
        RECT 103.310 89.005 103.920 90.205 ;
        RECT 103.690 88.975 103.920 89.005 ;
        RECT 104.130 90.925 104.360 90.975 ;
        RECT 104.130 89.045 104.670 90.925 ;
        RECT 104.890 90.905 105.060 93.885 ;
        RECT 105.260 93.835 105.490 93.885 ;
        RECT 105.700 93.915 106.190 99.835 ;
        RECT 106.840 99.755 107.070 99.835 ;
        RECT 105.700 93.835 105.930 93.915 ;
        RECT 106.430 93.875 107.070 99.755 ;
        RECT 105.450 93.625 105.740 93.630 ;
        RECT 105.440 92.985 105.780 93.625 ;
        RECT 105.270 91.955 106.270 92.985 ;
        RECT 105.440 91.145 105.780 91.955 ;
        RECT 105.460 91.135 105.750 91.145 ;
        RECT 105.270 90.905 105.500 90.975 ;
        RECT 104.890 90.865 105.500 90.905 ;
        RECT 104.870 89.065 105.500 90.865 ;
        RECT 104.900 89.045 105.500 89.065 ;
        RECT 104.130 88.975 104.360 89.045 ;
        RECT 80.995 88.705 81.285 88.750 ;
        RECT 82.185 88.705 82.475 88.750 ;
        RECT 84.705 88.705 84.995 88.750 ;
        RECT 100.000 88.635 101.000 88.645 ;
        RECT 101.280 88.635 101.530 88.775 ;
        RECT 102.910 88.635 103.090 88.855 ;
        RECT 104.500 88.805 104.670 89.045 ;
        RECT 105.270 88.975 105.500 89.045 ;
        RECT 105.710 90.905 105.940 90.975 ;
        RECT 105.710 89.025 106.250 90.905 ;
        RECT 106.440 90.895 106.630 93.875 ;
        RECT 106.840 93.835 107.070 93.875 ;
        RECT 107.270 93.865 107.710 100.195 ;
        RECT 108.890 99.835 109.330 100.195 ;
        RECT 110.480 99.835 110.920 100.195 ;
        RECT 112.060 99.835 112.500 100.195 ;
        RECT 108.420 99.815 108.650 99.835 ;
        RECT 107.970 93.885 108.650 99.815 ;
        RECT 107.280 93.835 107.510 93.865 ;
        RECT 107.030 93.625 107.320 93.630 ;
        RECT 107.010 92.955 107.370 93.625 ;
        RECT 106.820 91.925 107.820 92.955 ;
        RECT 107.010 91.135 107.370 91.925 ;
        RECT 106.850 90.895 107.080 90.975 ;
        RECT 106.440 89.045 107.080 90.895 ;
        RECT 105.710 88.975 105.940 89.025 ;
        RECT 104.490 88.635 104.670 88.805 ;
        RECT 106.080 88.635 106.250 89.025 ;
        RECT 106.850 88.975 107.080 89.045 ;
        RECT 107.290 90.925 107.520 90.975 ;
        RECT 107.980 90.935 108.240 93.885 ;
        RECT 108.420 93.835 108.650 93.885 ;
        RECT 108.860 93.895 109.330 99.835 ;
        RECT 110.000 99.795 110.230 99.835 ;
        RECT 108.860 93.835 109.090 93.895 ;
        RECT 109.550 93.885 110.230 99.795 ;
        RECT 108.610 93.625 108.900 93.630 ;
        RECT 108.580 92.985 108.920 93.625 ;
        RECT 108.440 91.955 109.440 92.985 ;
        RECT 108.580 91.135 108.920 91.955 ;
        RECT 108.430 90.935 108.660 90.975 ;
        RECT 107.290 89.045 107.830 90.925 ;
        RECT 107.290 88.975 107.520 89.045 ;
        RECT 107.660 88.635 107.830 89.045 ;
        RECT 107.980 89.015 108.660 90.935 ;
        RECT 108.430 88.975 108.660 89.015 ;
        RECT 108.870 90.915 109.100 90.975 ;
        RECT 108.870 89.035 109.420 90.915 ;
        RECT 109.600 90.895 109.860 93.885 ;
        RECT 110.000 93.835 110.230 93.885 ;
        RECT 110.440 93.875 110.920 99.835 ;
        RECT 111.580 99.795 111.810 99.835 ;
        RECT 111.150 93.905 111.810 99.795 ;
        RECT 111.150 93.885 111.410 93.905 ;
        RECT 110.440 93.835 110.670 93.875 ;
        RECT 111.160 93.675 111.410 93.885 ;
        RECT 111.580 93.835 111.810 93.905 ;
        RECT 112.020 93.925 112.500 99.835 ;
        RECT 112.020 93.835 112.250 93.925 ;
        RECT 110.190 93.625 110.480 93.630 ;
        RECT 110.180 92.955 110.510 93.625 ;
        RECT 110.010 91.925 111.010 92.955 ;
        RECT 110.180 91.135 110.510 91.925 ;
        RECT 111.160 91.575 111.460 93.675 ;
        RECT 111.770 93.625 112.060 93.630 ;
        RECT 111.750 92.975 112.110 93.625 ;
        RECT 111.670 91.945 112.670 92.975 ;
        RECT 111.240 91.125 111.460 91.575 ;
        RECT 111.750 91.135 112.110 91.945 ;
        RECT 110.010 90.895 110.240 90.975 ;
        RECT 109.580 89.045 110.240 90.895 ;
        RECT 108.870 88.975 109.100 89.035 ;
        RECT 109.260 88.635 109.420 89.035 ;
        RECT 110.010 88.975 110.240 89.045 ;
        RECT 110.450 90.915 110.680 90.975 ;
        RECT 110.450 89.025 111.000 90.915 ;
        RECT 111.240 90.885 111.420 91.125 ;
        RECT 111.590 90.885 111.820 90.975 ;
        RECT 111.240 90.735 111.820 90.885 ;
        RECT 111.210 89.065 111.820 90.735 ;
        RECT 111.220 89.035 111.820 89.065 ;
        RECT 110.450 88.975 110.680 89.025 ;
        RECT 110.830 88.635 111.000 89.025 ;
        RECT 111.590 88.975 111.820 89.035 ;
        RECT 112.030 90.915 112.260 90.975 ;
        RECT 112.030 89.065 112.720 90.915 ;
        RECT 112.030 88.975 112.260 89.065 ;
        RECT 112.410 88.815 112.720 89.065 ;
        RECT 112.390 88.775 112.720 88.815 ;
        RECT 112.390 88.635 112.880 88.775 ;
        RECT 70.455 88.410 71.590 88.550 ;
        RECT 80.600 88.550 80.890 88.595 ;
        RECT 82.700 88.550 82.990 88.595 ;
        RECT 84.270 88.550 84.560 88.595 ;
        RECT 80.600 88.410 84.560 88.550 ;
        RECT 70.455 88.365 70.745 88.410 ;
        RECT 80.600 88.365 80.890 88.410 ;
        RECT 82.700 88.365 82.990 88.410 ;
        RECT 84.270 88.365 84.560 88.410 ;
        RECT 88.380 88.350 88.700 88.610 ;
        RECT 100.000 88.605 112.880 88.635 ;
        RECT 99.980 88.550 112.880 88.605 ;
        RECT 113.070 88.550 113.700 101.660 ;
        RECT 119.900 101.650 120.990 101.675 ;
        RECT 134.480 99.950 135.430 101.710 ;
        RECT 136.630 99.960 138.450 102.060 ;
        RECT 139.570 99.960 141.390 102.060 ;
        RECT 142.470 99.960 144.300 102.090 ;
        RECT 145.440 99.960 147.270 102.090 ;
        RECT 148.420 99.970 150.250 102.100 ;
        RECT 136.630 99.955 136.880 99.960 ;
        RECT 138.110 99.955 138.360 99.960 ;
        RECT 139.590 99.955 139.840 99.960 ;
        RECT 141.070 99.955 141.320 99.960 ;
        RECT 142.550 99.955 142.800 99.960 ;
        RECT 144.030 99.955 144.280 99.960 ;
        RECT 145.510 99.955 145.760 99.960 ;
        RECT 146.990 99.955 147.240 99.960 ;
        RECT 148.470 99.955 148.720 99.970 ;
        RECT 149.950 99.955 150.200 99.970 ;
        RECT 151.370 99.960 153.200 102.090 ;
        RECT 151.430 99.955 151.680 99.960 ;
        RECT 152.910 99.955 153.160 99.960 ;
        RECT 154.340 99.950 156.170 102.080 ;
        RECT 157.270 99.980 158.460 103.930 ;
        RECT 157.350 99.955 157.600 99.980 ;
        RECT 135.150 99.340 135.400 99.365 ;
        RECT 136.630 99.340 136.880 99.365 ;
        RECT 135.100 99.300 136.910 99.340 ;
        RECT 135.100 97.270 136.940 99.300 ;
        RECT 138.090 97.270 139.910 99.370 ;
        RECT 141.030 97.280 142.850 99.380 ;
        RECT 144.030 99.360 144.280 99.365 ;
        RECT 145.510 99.360 145.760 99.365 ;
        RECT 135.100 97.240 136.910 97.270 ;
        RECT 138.110 97.260 138.360 97.270 ;
        RECT 139.590 97.260 139.840 97.270 ;
        RECT 141.070 97.260 141.320 97.280 ;
        RECT 142.550 97.260 142.800 97.280 ;
        RECT 143.960 97.230 145.790 99.360 ;
        RECT 146.940 97.240 148.770 99.370 ;
        RECT 149.930 97.240 151.760 99.370 ;
        RECT 152.910 99.360 153.160 99.365 ;
        RECT 154.390 99.360 154.640 99.365 ;
        RECT 152.850 97.230 154.680 99.360 ;
        RECT 155.820 97.240 157.650 99.370 ;
        RECT 117.600 93.110 130.450 93.240 ;
        RECT 117.600 92.280 130.480 93.110 ;
        RECT 118.410 91.720 119.370 91.950 ;
        RECT 118.130 91.480 118.360 91.515 ;
        RECT 17.170 88.070 25.220 88.210 ;
        RECT 21.680 88.010 22.000 88.070 ;
        RECT 24.900 88.010 25.220 88.070 ;
        RECT 26.295 88.025 26.585 88.255 ;
        RECT 27.215 88.210 27.505 88.255 ;
        RECT 29.500 88.210 29.820 88.270 ;
        RECT 27.215 88.070 29.820 88.210 ;
        RECT 27.215 88.025 27.505 88.070 ;
        RECT 29.500 88.010 29.820 88.070 ;
        RECT 48.820 88.010 49.140 88.270 ;
        RECT 63.540 88.210 63.860 88.270 ;
        RECT 67.220 88.210 67.540 88.270 ;
        RECT 63.540 88.070 67.540 88.210 ;
        RECT 63.540 88.010 63.860 88.070 ;
        RECT 67.220 88.010 67.540 88.070 ;
        RECT 72.740 88.210 73.060 88.270 ;
        RECT 74.120 88.210 74.440 88.270 ;
        RECT 72.740 88.070 74.440 88.210 ;
        RECT 72.740 88.010 73.060 88.070 ;
        RECT 74.120 88.010 74.440 88.070 ;
        RECT 79.195 88.210 79.485 88.255 ;
        RECT 83.320 88.210 83.640 88.270 ;
        RECT 79.195 88.070 83.640 88.210 ;
        RECT 79.195 88.025 79.485 88.070 ;
        RECT 83.320 88.010 83.640 88.070 ;
        RECT 11.950 87.390 90.610 87.870 ;
        RECT 99.980 87.685 113.700 88.550 ;
        RECT 99.980 87.645 113.630 87.685 ;
        RECT 99.980 87.615 112.880 87.645 ;
        RECT 100.000 87.575 112.880 87.615 ;
        RECT 20.760 86.990 21.080 87.250 ;
        RECT 23.995 87.190 24.285 87.235 ;
        RECT 25.820 87.190 26.140 87.250 ;
        RECT 23.995 87.050 26.140 87.190 ;
        RECT 23.995 87.005 24.285 87.050 ;
        RECT 25.820 86.990 26.140 87.050 ;
        RECT 43.760 87.190 44.080 87.250 ;
        RECT 44.235 87.190 44.525 87.235 ;
        RECT 48.820 87.190 49.140 87.250 ;
        RECT 43.760 87.050 49.140 87.190 ;
        RECT 43.760 86.990 44.080 87.050 ;
        RECT 44.235 87.005 44.525 87.050 ;
        RECT 48.820 86.990 49.140 87.050 ;
        RECT 66.315 87.190 66.605 87.235 ;
        RECT 66.760 87.190 67.080 87.250 ;
        RECT 68.140 87.190 68.460 87.250 ;
        RECT 71.835 87.190 72.125 87.235 ;
        RECT 74.120 87.190 74.440 87.250 ;
        RECT 81.480 87.190 81.800 87.250 ;
        RECT 81.955 87.190 82.245 87.235 ;
        RECT 66.315 87.050 72.125 87.190 ;
        RECT 66.315 87.005 66.605 87.050 ;
        RECT 66.760 86.990 67.080 87.050 ;
        RECT 68.140 86.990 68.460 87.050 ;
        RECT 71.835 87.005 72.125 87.050 ;
        RECT 72.470 87.050 79.410 87.190 ;
        RECT 22.140 86.650 22.460 86.910 ;
        RECT 26.780 86.850 27.070 86.895 ;
        RECT 28.880 86.850 29.170 86.895 ;
        RECT 30.450 86.850 30.740 86.895 ;
        RECT 26.780 86.710 30.740 86.850 ;
        RECT 26.780 86.665 27.070 86.710 ;
        RECT 28.880 86.665 29.170 86.710 ;
        RECT 30.450 86.665 30.740 86.710 ;
        RECT 42.395 86.850 42.685 86.895 ;
        RECT 42.840 86.850 43.160 86.910 ;
        RECT 42.395 86.710 43.160 86.850 ;
        RECT 42.395 86.665 42.685 86.710 ;
        RECT 42.840 86.650 43.160 86.710 ;
        RECT 46.980 86.650 47.300 86.910 ;
        RECT 47.900 86.850 48.220 86.910 ;
        RECT 49.740 86.850 50.060 86.910 ;
        RECT 47.900 86.710 50.060 86.850 ;
        RECT 47.900 86.650 48.220 86.710 ;
        RECT 49.740 86.650 50.060 86.710 ;
        RECT 56.220 86.850 56.510 86.895 ;
        RECT 58.320 86.850 58.610 86.895 ;
        RECT 59.890 86.850 60.180 86.895 ;
        RECT 56.220 86.710 60.180 86.850 ;
        RECT 56.220 86.665 56.510 86.710 ;
        RECT 58.320 86.665 58.610 86.710 ;
        RECT 59.890 86.665 60.180 86.710 ;
        RECT 62.635 86.850 62.925 86.895 ;
        RECT 72.470 86.850 72.610 87.050 ;
        RECT 74.120 86.990 74.440 87.050 ;
        RECT 76.420 86.850 76.740 86.910 ;
        RECT 62.635 86.710 64.690 86.850 ;
        RECT 62.635 86.665 62.925 86.710 ;
        RECT 20.315 86.510 20.605 86.555 ;
        RECT 22.230 86.510 22.370 86.650 ;
        RECT 23.980 86.510 24.300 86.570 ;
        RECT 20.315 86.370 21.910 86.510 ;
        RECT 22.230 86.370 24.300 86.510 ;
        RECT 20.315 86.325 20.605 86.370 ;
        RECT 21.770 86.215 21.910 86.370 ;
        RECT 21.695 85.985 21.985 86.215 ;
        RECT 22.140 85.970 22.460 86.230 ;
        RECT 23.610 86.215 23.750 86.370 ;
        RECT 23.980 86.310 24.300 86.370 ;
        RECT 25.360 86.510 25.680 86.570 ;
        RECT 26.295 86.510 26.585 86.555 ;
        RECT 25.360 86.370 26.585 86.510 ;
        RECT 25.360 86.310 25.680 86.370 ;
        RECT 26.295 86.325 26.585 86.370 ;
        RECT 27.175 86.510 27.465 86.555 ;
        RECT 28.365 86.510 28.655 86.555 ;
        RECT 30.885 86.510 31.175 86.555 ;
        RECT 27.175 86.370 31.175 86.510 ;
        RECT 27.175 86.325 27.465 86.370 ;
        RECT 28.365 86.325 28.655 86.370 ;
        RECT 30.885 86.325 31.175 86.370 ;
        RECT 54.340 86.310 54.660 86.570 ;
        RECT 55.720 86.310 56.040 86.570 ;
        RECT 56.615 86.510 56.905 86.555 ;
        RECT 57.805 86.510 58.095 86.555 ;
        RECT 60.325 86.510 60.615 86.555 ;
        RECT 63.095 86.510 63.385 86.555 ;
        RECT 56.615 86.370 60.615 86.510 ;
        RECT 56.615 86.325 56.905 86.370 ;
        RECT 57.805 86.325 58.095 86.370 ;
        RECT 60.325 86.325 60.615 86.370 ;
        RECT 60.870 86.370 63.385 86.510 ;
        RECT 23.535 85.985 23.825 86.215 ;
        RECT 41.935 85.985 42.225 86.215 ;
        RECT 57.070 86.170 57.360 86.215 ;
        RECT 60.870 86.170 61.010 86.370 ;
        RECT 63.095 86.325 63.385 86.370 ;
        RECT 57.070 86.030 61.010 86.170 ;
        RECT 57.070 85.985 57.360 86.030 ;
        RECT 18.475 85.830 18.765 85.875 ;
        RECT 19.395 85.830 19.685 85.875 ;
        RECT 20.760 85.830 21.080 85.890 ;
        RECT 18.475 85.690 19.150 85.830 ;
        RECT 18.475 85.645 18.765 85.690 ;
        RECT 19.010 85.550 19.150 85.690 ;
        RECT 19.395 85.690 21.080 85.830 ;
        RECT 19.395 85.645 19.685 85.690 ;
        RECT 20.760 85.630 21.080 85.690 ;
        RECT 26.740 85.830 27.060 85.890 ;
        RECT 27.520 85.830 27.810 85.875 ;
        RECT 26.740 85.690 27.810 85.830 ;
        RECT 42.010 85.830 42.150 85.985 ;
        RECT 64.000 85.970 64.320 86.230 ;
        RECT 64.550 86.215 64.690 86.710 ;
        RECT 71.910 86.710 72.610 86.850 ;
        RECT 72.830 86.710 76.740 86.850 ;
        RECT 71.910 86.570 72.050 86.710 ;
        RECT 68.230 86.370 69.290 86.510 ;
        RECT 64.475 86.170 64.765 86.215 ;
        RECT 64.920 86.170 65.240 86.230 ;
        RECT 64.475 86.030 65.240 86.170 ;
        RECT 64.475 85.985 64.765 86.030 ;
        RECT 64.920 85.970 65.240 86.030 ;
        RECT 65.395 85.985 65.685 86.215 ;
        RECT 65.855 86.170 66.145 86.215 ;
        RECT 66.300 86.170 66.620 86.230 ;
        RECT 65.855 86.030 66.620 86.170 ;
        RECT 65.855 85.985 66.145 86.030 ;
        RECT 44.220 85.830 44.540 85.890 ;
        RECT 42.010 85.690 44.540 85.830 ;
        RECT 26.740 85.630 27.060 85.690 ;
        RECT 27.520 85.645 27.810 85.690 ;
        RECT 44.220 85.630 44.540 85.690 ;
        RECT 48.820 85.830 49.140 85.890 ;
        RECT 51.580 85.830 51.900 85.890 ;
        RECT 48.820 85.690 51.900 85.830 ;
        RECT 48.820 85.630 49.140 85.690 ;
        RECT 51.580 85.630 51.900 85.690 ;
        RECT 18.920 85.490 19.240 85.550 ;
        RECT 21.220 85.490 21.540 85.550 ;
        RECT 18.920 85.350 21.540 85.490 ;
        RECT 18.920 85.290 19.240 85.350 ;
        RECT 21.220 85.290 21.540 85.350 ;
        RECT 33.180 85.290 33.500 85.550 ;
        RECT 38.700 85.290 39.020 85.550 ;
        RECT 45.140 85.290 45.460 85.550 ;
        RECT 46.535 85.490 46.825 85.535 ;
        RECT 47.900 85.490 48.220 85.550 ;
        RECT 46.535 85.350 48.220 85.490 ;
        RECT 46.535 85.305 46.825 85.350 ;
        RECT 47.900 85.290 48.220 85.350 ;
        RECT 51.120 85.290 51.440 85.550 ;
        RECT 52.960 85.290 53.280 85.550 ;
        RECT 53.435 85.490 53.725 85.535 ;
        RECT 56.180 85.490 56.500 85.550 ;
        RECT 53.435 85.350 56.500 85.490 ;
        RECT 53.435 85.305 53.725 85.350 ;
        RECT 56.180 85.290 56.500 85.350 ;
        RECT 64.460 85.490 64.780 85.550 ;
        RECT 65.470 85.490 65.610 85.985 ;
        RECT 66.300 85.970 66.620 86.030 ;
        RECT 67.220 85.970 67.540 86.230 ;
        RECT 68.230 86.215 68.370 86.370 ;
        RECT 69.150 86.230 69.290 86.370 ;
        RECT 71.820 86.310 72.140 86.570 ;
        RECT 72.830 86.555 72.970 86.710 ;
        RECT 76.420 86.650 76.740 86.710 ;
        RECT 72.755 86.325 73.045 86.555 ;
        RECT 75.500 86.510 75.820 86.570 ;
        RECT 75.975 86.510 76.265 86.555 ;
        RECT 78.735 86.510 79.025 86.555 ;
        RECT 75.500 86.370 79.025 86.510 ;
        RECT 75.500 86.310 75.820 86.370 ;
        RECT 75.975 86.325 76.265 86.370 ;
        RECT 78.735 86.325 79.025 86.370 ;
        RECT 68.155 85.985 68.445 86.215 ;
        RECT 68.615 85.985 68.905 86.215 ;
        RECT 69.060 86.170 69.380 86.230 ;
        RECT 69.535 86.170 69.825 86.215 ;
        RECT 69.060 86.030 69.825 86.170 ;
        RECT 64.460 85.350 65.610 85.490 ;
        RECT 67.310 85.490 67.450 85.970 ;
        RECT 68.690 85.490 68.830 85.985 ;
        RECT 69.060 85.970 69.380 86.030 ;
        RECT 69.535 85.985 69.825 86.030 ;
        RECT 71.360 85.970 71.680 86.230 ;
        RECT 73.200 86.170 73.520 86.230 ;
        RECT 74.135 86.170 74.425 86.215 ;
        RECT 73.200 86.030 74.425 86.170 ;
        RECT 73.200 85.970 73.520 86.030 ;
        RECT 74.135 85.985 74.425 86.030 ;
        RECT 76.895 85.985 77.185 86.215 ;
        RECT 77.815 85.985 78.105 86.215 ;
        RECT 78.275 86.170 78.565 86.215 ;
        RECT 79.270 86.170 79.410 87.050 ;
        RECT 81.480 87.050 82.245 87.190 ;
        RECT 81.480 86.990 81.800 87.050 ;
        RECT 81.955 87.005 82.245 87.050 ;
        RECT 87.015 87.190 87.305 87.235 ;
        RECT 87.460 87.190 87.780 87.250 ;
        RECT 87.015 87.050 87.780 87.190 ;
        RECT 87.015 87.005 87.305 87.050 ;
        RECT 87.460 86.990 87.780 87.050 ;
        RECT 80.575 86.510 80.865 86.555 ;
        RECT 84.715 86.510 85.005 86.555 ;
        RECT 80.575 86.370 85.005 86.510 ;
        RECT 80.575 86.325 80.865 86.370 ;
        RECT 84.715 86.325 85.005 86.370 ;
        RECT 78.275 86.030 79.410 86.170 ;
        RECT 79.655 86.170 79.945 86.215 ;
        RECT 80.100 86.170 80.420 86.230 ;
        RECT 79.655 86.030 80.420 86.170 ;
        RECT 78.275 85.985 78.565 86.030 ;
        RECT 79.655 85.985 79.945 86.030 ;
        RECT 75.040 85.630 75.360 85.890 ;
        RECT 75.960 85.830 76.280 85.890 ;
        RECT 76.970 85.830 77.110 85.985 ;
        RECT 75.960 85.690 77.110 85.830 ;
        RECT 75.960 85.630 76.280 85.690 ;
        RECT 67.310 85.350 68.830 85.490 ;
        RECT 64.460 85.290 64.780 85.350 ;
        RECT 69.060 85.290 69.380 85.550 ;
        RECT 72.755 85.490 73.045 85.535 ;
        RECT 74.580 85.490 74.900 85.550 ;
        RECT 77.890 85.490 78.030 85.985 ;
        RECT 80.100 85.970 80.420 86.030 ;
        RECT 83.795 86.170 84.085 86.215 ;
        RECT 85.620 86.170 85.940 86.230 ;
        RECT 83.795 86.030 85.940 86.170 ;
        RECT 83.795 85.985 84.085 86.030 ;
        RECT 85.620 85.970 85.940 86.030 ;
        RECT 86.080 85.970 86.400 86.230 ;
        RECT 83.320 85.830 83.640 85.890 ;
        RECT 84.255 85.830 84.545 85.875 ;
        RECT 83.320 85.690 84.545 85.830 ;
        RECT 83.320 85.630 83.640 85.690 ;
        RECT 84.255 85.645 84.545 85.690 ;
        RECT 72.755 85.350 78.030 85.490 ;
        RECT 72.755 85.305 73.045 85.350 ;
        RECT 74.580 85.290 74.900 85.350 ;
        RECT 11.950 84.670 90.610 85.150 ;
        RECT 100.540 84.895 101.150 87.235 ;
        RECT 101.980 87.045 102.640 87.365 ;
        RECT 102.030 84.925 102.640 87.045 ;
        RECT 102.480 84.895 102.640 84.925 ;
        RECT 103.500 84.885 104.050 87.235 ;
        RECT 105.010 84.865 105.560 87.215 ;
        RECT 106.470 84.895 107.020 87.245 ;
        RECT 107.950 84.925 108.500 87.275 ;
        RECT 109.400 84.915 109.950 87.265 ;
        RECT 110.900 84.925 111.450 87.275 ;
        RECT 112.320 87.135 112.880 87.575 ;
        RECT 112.320 84.975 112.890 87.135 ;
        RECT 112.320 84.965 112.880 84.975 ;
        RECT 26.740 84.270 27.060 84.530 ;
        RECT 44.220 84.470 44.540 84.530 ;
        RECT 45.155 84.470 45.445 84.515 ;
        RECT 44.220 84.330 45.445 84.470 ;
        RECT 44.220 84.270 44.540 84.330 ;
        RECT 45.155 84.285 45.445 84.330 ;
        RECT 45.615 84.470 45.905 84.515 ;
        RECT 46.520 84.470 46.840 84.530 ;
        RECT 45.615 84.330 46.840 84.470 ;
        RECT 45.615 84.285 45.905 84.330 ;
        RECT 46.520 84.270 46.840 84.330 ;
        RECT 55.260 84.470 55.580 84.530 ;
        RECT 55.735 84.470 56.025 84.515 ;
        RECT 55.260 84.330 56.025 84.470 ;
        RECT 55.260 84.270 55.580 84.330 ;
        RECT 55.735 84.285 56.025 84.330 ;
        RECT 26.280 84.130 26.600 84.190 ;
        RECT 29.055 84.130 29.345 84.175 ;
        RECT 41.000 84.130 41.320 84.190 ;
        RECT 47.440 84.130 47.760 84.190 ;
        RECT 26.280 83.990 29.345 84.130 ;
        RECT 26.280 83.930 26.600 83.990 ;
        RECT 29.055 83.945 29.345 83.990 ;
        RECT 38.330 83.990 47.760 84.130 ;
        RECT 28.595 83.790 28.885 83.835 ;
        RECT 29.960 83.790 30.280 83.850 ;
        RECT 33.180 83.790 33.500 83.850 ;
        RECT 38.330 83.835 38.470 83.990 ;
        RECT 41.000 83.930 41.320 83.990 ;
        RECT 47.440 83.930 47.760 83.990 ;
        RECT 47.900 83.930 48.220 84.190 ;
        RECT 50.170 84.130 50.460 84.175 ;
        RECT 51.120 84.130 51.440 84.190 ;
        RECT 50.170 83.990 51.440 84.130 ;
        RECT 50.170 83.945 50.460 83.990 ;
        RECT 51.120 83.930 51.440 83.990 ;
        RECT 39.620 83.835 39.940 83.850 ;
        RECT 28.595 83.650 33.500 83.790 ;
        RECT 28.595 83.605 28.885 83.650 ;
        RECT 29.960 83.590 30.280 83.650 ;
        RECT 33.180 83.590 33.500 83.650 ;
        RECT 38.255 83.605 38.545 83.835 ;
        RECT 39.590 83.605 39.940 83.835 ;
        RECT 39.620 83.590 39.940 83.605 ;
        RECT 45.600 83.790 45.920 83.850 ;
        RECT 46.535 83.790 46.825 83.835 ;
        RECT 45.600 83.650 46.825 83.790 ;
        RECT 55.810 83.790 55.950 84.285 ;
        RECT 56.180 84.270 56.500 84.530 ;
        RECT 65.380 84.470 65.700 84.530 ;
        RECT 66.775 84.470 67.065 84.515 ;
        RECT 67.680 84.470 68.000 84.530 ;
        RECT 69.060 84.470 69.380 84.530 ;
        RECT 65.380 84.330 69.380 84.470 ;
        RECT 65.380 84.270 65.700 84.330 ;
        RECT 66.775 84.285 67.065 84.330 ;
        RECT 67.680 84.270 68.000 84.330 ;
        RECT 69.060 84.270 69.380 84.330 ;
        RECT 69.980 84.470 70.300 84.530 ;
        RECT 72.740 84.470 73.060 84.530 ;
        RECT 74.465 84.470 74.755 84.515 ;
        RECT 69.980 84.330 74.755 84.470 ;
        RECT 118.030 84.370 118.360 91.480 ;
        RECT 69.980 84.270 70.300 84.330 ;
        RECT 72.740 84.270 73.060 84.330 ;
        RECT 74.465 84.285 74.755 84.330 ;
        RECT 70.455 84.130 70.745 84.175 ;
        RECT 71.360 84.130 71.680 84.190 ;
        RECT 65.055 83.990 71.680 84.130 ;
        RECT 65.055 83.850 65.195 83.990 ;
        RECT 70.455 83.945 70.745 83.990 ;
        RECT 71.360 83.930 71.680 83.990 ;
        RECT 75.500 83.930 75.820 84.190 ;
        RECT 58.955 83.790 59.245 83.835 ;
        RECT 55.810 83.650 59.245 83.790 ;
        RECT 45.600 83.590 45.920 83.650 ;
        RECT 46.535 83.605 46.825 83.650 ;
        RECT 58.955 83.605 59.245 83.650 ;
        RECT 64.920 83.590 65.240 83.850 ;
        RECT 77.800 83.790 78.120 83.850 ;
        RECT 65.470 83.650 78.120 83.790 ;
        RECT 29.500 83.250 29.820 83.510 ;
        RECT 39.135 83.450 39.425 83.495 ;
        RECT 40.325 83.450 40.615 83.495 ;
        RECT 42.845 83.450 43.135 83.495 ;
        RECT 39.135 83.310 43.135 83.450 ;
        RECT 39.135 83.265 39.425 83.310 ;
        RECT 40.325 83.265 40.615 83.310 ;
        RECT 42.845 83.265 43.135 83.310 ;
        RECT 45.140 83.450 45.460 83.510 ;
        RECT 46.995 83.450 47.285 83.495 ;
        RECT 45.140 83.310 47.285 83.450 ;
        RECT 45.140 83.250 45.460 83.310 ;
        RECT 46.995 83.265 47.285 83.310 ;
        RECT 47.440 83.450 47.760 83.510 ;
        RECT 48.835 83.450 49.125 83.495 ;
        RECT 47.440 83.310 49.125 83.450 ;
        RECT 47.440 83.250 47.760 83.310 ;
        RECT 48.835 83.265 49.125 83.310 ;
        RECT 49.715 83.450 50.005 83.495 ;
        RECT 50.905 83.450 51.195 83.495 ;
        RECT 53.425 83.450 53.715 83.495 ;
        RECT 49.715 83.310 53.715 83.450 ;
        RECT 49.715 83.265 50.005 83.310 ;
        RECT 50.905 83.265 51.195 83.310 ;
        RECT 53.425 83.265 53.715 83.310 ;
        RECT 38.740 83.110 39.030 83.155 ;
        RECT 40.840 83.110 41.130 83.155 ;
        RECT 42.410 83.110 42.700 83.155 ;
        RECT 49.320 83.110 49.610 83.155 ;
        RECT 51.420 83.110 51.710 83.155 ;
        RECT 52.990 83.110 53.280 83.155 ;
        RECT 38.740 82.970 42.700 83.110 ;
        RECT 38.740 82.925 39.030 82.970 ;
        RECT 40.840 82.925 41.130 82.970 ;
        RECT 42.410 82.925 42.700 82.970 ;
        RECT 42.930 82.970 48.545 83.110 ;
        RECT 33.180 82.770 33.500 82.830 ;
        RECT 42.930 82.770 43.070 82.970 ;
        RECT 33.180 82.630 43.070 82.770 ;
        RECT 33.180 82.570 33.500 82.630 ;
        RECT 47.900 82.570 48.220 82.830 ;
        RECT 48.405 82.770 48.545 82.970 ;
        RECT 49.320 82.970 53.280 83.110 ;
        RECT 49.320 82.925 49.610 82.970 ;
        RECT 51.420 82.925 51.710 82.970 ;
        RECT 52.990 82.925 53.280 82.970 ;
        RECT 65.470 82.770 65.610 83.650 ;
        RECT 77.800 83.590 78.120 83.650 ;
        RECT 84.255 83.790 84.545 83.835 ;
        RECT 87.000 83.790 87.320 83.850 ;
        RECT 88.395 83.790 88.685 83.835 ;
        RECT 84.255 83.650 88.685 83.790 ;
        RECT 84.255 83.605 84.545 83.650 ;
        RECT 87.000 83.590 87.320 83.650 ;
        RECT 88.395 83.605 88.685 83.650 ;
        RECT 99.980 83.715 100.370 83.725 ;
        RECT 70.900 83.450 71.220 83.510 ;
        RECT 67.770 83.310 71.220 83.450 ;
        RECT 67.770 83.155 67.910 83.310 ;
        RECT 70.900 83.250 71.220 83.310 ;
        RECT 67.695 82.925 67.985 83.155 ;
        RECT 68.600 82.910 68.920 83.170 ;
        RECT 73.200 83.110 73.520 83.170 ;
        RECT 71.070 82.970 73.520 83.110 ;
        RECT 48.405 82.630 65.610 82.770 ;
        RECT 66.760 82.570 67.080 82.830 ;
        RECT 68.155 82.770 68.445 82.815 ;
        RECT 71.070 82.770 71.210 82.970 ;
        RECT 73.200 82.910 73.520 82.970 ;
        RECT 68.155 82.630 71.210 82.770 ;
        RECT 71.360 82.770 71.680 82.830 ;
        RECT 73.675 82.770 73.965 82.815 ;
        RECT 71.360 82.630 73.965 82.770 ;
        RECT 68.155 82.585 68.445 82.630 ;
        RECT 71.360 82.570 71.680 82.630 ;
        RECT 73.675 82.585 73.965 82.630 ;
        RECT 74.580 82.570 74.900 82.830 ;
        RECT 85.160 82.570 85.480 82.830 ;
        RECT 85.620 82.570 85.940 82.830 ;
        RECT 11.950 81.950 90.610 82.430 ;
        RECT 21.220 81.750 21.540 81.810 ;
        RECT 22.155 81.750 22.445 81.795 ;
        RECT 23.060 81.750 23.380 81.810 ;
        RECT 17.630 81.610 23.380 81.750 ;
        RECT 17.630 81.115 17.770 81.610 ;
        RECT 21.220 81.550 21.540 81.610 ;
        RECT 22.155 81.565 22.445 81.610 ;
        RECT 23.060 81.550 23.380 81.610 ;
        RECT 39.620 81.750 39.940 81.810 ;
        RECT 41.015 81.750 41.305 81.795 ;
        RECT 39.620 81.610 41.305 81.750 ;
        RECT 39.620 81.550 39.940 81.610 ;
        RECT 41.015 81.565 41.305 81.610 ;
        RECT 47.900 81.750 48.220 81.810 ;
        RECT 51.135 81.750 51.425 81.795 ;
        RECT 47.900 81.610 51.425 81.750 ;
        RECT 47.900 81.550 48.220 81.610 ;
        RECT 51.135 81.565 51.425 81.610 ;
        RECT 51.580 81.750 51.900 81.810 ;
        RECT 52.055 81.750 52.345 81.795 ;
        RECT 51.580 81.610 52.345 81.750 ;
        RECT 51.580 81.550 51.900 81.610 ;
        RECT 52.055 81.565 52.345 81.610 ;
        RECT 52.960 81.750 53.280 81.810 ;
        RECT 53.435 81.750 53.725 81.795 ;
        RECT 52.960 81.610 53.725 81.750 ;
        RECT 52.960 81.550 53.280 81.610 ;
        RECT 53.435 81.565 53.725 81.610 ;
        RECT 66.760 81.750 67.080 81.810 ;
        RECT 67.695 81.750 67.985 81.795 ;
        RECT 66.760 81.610 67.985 81.750 ;
        RECT 66.760 81.550 67.080 81.610 ;
        RECT 67.695 81.565 67.985 81.610 ;
        RECT 75.975 81.750 76.265 81.795 ;
        RECT 84.700 81.750 85.020 81.810 ;
        RECT 75.975 81.610 85.020 81.750 ;
        RECT 75.975 81.565 76.265 81.610 ;
        RECT 84.700 81.550 85.020 81.610 ;
        RECT 87.000 81.550 87.320 81.810 ;
        RECT 88.380 81.550 88.700 81.810 ;
        RECT 99.980 81.555 101.000 83.715 ;
        RECT 20.760 81.410 21.080 81.470 ;
        RECT 24.455 81.410 24.745 81.455 ;
        RECT 34.100 81.410 34.420 81.470 ;
        RECT 72.280 81.410 72.600 81.470 ;
        RECT 75.500 81.410 75.820 81.470 ;
        RECT 18.090 81.270 23.290 81.410 ;
        RECT 17.555 80.885 17.845 81.115 ;
        RECT 18.090 80.775 18.230 81.270 ;
        RECT 20.760 81.210 21.080 81.270 ;
        RECT 18.475 81.070 18.765 81.115 ;
        RECT 22.140 81.070 22.460 81.130 ;
        RECT 18.475 80.930 22.460 81.070 ;
        RECT 18.475 80.885 18.765 80.930 ;
        RECT 16.635 80.545 16.925 80.775 ;
        RECT 18.015 80.545 18.305 80.775 ;
        RECT 16.710 80.390 16.850 80.545 ;
        RECT 18.920 80.530 19.240 80.790 ;
        RECT 19.470 80.775 19.610 80.930 ;
        RECT 22.140 80.870 22.460 80.930 ;
        RECT 19.395 80.545 19.685 80.775 ;
        RECT 20.315 80.730 20.605 80.775 ;
        RECT 21.220 80.730 21.540 80.790 ;
        RECT 23.150 80.775 23.290 81.270 ;
        RECT 24.455 81.270 29.730 81.410 ;
        RECT 24.455 81.225 24.745 81.270 ;
        RECT 29.590 81.115 29.730 81.270 ;
        RECT 34.100 81.270 68.600 81.410 ;
        RECT 34.100 81.210 34.420 81.270 ;
        RECT 29.515 80.885 29.805 81.115 ;
        RECT 36.860 81.070 37.180 81.130 ;
        RECT 37.795 81.070 38.085 81.115 ;
        RECT 36.860 80.930 38.085 81.070 ;
        RECT 36.860 80.870 37.180 80.930 ;
        RECT 37.795 80.885 38.085 80.930 ;
        RECT 20.315 80.590 21.540 80.730 ;
        RECT 20.315 80.545 20.605 80.590 ;
        RECT 19.470 80.390 19.610 80.545 ;
        RECT 21.220 80.530 21.540 80.590 ;
        RECT 21.695 80.545 21.985 80.775 ;
        RECT 23.075 80.545 23.365 80.775 ;
        RECT 26.280 80.730 26.600 80.790 ;
        RECT 28.595 80.730 28.885 80.775 ;
        RECT 26.280 80.590 28.885 80.730 ;
        RECT 37.870 80.730 38.010 80.885 ;
        RECT 38.700 80.870 39.020 81.130 ;
        RECT 44.680 81.070 45.000 81.130 ;
        RECT 46.075 81.070 46.365 81.115 ;
        RECT 44.680 80.930 46.365 81.070 ;
        RECT 44.680 80.870 45.000 80.930 ;
        RECT 46.075 80.885 46.365 80.930 ;
        RECT 46.980 80.870 47.300 81.130 ;
        RECT 56.195 81.070 56.485 81.115 ;
        RECT 57.100 81.070 57.420 81.130 ;
        RECT 56.195 80.930 57.420 81.070 ;
        RECT 68.460 81.070 68.600 81.270 ;
        RECT 72.280 81.270 75.820 81.410 ;
        RECT 72.280 81.210 72.600 81.270 ;
        RECT 75.500 81.210 75.820 81.270 ;
        RECT 80.600 81.410 80.890 81.455 ;
        RECT 82.700 81.410 82.990 81.455 ;
        RECT 84.270 81.410 84.560 81.455 ;
        RECT 80.600 81.270 84.560 81.410 ;
        RECT 80.600 81.225 80.890 81.270 ;
        RECT 82.700 81.225 82.990 81.270 ;
        RECT 84.270 81.225 84.560 81.270 ;
        RECT 79.180 81.070 79.500 81.130 ;
        RECT 80.115 81.070 80.405 81.115 ;
        RECT 68.460 80.930 78.490 81.070 ;
        RECT 56.195 80.885 56.485 80.930 ;
        RECT 57.100 80.870 57.420 80.930 ;
        RECT 40.540 80.730 40.860 80.790 ;
        RECT 37.870 80.590 40.860 80.730 ;
        RECT 16.710 80.250 19.610 80.390 ;
        RECT 19.840 80.190 20.160 80.450 ;
        RECT 15.715 80.050 16.005 80.095 ;
        RECT 17.080 80.050 17.400 80.110 ;
        RECT 15.715 79.910 17.400 80.050 ;
        RECT 15.715 79.865 16.005 79.910 ;
        RECT 17.080 79.850 17.400 79.910 ;
        RECT 19.380 80.050 19.700 80.110 ;
        RECT 21.770 80.050 21.910 80.545 ;
        RECT 22.140 80.390 22.460 80.450 ;
        RECT 23.150 80.390 23.290 80.545 ;
        RECT 26.280 80.530 26.600 80.590 ;
        RECT 28.595 80.545 28.885 80.590 ;
        RECT 40.540 80.530 40.860 80.590 ;
        RECT 55.735 80.730 56.025 80.775 ;
        RECT 56.640 80.730 56.960 80.790 ;
        RECT 63.095 80.730 63.385 80.775 ;
        RECT 55.735 80.590 63.385 80.730 ;
        RECT 55.735 80.545 56.025 80.590 ;
        RECT 56.640 80.530 56.960 80.590 ;
        RECT 63.095 80.545 63.385 80.590 ;
        RECT 66.315 80.730 66.605 80.775 ;
        RECT 69.520 80.730 69.840 80.790 ;
        RECT 66.315 80.590 69.840 80.730 ;
        RECT 66.315 80.545 66.605 80.590 ;
        RECT 69.520 80.530 69.840 80.590 ;
        RECT 72.280 80.530 72.600 80.790 ;
        RECT 73.215 80.545 73.505 80.775 ;
        RECT 73.675 80.545 73.965 80.775 ;
        RECT 22.140 80.250 23.290 80.390 ;
        RECT 50.660 80.390 50.980 80.450 ;
        RECT 52.975 80.390 53.265 80.435 ;
        RECT 50.660 80.250 53.265 80.390 ;
        RECT 22.140 80.190 22.460 80.250 ;
        RECT 50.660 80.190 50.980 80.250 ;
        RECT 52.975 80.205 53.265 80.250 ;
        RECT 64.920 80.390 65.240 80.450 ;
        RECT 67.680 80.435 68.000 80.450 ;
        RECT 66.775 80.390 67.065 80.435 ;
        RECT 64.920 80.250 67.065 80.390 ;
        RECT 64.920 80.190 65.240 80.250 ;
        RECT 66.775 80.205 67.065 80.250 ;
        RECT 67.680 80.205 68.065 80.435 ;
        RECT 67.680 80.190 68.000 80.205 ;
        RECT 19.380 79.910 21.910 80.050 ;
        RECT 26.755 80.050 27.045 80.095 ;
        RECT 27.660 80.050 27.980 80.110 ;
        RECT 26.755 79.910 27.980 80.050 ;
        RECT 19.380 79.850 19.700 79.910 ;
        RECT 26.755 79.865 27.045 79.910 ;
        RECT 27.660 79.850 27.980 79.910 ;
        RECT 29.055 80.050 29.345 80.095 ;
        RECT 34.100 80.050 34.420 80.110 ;
        RECT 29.055 79.910 34.420 80.050 ;
        RECT 29.055 79.865 29.345 79.910 ;
        RECT 34.100 79.850 34.420 79.910 ;
        RECT 39.175 80.050 39.465 80.095 ;
        RECT 41.460 80.050 41.780 80.110 ;
        RECT 39.175 79.910 41.780 80.050 ;
        RECT 39.175 79.865 39.465 79.910 ;
        RECT 41.460 79.850 41.780 79.910 ;
        RECT 43.300 79.850 43.620 80.110 ;
        RECT 50.200 79.850 50.520 80.110 ;
        RECT 51.975 80.050 52.265 80.095 ;
        RECT 53.880 80.050 54.200 80.110 ;
        RECT 51.975 79.910 54.200 80.050 ;
        RECT 51.975 79.865 52.265 79.910 ;
        RECT 53.880 79.850 54.200 79.910 ;
        RECT 55.275 80.050 55.565 80.095 ;
        RECT 58.020 80.050 58.340 80.110 ;
        RECT 55.275 79.910 58.340 80.050 ;
        RECT 55.275 79.865 55.565 79.910 ;
        RECT 58.020 79.850 58.340 79.910 ;
        RECT 68.600 80.050 68.920 80.110 ;
        RECT 73.290 80.050 73.430 80.545 ;
        RECT 73.750 80.390 73.890 80.545 ;
        RECT 74.120 80.530 74.440 80.790 ;
        RECT 74.580 80.730 74.900 80.790 ;
        RECT 75.055 80.730 75.345 80.775 ;
        RECT 74.580 80.590 75.345 80.730 ;
        RECT 74.580 80.530 74.900 80.590 ;
        RECT 75.055 80.545 75.345 80.590 ;
        RECT 76.880 80.530 77.200 80.790 ;
        RECT 77.340 80.730 77.660 80.790 ;
        RECT 78.350 80.775 78.490 80.930 ;
        RECT 79.180 80.930 80.405 81.070 ;
        RECT 79.180 80.870 79.500 80.930 ;
        RECT 80.115 80.885 80.405 80.930 ;
        RECT 80.995 81.070 81.285 81.115 ;
        RECT 82.185 81.070 82.475 81.115 ;
        RECT 84.705 81.070 84.995 81.115 ;
        RECT 80.995 80.930 84.995 81.070 ;
        RECT 80.995 80.885 81.285 80.930 ;
        RECT 82.185 80.885 82.475 80.930 ;
        RECT 84.705 80.885 84.995 80.930 ;
        RECT 77.815 80.730 78.105 80.775 ;
        RECT 77.340 80.590 78.105 80.730 ;
        RECT 77.340 80.530 77.660 80.590 ;
        RECT 77.815 80.545 78.105 80.590 ;
        RECT 78.275 80.545 78.565 80.775 ;
        RECT 78.720 80.530 79.040 80.790 ;
        RECT 85.160 80.730 85.480 80.790 ;
        RECT 87.475 80.730 87.765 80.775 ;
        RECT 85.160 80.590 87.765 80.730 ;
        RECT 85.160 80.530 85.480 80.590 ;
        RECT 87.475 80.545 87.765 80.590 ;
        RECT 80.100 80.390 80.420 80.450 ;
        RECT 73.750 80.250 80.420 80.390 ;
        RECT 77.890 80.110 78.030 80.250 ;
        RECT 80.100 80.190 80.420 80.250 ;
        RECT 81.450 80.390 81.740 80.435 ;
        RECT 81.940 80.390 82.260 80.450 ;
        RECT 81.450 80.250 82.260 80.390 ;
        RECT 81.450 80.205 81.740 80.250 ;
        RECT 81.940 80.190 82.260 80.250 ;
        RECT 68.600 79.910 73.430 80.050 ;
        RECT 68.600 79.850 68.920 79.910 ;
        RECT 77.800 79.850 78.120 80.110 ;
        RECT 79.655 80.050 79.945 80.095 ;
        RECT 84.240 80.050 84.560 80.110 ;
        RECT 79.655 79.910 84.560 80.050 ;
        RECT 79.655 79.865 79.945 79.910 ;
        RECT 84.240 79.850 84.560 79.910 ;
        RECT 11.950 79.230 90.610 79.710 ;
        RECT 21.220 78.830 21.540 79.090 ;
        RECT 34.100 78.830 34.420 79.090 ;
        RECT 44.680 79.030 45.000 79.090 ;
        RECT 45.155 79.030 45.445 79.075 ;
        RECT 44.680 78.890 45.445 79.030 ;
        RECT 44.680 78.830 45.000 78.890 ;
        RECT 45.155 78.845 45.445 78.890 ;
        RECT 46.075 79.030 46.365 79.075 ;
        RECT 46.980 79.030 47.300 79.090 ;
        RECT 46.075 78.890 47.300 79.030 ;
        RECT 46.075 78.845 46.365 78.890 ;
        RECT 46.980 78.830 47.300 78.890 ;
        RECT 56.195 79.030 56.485 79.075 ;
        RECT 56.640 79.030 56.960 79.090 ;
        RECT 69.060 79.030 69.380 79.090 ;
        RECT 71.820 79.030 72.140 79.090 ;
        RECT 76.435 79.030 76.725 79.075 ;
        RECT 76.880 79.030 77.200 79.090 ;
        RECT 56.195 78.890 56.960 79.030 ;
        RECT 56.195 78.845 56.485 78.890 ;
        RECT 56.640 78.830 56.960 78.890 ;
        RECT 65.010 78.890 74.350 79.030 ;
        RECT 20.300 78.690 20.620 78.750 ;
        RECT 14.410 78.550 20.620 78.690 ;
        RECT 21.310 78.690 21.450 78.830 ;
        RECT 41.000 78.690 41.320 78.750 ;
        RECT 21.310 78.550 25.130 78.690 ;
        RECT 14.410 78.395 14.550 78.550 ;
        RECT 20.300 78.490 20.620 78.550 ;
        RECT 15.700 78.395 16.020 78.410 ;
        RECT 14.335 78.165 14.625 78.395 ;
        RECT 15.670 78.165 16.020 78.395 ;
        RECT 15.700 78.150 16.020 78.165 ;
        RECT 22.140 78.350 22.460 78.410 ;
        RECT 24.990 78.395 25.130 78.550 ;
        RECT 27.290 78.550 41.320 78.690 ;
        RECT 27.290 78.395 27.430 78.550 ;
        RECT 23.535 78.350 23.825 78.395 ;
        RECT 22.140 78.210 23.825 78.350 ;
        RECT 22.140 78.150 22.460 78.210 ;
        RECT 23.535 78.165 23.825 78.210 ;
        RECT 24.915 78.165 25.205 78.395 ;
        RECT 27.215 78.165 27.505 78.395 ;
        RECT 27.660 78.350 27.980 78.410 ;
        RECT 38.330 78.395 38.470 78.550 ;
        RECT 41.000 78.490 41.320 78.550 ;
        RECT 50.660 78.690 50.980 78.750 ;
        RECT 54.340 78.690 54.660 78.750 ;
        RECT 50.660 78.550 54.660 78.690 ;
        RECT 50.660 78.490 50.980 78.550 ;
        RECT 54.340 78.490 54.660 78.550 ;
        RECT 61.870 78.690 62.160 78.735 ;
        RECT 64.015 78.690 64.305 78.735 ;
        RECT 61.870 78.550 64.305 78.690 ;
        RECT 61.870 78.505 62.160 78.550 ;
        RECT 64.015 78.505 64.305 78.550 ;
        RECT 39.620 78.395 39.940 78.410 ;
        RECT 28.495 78.350 28.785 78.395 ;
        RECT 27.660 78.210 28.785 78.350 ;
        RECT 27.660 78.150 27.980 78.210 ;
        RECT 28.495 78.165 28.785 78.210 ;
        RECT 38.255 78.165 38.545 78.395 ;
        RECT 39.590 78.165 39.940 78.395 ;
        RECT 39.620 78.150 39.940 78.165 ;
        RECT 51.580 78.395 51.900 78.410 ;
        RECT 51.580 78.165 51.930 78.395 ;
        RECT 62.620 78.350 62.940 78.410 ;
        RECT 65.010 78.395 65.150 78.890 ;
        RECT 69.060 78.830 69.380 78.890 ;
        RECT 71.820 78.830 72.140 78.890 ;
        RECT 68.600 78.690 68.920 78.750 ;
        RECT 72.280 78.690 72.600 78.750 ;
        RECT 73.675 78.690 73.965 78.735 ;
        RECT 68.230 78.550 68.920 78.690 ;
        RECT 63.095 78.350 63.385 78.395 ;
        RECT 62.620 78.210 63.385 78.350 ;
        RECT 51.580 78.150 51.900 78.165 ;
        RECT 62.620 78.150 62.940 78.210 ;
        RECT 63.095 78.165 63.385 78.210 ;
        RECT 64.935 78.165 65.225 78.395 ;
        RECT 65.395 78.350 65.685 78.395 ;
        RECT 65.840 78.350 66.160 78.410 ;
        RECT 68.230 78.395 68.370 78.550 ;
        RECT 68.600 78.490 68.920 78.550 ;
        RECT 69.150 78.550 73.965 78.690 ;
        RECT 74.210 78.690 74.350 78.890 ;
        RECT 76.435 78.890 77.200 79.030 ;
        RECT 76.435 78.845 76.725 78.890 ;
        RECT 76.880 78.830 77.200 78.890 ;
        RECT 81.940 78.830 82.260 79.090 ;
        RECT 83.795 79.030 84.085 79.075 ;
        RECT 85.620 79.030 85.940 79.090 ;
        RECT 83.795 78.890 85.940 79.030 ;
        RECT 83.795 78.845 84.085 78.890 ;
        RECT 85.620 78.830 85.940 78.890 ;
        RECT 74.595 78.690 74.885 78.735 ;
        RECT 74.210 78.550 74.885 78.690 ;
        RECT 65.395 78.210 66.160 78.350 ;
        RECT 65.395 78.165 65.685 78.210 ;
        RECT 65.840 78.150 66.160 78.210 ;
        RECT 66.315 78.165 66.605 78.395 ;
        RECT 68.155 78.165 68.445 78.395 ;
        RECT 69.150 78.350 69.290 78.550 ;
        RECT 72.280 78.490 72.600 78.550 ;
        RECT 73.675 78.505 73.965 78.550 ;
        RECT 74.595 78.505 74.885 78.550 ;
        RECT 84.240 78.490 84.560 78.750 ;
        RECT 68.690 78.210 69.290 78.350 ;
        RECT 15.215 78.010 15.505 78.055 ;
        RECT 16.405 78.010 16.695 78.055 ;
        RECT 18.925 78.010 19.215 78.055 ;
        RECT 15.215 77.870 19.215 78.010 ;
        RECT 15.215 77.825 15.505 77.870 ;
        RECT 16.405 77.825 16.695 77.870 ;
        RECT 18.925 77.825 19.215 77.870 ;
        RECT 28.095 78.010 28.385 78.055 ;
        RECT 29.285 78.010 29.575 78.055 ;
        RECT 31.805 78.010 32.095 78.055 ;
        RECT 28.095 77.870 32.095 78.010 ;
        RECT 28.095 77.825 28.385 77.870 ;
        RECT 29.285 77.825 29.575 77.870 ;
        RECT 31.805 77.825 32.095 77.870 ;
        RECT 39.135 78.010 39.425 78.055 ;
        RECT 40.325 78.010 40.615 78.055 ;
        RECT 42.845 78.010 43.135 78.055 ;
        RECT 39.135 77.870 43.135 78.010 ;
        RECT 39.135 77.825 39.425 77.870 ;
        RECT 40.325 77.825 40.615 77.870 ;
        RECT 42.845 77.825 43.135 77.870 ;
        RECT 48.385 78.010 48.675 78.055 ;
        RECT 50.905 78.010 51.195 78.055 ;
        RECT 52.095 78.010 52.385 78.055 ;
        RECT 48.385 77.870 52.385 78.010 ;
        RECT 48.385 77.825 48.675 77.870 ;
        RECT 50.905 77.825 51.195 77.870 ;
        RECT 52.095 77.825 52.385 77.870 ;
        RECT 52.975 77.825 53.265 78.055 ;
        RECT 58.505 78.010 58.795 78.055 ;
        RECT 61.025 78.010 61.315 78.055 ;
        RECT 62.215 78.010 62.505 78.055 ;
        RECT 58.505 77.870 62.505 78.010 ;
        RECT 66.390 78.010 66.530 78.165 ;
        RECT 68.690 78.055 68.830 78.210 ;
        RECT 69.520 78.150 69.840 78.410 ;
        RECT 70.440 78.350 70.760 78.410 ;
        RECT 71.375 78.350 71.665 78.395 ;
        RECT 70.440 78.210 71.665 78.350 ;
        RECT 70.440 78.150 70.760 78.210 ;
        RECT 71.375 78.165 71.665 78.210 ;
        RECT 67.235 78.010 67.525 78.055 ;
        RECT 66.390 77.870 67.525 78.010 ;
        RECT 58.505 77.825 58.795 77.870 ;
        RECT 61.025 77.825 61.315 77.870 ;
        RECT 62.215 77.825 62.505 77.870 ;
        RECT 67.235 77.825 67.525 77.870 ;
        RECT 68.615 77.825 68.905 78.055 ;
        RECT 69.060 78.010 69.380 78.070 ;
        RECT 69.980 78.010 70.300 78.070 ;
        RECT 69.060 77.870 70.300 78.010 ;
        RECT 71.450 78.010 71.590 78.165 ;
        RECT 72.740 78.150 73.060 78.410 ;
        RECT 74.135 78.165 74.425 78.395 ;
        RECT 75.515 78.350 75.805 78.395 ;
        RECT 76.880 78.350 77.200 78.410 ;
        RECT 75.515 78.210 77.200 78.350 ;
        RECT 75.515 78.165 75.805 78.210 ;
        RECT 74.210 78.010 74.350 78.165 ;
        RECT 76.880 78.150 77.200 78.210 ;
        RECT 86.095 78.350 86.385 78.395 ;
        RECT 87.000 78.350 87.320 78.410 ;
        RECT 86.095 78.210 87.320 78.350 ;
        RECT 86.095 78.165 86.385 78.210 ;
        RECT 87.000 78.150 87.320 78.210 ;
        RECT 78.260 78.010 78.580 78.070 ;
        RECT 71.450 77.870 78.580 78.010 ;
        RECT 14.820 77.670 15.110 77.715 ;
        RECT 16.920 77.670 17.210 77.715 ;
        RECT 18.490 77.670 18.780 77.715 ;
        RECT 14.820 77.530 18.780 77.670 ;
        RECT 14.820 77.485 15.110 77.530 ;
        RECT 16.920 77.485 17.210 77.530 ;
        RECT 18.490 77.485 18.780 77.530 ;
        RECT 23.520 77.670 23.840 77.730 ;
        RECT 26.295 77.670 26.585 77.715 ;
        RECT 23.520 77.530 26.585 77.670 ;
        RECT 23.520 77.470 23.840 77.530 ;
        RECT 26.295 77.485 26.585 77.530 ;
        RECT 27.700 77.670 27.990 77.715 ;
        RECT 29.800 77.670 30.090 77.715 ;
        RECT 31.370 77.670 31.660 77.715 ;
        RECT 27.700 77.530 31.660 77.670 ;
        RECT 27.700 77.485 27.990 77.530 ;
        RECT 29.800 77.485 30.090 77.530 ;
        RECT 31.370 77.485 31.660 77.530 ;
        RECT 38.740 77.670 39.030 77.715 ;
        RECT 40.840 77.670 41.130 77.715 ;
        RECT 42.410 77.670 42.700 77.715 ;
        RECT 38.740 77.530 42.700 77.670 ;
        RECT 38.740 77.485 39.030 77.530 ;
        RECT 40.840 77.485 41.130 77.530 ;
        RECT 42.410 77.485 42.700 77.530 ;
        RECT 48.820 77.670 49.110 77.715 ;
        RECT 50.390 77.670 50.680 77.715 ;
        RECT 52.490 77.670 52.780 77.715 ;
        RECT 48.820 77.530 52.780 77.670 ;
        RECT 48.820 77.485 49.110 77.530 ;
        RECT 50.390 77.485 50.680 77.530 ;
        RECT 52.490 77.485 52.780 77.530 ;
        RECT 23.980 77.130 24.300 77.390 ;
        RECT 51.120 77.330 51.440 77.390 ;
        RECT 53.050 77.330 53.190 77.825 ;
        RECT 69.060 77.810 69.380 77.870 ;
        RECT 69.980 77.810 70.300 77.870 ;
        RECT 78.260 77.810 78.580 77.870 ;
        RECT 84.700 77.810 85.020 78.070 ;
        RECT 99.980 77.735 100.370 81.555 ;
        RECT 101.460 81.315 102.460 83.715 ;
        RECT 102.950 81.585 103.950 83.735 ;
        RECT 101.210 81.085 102.460 81.315 ;
        RECT 100.650 80.925 102.460 81.085 ;
        RECT 102.720 80.945 103.950 81.585 ;
        RECT 104.430 81.575 105.430 83.725 ;
        RECT 105.890 81.575 106.890 83.715 ;
        RECT 100.650 80.625 101.930 80.925 ;
        RECT 100.650 78.745 101.650 80.625 ;
        RECT 102.720 80.475 103.400 80.945 ;
        RECT 104.210 80.935 105.430 81.575 ;
        RECT 104.210 80.475 104.890 80.935 ;
        RECT 105.700 80.925 106.890 81.575 ;
        RECT 107.390 81.545 108.390 83.735 ;
        RECT 110.330 83.715 112.640 83.725 ;
        RECT 107.150 80.945 108.390 81.545 ;
        RECT 108.900 81.535 109.900 83.715 ;
        RECT 110.330 81.545 112.810 83.715 ;
        RECT 118.020 83.515 118.360 84.370 ;
        RECT 118.020 83.510 118.340 83.515 ;
        RECT 118.020 82.930 118.260 83.510 ;
        RECT 118.670 83.310 119.140 91.720 ;
        RECT 119.640 91.515 119.860 92.280 ;
        RECT 120.840 91.720 122.800 91.950 ;
        RECT 124.270 91.720 126.230 91.950 ;
        RECT 127.700 91.720 128.660 91.950 ;
        RECT 119.420 91.310 119.860 91.515 ;
        RECT 120.560 91.490 120.790 91.515 ;
        RECT 120.560 91.480 120.800 91.490 ;
        RECT 119.420 83.570 119.810 91.310 ;
        RECT 120.390 84.420 120.800 91.480 ;
        RECT 121.380 85.130 122.280 91.720 ;
        RECT 122.850 91.470 123.080 91.515 ;
        RECT 123.990 91.490 124.220 91.515 ;
        RECT 120.380 83.600 120.800 84.420 ;
        RECT 121.350 84.120 122.350 85.130 ;
        RECT 119.420 83.515 119.650 83.570 ;
        RECT 120.380 83.515 120.790 83.600 ;
        RECT 118.410 83.080 119.370 83.310 ;
        RECT 118.020 82.440 118.340 82.930 ;
        RECT 105.700 80.475 106.380 80.925 ;
        RECT 107.150 80.475 107.830 80.945 ;
        RECT 102.100 80.005 103.400 80.475 ;
        RECT 102.100 78.835 103.140 80.005 ;
        RECT 103.610 79.995 104.890 80.475 ;
        RECT 105.080 79.995 106.380 80.475 ;
        RECT 103.610 78.835 104.650 79.995 ;
        RECT 105.080 78.835 106.120 79.995 ;
        RECT 106.570 79.965 107.830 80.475 ;
        RECT 108.650 80.925 109.900 81.535 ;
        RECT 110.160 80.935 112.810 81.545 ;
        RECT 117.580 81.190 118.420 82.440 ;
        RECT 108.650 80.465 109.330 80.925 ;
        RECT 110.160 80.475 110.840 80.935 ;
        RECT 111.810 80.925 112.810 80.935 ;
        RECT 100.650 78.295 101.880 78.745 ;
        RECT 102.100 78.295 103.430 78.835 ;
        RECT 103.610 78.295 104.920 78.835 ;
        RECT 105.080 78.295 106.410 78.835 ;
        RECT 106.570 78.825 107.610 79.965 ;
        RECT 108.050 79.955 109.330 80.465 ;
        RECT 109.530 79.965 110.840 80.475 ;
        RECT 118.020 80.140 118.260 81.190 ;
        RECT 118.560 80.530 119.230 83.080 ;
        RECT 120.380 81.300 120.700 83.515 ;
        RECT 121.380 83.310 122.280 84.120 ;
        RECT 122.850 83.580 123.370 91.470 ;
        RECT 122.850 83.515 123.080 83.580 ;
        RECT 123.850 83.570 124.230 91.490 ;
        RECT 124.930 85.090 125.750 91.720 ;
        RECT 126.280 91.470 126.510 91.515 ;
        RECT 127.420 91.470 127.650 91.515 ;
        RECT 124.840 84.090 125.840 85.090 ;
        RECT 123.860 83.515 124.220 83.570 ;
        RECT 120.840 83.080 122.800 83.310 ;
        RECT 123.860 81.950 124.120 83.515 ;
        RECT 124.930 83.310 125.750 84.090 ;
        RECT 126.280 83.600 127.660 91.470 ;
        RECT 128.010 91.350 128.430 91.720 ;
        RECT 128.710 91.470 128.940 91.515 ;
        RECT 129.340 91.470 130.480 92.280 ;
        RECT 128.710 87.490 130.480 91.470 ;
        RECT 128.710 86.490 130.470 87.490 ;
        RECT 126.280 83.515 126.510 83.600 ;
        RECT 127.420 83.515 127.650 83.600 ;
        RECT 128.010 83.310 128.430 83.980 ;
        RECT 128.710 83.610 130.480 86.490 ;
        RECT 128.710 83.515 128.940 83.610 ;
        RECT 124.270 83.080 126.230 83.310 ;
        RECT 127.700 83.080 128.660 83.310 ;
        RECT 127.800 82.200 128.590 83.080 ;
        RECT 129.340 82.600 130.480 83.610 ;
        RECT 123.860 81.330 127.480 81.950 ;
        RECT 127.750 81.440 128.640 82.200 ;
        RECT 118.420 80.300 119.380 80.530 ;
        RECT 108.050 78.825 109.090 79.955 ;
        RECT 106.570 78.295 107.840 78.825 ;
        RECT 101.200 77.735 101.880 78.295 ;
        RECT 102.750 77.745 103.430 78.295 ;
        RECT 104.240 77.755 104.920 78.295 ;
        RECT 105.730 77.755 106.410 78.295 ;
        RECT 107.160 77.755 107.840 78.295 ;
        RECT 108.050 78.285 109.350 78.825 ;
        RECT 109.530 78.295 110.570 79.965 ;
        RECT 118.020 79.130 118.370 80.140 ;
        RECT 108.670 77.755 109.350 78.285 ;
        RECT 58.940 77.670 59.230 77.715 ;
        RECT 60.510 77.670 60.800 77.715 ;
        RECT 62.610 77.670 62.900 77.715 ;
        RECT 58.940 77.530 62.900 77.670 ;
        RECT 58.940 77.485 59.230 77.530 ;
        RECT 60.510 77.485 60.800 77.530 ;
        RECT 62.610 77.485 62.900 77.530 ;
        RECT 65.840 77.470 66.160 77.730 ;
        RECT 72.740 77.670 73.060 77.730 ;
        RECT 74.120 77.670 74.440 77.730 ;
        RECT 72.740 77.530 74.440 77.670 ;
        RECT 72.740 77.470 73.060 77.530 ;
        RECT 74.120 77.470 74.440 77.530 ;
        RECT 51.120 77.190 53.190 77.330 ;
        RECT 87.015 77.330 87.305 77.375 ;
        RECT 87.460 77.330 87.780 77.390 ;
        RECT 87.015 77.190 87.780 77.330 ;
        RECT 51.120 77.130 51.440 77.190 ;
        RECT 87.015 77.145 87.305 77.190 ;
        RECT 87.460 77.130 87.780 77.190 ;
        RECT 11.950 76.510 90.610 76.990 ;
        RECT 15.255 76.310 15.545 76.355 ;
        RECT 15.700 76.310 16.020 76.370 ;
        RECT 15.255 76.170 16.020 76.310 ;
        RECT 15.255 76.125 15.545 76.170 ;
        RECT 15.700 76.110 16.020 76.170 ;
        RECT 19.855 76.310 20.145 76.355 ;
        RECT 21.220 76.310 21.540 76.370 ;
        RECT 19.855 76.170 21.540 76.310 ;
        RECT 19.855 76.125 20.145 76.170 ;
        RECT 21.220 76.110 21.540 76.170 ;
        RECT 22.140 76.110 22.460 76.370 ;
        RECT 39.620 76.310 39.940 76.370 ;
        RECT 41.015 76.310 41.305 76.355 ;
        RECT 50.660 76.310 50.980 76.370 ;
        RECT 39.620 76.170 41.305 76.310 ;
        RECT 39.620 76.110 39.940 76.170 ;
        RECT 41.015 76.125 41.305 76.170 ;
        RECT 43.850 76.170 50.980 76.310 ;
        RECT 18.015 75.970 18.305 76.015 ;
        RECT 22.230 75.970 22.370 76.110 ;
        RECT 18.015 75.830 22.370 75.970 ;
        RECT 28.160 75.970 28.450 76.015 ;
        RECT 30.260 75.970 30.550 76.015 ;
        RECT 31.830 75.970 32.120 76.015 ;
        RECT 28.160 75.830 32.120 75.970 ;
        RECT 18.015 75.785 18.305 75.830 ;
        RECT 28.160 75.785 28.450 75.830 ;
        RECT 30.260 75.785 30.550 75.830 ;
        RECT 31.830 75.785 32.120 75.830 ;
        RECT 40.540 75.970 40.860 76.030 ;
        RECT 43.850 75.970 43.990 76.170 ;
        RECT 50.660 76.110 50.980 76.170 ;
        RECT 51.135 76.310 51.425 76.355 ;
        RECT 51.580 76.310 51.900 76.370 ;
        RECT 51.135 76.170 51.900 76.310 ;
        RECT 51.135 76.125 51.425 76.170 ;
        RECT 51.580 76.110 51.900 76.170 ;
        RECT 55.735 76.310 56.025 76.355 ;
        RECT 71.360 76.310 71.680 76.370 ;
        RECT 71.835 76.310 72.125 76.355 ;
        RECT 75.040 76.310 75.360 76.370 ;
        RECT 55.735 76.170 63.310 76.310 ;
        RECT 55.735 76.125 56.025 76.170 ;
        RECT 55.810 75.970 55.950 76.125 ;
        RECT 40.540 75.830 43.990 75.970 ;
        RECT 40.540 75.770 40.860 75.830 ;
        RECT 16.620 75.630 16.940 75.690 ;
        RECT 19.840 75.630 20.160 75.690 ;
        RECT 16.250 75.490 20.160 75.630 ;
        RECT 16.250 75.335 16.390 75.490 ;
        RECT 16.620 75.430 16.940 75.490 ;
        RECT 19.840 75.430 20.160 75.490 ;
        RECT 28.555 75.630 28.845 75.675 ;
        RECT 29.745 75.630 30.035 75.675 ;
        RECT 32.265 75.630 32.555 75.675 ;
        RECT 28.555 75.490 32.555 75.630 ;
        RECT 28.555 75.445 28.845 75.490 ;
        RECT 29.745 75.445 30.035 75.490 ;
        RECT 32.265 75.445 32.555 75.490 ;
        RECT 43.300 75.430 43.620 75.690 ;
        RECT 43.850 75.675 43.990 75.830 ;
        RECT 47.530 75.830 55.950 75.970 ;
        RECT 58.480 75.970 58.770 76.015 ;
        RECT 60.050 75.970 60.340 76.015 ;
        RECT 62.150 75.970 62.440 76.015 ;
        RECT 58.480 75.830 62.440 75.970 ;
        RECT 47.530 75.675 47.670 75.830 ;
        RECT 58.480 75.785 58.770 75.830 ;
        RECT 60.050 75.785 60.340 75.830 ;
        RECT 62.150 75.785 62.440 75.830 ;
        RECT 43.775 75.445 44.065 75.675 ;
        RECT 47.455 75.445 47.745 75.675 ;
        RECT 47.915 75.445 48.205 75.675 ;
        RECT 50.200 75.630 50.520 75.690 ;
        RECT 53.435 75.630 53.725 75.675 ;
        RECT 50.200 75.490 53.725 75.630 ;
        RECT 16.175 75.105 16.465 75.335 ;
        RECT 17.080 75.090 17.400 75.350 ;
        RECT 21.220 75.290 21.540 75.350 ;
        RECT 21.695 75.290 21.985 75.335 ;
        RECT 21.220 75.150 21.985 75.290 ;
        RECT 21.220 75.090 21.540 75.150 ;
        RECT 21.695 75.105 21.985 75.150 ;
        RECT 23.535 75.290 23.825 75.335 ;
        RECT 23.980 75.290 24.300 75.350 ;
        RECT 23.535 75.150 24.300 75.290 ;
        RECT 23.535 75.105 23.825 75.150 ;
        RECT 23.980 75.090 24.300 75.150 ;
        RECT 27.675 75.290 27.965 75.335 ;
        RECT 40.095 75.290 40.385 75.335 ;
        RECT 41.000 75.290 41.320 75.350 ;
        RECT 27.675 75.150 41.320 75.290 ;
        RECT 27.675 75.105 27.965 75.150 ;
        RECT 40.095 75.105 40.385 75.150 ;
        RECT 41.000 75.090 41.320 75.150 ;
        RECT 46.060 75.290 46.380 75.350 ;
        RECT 47.990 75.290 48.130 75.445 ;
        RECT 50.200 75.430 50.520 75.490 ;
        RECT 53.435 75.445 53.725 75.490 ;
        RECT 54.340 75.430 54.660 75.690 ;
        RECT 63.170 75.675 63.310 76.170 ;
        RECT 71.360 76.170 75.360 76.310 ;
        RECT 71.360 76.110 71.680 76.170 ;
        RECT 71.835 76.125 72.125 76.170 ;
        RECT 75.040 76.110 75.360 76.170 ;
        RECT 87.000 76.110 87.320 76.370 ;
        RECT 65.840 75.970 66.160 76.030 ;
        RECT 80.600 75.970 80.890 76.015 ;
        RECT 82.700 75.970 82.990 76.015 ;
        RECT 84.270 75.970 84.560 76.015 ;
        RECT 65.840 75.830 69.750 75.970 ;
        RECT 65.840 75.770 66.160 75.830 ;
        RECT 58.045 75.630 58.335 75.675 ;
        RECT 60.565 75.630 60.855 75.675 ;
        RECT 61.755 75.630 62.045 75.675 ;
        RECT 58.045 75.490 62.045 75.630 ;
        RECT 58.045 75.445 58.335 75.490 ;
        RECT 60.565 75.445 60.855 75.490 ;
        RECT 61.755 75.445 62.045 75.490 ;
        RECT 63.095 75.445 63.385 75.675 ;
        RECT 66.315 75.630 66.605 75.675 ;
        RECT 66.315 75.490 68.370 75.630 ;
        RECT 66.315 75.445 66.605 75.490 ;
        RECT 46.060 75.150 48.130 75.290 ;
        RECT 51.120 75.290 51.440 75.350 ;
        RECT 55.720 75.290 56.040 75.350 ;
        RECT 62.620 75.290 62.940 75.350 ;
        RECT 51.120 75.150 62.940 75.290 ;
        RECT 46.060 75.090 46.380 75.150 ;
        RECT 51.120 75.090 51.440 75.150 ;
        RECT 55.720 75.090 56.040 75.150 ;
        RECT 62.620 75.090 62.940 75.150 ;
        RECT 64.460 75.290 64.780 75.350 ;
        RECT 67.680 75.290 68.000 75.350 ;
        RECT 68.230 75.335 68.370 75.490 ;
        RECT 69.060 75.430 69.380 75.690 ;
        RECT 69.610 75.335 69.750 75.830 ;
        RECT 80.600 75.830 84.560 75.970 ;
        RECT 80.600 75.785 80.890 75.830 ;
        RECT 82.700 75.785 82.990 75.830 ;
        RECT 84.270 75.785 84.560 75.830 ;
        RECT 69.980 75.630 70.300 75.690 ;
        RECT 71.820 75.630 72.140 75.690 ;
        RECT 69.980 75.490 72.140 75.630 ;
        RECT 69.980 75.430 70.300 75.490 ;
        RECT 71.820 75.430 72.140 75.490 ;
        RECT 75.500 75.630 75.820 75.690 ;
        RECT 77.340 75.630 77.660 75.690 ;
        RECT 75.500 75.490 77.660 75.630 ;
        RECT 75.500 75.430 75.820 75.490 ;
        RECT 77.340 75.430 77.660 75.490 ;
        RECT 79.180 75.630 79.500 75.690 ;
        RECT 80.100 75.630 80.420 75.690 ;
        RECT 79.180 75.490 80.420 75.630 ;
        RECT 79.180 75.430 79.500 75.490 ;
        RECT 80.100 75.430 80.420 75.490 ;
        RECT 80.995 75.630 81.285 75.675 ;
        RECT 82.185 75.630 82.475 75.675 ;
        RECT 84.705 75.630 84.995 75.675 ;
        RECT 80.995 75.490 84.995 75.630 ;
        RECT 99.980 75.585 101.000 77.735 ;
        RECT 101.200 77.165 102.510 77.735 ;
        RECT 102.750 77.255 103.960 77.745 ;
        RECT 104.240 77.255 105.470 77.755 ;
        RECT 105.730 77.255 106.940 77.755 ;
        RECT 101.470 75.575 102.510 77.165 ;
        RECT 102.920 75.565 103.960 77.255 ;
        RECT 104.430 75.575 105.470 77.255 ;
        RECT 105.900 75.575 106.940 77.255 ;
        RECT 107.160 77.245 108.430 77.755 ;
        RECT 108.670 77.245 109.900 77.755 ;
        RECT 107.390 75.575 108.430 77.245 ;
        RECT 108.860 75.575 109.900 77.245 ;
        RECT 118.030 76.180 118.370 79.130 ;
        RECT 118.140 76.140 118.370 76.180 ;
        RECT 118.670 75.980 119.110 80.300 ;
        RECT 120.380 80.140 120.710 81.300 ;
        RECT 120.850 80.300 122.810 80.530 ;
        RECT 119.430 80.130 119.660 80.140 ;
        RECT 119.430 77.820 119.840 80.130 ;
        RECT 120.380 80.100 120.800 80.140 ;
        RECT 121.160 80.100 122.500 80.300 ;
        RECT 123.860 80.140 124.120 81.330 ;
        RECT 127.070 80.680 127.470 81.330 ;
        RECT 129.410 81.250 130.480 82.600 ;
        RECT 134.410 84.950 139.730 85.560 ;
        RECT 134.410 84.870 136.330 84.950 ;
        RECT 134.410 84.540 136.160 84.870 ;
        RECT 134.410 83.750 134.760 84.540 ;
        RECT 136.910 84.520 139.710 84.770 ;
        RECT 135.150 84.300 135.440 84.330 ;
        RECT 135.140 84.050 135.460 84.300 ;
        RECT 136.910 83.895 137.070 84.520 ;
        RECT 137.210 84.050 137.540 84.380 ;
        RECT 137.820 84.250 138.030 84.520 ;
        RECT 137.890 83.910 138.030 84.250 ;
        RECT 138.170 84.050 138.500 84.380 ;
        RECT 138.970 84.040 139.710 84.520 ;
        RECT 137.890 83.895 138.180 83.910 ;
        RECT 138.970 83.895 139.140 84.040 ;
        RECT 139.320 83.960 139.710 84.040 ;
        RECT 134.960 83.750 135.190 83.895 ;
        RECT 129.410 80.820 131.250 81.250 ;
        RECT 129.410 80.780 130.470 80.820 ;
        RECT 128.470 80.680 129.220 80.690 ;
        RECT 127.070 80.630 129.220 80.680 ;
        RECT 127.070 80.590 129.400 80.630 ;
        RECT 124.280 80.300 126.240 80.530 ;
        RECT 127.070 80.340 130.630 80.590 ;
        RECT 127.070 80.330 128.410 80.340 ;
        RECT 128.120 80.310 128.410 80.330 ;
        RECT 120.380 79.170 122.500 80.100 ;
        RECT 119.430 76.140 119.930 77.820 ;
        RECT 120.500 76.200 122.500 79.170 ;
        RECT 120.570 76.140 120.800 76.200 ;
        RECT 118.420 75.750 119.380 75.980 ;
        RECT 119.730 75.520 119.930 76.140 ;
        RECT 121.160 75.980 122.500 76.200 ;
        RECT 122.860 80.090 123.090 80.140 ;
        RECT 123.860 80.090 124.230 80.140 ;
        RECT 124.570 80.090 125.940 80.300 ;
        RECT 129.280 80.250 130.630 80.340 ;
        RECT 130.230 80.245 130.520 80.250 ;
        RECT 122.860 77.870 123.310 80.090 ;
        RECT 123.860 79.800 125.940 80.090 ;
        RECT 122.860 77.380 123.360 77.870 ;
        RECT 122.860 76.710 123.450 77.380 ;
        RECT 122.860 76.460 123.510 76.710 ;
        RECT 122.860 76.430 123.560 76.460 ;
        RECT 122.860 76.140 123.090 76.430 ;
        RECT 123.320 76.060 123.560 76.430 ;
        RECT 123.870 76.200 125.940 79.800 ;
        RECT 123.870 76.180 124.230 76.200 ;
        RECT 124.000 76.140 124.230 76.180 ;
        RECT 120.850 75.750 122.810 75.980 ;
        RECT 123.240 75.820 123.560 76.060 ;
        RECT 124.570 75.980 125.940 76.200 ;
        RECT 126.290 79.960 126.520 80.140 ;
        RECT 127.930 80.090 128.160 80.150 ;
        RECT 128.370 80.090 128.600 80.150 ;
        RECT 127.180 80.080 128.160 80.090 ;
        RECT 126.750 79.960 128.160 80.080 ;
        RECT 126.290 79.210 128.160 79.960 ;
        RECT 128.350 79.950 128.750 80.090 ;
        RECT 130.040 79.950 130.270 80.040 ;
        RECT 130.480 79.990 130.710 80.040 ;
        RECT 130.880 79.990 131.250 80.820 ;
        RECT 128.350 79.220 130.310 79.950 ;
        RECT 128.350 79.210 128.750 79.220 ;
        RECT 126.290 78.750 127.650 79.210 ;
        RECT 127.930 79.150 128.160 79.210 ;
        RECT 128.370 79.150 128.600 79.210 ;
        RECT 126.290 78.480 128.750 78.750 ;
        RECT 126.290 78.440 128.460 78.480 ;
        RECT 126.290 76.690 127.640 78.440 ;
        RECT 128.920 78.260 130.300 79.220 ;
        RECT 128.920 78.130 130.320 78.260 ;
        RECT 128.200 77.130 130.320 78.130 ;
        RECT 128.920 77.100 130.320 77.130 ;
        RECT 130.040 77.090 130.320 77.100 ;
        RECT 130.480 77.130 131.250 79.990 ;
        RECT 134.410 79.895 135.190 83.750 ;
        RECT 135.400 83.840 135.630 83.895 ;
        RECT 135.400 80.660 136.040 83.840 ;
        RECT 135.400 79.950 136.050 80.660 ;
        RECT 136.540 80.130 136.770 83.895 ;
        RECT 136.910 83.750 137.250 83.895 ;
        RECT 135.400 79.895 135.630 79.950 ;
        RECT 134.410 79.880 135.160 79.895 ;
        RECT 134.410 79.870 134.760 79.880 ;
        RECT 135.150 79.590 135.440 79.690 ;
        RECT 134.910 79.080 135.590 79.590 ;
        RECT 134.410 78.080 135.590 79.080 ;
        RECT 134.910 77.590 135.590 78.080 ;
        RECT 135.140 77.550 135.430 77.590 ;
        RECT 134.950 77.340 135.180 77.390 ;
        RECT 130.040 77.040 130.270 77.090 ;
        RECT 130.480 77.040 130.710 77.130 ;
        RECT 130.880 77.100 131.250 77.130 ;
        RECT 126.290 76.390 128.990 76.690 ;
        RECT 126.290 76.140 126.520 76.390 ;
        RECT 123.200 75.520 123.560 75.820 ;
        RECT 124.280 75.750 126.240 75.980 ;
        RECT 126.900 75.520 128.990 76.390 ;
        RECT 80.995 75.445 81.285 75.490 ;
        RECT 82.185 75.445 82.475 75.490 ;
        RECT 84.705 75.445 84.995 75.490 ;
        RECT 64.460 75.150 68.000 75.290 ;
        RECT 64.460 75.090 64.780 75.150 ;
        RECT 67.680 75.090 68.000 75.150 ;
        RECT 68.155 75.105 68.445 75.335 ;
        RECT 69.535 75.105 69.825 75.335 ;
        RECT 70.900 75.090 71.220 75.350 ;
        RECT 71.910 75.290 72.050 75.430 ;
        RECT 72.295 75.290 72.585 75.335 ;
        RECT 71.910 75.150 72.585 75.290 ;
        RECT 72.295 75.105 72.585 75.150 ;
        RECT 73.200 75.090 73.520 75.350 ;
        RECT 73.660 75.290 73.980 75.350 ;
        RECT 74.135 75.290 74.425 75.335 ;
        RECT 86.540 75.290 86.860 75.350 ;
        RECT 73.660 75.150 86.860 75.290 ;
        RECT 73.660 75.090 73.980 75.150 ;
        RECT 74.135 75.105 74.425 75.150 ;
        RECT 86.540 75.090 86.860 75.150 ;
        RECT 87.460 75.090 87.780 75.350 ;
        RECT 19.380 74.950 19.700 75.010 ;
        RECT 19.855 74.950 20.145 74.995 ;
        RECT 19.380 74.810 20.145 74.950 ;
        RECT 19.380 74.750 19.700 74.810 ;
        RECT 19.855 74.765 20.145 74.810 ;
        RECT 26.740 74.950 27.060 75.010 ;
        RECT 28.900 74.950 29.190 74.995 ;
        RECT 36.400 74.950 36.720 75.010 ;
        RECT 61.410 74.950 61.700 74.995 ;
        RECT 66.775 74.950 67.065 74.995 ;
        RECT 26.740 74.810 29.190 74.950 ;
        RECT 26.740 74.750 27.060 74.810 ;
        RECT 28.900 74.765 29.190 74.810 ;
        RECT 34.650 74.810 54.800 74.950 ;
        RECT 20.760 74.410 21.080 74.670 ;
        RECT 24.440 74.410 24.760 74.670 ;
        RECT 34.650 74.655 34.790 74.810 ;
        RECT 36.400 74.750 36.720 74.810 ;
        RECT 34.575 74.425 34.865 74.655 ;
        RECT 42.855 74.610 43.145 74.655 ;
        RECT 45.155 74.610 45.445 74.655 ;
        RECT 42.855 74.470 45.445 74.610 ;
        RECT 42.855 74.425 43.145 74.470 ;
        RECT 45.155 74.425 45.445 74.470 ;
        RECT 46.980 74.410 47.300 74.670 ;
        RECT 52.960 74.410 53.280 74.670 ;
        RECT 54.660 74.610 54.800 74.810 ;
        RECT 61.410 74.810 67.065 74.950 ;
        RECT 61.410 74.765 61.700 74.810 ;
        RECT 66.775 74.765 67.065 74.810 ;
        RECT 69.060 74.950 69.380 75.010 ;
        RECT 71.820 74.950 72.140 75.010 ;
        RECT 79.640 74.950 79.960 75.010 ;
        RECT 81.480 74.995 81.800 75.010 ;
        RECT 69.060 74.810 72.140 74.950 ;
        RECT 69.060 74.750 69.380 74.810 ;
        RECT 71.820 74.750 72.140 74.810 ;
        RECT 72.830 74.810 79.960 74.950 ;
        RECT 72.830 74.670 72.970 74.810 ;
        RECT 79.640 74.750 79.960 74.810 ;
        RECT 81.450 74.765 81.800 74.995 ;
        RECT 117.630 74.950 128.990 75.520 ;
        RECT 81.480 74.750 81.800 74.765 ;
        RECT 117.600 74.770 128.990 74.950 ;
        RECT 134.410 76.460 135.180 77.340 ;
        RECT 134.410 76.240 134.810 76.460 ;
        RECT 134.950 76.390 135.180 76.460 ;
        RECT 135.390 77.330 135.620 77.390 ;
        RECT 135.830 77.330 136.050 79.950 ;
        RECT 136.330 79.895 136.770 80.130 ;
        RECT 137.020 79.895 137.250 83.750 ;
        RECT 137.500 80.070 137.730 83.895 ;
        RECT 137.890 83.760 138.210 83.895 ;
        RECT 137.390 79.895 137.730 80.070 ;
        RECT 137.980 79.895 138.210 83.760 ;
        RECT 138.460 80.090 138.690 83.895 ;
        RECT 138.380 80.040 138.690 80.090 ;
        RECT 138.350 79.895 138.690 80.040 ;
        RECT 138.940 79.895 139.170 83.895 ;
        RECT 136.330 79.880 136.620 79.895 ;
        RECT 137.390 79.890 137.600 79.895 ;
        RECT 138.350 79.890 138.550 79.895 ;
        RECT 136.330 79.200 136.590 79.880 ;
        RECT 136.730 79.410 137.060 79.740 ;
        RECT 137.390 79.230 137.550 79.890 ;
        RECT 137.690 79.410 138.020 79.740 ;
        RECT 138.350 79.260 138.510 79.890 ;
        RECT 138.650 79.410 138.980 79.740 ;
        RECT 136.330 79.190 136.620 79.200 ;
        RECT 137.390 79.190 137.600 79.230 ;
        RECT 138.350 79.190 138.550 79.260 ;
        RECT 136.330 79.050 138.550 79.190 ;
        RECT 139.410 79.140 139.700 83.960 ;
        RECT 135.390 77.050 136.050 77.330 ;
        RECT 136.320 79.020 138.550 79.050 ;
        RECT 136.320 78.540 138.520 79.020 ;
        RECT 136.320 78.190 138.790 78.540 ;
        RECT 136.320 78.100 138.800 78.190 ;
        RECT 138.940 78.140 139.940 79.140 ;
        RECT 136.320 77.390 136.730 78.100 ;
        RECT 137.200 77.550 137.530 77.880 ;
        RECT 137.680 77.530 137.850 78.100 ;
        RECT 138.470 78.090 138.800 78.100 ;
        RECT 138.160 77.550 138.490 77.880 ;
        RECT 138.650 77.530 138.800 78.090 ;
        RECT 137.680 77.390 137.820 77.530 ;
        RECT 138.650 77.390 138.790 77.530 ;
        RECT 136.320 77.150 136.760 77.390 ;
        RECT 135.390 76.450 136.020 77.050 ;
        RECT 135.390 76.390 135.620 76.450 ;
        RECT 136.530 76.390 136.760 77.150 ;
        RECT 137.010 76.560 137.240 77.390 ;
        RECT 137.490 77.160 137.820 77.390 ;
        RECT 137.010 76.390 137.340 76.560 ;
        RECT 137.490 76.390 137.720 77.160 ;
        RECT 137.970 76.620 138.200 77.390 ;
        RECT 138.450 77.170 138.790 77.390 ;
        RECT 138.930 77.310 139.160 77.390 ;
        RECT 139.410 77.310 139.700 78.140 ;
        RECT 137.970 76.390 138.310 76.620 ;
        RECT 138.450 76.390 138.680 77.170 ;
        RECT 138.930 76.390 139.700 77.310 ;
        RECT 134.410 75.700 134.900 76.240 ;
        RECT 135.110 76.020 135.460 76.230 ;
        RECT 135.120 75.960 135.460 76.020 ;
        RECT 136.720 75.910 137.050 76.240 ;
        RECT 137.200 75.750 137.340 76.390 ;
        RECT 138.150 76.240 138.310 76.390 ;
        RECT 137.680 75.910 138.010 76.240 ;
        RECT 138.150 75.750 138.320 76.240 ;
        RECT 138.640 75.910 138.970 76.240 ;
        RECT 139.110 75.750 139.700 76.390 ;
        RECT 134.410 75.680 135.410 75.700 ;
        RECT 134.410 75.250 136.210 75.680 ;
        RECT 136.430 75.550 139.700 75.750 ;
        RECT 136.430 75.540 139.260 75.550 ;
        RECT 136.430 75.390 139.180 75.540 ;
        RECT 139.440 75.250 139.700 75.290 ;
        RECT 117.600 74.690 128.980 74.770 ;
        RECT 134.410 74.700 139.700 75.250 ;
        RECT 134.420 74.690 139.700 74.700 ;
        RECT 72.280 74.610 72.600 74.670 ;
        RECT 54.660 74.470 72.600 74.610 ;
        RECT 72.280 74.410 72.600 74.470 ;
        RECT 72.740 74.410 73.060 74.670 ;
        RECT 74.120 74.610 74.440 74.670 ;
        RECT 75.055 74.610 75.345 74.655 ;
        RECT 80.560 74.610 80.880 74.670 ;
        RECT 74.120 74.470 80.880 74.610 ;
        RECT 74.120 74.410 74.440 74.470 ;
        RECT 75.055 74.425 75.345 74.470 ;
        RECT 80.560 74.410 80.880 74.470 ;
        RECT 88.380 74.410 88.700 74.670 ;
        RECT 11.950 73.790 90.610 74.270 ;
        RECT 16.175 73.590 16.465 73.635 ;
        RECT 21.220 73.590 21.540 73.650 ;
        RECT 24.915 73.590 25.205 73.635 ;
        RECT 26.280 73.590 26.600 73.650 ;
        RECT 16.175 73.450 26.600 73.590 ;
        RECT 16.175 73.405 16.465 73.450 ;
        RECT 21.220 73.390 21.540 73.450 ;
        RECT 24.915 73.405 25.205 73.450 ;
        RECT 26.280 73.390 26.600 73.450 ;
        RECT 26.740 73.390 27.060 73.650 ;
        RECT 57.560 73.590 57.880 73.650 ;
        RECT 39.250 73.450 57.880 73.590 ;
        RECT 20.300 73.250 20.620 73.310 ;
        RECT 25.360 73.250 25.680 73.310 ;
        RECT 30.895 73.250 31.185 73.295 ;
        RECT 20.300 73.110 31.185 73.250 ;
        RECT 20.300 73.050 20.620 73.110 ;
        RECT 25.360 73.050 25.680 73.110 ;
        RECT 30.895 73.065 31.185 73.110 ;
        RECT 38.240 73.250 38.560 73.310 ;
        RECT 39.250 73.295 39.390 73.450 ;
        RECT 57.560 73.390 57.880 73.450 ;
        RECT 65.840 73.590 66.160 73.650 ;
        RECT 67.235 73.590 67.525 73.635 ;
        RECT 65.840 73.450 67.525 73.590 ;
        RECT 65.840 73.390 66.160 73.450 ;
        RECT 67.235 73.405 67.525 73.450 ;
        RECT 68.600 73.390 68.920 73.650 ;
        RECT 69.060 73.390 69.380 73.650 ;
        RECT 69.520 73.390 69.840 73.650 ;
        RECT 72.280 73.590 72.600 73.650 ;
        RECT 72.280 73.450 72.970 73.590 ;
        RECT 72.280 73.390 72.600 73.450 ;
        RECT 39.175 73.250 39.465 73.295 ;
        RECT 38.240 73.110 39.465 73.250 ;
        RECT 38.240 73.050 38.560 73.110 ;
        RECT 39.175 73.065 39.465 73.110 ;
        RECT 39.620 73.250 39.940 73.310 ;
        RECT 41.000 73.250 41.320 73.310 ;
        RECT 42.855 73.250 43.145 73.295 ;
        RECT 39.620 73.110 43.145 73.250 ;
        RECT 39.620 73.050 39.940 73.110 ;
        RECT 41.000 73.050 41.320 73.110 ;
        RECT 42.855 73.065 43.145 73.110 ;
        RECT 52.040 73.250 52.360 73.310 ;
        RECT 64.920 73.250 65.240 73.310 ;
        RECT 68.690 73.250 68.830 73.390 ;
        RECT 52.040 73.110 61.930 73.250 ;
        RECT 15.715 72.725 16.005 72.955 ;
        RECT 15.790 72.230 15.930 72.725 ;
        RECT 19.840 72.710 20.160 72.970 ;
        RECT 21.220 72.910 21.540 72.970 ;
        RECT 20.390 72.770 21.540 72.910 ;
        RECT 16.620 72.370 16.940 72.630 ;
        RECT 20.390 72.615 20.530 72.770 ;
        RECT 21.220 72.710 21.540 72.770 ;
        RECT 27.215 72.910 27.505 72.955 ;
        RECT 38.330 72.910 38.470 73.050 ;
        RECT 27.215 72.770 38.470 72.910 ;
        RECT 42.930 72.910 43.070 73.065 ;
        RECT 52.040 73.050 52.360 73.110 ;
        RECT 46.995 72.910 47.285 72.955 ;
        RECT 42.930 72.770 47.285 72.910 ;
        RECT 27.215 72.725 27.505 72.770 ;
        RECT 46.995 72.725 47.285 72.770 ;
        RECT 48.330 72.910 48.620 72.955 ;
        RECT 48.330 72.770 54.570 72.910 ;
        RECT 48.330 72.725 48.620 72.770 ;
        RECT 20.315 72.385 20.605 72.615 ;
        RECT 20.760 72.370 21.080 72.630 ;
        RECT 23.520 72.370 23.840 72.630 ;
        RECT 24.455 72.570 24.745 72.615 ;
        RECT 36.400 72.570 36.720 72.630 ;
        RECT 24.455 72.430 36.720 72.570 ;
        RECT 24.455 72.385 24.745 72.430 ;
        RECT 36.400 72.370 36.720 72.430 ;
        RECT 47.875 72.570 48.165 72.615 ;
        RECT 49.065 72.570 49.355 72.615 ;
        RECT 51.585 72.570 51.875 72.615 ;
        RECT 47.875 72.430 51.875 72.570 ;
        RECT 47.875 72.385 48.165 72.430 ;
        RECT 49.065 72.385 49.355 72.430 ;
        RECT 51.585 72.385 51.875 72.430 ;
        RECT 52.040 72.570 52.360 72.630 ;
        RECT 52.040 72.430 54.110 72.570 ;
        RECT 52.040 72.370 52.360 72.430 ;
        RECT 19.380 72.230 19.700 72.290 ;
        RECT 53.970 72.275 54.110 72.430 ;
        RECT 54.430 72.275 54.570 72.770 ;
        RECT 56.180 72.710 56.500 72.970 ;
        RECT 61.790 72.955 61.930 73.110 ;
        RECT 64.920 73.110 68.830 73.250 ;
        RECT 64.920 73.050 65.240 73.110 ;
        RECT 56.655 72.910 56.945 72.955 ;
        RECT 58.495 72.910 58.785 72.955 ;
        RECT 56.655 72.770 58.785 72.910 ;
        RECT 56.655 72.725 56.945 72.770 ;
        RECT 58.495 72.725 58.785 72.770 ;
        RECT 61.715 72.725 62.005 72.955 ;
        RECT 62.620 72.910 62.940 72.970 ;
        RECT 64.475 72.910 64.765 72.955 ;
        RECT 62.620 72.770 64.765 72.910 ;
        RECT 62.620 72.710 62.940 72.770 ;
        RECT 64.475 72.725 64.765 72.770 ;
        RECT 67.220 72.710 67.540 72.970 ;
        RECT 68.230 72.955 68.370 73.110 ;
        RECT 68.155 72.725 68.445 72.955 ;
        RECT 68.600 72.710 68.920 72.970 ;
        RECT 69.610 72.955 69.750 73.390 ;
        RECT 70.960 73.110 71.590 73.250 ;
        RECT 70.960 72.955 71.100 73.110 ;
        RECT 69.535 72.910 69.825 72.955 ;
        RECT 69.150 72.770 69.825 72.910 ;
        RECT 57.115 72.385 57.405 72.615 ;
        RECT 47.480 72.230 47.770 72.275 ;
        RECT 49.580 72.230 49.870 72.275 ;
        RECT 51.150 72.230 51.440 72.275 ;
        RECT 15.790 72.090 20.300 72.230 ;
        RECT 19.380 72.030 19.700 72.090 ;
        RECT 13.860 71.690 14.180 71.950 ;
        RECT 17.540 71.890 17.860 71.950 ;
        RECT 18.015 71.890 18.305 71.935 ;
        RECT 17.540 71.750 18.305 71.890 ;
        RECT 20.160 71.890 20.300 72.090 ;
        RECT 47.480 72.090 51.440 72.230 ;
        RECT 47.480 72.045 47.770 72.090 ;
        RECT 49.580 72.045 49.870 72.090 ;
        RECT 51.150 72.045 51.440 72.090 ;
        RECT 53.895 72.045 54.185 72.275 ;
        RECT 54.355 72.045 54.645 72.275 ;
        RECT 54.800 72.230 55.120 72.290 ;
        RECT 57.190 72.230 57.330 72.385 ;
        RECT 69.150 72.290 69.290 72.770 ;
        RECT 69.535 72.725 69.825 72.770 ;
        RECT 70.025 72.725 70.315 72.955 ;
        RECT 70.885 72.725 71.175 72.955 ;
        RECT 54.800 72.090 57.330 72.230 ;
        RECT 54.800 72.030 55.120 72.090 ;
        RECT 69.060 72.030 69.380 72.290 ;
        RECT 70.075 72.230 70.215 72.725 ;
        RECT 71.450 72.570 71.590 73.110 ;
        RECT 72.280 72.710 72.600 72.970 ;
        RECT 72.830 72.925 72.970 73.450 ;
        RECT 75.055 73.405 75.345 73.635 ;
        RECT 75.500 73.590 75.820 73.650 ;
        RECT 78.720 73.590 79.040 73.650 ;
        RECT 75.500 73.450 79.040 73.590 ;
        RECT 73.215 73.250 73.505 73.295 ;
        RECT 74.580 73.250 74.900 73.310 ;
        RECT 73.215 73.110 74.900 73.250 ;
        RECT 75.130 73.250 75.270 73.405 ;
        RECT 75.500 73.390 75.820 73.450 ;
        RECT 78.720 73.390 79.040 73.450 ;
        RECT 81.480 73.390 81.800 73.650 ;
        RECT 83.795 73.250 84.085 73.295 ;
        RECT 75.130 73.110 84.085 73.250 ;
        RECT 73.215 73.065 73.505 73.110 ;
        RECT 74.580 73.050 74.900 73.110 ;
        RECT 83.795 73.065 84.085 73.110 ;
        RECT 72.830 72.910 73.430 72.925 ;
        RECT 73.675 72.910 73.965 72.955 ;
        RECT 72.830 72.785 73.965 72.910 ;
        RECT 73.290 72.770 73.965 72.785 ;
        RECT 73.675 72.725 73.965 72.770 ;
        RECT 74.135 72.725 74.425 72.955 ;
        RECT 75.515 72.910 75.805 72.955 ;
        RECT 75.960 72.910 76.280 72.970 ;
        RECT 75.515 72.770 76.280 72.910 ;
        RECT 75.515 72.725 75.805 72.770 ;
        RECT 72.740 72.570 73.060 72.630 ;
        RECT 71.450 72.430 73.060 72.570 ;
        RECT 74.210 72.570 74.350 72.725 ;
        RECT 75.960 72.710 76.280 72.770 ;
        RECT 76.420 72.710 76.740 72.970 ;
        RECT 76.895 72.725 77.185 72.955 ;
        RECT 77.355 72.910 77.645 72.955 ;
        RECT 77.800 72.910 78.120 72.970 ;
        RECT 77.355 72.770 78.120 72.910 ;
        RECT 77.355 72.725 77.645 72.770 ;
        RECT 74.580 72.570 74.900 72.630 ;
        RECT 74.210 72.430 74.900 72.570 ;
        RECT 76.970 72.570 77.110 72.725 ;
        RECT 77.800 72.710 78.120 72.770 ;
        RECT 83.335 72.910 83.625 72.955 ;
        RECT 85.635 72.910 85.925 72.955 ;
        RECT 83.335 72.770 85.925 72.910 ;
        RECT 83.335 72.725 83.625 72.770 ;
        RECT 85.635 72.725 85.925 72.770 ;
        RECT 87.000 72.910 87.320 72.970 ;
        RECT 88.395 72.910 88.685 72.955 ;
        RECT 87.000 72.770 88.685 72.910 ;
        RECT 87.000 72.710 87.320 72.770 ;
        RECT 88.395 72.725 88.685 72.770 ;
        RECT 78.260 72.570 78.580 72.630 ;
        RECT 76.970 72.430 78.580 72.570 ;
        RECT 72.740 72.370 73.060 72.430 ;
        RECT 74.580 72.370 74.900 72.430 ;
        RECT 78.260 72.370 78.580 72.430 ;
        RECT 84.255 72.385 84.545 72.615 ;
        RECT 78.735 72.230 79.025 72.275 ;
        RECT 84.330 72.230 84.470 72.385 ;
        RECT 70.075 72.090 71.590 72.230 ;
        RECT 65.380 71.890 65.700 71.950 ;
        RECT 20.160 71.750 65.700 71.890 ;
        RECT 17.540 71.690 17.860 71.750 ;
        RECT 18.015 71.705 18.305 71.750 ;
        RECT 65.380 71.690 65.700 71.750 ;
        RECT 70.900 71.690 71.220 71.950 ;
        RECT 71.450 71.890 71.590 72.090 ;
        RECT 78.735 72.090 84.470 72.230 ;
        RECT 78.735 72.045 79.025 72.090 ;
        RECT 74.120 71.890 74.440 71.950 ;
        RECT 71.450 71.750 74.440 71.890 ;
        RECT 74.120 71.690 74.440 71.750 ;
        RECT 11.950 71.070 90.610 71.550 ;
        RECT 18.000 70.870 18.320 70.930 ;
        RECT 19.380 70.870 19.700 70.930 ;
        RECT 20.315 70.870 20.605 70.915 ;
        RECT 18.000 70.730 20.605 70.870 ;
        RECT 18.000 70.670 18.320 70.730 ;
        RECT 19.380 70.670 19.700 70.730 ;
        RECT 20.315 70.685 20.605 70.730 ;
        RECT 72.280 70.670 72.600 70.930 ;
        RECT 74.120 70.670 74.440 70.930 ;
        RECT 75.055 70.870 75.345 70.915 ;
        RECT 76.420 70.870 76.740 70.930 ;
        RECT 75.055 70.730 76.740 70.870 ;
        RECT 75.055 70.685 75.345 70.730 ;
        RECT 76.420 70.670 76.740 70.730 ;
        RECT 13.900 70.530 14.190 70.575 ;
        RECT 16.000 70.530 16.290 70.575 ;
        RECT 17.570 70.530 17.860 70.575 ;
        RECT 13.900 70.390 17.860 70.530 ;
        RECT 13.900 70.345 14.190 70.390 ;
        RECT 16.000 70.345 16.290 70.390 ;
        RECT 17.570 70.345 17.860 70.390 ;
        RECT 19.840 70.530 20.160 70.590 ;
        RECT 23.520 70.530 23.840 70.590 ;
        RECT 19.840 70.390 23.840 70.530 ;
        RECT 19.840 70.330 20.160 70.390 ;
        RECT 23.520 70.330 23.840 70.390 ;
        RECT 25.860 70.530 26.150 70.575 ;
        RECT 27.960 70.530 28.250 70.575 ;
        RECT 29.530 70.530 29.820 70.575 ;
        RECT 25.860 70.390 29.820 70.530 ;
        RECT 25.860 70.345 26.150 70.390 ;
        RECT 27.960 70.345 28.250 70.390 ;
        RECT 29.530 70.345 29.820 70.390 ;
        RECT 39.660 70.530 39.950 70.575 ;
        RECT 41.760 70.530 42.050 70.575 ;
        RECT 43.330 70.530 43.620 70.575 ;
        RECT 39.660 70.390 43.620 70.530 ;
        RECT 39.660 70.345 39.950 70.390 ;
        RECT 41.760 70.345 42.050 70.390 ;
        RECT 43.330 70.345 43.620 70.390 ;
        RECT 46.075 70.530 46.365 70.575 ;
        RECT 70.900 70.530 71.220 70.590 ;
        RECT 72.740 70.530 73.060 70.590 ;
        RECT 74.210 70.530 74.350 70.670 ;
        RECT 46.075 70.390 54.110 70.530 ;
        RECT 46.075 70.345 46.365 70.390 ;
        RECT 53.970 70.250 54.110 70.390 ;
        RECT 70.900 70.390 74.350 70.530 ;
        RECT 75.500 70.530 75.820 70.590 ;
        RECT 77.800 70.530 78.120 70.590 ;
        RECT 75.500 70.390 78.120 70.530 ;
        RECT 70.900 70.330 71.220 70.390 ;
        RECT 72.740 70.330 73.060 70.390 ;
        RECT 75.500 70.330 75.820 70.390 ;
        RECT 77.800 70.330 78.120 70.390 ;
        RECT 14.295 70.190 14.585 70.235 ;
        RECT 15.485 70.190 15.775 70.235 ;
        RECT 18.005 70.190 18.295 70.235 ;
        RECT 14.295 70.050 18.295 70.190 ;
        RECT 14.295 70.005 14.585 70.050 ;
        RECT 15.485 70.005 15.775 70.050 ;
        RECT 18.005 70.005 18.295 70.050 ;
        RECT 25.360 69.990 25.680 70.250 ;
        RECT 26.255 70.190 26.545 70.235 ;
        RECT 27.445 70.190 27.735 70.235 ;
        RECT 29.965 70.190 30.255 70.235 ;
        RECT 26.255 70.050 30.255 70.190 ;
        RECT 26.255 70.005 26.545 70.050 ;
        RECT 27.445 70.005 27.735 70.050 ;
        RECT 29.965 70.005 30.255 70.050 ;
        RECT 38.255 70.190 38.545 70.235 ;
        RECT 40.055 70.190 40.345 70.235 ;
        RECT 41.245 70.190 41.535 70.235 ;
        RECT 43.765 70.190 44.055 70.235 ;
        RECT 38.255 70.050 38.930 70.190 ;
        RECT 38.255 70.005 38.545 70.050 ;
        RECT 13.415 69.850 13.705 69.895 ;
        RECT 20.300 69.850 20.620 69.910 ;
        RECT 13.415 69.710 20.620 69.850 ;
        RECT 13.415 69.665 13.705 69.710 ;
        RECT 20.300 69.650 20.620 69.710 ;
        RECT 13.860 69.510 14.180 69.570 ;
        RECT 14.640 69.510 14.930 69.555 ;
        RECT 13.860 69.370 14.930 69.510 ;
        RECT 13.860 69.310 14.180 69.370 ;
        RECT 14.640 69.325 14.930 69.370 ;
        RECT 26.710 69.510 27.000 69.555 ;
        RECT 27.660 69.510 27.980 69.570 ;
        RECT 26.710 69.370 27.980 69.510 ;
        RECT 38.790 69.510 38.930 70.050 ;
        RECT 40.055 70.050 44.055 70.190 ;
        RECT 40.055 70.005 40.345 70.050 ;
        RECT 41.245 70.005 41.535 70.050 ;
        RECT 43.765 70.005 44.055 70.050 ;
        RECT 49.755 70.190 50.045 70.235 ;
        RECT 50.660 70.190 50.980 70.250 ;
        RECT 49.755 70.050 50.980 70.190 ;
        RECT 49.755 70.005 50.045 70.050 ;
        RECT 50.660 69.990 50.980 70.050 ;
        RECT 53.880 69.990 54.200 70.250 ;
        RECT 62.620 70.190 62.940 70.250 ;
        RECT 63.095 70.190 63.385 70.235 ;
        RECT 62.620 70.050 63.385 70.190 ;
        RECT 62.620 69.990 62.940 70.050 ;
        RECT 63.095 70.005 63.385 70.050 ;
        RECT 66.760 70.190 67.080 70.250 ;
        RECT 68.155 70.190 68.445 70.235 ;
        RECT 66.760 70.050 73.430 70.190 ;
        RECT 66.760 69.990 67.080 70.050 ;
        RECT 68.155 70.005 68.445 70.050 ;
        RECT 39.175 69.850 39.465 69.895 ;
        RECT 39.620 69.850 39.940 69.910 ;
        RECT 47.440 69.850 47.760 69.910 ;
        RECT 39.175 69.710 39.940 69.850 ;
        RECT 39.175 69.665 39.465 69.710 ;
        RECT 39.620 69.650 39.940 69.710 ;
        RECT 40.170 69.710 47.760 69.850 ;
        RECT 40.170 69.510 40.310 69.710 ;
        RECT 47.440 69.650 47.760 69.710 ;
        RECT 57.560 69.850 57.880 69.910 ;
        RECT 59.415 69.850 59.705 69.895 ;
        RECT 64.000 69.850 64.320 69.910 ;
        RECT 57.560 69.710 64.320 69.850 ;
        RECT 57.560 69.650 57.880 69.710 ;
        RECT 59.415 69.665 59.705 69.710 ;
        RECT 64.000 69.650 64.320 69.710 ;
        RECT 64.475 69.665 64.765 69.895 ;
        RECT 38.790 69.370 40.310 69.510 ;
        RECT 40.510 69.510 40.800 69.555 ;
        RECT 55.720 69.510 56.040 69.570 ;
        RECT 64.550 69.510 64.690 69.665 ;
        RECT 69.060 69.650 69.380 69.910 ;
        RECT 69.520 69.850 69.840 69.910 ;
        RECT 70.915 69.850 71.205 69.895 ;
        RECT 69.520 69.710 71.205 69.850 ;
        RECT 69.520 69.650 69.840 69.710 ;
        RECT 70.915 69.665 71.205 69.710 ;
        RECT 71.375 69.665 71.665 69.895 ;
        RECT 40.510 69.370 46.750 69.510 ;
        RECT 26.710 69.325 27.000 69.370 ;
        RECT 27.660 69.310 27.980 69.370 ;
        RECT 40.510 69.325 40.800 69.370 ;
        RECT 32.275 69.170 32.565 69.215 ;
        RECT 32.720 69.170 33.040 69.230 ;
        RECT 32.275 69.030 33.040 69.170 ;
        RECT 32.275 68.985 32.565 69.030 ;
        RECT 32.720 68.970 33.040 69.030 ;
        RECT 35.020 68.970 35.340 69.230 ;
        RECT 36.860 68.970 37.180 69.230 ;
        RECT 37.320 68.970 37.640 69.230 ;
        RECT 46.610 69.215 46.750 69.370 ;
        RECT 55.720 69.370 64.690 69.510 ;
        RECT 65.380 69.510 65.700 69.570 ;
        RECT 69.980 69.510 70.300 69.570 ;
        RECT 71.450 69.510 71.590 69.665 ;
        RECT 71.820 69.650 72.140 69.910 ;
        RECT 73.290 69.895 73.430 70.050 ;
        RECT 73.660 69.990 73.980 70.250 ;
        RECT 78.720 70.190 79.040 70.250 ;
        RECT 78.720 70.050 79.870 70.190 ;
        RECT 78.720 69.990 79.040 70.050 ;
        RECT 72.755 69.665 73.045 69.895 ;
        RECT 73.215 69.665 73.505 69.895 ;
        RECT 65.380 69.370 68.600 69.510 ;
        RECT 55.720 69.310 56.040 69.370 ;
        RECT 65.380 69.310 65.700 69.370 ;
        RECT 46.535 68.985 46.825 69.215 ;
        RECT 48.360 68.970 48.680 69.230 ;
        RECT 48.835 69.170 49.125 69.215 ;
        RECT 51.135 69.170 51.425 69.215 ;
        RECT 48.835 69.030 51.425 69.170 ;
        RECT 48.835 68.985 49.125 69.030 ;
        RECT 51.135 68.985 51.425 69.030 ;
        RECT 65.840 69.170 66.160 69.230 ;
        RECT 67.695 69.170 67.985 69.215 ;
        RECT 65.840 69.030 67.985 69.170 ;
        RECT 68.460 69.170 68.600 69.370 ;
        RECT 69.980 69.370 71.590 69.510 ;
        RECT 72.280 69.510 72.600 69.570 ;
        RECT 72.830 69.510 72.970 69.665 ;
        RECT 73.750 69.510 73.890 69.990 ;
        RECT 77.800 69.650 78.120 69.910 ;
        RECT 79.730 69.895 79.870 70.050 ;
        RECT 79.655 69.665 79.945 69.895 ;
        RECT 85.175 69.850 85.465 69.895 ;
        RECT 86.080 69.850 86.400 69.910 ;
        RECT 85.175 69.710 86.400 69.850 ;
        RECT 85.175 69.665 85.465 69.710 ;
        RECT 86.080 69.650 86.400 69.710 ;
        RECT 88.380 69.650 88.700 69.910 ;
        RECT 72.280 69.370 73.890 69.510 ;
        RECT 77.340 69.510 77.660 69.570 ;
        RECT 78.260 69.510 78.580 69.570 ;
        RECT 78.735 69.510 79.025 69.555 ;
        RECT 77.340 69.370 79.025 69.510 ;
        RECT 69.980 69.310 70.300 69.370 ;
        RECT 72.280 69.310 72.600 69.370 ;
        RECT 77.340 69.310 77.660 69.370 ;
        RECT 78.260 69.310 78.580 69.370 ;
        RECT 78.735 69.325 79.025 69.370 ;
        RECT 79.195 69.510 79.485 69.555 ;
        RECT 81.480 69.510 81.800 69.570 ;
        RECT 79.195 69.370 81.800 69.510 ;
        RECT 79.195 69.325 79.485 69.370 ;
        RECT 79.270 69.170 79.410 69.325 ;
        RECT 81.480 69.310 81.800 69.370 ;
        RECT 68.460 69.030 79.410 69.170 ;
        RECT 80.575 69.170 80.865 69.215 ;
        RECT 83.320 69.170 83.640 69.230 ;
        RECT 80.575 69.030 83.640 69.170 ;
        RECT 65.840 68.970 66.160 69.030 ;
        RECT 67.695 68.985 67.985 69.030 ;
        RECT 80.575 68.985 80.865 69.030 ;
        RECT 83.320 68.970 83.640 69.030 ;
        RECT 84.240 68.970 84.560 69.230 ;
        RECT 85.620 68.970 85.940 69.230 ;
        RECT 11.950 68.350 90.610 68.830 ;
        RECT 12.940 68.150 13.260 68.210 ;
        RECT 13.875 68.150 14.165 68.195 ;
        RECT 12.940 68.010 14.165 68.150 ;
        RECT 12.940 67.950 13.260 68.010 ;
        RECT 13.875 67.965 14.165 68.010 ;
        RECT 14.870 68.010 22.370 68.150 ;
        RECT 14.870 67.515 15.010 68.010 ;
        RECT 20.300 67.810 20.620 67.870 ;
        RECT 16.250 67.670 20.620 67.810 ;
        RECT 16.250 67.515 16.390 67.670 ;
        RECT 20.300 67.610 20.620 67.670 ;
        RECT 17.540 67.515 17.860 67.530 ;
        RECT 14.795 67.285 15.085 67.515 ;
        RECT 16.175 67.285 16.465 67.515 ;
        RECT 17.510 67.470 17.860 67.515 ;
        RECT 17.345 67.330 17.860 67.470 ;
        RECT 22.230 67.470 22.370 68.010 ;
        RECT 23.075 67.965 23.365 68.195 ;
        RECT 25.835 68.150 26.125 68.195 ;
        RECT 26.280 68.150 26.600 68.210 ;
        RECT 25.835 68.010 26.600 68.150 ;
        RECT 25.835 67.965 26.125 68.010 ;
        RECT 23.150 67.810 23.290 67.965 ;
        RECT 26.280 67.950 26.600 68.010 ;
        RECT 27.660 67.950 27.980 68.210 ;
        RECT 36.860 68.150 37.180 68.210 ;
        RECT 38.715 68.150 39.005 68.195 ;
        RECT 36.860 68.010 39.005 68.150 ;
        RECT 36.860 67.950 37.180 68.010 ;
        RECT 38.715 67.965 39.005 68.010 ;
        RECT 41.920 68.150 42.240 68.210 ;
        RECT 46.980 68.150 47.300 68.210 ;
        RECT 41.920 68.010 47.300 68.150 ;
        RECT 41.920 67.950 42.240 68.010 ;
        RECT 46.980 67.950 47.300 68.010 ;
        RECT 51.595 68.150 51.885 68.195 ;
        RECT 52.960 68.150 53.280 68.210 ;
        RECT 51.595 68.010 53.280 68.150 ;
        RECT 51.595 67.965 51.885 68.010 ;
        RECT 52.960 67.950 53.280 68.010 ;
        RECT 53.895 68.150 54.185 68.195 ;
        RECT 55.720 68.150 56.040 68.210 ;
        RECT 53.895 68.010 56.040 68.150 ;
        RECT 53.895 67.965 54.185 68.010 ;
        RECT 55.720 67.950 56.040 68.010 ;
        RECT 64.015 67.965 64.305 68.195 ;
        RECT 23.520 67.810 23.840 67.870 ;
        RECT 61.410 67.810 61.700 67.855 ;
        RECT 64.090 67.810 64.230 67.965 ;
        RECT 65.840 67.950 66.160 68.210 ;
        RECT 73.215 67.965 73.505 68.195 ;
        RECT 76.895 68.150 77.185 68.195 ;
        RECT 85.160 68.150 85.480 68.210 ;
        RECT 76.895 68.010 85.480 68.150 ;
        RECT 76.895 67.965 77.185 68.010 ;
        RECT 23.150 67.670 58.250 67.810 ;
        RECT 23.520 67.610 23.840 67.670 ;
        RECT 22.230 67.330 29.730 67.470 ;
        RECT 17.510 67.285 17.860 67.330 ;
        RECT 17.540 67.270 17.860 67.285 ;
        RECT 17.055 67.130 17.345 67.175 ;
        RECT 18.245 67.130 18.535 67.175 ;
        RECT 20.765 67.130 21.055 67.175 ;
        RECT 17.055 66.990 21.055 67.130 ;
        RECT 17.055 66.945 17.345 66.990 ;
        RECT 18.245 66.945 18.535 66.990 ;
        RECT 20.765 66.945 21.055 66.990 ;
        RECT 24.440 66.930 24.760 67.190 ;
        RECT 25.375 67.130 25.665 67.175 ;
        RECT 26.740 67.130 27.060 67.190 ;
        RECT 25.375 66.990 27.060 67.130 ;
        RECT 29.590 67.130 29.730 67.330 ;
        RECT 41.920 67.270 42.240 67.530 ;
        RECT 42.380 67.270 42.700 67.530 ;
        RECT 42.855 67.470 43.145 67.515 ;
        RECT 43.300 67.470 43.620 67.530 ;
        RECT 42.855 67.330 43.620 67.470 ;
        RECT 42.855 67.285 43.145 67.330 ;
        RECT 43.300 67.270 43.620 67.330 ;
        RECT 43.775 67.285 44.065 67.515 ;
        RECT 44.235 67.470 44.525 67.515 ;
        RECT 47.900 67.470 48.220 67.530 ;
        RECT 44.235 67.330 48.220 67.470 ;
        RECT 44.235 67.285 44.525 67.330 ;
        RECT 29.960 67.130 30.280 67.190 ;
        RECT 43.850 67.130 43.990 67.285 ;
        RECT 47.900 67.270 48.220 67.330 ;
        RECT 53.435 67.470 53.725 67.515 ;
        RECT 57.560 67.470 57.880 67.530 ;
        RECT 53.435 67.330 57.880 67.470 ;
        RECT 58.110 67.470 58.250 67.670 ;
        RECT 61.410 67.670 64.230 67.810 ;
        RECT 64.550 67.670 72.970 67.810 ;
        RECT 61.410 67.625 61.700 67.670 ;
        RECT 64.550 67.470 64.690 67.670 ;
        RECT 58.110 67.330 64.690 67.470 ;
        RECT 66.315 67.470 66.605 67.515 ;
        RECT 67.220 67.470 67.540 67.530 ;
        RECT 69.520 67.470 69.840 67.530 ;
        RECT 66.315 67.330 69.840 67.470 ;
        RECT 53.435 67.285 53.725 67.330 ;
        RECT 57.560 67.270 57.880 67.330 ;
        RECT 66.315 67.285 66.605 67.330 ;
        RECT 67.220 67.270 67.540 67.330 ;
        RECT 69.520 67.270 69.840 67.330 ;
        RECT 70.900 67.470 71.220 67.530 ;
        RECT 71.375 67.470 71.665 67.515 ;
        RECT 70.900 67.330 71.665 67.470 ;
        RECT 70.900 67.270 71.220 67.330 ;
        RECT 71.375 67.285 71.665 67.330 ;
        RECT 72.280 67.270 72.600 67.530 ;
        RECT 29.590 66.990 43.990 67.130 ;
        RECT 25.375 66.945 25.665 66.990 ;
        RECT 26.740 66.930 27.060 66.990 ;
        RECT 29.960 66.930 30.280 66.990 ;
        RECT 46.980 66.930 47.300 67.190 ;
        RECT 49.740 66.930 50.060 67.190 ;
        RECT 54.355 66.945 54.645 67.175 ;
        RECT 58.045 67.130 58.335 67.175 ;
        RECT 60.565 67.130 60.855 67.175 ;
        RECT 61.755 67.130 62.045 67.175 ;
        RECT 58.045 66.990 62.045 67.130 ;
        RECT 58.045 66.945 58.335 66.990 ;
        RECT 60.565 66.945 60.855 66.990 ;
        RECT 61.755 66.945 62.045 66.990 ;
        RECT 62.635 67.130 62.925 67.175 ;
        RECT 63.080 67.130 63.400 67.190 ;
        RECT 62.635 66.990 63.400 67.130 ;
        RECT 62.635 66.945 62.925 66.990 ;
        RECT 16.660 66.790 16.950 66.835 ;
        RECT 18.760 66.790 19.050 66.835 ;
        RECT 20.330 66.790 20.620 66.835 ;
        RECT 16.660 66.650 20.620 66.790 ;
        RECT 16.660 66.605 16.950 66.650 ;
        RECT 18.760 66.605 19.050 66.650 ;
        RECT 20.330 66.605 20.620 66.650 ;
        RECT 45.155 66.790 45.445 66.835 ;
        RECT 51.580 66.790 51.900 66.850 ;
        RECT 45.155 66.650 51.900 66.790 ;
        RECT 45.155 66.605 45.445 66.650 ;
        RECT 51.580 66.590 51.900 66.650 ;
        RECT 18.000 66.450 18.320 66.510 ;
        RECT 19.840 66.450 20.160 66.510 ;
        RECT 18.000 66.310 20.160 66.450 ;
        RECT 18.000 66.250 18.320 66.310 ;
        RECT 19.840 66.250 20.160 66.310 ;
        RECT 46.060 66.450 46.380 66.510 ;
        RECT 54.430 66.450 54.570 66.945 ;
        RECT 63.080 66.930 63.400 66.990 ;
        RECT 66.775 67.130 67.065 67.175 ;
        RECT 68.140 67.130 68.460 67.190 ;
        RECT 66.775 66.990 68.460 67.130 ;
        RECT 72.830 67.130 72.970 67.670 ;
        RECT 73.290 67.470 73.430 67.965 ;
        RECT 85.160 67.950 85.480 68.010 ;
        RECT 87.000 68.150 87.320 68.210 ;
        RECT 87.475 68.150 87.765 68.195 ;
        RECT 88.380 68.150 88.700 68.210 ;
        RECT 87.000 68.010 88.700 68.150 ;
        RECT 87.000 67.950 87.320 68.010 ;
        RECT 87.475 67.965 87.765 68.010 ;
        RECT 88.380 67.950 88.700 68.010 ;
        RECT 75.960 67.810 76.280 67.870 ;
        RECT 74.670 67.670 76.280 67.810 ;
        RECT 74.670 67.515 74.810 67.670 ;
        RECT 75.960 67.610 76.280 67.670 ;
        RECT 78.260 67.610 78.580 67.870 ;
        RECT 81.910 67.810 82.200 67.855 ;
        RECT 82.400 67.810 82.720 67.870 ;
        RECT 81.910 67.670 82.720 67.810 ;
        RECT 81.910 67.625 82.200 67.670 ;
        RECT 82.400 67.610 82.720 67.670 ;
        RECT 73.675 67.470 73.965 67.515 ;
        RECT 73.290 67.330 73.965 67.470 ;
        RECT 73.675 67.285 73.965 67.330 ;
        RECT 74.595 67.285 74.885 67.515 ;
        RECT 75.040 67.270 75.360 67.530 ;
        RECT 75.500 67.270 75.820 67.530 ;
        RECT 77.340 67.270 77.660 67.530 ;
        RECT 78.735 67.285 79.025 67.515 ;
        RECT 78.810 67.130 78.950 67.285 ;
        RECT 79.180 67.270 79.500 67.530 ;
        RECT 80.100 67.470 80.420 67.530 ;
        RECT 80.575 67.470 80.865 67.515 ;
        RECT 80.100 67.330 80.865 67.470 ;
        RECT 80.100 67.270 80.420 67.330 ;
        RECT 80.575 67.285 80.865 67.330 ;
        RECT 81.020 67.270 81.340 67.530 ;
        RECT 88.840 67.270 89.160 67.530 ;
        RECT 81.110 67.130 81.250 67.270 ;
        RECT 72.830 66.990 81.250 67.130 ;
        RECT 81.455 67.130 81.745 67.175 ;
        RECT 82.645 67.130 82.935 67.175 ;
        RECT 85.165 67.130 85.455 67.175 ;
        RECT 81.455 66.990 85.455 67.130 ;
        RECT 66.775 66.945 67.065 66.990 ;
        RECT 68.140 66.930 68.460 66.990 ;
        RECT 81.455 66.945 81.745 66.990 ;
        RECT 82.645 66.945 82.935 66.990 ;
        RECT 85.165 66.945 85.455 66.990 ;
        RECT 58.480 66.790 58.770 66.835 ;
        RECT 60.050 66.790 60.340 66.835 ;
        RECT 62.150 66.790 62.440 66.835 ;
        RECT 58.480 66.650 62.440 66.790 ;
        RECT 58.480 66.605 58.770 66.650 ;
        RECT 60.050 66.605 60.340 66.650 ;
        RECT 62.150 66.605 62.440 66.650 ;
        RECT 70.440 66.790 70.760 66.850 ;
        RECT 75.040 66.790 75.360 66.850 ;
        RECT 70.440 66.650 75.360 66.790 ;
        RECT 70.440 66.590 70.760 66.650 ;
        RECT 75.040 66.590 75.360 66.650 ;
        RECT 75.960 66.790 76.280 66.850 ;
        RECT 79.180 66.790 79.500 66.850 ;
        RECT 75.960 66.650 79.500 66.790 ;
        RECT 75.960 66.590 76.280 66.650 ;
        RECT 79.180 66.590 79.500 66.650 ;
        RECT 81.060 66.790 81.350 66.835 ;
        RECT 83.160 66.790 83.450 66.835 ;
        RECT 84.730 66.790 85.020 66.835 ;
        RECT 81.060 66.650 85.020 66.790 ;
        RECT 81.060 66.605 81.350 66.650 ;
        RECT 83.160 66.605 83.450 66.650 ;
        RECT 84.730 66.605 85.020 66.650 ;
        RECT 86.540 66.790 86.860 66.850 ;
        RECT 87.935 66.790 88.225 66.835 ;
        RECT 86.540 66.650 88.225 66.790 ;
        RECT 86.540 66.590 86.860 66.650 ;
        RECT 87.935 66.605 88.225 66.650 ;
        RECT 57.100 66.450 57.420 66.510 ;
        RECT 58.940 66.450 59.260 66.510 ;
        RECT 46.060 66.310 59.260 66.450 ;
        RECT 46.060 66.250 46.380 66.310 ;
        RECT 57.100 66.250 57.420 66.310 ;
        RECT 58.940 66.250 59.260 66.310 ;
        RECT 71.360 66.250 71.680 66.510 ;
        RECT 80.115 66.450 80.405 66.495 ;
        RECT 84.240 66.450 84.560 66.510 ;
        RECT 80.115 66.310 84.560 66.450 ;
        RECT 80.115 66.265 80.405 66.310 ;
        RECT 84.240 66.250 84.560 66.310 ;
        RECT 11.950 65.630 90.610 66.110 ;
        RECT 26.740 65.430 27.060 65.490 ;
        RECT 32.720 65.430 33.040 65.490 ;
        RECT 39.160 65.430 39.480 65.490 ;
        RECT 26.740 65.290 39.480 65.430 ;
        RECT 26.740 65.230 27.060 65.290 ;
        RECT 32.720 65.230 33.040 65.290 ;
        RECT 39.160 65.230 39.480 65.290 ;
        RECT 40.095 65.430 40.385 65.475 ;
        RECT 41.920 65.430 42.240 65.490 ;
        RECT 40.095 65.290 42.240 65.430 ;
        RECT 40.095 65.245 40.385 65.290 ;
        RECT 41.920 65.230 42.240 65.290 ;
        RECT 47.900 65.430 48.220 65.490 ;
        RECT 48.820 65.430 49.140 65.490 ;
        RECT 47.900 65.290 49.140 65.430 ;
        RECT 47.900 65.230 48.220 65.290 ;
        RECT 48.820 65.230 49.140 65.290 ;
        RECT 58.020 65.230 58.340 65.490 ;
        RECT 75.975 65.430 76.265 65.475 ;
        RECT 77.340 65.430 77.660 65.490 ;
        RECT 75.975 65.290 77.660 65.430 ;
        RECT 75.975 65.245 76.265 65.290 ;
        RECT 77.340 65.230 77.660 65.290 ;
        RECT 82.400 65.230 82.720 65.490 ;
        RECT 33.180 65.090 33.500 65.150 ;
        RECT 16.710 64.950 33.500 65.090 ;
        RECT 14.780 64.210 15.100 64.470 ;
        RECT 16.710 64.455 16.850 64.950 ;
        RECT 33.180 64.890 33.500 64.950 ;
        RECT 33.680 65.090 33.970 65.135 ;
        RECT 35.780 65.090 36.070 65.135 ;
        RECT 37.350 65.090 37.640 65.135 ;
        RECT 33.680 64.950 37.640 65.090 ;
        RECT 33.680 64.905 33.970 64.950 ;
        RECT 35.780 64.905 36.070 64.950 ;
        RECT 37.350 64.905 37.640 64.950 ;
        RECT 51.620 65.090 51.910 65.135 ;
        RECT 53.720 65.090 54.010 65.135 ;
        RECT 55.290 65.090 55.580 65.135 ;
        RECT 51.620 64.950 55.580 65.090 ;
        RECT 51.620 64.905 51.910 64.950 ;
        RECT 53.720 64.905 54.010 64.950 ;
        RECT 55.290 64.905 55.580 64.950 ;
        RECT 25.820 64.750 26.140 64.810 ;
        RECT 34.075 64.750 34.365 64.795 ;
        RECT 35.265 64.750 35.555 64.795 ;
        RECT 37.785 64.750 38.075 64.795 ;
        RECT 25.820 64.610 26.970 64.750 ;
        RECT 25.820 64.550 26.140 64.610 ;
        RECT 16.635 64.225 16.925 64.455 ;
        RECT 19.855 64.410 20.145 64.455 ;
        RECT 21.220 64.410 21.540 64.470 ;
        RECT 26.830 64.455 26.970 64.610 ;
        RECT 34.075 64.610 38.075 64.750 ;
        RECT 34.075 64.565 34.365 64.610 ;
        RECT 35.265 64.565 35.555 64.610 ;
        RECT 37.785 64.565 38.075 64.610 ;
        RECT 46.535 64.750 46.825 64.795 ;
        RECT 47.440 64.750 47.760 64.810 ;
        RECT 46.535 64.610 47.760 64.750 ;
        RECT 46.535 64.565 46.825 64.610 ;
        RECT 47.440 64.550 47.760 64.610 ;
        RECT 51.120 64.550 51.440 64.810 ;
        RECT 52.015 64.750 52.305 64.795 ;
        RECT 53.205 64.750 53.495 64.795 ;
        RECT 55.725 64.750 56.015 64.795 ;
        RECT 52.015 64.610 56.015 64.750 ;
        RECT 58.110 64.750 58.250 65.230 ;
        RECT 88.380 64.890 88.700 65.150 ;
        RECT 61.255 64.750 61.545 64.795 ;
        RECT 58.110 64.610 61.545 64.750 ;
        RECT 52.015 64.565 52.305 64.610 ;
        RECT 53.205 64.565 53.495 64.610 ;
        RECT 55.725 64.565 56.015 64.610 ;
        RECT 61.255 64.565 61.545 64.610 ;
        RECT 65.855 64.750 66.145 64.795 ;
        RECT 66.300 64.750 66.620 64.810 ;
        RECT 69.060 64.750 69.380 64.810 ;
        RECT 72.280 64.750 72.600 64.810 ;
        RECT 65.855 64.610 66.620 64.750 ;
        RECT 65.855 64.565 66.145 64.610 ;
        RECT 66.300 64.550 66.620 64.610 ;
        RECT 67.310 64.610 72.600 64.750 ;
        RECT 19.855 64.270 21.540 64.410 ;
        RECT 19.855 64.225 20.145 64.270 ;
        RECT 21.220 64.210 21.540 64.270 ;
        RECT 26.755 64.225 27.045 64.455 ;
        RECT 27.215 64.225 27.505 64.455 ;
        RECT 27.675 64.225 27.965 64.455 ;
        RECT 25.820 64.070 26.140 64.130 ;
        RECT 27.290 64.070 27.430 64.225 ;
        RECT 25.820 63.930 27.430 64.070 ;
        RECT 25.820 63.870 26.140 63.930 ;
        RECT 10.640 63.730 10.960 63.790 ;
        RECT 13.875 63.730 14.165 63.775 ;
        RECT 10.640 63.590 14.165 63.730 ;
        RECT 10.640 63.530 10.960 63.590 ;
        RECT 13.875 63.545 14.165 63.590 ;
        RECT 15.700 63.530 16.020 63.790 ;
        RECT 18.935 63.730 19.225 63.775 ;
        RECT 21.680 63.730 22.000 63.790 ;
        RECT 18.935 63.590 22.000 63.730 ;
        RECT 18.935 63.545 19.225 63.590 ;
        RECT 21.680 63.530 22.000 63.590 ;
        RECT 24.440 63.730 24.760 63.790 ;
        RECT 25.375 63.730 25.665 63.775 ;
        RECT 24.440 63.590 25.665 63.730 ;
        RECT 24.440 63.530 24.760 63.590 ;
        RECT 25.375 63.545 25.665 63.590 ;
        RECT 26.740 63.730 27.060 63.790 ;
        RECT 27.750 63.730 27.890 64.225 ;
        RECT 28.580 64.210 28.900 64.470 ;
        RECT 29.960 64.210 30.280 64.470 ;
        RECT 33.195 64.410 33.485 64.455 ;
        RECT 39.620 64.410 39.940 64.470 ;
        RECT 33.195 64.270 39.940 64.410 ;
        RECT 33.195 64.225 33.485 64.270 ;
        RECT 39.620 64.210 39.940 64.270 ;
        RECT 45.155 64.410 45.445 64.455 ;
        RECT 46.980 64.410 47.300 64.470 ;
        RECT 45.155 64.270 47.300 64.410 ;
        RECT 45.155 64.225 45.445 64.270 ;
        RECT 46.980 64.210 47.300 64.270 ;
        RECT 49.755 64.410 50.045 64.455 ;
        RECT 50.200 64.410 50.520 64.470 ;
        RECT 49.755 64.270 50.520 64.410 ;
        RECT 49.755 64.225 50.045 64.270 ;
        RECT 50.200 64.210 50.520 64.270 ;
        RECT 56.640 64.410 56.960 64.470 ;
        RECT 62.175 64.410 62.465 64.455 ;
        RECT 56.640 64.270 62.465 64.410 ;
        RECT 56.640 64.210 56.960 64.270 ;
        RECT 62.175 64.225 62.465 64.270 ;
        RECT 64.460 64.410 64.780 64.470 ;
        RECT 66.760 64.410 67.080 64.470 ;
        RECT 67.310 64.455 67.450 64.610 ;
        RECT 69.060 64.550 69.380 64.610 ;
        RECT 72.280 64.550 72.600 64.610 ;
        RECT 72.755 64.750 73.045 64.795 ;
        RECT 75.500 64.750 75.820 64.810 ;
        RECT 80.100 64.750 80.420 64.810 ;
        RECT 72.755 64.610 80.420 64.750 ;
        RECT 72.755 64.565 73.045 64.610 ;
        RECT 75.500 64.550 75.820 64.610 ;
        RECT 80.100 64.550 80.420 64.610 ;
        RECT 84.240 64.750 84.560 64.810 ;
        RECT 84.715 64.750 85.005 64.795 ;
        RECT 84.240 64.610 85.005 64.750 ;
        RECT 84.240 64.550 84.560 64.610 ;
        RECT 84.715 64.565 85.005 64.610 ;
        RECT 85.160 64.550 85.480 64.810 ;
        RECT 64.460 64.270 67.080 64.410 ;
        RECT 64.460 64.210 64.780 64.270 ;
        RECT 66.760 64.210 67.080 64.270 ;
        RECT 67.235 64.225 67.525 64.455 ;
        RECT 71.360 64.410 71.680 64.470 ;
        RECT 74.135 64.410 74.425 64.455 ;
        RECT 71.360 64.270 74.425 64.410 ;
        RECT 71.360 64.210 71.680 64.270 ;
        RECT 74.135 64.225 74.425 64.270 ;
        RECT 75.055 64.410 75.345 64.455 ;
        RECT 76.420 64.410 76.740 64.470 ;
        RECT 78.260 64.410 78.580 64.470 ;
        RECT 75.055 64.270 78.580 64.410 ;
        RECT 75.055 64.225 75.345 64.270 ;
        RECT 76.420 64.210 76.740 64.270 ;
        RECT 78.260 64.210 78.580 64.270 ;
        RECT 79.195 64.410 79.485 64.455 ;
        RECT 86.540 64.410 86.860 64.470 ;
        RECT 79.195 64.270 86.860 64.410 ;
        RECT 79.195 64.225 79.485 64.270 ;
        RECT 86.540 64.210 86.860 64.270 ;
        RECT 87.475 64.410 87.765 64.455 ;
        RECT 87.920 64.410 88.240 64.470 ;
        RECT 87.475 64.270 88.240 64.410 ;
        RECT 87.475 64.225 87.765 64.270 ;
        RECT 87.920 64.210 88.240 64.270 ;
        RECT 29.055 63.885 29.345 64.115 ;
        RECT 34.530 64.070 34.820 64.115 ;
        RECT 35.020 64.070 35.340 64.130 ;
        RECT 34.530 63.930 35.340 64.070 ;
        RECT 34.530 63.885 34.820 63.930 ;
        RECT 26.740 63.590 27.890 63.730 ;
        RECT 28.120 63.730 28.440 63.790 ;
        RECT 29.130 63.730 29.270 63.885 ;
        RECT 35.020 63.870 35.340 63.930 ;
        RECT 52.470 64.070 52.760 64.115 ;
        RECT 53.880 64.070 54.200 64.130 ;
        RECT 52.470 63.930 54.200 64.070 ;
        RECT 52.470 63.885 52.760 63.930 ;
        RECT 53.880 63.870 54.200 63.930 ;
        RECT 64.000 64.070 64.320 64.130 ;
        RECT 66.300 64.070 66.620 64.130 ;
        RECT 68.615 64.070 68.905 64.115 ;
        RECT 64.000 63.930 68.905 64.070 ;
        RECT 64.000 63.870 64.320 63.930 ;
        RECT 66.300 63.870 66.620 63.930 ;
        RECT 68.615 63.885 68.905 63.930 ;
        RECT 84.255 64.070 84.545 64.115 ;
        RECT 85.620 64.070 85.940 64.130 ;
        RECT 84.255 63.930 85.940 64.070 ;
        RECT 84.255 63.885 84.545 63.930 ;
        RECT 85.620 63.870 85.940 63.930 ;
        RECT 28.120 63.590 29.270 63.730 ;
        RECT 30.420 63.730 30.740 63.790 ;
        RECT 30.895 63.730 31.185 63.775 ;
        RECT 30.420 63.590 31.185 63.730 ;
        RECT 26.740 63.530 27.060 63.590 ;
        RECT 28.120 63.530 28.440 63.590 ;
        RECT 30.420 63.530 30.740 63.590 ;
        RECT 30.895 63.545 31.185 63.590 ;
        RECT 43.300 63.530 43.620 63.790 ;
        RECT 45.600 63.530 45.920 63.790 ;
        RECT 47.900 63.730 48.220 63.790 ;
        RECT 49.295 63.730 49.585 63.775 ;
        RECT 51.120 63.730 51.440 63.790 ;
        RECT 47.900 63.590 51.440 63.730 ;
        RECT 47.900 63.530 48.220 63.590 ;
        RECT 49.295 63.545 49.585 63.590 ;
        RECT 51.120 63.530 51.440 63.590 ;
        RECT 58.480 63.530 58.800 63.790 ;
        RECT 65.380 63.530 65.700 63.790 ;
        RECT 65.840 63.530 66.160 63.790 ;
        RECT 81.955 63.730 82.245 63.775 ;
        RECT 83.780 63.730 84.100 63.790 ;
        RECT 81.955 63.590 84.100 63.730 ;
        RECT 81.955 63.545 82.245 63.590 ;
        RECT 83.780 63.530 84.100 63.590 ;
        RECT 11.950 62.910 90.610 63.390 ;
        RECT 25.360 62.710 25.680 62.770 ;
        RECT 28.120 62.710 28.440 62.770 ;
        RECT 14.870 62.570 28.440 62.710 ;
        RECT 14.870 62.415 15.010 62.570 ;
        RECT 25.360 62.510 25.680 62.570 ;
        RECT 28.120 62.510 28.440 62.570 ;
        RECT 29.960 62.710 30.280 62.770 ;
        RECT 37.335 62.710 37.625 62.755 ;
        RECT 29.960 62.570 37.625 62.710 ;
        RECT 29.960 62.510 30.280 62.570 ;
        RECT 37.335 62.525 37.625 62.570 ;
        RECT 47.915 62.710 48.205 62.755 ;
        RECT 49.740 62.710 50.060 62.770 ;
        RECT 47.915 62.570 50.060 62.710 ;
        RECT 47.915 62.525 48.205 62.570 ;
        RECT 49.740 62.510 50.060 62.570 ;
        RECT 51.580 62.510 51.900 62.770 ;
        RECT 53.880 62.510 54.200 62.770 ;
        RECT 56.195 62.710 56.485 62.755 ;
        RECT 56.640 62.710 56.960 62.770 ;
        RECT 56.195 62.570 56.960 62.710 ;
        RECT 56.195 62.525 56.485 62.570 ;
        RECT 56.640 62.510 56.960 62.570 ;
        RECT 64.015 62.525 64.305 62.755 ;
        RECT 65.380 62.710 65.700 62.770 ;
        RECT 65.380 62.570 66.990 62.710 ;
        RECT 14.795 62.185 15.085 62.415 ;
        RECT 15.715 62.370 16.005 62.415 ;
        RECT 20.760 62.370 21.080 62.430 ;
        RECT 30.880 62.370 31.200 62.430 ;
        RECT 34.100 62.370 34.420 62.430 ;
        RECT 15.715 62.230 21.080 62.370 ;
        RECT 15.715 62.185 16.005 62.230 ;
        RECT 20.760 62.170 21.080 62.230 ;
        RECT 23.150 62.230 30.650 62.370 ;
        RECT 20.300 62.030 20.620 62.090 ;
        RECT 23.150 62.075 23.290 62.230 ;
        RECT 24.440 62.075 24.760 62.090 ;
        RECT 30.510 62.075 30.650 62.230 ;
        RECT 30.880 62.230 34.420 62.370 ;
        RECT 30.880 62.170 31.200 62.230 ;
        RECT 34.100 62.170 34.420 62.230 ;
        RECT 42.350 62.370 42.640 62.415 ;
        RECT 43.300 62.370 43.620 62.430 ;
        RECT 42.350 62.230 43.620 62.370 ;
        RECT 42.350 62.185 42.640 62.230 ;
        RECT 43.300 62.170 43.620 62.230 ;
        RECT 52.055 62.370 52.345 62.415 ;
        RECT 58.480 62.370 58.800 62.430 ;
        RECT 52.055 62.230 58.800 62.370 ;
        RECT 52.055 62.185 52.345 62.230 ;
        RECT 58.480 62.170 58.800 62.230 ;
        RECT 61.870 62.370 62.160 62.415 ;
        RECT 64.090 62.370 64.230 62.525 ;
        RECT 65.380 62.510 65.700 62.570 ;
        RECT 61.870 62.230 64.230 62.370 ;
        RECT 61.870 62.185 62.160 62.230 ;
        RECT 65.840 62.170 66.160 62.430 ;
        RECT 31.800 62.075 32.120 62.090 ;
        RECT 23.075 62.030 23.365 62.075 ;
        RECT 24.410 62.030 24.760 62.075 ;
        RECT 20.300 61.890 23.365 62.030 ;
        RECT 24.245 61.890 24.760 62.030 ;
        RECT 20.300 61.830 20.620 61.890 ;
        RECT 23.075 61.845 23.365 61.890 ;
        RECT 24.410 61.845 24.760 61.890 ;
        RECT 30.435 61.845 30.725 62.075 ;
        RECT 31.770 61.845 32.120 62.075 ;
        RECT 24.440 61.830 24.760 61.845 ;
        RECT 31.800 61.830 32.120 61.845 ;
        RECT 39.620 62.030 39.940 62.090 ;
        RECT 41.015 62.030 41.305 62.075 ;
        RECT 39.620 61.890 41.305 62.030 ;
        RECT 39.620 61.830 39.940 61.890 ;
        RECT 41.015 61.845 41.305 61.890 ;
        RECT 63.080 61.830 63.400 62.090 ;
        RECT 64.460 62.030 64.780 62.090 ;
        RECT 64.935 62.030 65.225 62.075 ;
        RECT 64.460 61.890 65.225 62.030 ;
        RECT 64.460 61.830 64.780 61.890 ;
        RECT 64.935 61.845 65.225 61.890 ;
        RECT 65.380 61.830 65.700 62.090 ;
        RECT 66.850 62.075 66.990 62.570 ;
        RECT 69.520 62.510 69.840 62.770 ;
        RECT 77.800 62.710 78.120 62.770 ;
        RECT 80.115 62.710 80.405 62.755 ;
        RECT 77.800 62.570 80.405 62.710 ;
        RECT 77.800 62.510 78.120 62.570 ;
        RECT 80.115 62.525 80.405 62.570 ;
        RECT 83.780 62.510 84.100 62.770 ;
        RECT 86.080 62.510 86.400 62.770 ;
        RECT 69.610 62.370 69.750 62.510 ;
        RECT 73.200 62.370 73.520 62.430 ;
        RECT 68.230 62.230 73.520 62.370 ;
        RECT 66.775 61.845 67.065 62.075 ;
        RECT 67.220 61.830 67.540 62.090 ;
        RECT 68.230 62.075 68.370 62.230 ;
        RECT 73.200 62.170 73.520 62.230 ;
        RECT 68.155 61.845 68.445 62.075 ;
        RECT 69.535 62.030 69.825 62.075 ;
        RECT 75.500 62.030 75.820 62.090 ;
        RECT 69.535 61.890 75.820 62.030 ;
        RECT 69.535 61.845 69.825 61.890 ;
        RECT 21.220 61.490 21.540 61.750 ;
        RECT 22.600 61.490 22.920 61.750 ;
        RECT 23.955 61.690 24.245 61.735 ;
        RECT 25.145 61.690 25.435 61.735 ;
        RECT 27.665 61.690 27.955 61.735 ;
        RECT 23.955 61.550 27.955 61.690 ;
        RECT 23.955 61.505 24.245 61.550 ;
        RECT 25.145 61.505 25.435 61.550 ;
        RECT 27.665 61.505 27.955 61.550 ;
        RECT 31.315 61.690 31.605 61.735 ;
        RECT 32.505 61.690 32.795 61.735 ;
        RECT 35.025 61.690 35.315 61.735 ;
        RECT 31.315 61.550 35.315 61.690 ;
        RECT 31.315 61.505 31.605 61.550 ;
        RECT 32.505 61.505 32.795 61.550 ;
        RECT 35.025 61.505 35.315 61.550 ;
        RECT 41.895 61.690 42.185 61.735 ;
        RECT 43.085 61.690 43.375 61.735 ;
        RECT 45.605 61.690 45.895 61.735 ;
        RECT 41.895 61.550 45.895 61.690 ;
        RECT 41.895 61.505 42.185 61.550 ;
        RECT 43.085 61.505 43.375 61.550 ;
        RECT 45.605 61.505 45.895 61.550 ;
        RECT 51.120 61.690 51.440 61.750 ;
        RECT 54.340 61.690 54.660 61.750 ;
        RECT 51.120 61.550 54.660 61.690 ;
        RECT 51.120 61.490 51.440 61.550 ;
        RECT 54.340 61.490 54.660 61.550 ;
        RECT 58.505 61.690 58.795 61.735 ;
        RECT 61.025 61.690 61.315 61.735 ;
        RECT 62.215 61.690 62.505 61.735 ;
        RECT 58.505 61.550 62.505 61.690 ;
        RECT 63.170 61.690 63.310 61.830 ;
        RECT 69.610 61.690 69.750 61.845 ;
        RECT 75.500 61.830 75.820 61.890 ;
        RECT 76.420 62.030 76.740 62.090 ;
        RECT 79.640 62.030 79.960 62.090 ;
        RECT 76.420 61.890 79.960 62.030 ;
        RECT 76.420 61.830 76.740 61.890 ;
        RECT 79.640 61.830 79.960 61.890 ;
        RECT 80.575 61.845 80.865 62.075 ;
        RECT 63.170 61.550 69.750 61.690 ;
        RECT 72.280 61.690 72.600 61.750 ;
        RECT 80.650 61.690 80.790 61.845 ;
        RECT 87.000 61.830 87.320 62.090 ;
        RECT 87.460 61.830 87.780 62.090 ;
        RECT 72.280 61.550 80.790 61.690 ;
        RECT 58.505 61.505 58.795 61.550 ;
        RECT 61.025 61.505 61.315 61.550 ;
        RECT 62.215 61.505 62.505 61.550 ;
        RECT 72.280 61.490 72.600 61.550 ;
        RECT 84.240 61.490 84.560 61.750 ;
        RECT 84.715 61.505 85.005 61.735 ;
        RECT 14.780 61.350 15.100 61.410 ;
        RECT 23.560 61.350 23.850 61.395 ;
        RECT 25.660 61.350 25.950 61.395 ;
        RECT 27.230 61.350 27.520 61.395 ;
        RECT 14.780 61.210 20.300 61.350 ;
        RECT 14.780 61.150 15.100 61.210 ;
        RECT 16.635 61.010 16.925 61.055 ;
        RECT 17.080 61.010 17.400 61.070 ;
        RECT 16.635 60.870 17.400 61.010 ;
        RECT 20.160 61.010 20.300 61.210 ;
        RECT 23.560 61.210 27.520 61.350 ;
        RECT 23.560 61.165 23.850 61.210 ;
        RECT 25.660 61.165 25.950 61.210 ;
        RECT 27.230 61.165 27.520 61.210 ;
        RECT 30.920 61.350 31.210 61.395 ;
        RECT 33.020 61.350 33.310 61.395 ;
        RECT 34.590 61.350 34.880 61.395 ;
        RECT 30.920 61.210 34.880 61.350 ;
        RECT 30.920 61.165 31.210 61.210 ;
        RECT 33.020 61.165 33.310 61.210 ;
        RECT 34.590 61.165 34.880 61.210 ;
        RECT 41.500 61.350 41.790 61.395 ;
        RECT 43.600 61.350 43.890 61.395 ;
        RECT 45.170 61.350 45.460 61.395 ;
        RECT 41.500 61.210 45.460 61.350 ;
        RECT 41.500 61.165 41.790 61.210 ;
        RECT 43.600 61.165 43.890 61.210 ;
        RECT 45.170 61.165 45.460 61.210 ;
        RECT 58.940 61.350 59.230 61.395 ;
        RECT 60.510 61.350 60.800 61.395 ;
        RECT 62.610 61.350 62.900 61.395 ;
        RECT 58.940 61.210 62.900 61.350 ;
        RECT 58.940 61.165 59.230 61.210 ;
        RECT 60.510 61.165 60.800 61.210 ;
        RECT 62.610 61.165 62.900 61.210 ;
        RECT 75.960 61.350 76.280 61.410 ;
        RECT 84.790 61.350 84.930 61.505 ;
        RECT 75.960 61.210 84.930 61.350 ;
        RECT 75.960 61.150 76.280 61.210 ;
        RECT 88.380 61.150 88.700 61.410 ;
        RECT 26.280 61.010 26.600 61.070 ;
        RECT 29.975 61.010 30.265 61.055 ;
        RECT 34.100 61.010 34.420 61.070 ;
        RECT 20.160 60.870 34.420 61.010 ;
        RECT 16.635 60.825 16.925 60.870 ;
        RECT 17.080 60.810 17.400 60.870 ;
        RECT 26.280 60.810 26.600 60.870 ;
        RECT 29.975 60.825 30.265 60.870 ;
        RECT 34.100 60.810 34.420 60.870 ;
        RECT 67.695 61.010 67.985 61.055 ;
        RECT 68.600 61.010 68.920 61.070 ;
        RECT 67.695 60.870 68.920 61.010 ;
        RECT 67.695 60.825 67.985 60.870 ;
        RECT 68.600 60.810 68.920 60.870 ;
        RECT 72.280 61.010 72.600 61.070 ;
        RECT 79.180 61.010 79.500 61.070 ;
        RECT 72.280 60.870 79.500 61.010 ;
        RECT 72.280 60.810 72.600 60.870 ;
        RECT 79.180 60.810 79.500 60.870 ;
        RECT 81.940 60.810 82.260 61.070 ;
        RECT 11.950 60.190 90.610 60.670 ;
        RECT 12.020 59.990 12.340 60.050 ;
        RECT 13.875 59.990 14.165 60.035 ;
        RECT 12.020 59.850 14.165 59.990 ;
        RECT 12.020 59.790 12.340 59.850 ;
        RECT 13.875 59.805 14.165 59.850 ;
        RECT 21.220 59.990 21.540 60.050 ;
        RECT 24.900 59.990 25.220 60.050 ;
        RECT 21.220 59.850 25.220 59.990 ;
        RECT 21.220 59.790 21.540 59.850 ;
        RECT 24.900 59.790 25.220 59.850 ;
        RECT 26.740 59.990 27.060 60.050 ;
        RECT 27.215 59.990 27.505 60.035 ;
        RECT 26.740 59.850 27.505 59.990 ;
        RECT 26.740 59.790 27.060 59.850 ;
        RECT 27.215 59.805 27.505 59.850 ;
        RECT 31.355 59.990 31.645 60.035 ;
        RECT 31.800 59.990 32.120 60.050 ;
        RECT 31.355 59.850 32.120 59.990 ;
        RECT 31.355 59.805 31.645 59.850 ;
        RECT 31.800 59.790 32.120 59.850 ;
        RECT 41.015 59.990 41.305 60.035 ;
        RECT 41.460 59.990 41.780 60.050 ;
        RECT 41.015 59.850 41.780 59.990 ;
        RECT 41.015 59.805 41.305 59.850 ;
        RECT 41.460 59.790 41.780 59.850 ;
        RECT 48.360 59.990 48.680 60.050 ;
        RECT 49.295 59.990 49.585 60.035 ;
        RECT 48.360 59.850 49.585 59.990 ;
        RECT 48.360 59.790 48.680 59.850 ;
        RECT 49.295 59.805 49.585 59.850 ;
        RECT 54.815 59.990 55.105 60.035 ;
        RECT 56.180 59.990 56.500 60.050 ;
        RECT 54.815 59.850 56.500 59.990 ;
        RECT 54.815 59.805 55.105 59.850 ;
        RECT 56.180 59.790 56.500 59.850 ;
        RECT 65.380 59.990 65.700 60.050 ;
        RECT 70.900 59.990 71.220 60.050 ;
        RECT 65.380 59.850 71.220 59.990 ;
        RECT 65.380 59.790 65.700 59.850 ;
        RECT 70.900 59.790 71.220 59.850 ;
        RECT 71.360 59.990 71.680 60.050 ;
        RECT 75.500 59.990 75.820 60.050 ;
        RECT 71.360 59.850 75.820 59.990 ;
        RECT 71.360 59.790 71.680 59.850 ;
        RECT 75.500 59.790 75.820 59.850 ;
        RECT 75.960 59.790 76.280 60.050 ;
        RECT 79.655 59.990 79.945 60.035 ;
        RECT 84.240 59.990 84.560 60.050 ;
        RECT 79.655 59.850 84.560 59.990 ;
        RECT 79.655 59.805 79.945 59.850 ;
        RECT 84.240 59.790 84.560 59.850 ;
        RECT 86.540 59.990 86.860 60.050 ;
        RECT 87.475 59.990 87.765 60.035 ;
        RECT 86.540 59.850 87.765 59.990 ;
        RECT 86.540 59.790 86.860 59.850 ;
        RECT 87.475 59.805 87.765 59.850 ;
        RECT 15.740 59.650 16.030 59.695 ;
        RECT 17.840 59.650 18.130 59.695 ;
        RECT 19.410 59.650 19.700 59.695 ;
        RECT 15.740 59.510 19.700 59.650 ;
        RECT 15.740 59.465 16.030 59.510 ;
        RECT 17.840 59.465 18.130 59.510 ;
        RECT 19.410 59.465 19.700 59.510 ;
        RECT 20.760 59.650 21.080 59.710 ;
        RECT 22.155 59.650 22.445 59.695 ;
        RECT 23.520 59.650 23.840 59.710 ;
        RECT 29.500 59.650 29.820 59.710 ;
        RECT 20.760 59.510 23.840 59.650 ;
        RECT 20.760 59.450 21.080 59.510 ;
        RECT 22.155 59.465 22.445 59.510 ;
        RECT 23.520 59.450 23.840 59.510 ;
        RECT 28.570 59.510 29.820 59.650 ;
        RECT 16.135 59.310 16.425 59.355 ;
        RECT 17.325 59.310 17.615 59.355 ;
        RECT 19.845 59.310 20.135 59.355 ;
        RECT 16.135 59.170 20.135 59.310 ;
        RECT 16.135 59.125 16.425 59.170 ;
        RECT 17.325 59.125 17.615 59.170 ;
        RECT 19.845 59.125 20.135 59.170 ;
        RECT 14.795 58.785 15.085 59.015 ;
        RECT 14.870 58.630 15.010 58.785 ;
        RECT 15.240 58.770 15.560 59.030 ;
        RECT 20.760 58.970 21.080 59.030 ;
        RECT 16.250 58.830 21.080 58.970 ;
        RECT 16.250 58.630 16.390 58.830 ;
        RECT 20.760 58.770 21.080 58.830 ;
        RECT 25.360 58.770 25.680 59.030 ;
        RECT 26.280 58.770 26.600 59.030 ;
        RECT 28.135 58.970 28.425 59.015 ;
        RECT 28.570 58.970 28.710 59.510 ;
        RECT 29.500 59.450 29.820 59.510 ;
        RECT 34.140 59.650 34.430 59.695 ;
        RECT 36.240 59.650 36.530 59.695 ;
        RECT 37.810 59.650 38.100 59.695 ;
        RECT 34.140 59.510 38.100 59.650 ;
        RECT 34.140 59.465 34.430 59.510 ;
        RECT 36.240 59.465 36.530 59.510 ;
        RECT 37.810 59.465 38.100 59.510 ;
        RECT 39.160 59.650 39.480 59.710 ;
        RECT 64.000 59.650 64.320 59.710 ;
        RECT 71.820 59.650 72.140 59.710 ;
        RECT 81.060 59.650 81.350 59.695 ;
        RECT 83.160 59.650 83.450 59.695 ;
        RECT 84.730 59.650 85.020 59.695 ;
        RECT 39.160 59.510 66.990 59.650 ;
        RECT 39.160 59.450 39.480 59.510 ;
        RECT 64.000 59.450 64.320 59.510 ;
        RECT 30.420 59.310 30.740 59.370 ;
        RECT 29.130 59.170 30.740 59.310 ;
        RECT 29.130 59.015 29.270 59.170 ;
        RECT 30.420 59.110 30.740 59.170 ;
        RECT 34.535 59.310 34.825 59.355 ;
        RECT 35.725 59.310 36.015 59.355 ;
        RECT 38.245 59.310 38.535 59.355 ;
        RECT 34.535 59.170 38.535 59.310 ;
        RECT 34.535 59.125 34.825 59.170 ;
        RECT 35.725 59.125 36.015 59.170 ;
        RECT 38.245 59.125 38.535 59.170 ;
        RECT 44.235 59.310 44.525 59.355 ;
        RECT 46.060 59.310 46.380 59.370 ;
        RECT 44.235 59.170 46.380 59.310 ;
        RECT 44.235 59.125 44.525 59.170 ;
        RECT 46.060 59.110 46.380 59.170 ;
        RECT 46.995 59.310 47.285 59.355 ;
        RECT 56.640 59.310 56.960 59.370 ;
        RECT 57.115 59.310 57.405 59.355 ;
        RECT 46.995 59.170 56.410 59.310 ;
        RECT 46.995 59.125 47.285 59.170 ;
        RECT 26.785 58.830 28.710 58.970 ;
        RECT 16.620 58.675 16.940 58.690 ;
        RECT 14.870 58.490 16.390 58.630 ;
        RECT 16.590 58.445 16.940 58.675 ;
        RECT 16.620 58.430 16.940 58.445 ;
        RECT 17.540 58.630 17.860 58.690 ;
        RECT 21.680 58.630 22.000 58.690 ;
        RECT 26.785 58.630 26.925 58.830 ;
        RECT 28.135 58.785 28.425 58.830 ;
        RECT 29.055 58.785 29.345 59.015 ;
        RECT 29.515 58.785 29.805 59.015 ;
        RECT 29.975 58.970 30.265 59.015 ;
        RECT 30.880 58.970 31.200 59.030 ;
        RECT 29.975 58.830 31.200 58.970 ;
        RECT 29.975 58.785 30.265 58.830 ;
        RECT 17.540 58.490 26.925 58.630 ;
        RECT 27.660 58.630 27.980 58.690 ;
        RECT 29.590 58.630 29.730 58.785 ;
        RECT 30.880 58.770 31.200 58.830 ;
        RECT 33.655 58.970 33.945 59.015 ;
        RECT 39.620 58.970 39.940 59.030 ;
        RECT 33.655 58.830 39.940 58.970 ;
        RECT 33.655 58.785 33.945 58.830 ;
        RECT 39.620 58.770 39.940 58.830 ;
        RECT 47.455 58.970 47.745 59.015 ;
        RECT 49.740 58.970 50.060 59.030 ;
        RECT 47.455 58.830 50.060 58.970 ;
        RECT 56.270 58.970 56.410 59.170 ;
        RECT 56.640 59.170 57.405 59.310 ;
        RECT 56.640 59.110 56.960 59.170 ;
        RECT 57.115 59.125 57.405 59.170 ;
        RECT 58.035 59.310 58.325 59.355 ;
        RECT 58.940 59.310 59.260 59.370 ;
        RECT 66.300 59.310 66.620 59.370 ;
        RECT 58.035 59.170 59.260 59.310 ;
        RECT 58.035 59.125 58.325 59.170 ;
        RECT 58.940 59.110 59.260 59.170 ;
        RECT 65.930 59.170 66.620 59.310 ;
        RECT 66.850 59.310 66.990 59.510 ;
        RECT 67.770 59.510 72.140 59.650 ;
        RECT 67.770 59.310 67.910 59.510 ;
        RECT 71.820 59.450 72.140 59.510 ;
        RECT 72.370 59.510 77.110 59.650 ;
        RECT 66.850 59.170 67.910 59.310 ;
        RECT 68.155 59.310 68.445 59.355 ;
        RECT 72.370 59.310 72.510 59.510 ;
        RECT 68.155 59.170 72.510 59.310 ;
        RECT 72.740 59.310 73.060 59.370 ;
        RECT 73.675 59.310 73.965 59.355 ;
        RECT 72.740 59.170 73.965 59.310 ;
        RECT 63.080 58.970 63.400 59.030 ;
        RECT 56.270 58.830 63.400 58.970 ;
        RECT 47.455 58.785 47.745 58.830 ;
        RECT 49.740 58.770 50.060 58.830 ;
        RECT 63.080 58.770 63.400 58.830 ;
        RECT 65.380 58.770 65.700 59.030 ;
        RECT 65.930 59.015 66.070 59.170 ;
        RECT 66.300 59.110 66.620 59.170 ;
        RECT 68.155 59.125 68.445 59.170 ;
        RECT 72.740 59.110 73.060 59.170 ;
        RECT 73.675 59.125 73.965 59.170 ;
        RECT 74.120 59.110 74.440 59.370 ;
        RECT 65.855 58.785 66.145 59.015 ;
        RECT 67.220 58.770 67.540 59.030 ;
        RECT 67.680 58.770 68.000 59.030 ;
        RECT 68.615 58.970 68.905 59.015 ;
        RECT 69.060 58.970 69.380 59.030 ;
        RECT 68.615 58.830 69.380 58.970 ;
        RECT 68.615 58.785 68.905 58.830 ;
        RECT 27.660 58.490 29.730 58.630 ;
        RECT 34.990 58.630 35.280 58.675 ;
        RECT 37.780 58.630 38.100 58.690 ;
        RECT 34.990 58.490 38.100 58.630 ;
        RECT 17.540 58.430 17.860 58.490 ;
        RECT 21.680 58.430 22.000 58.490 ;
        RECT 27.660 58.430 27.980 58.490 ;
        RECT 34.990 58.445 35.280 58.490 ;
        RECT 37.780 58.430 38.100 58.490 ;
        RECT 43.315 58.630 43.605 58.675 ;
        RECT 53.880 58.630 54.200 58.690 ;
        RECT 43.315 58.490 54.200 58.630 ;
        RECT 43.315 58.445 43.605 58.490 ;
        RECT 53.880 58.430 54.200 58.490 ;
        RECT 66.300 58.430 66.620 58.690 ;
        RECT 18.000 58.290 18.320 58.350 ;
        RECT 19.840 58.290 20.160 58.350 ;
        RECT 18.000 58.150 20.160 58.290 ;
        RECT 18.000 58.090 18.320 58.150 ;
        RECT 19.840 58.090 20.160 58.150 ;
        RECT 27.200 58.290 27.520 58.350 ;
        RECT 29.960 58.290 30.280 58.350 ;
        RECT 27.200 58.150 30.280 58.290 ;
        RECT 27.200 58.090 27.520 58.150 ;
        RECT 29.960 58.090 30.280 58.150 ;
        RECT 40.555 58.290 40.845 58.335 ;
        RECT 42.840 58.290 43.160 58.350 ;
        RECT 40.555 58.150 43.160 58.290 ;
        RECT 40.555 58.105 40.845 58.150 ;
        RECT 42.840 58.090 43.160 58.150 ;
        RECT 56.655 58.290 56.945 58.335 ;
        RECT 58.940 58.290 59.260 58.350 ;
        RECT 56.655 58.150 59.260 58.290 ;
        RECT 56.655 58.105 56.945 58.150 ;
        RECT 58.940 58.090 59.260 58.150 ;
        RECT 64.475 58.290 64.765 58.335 ;
        RECT 64.920 58.290 65.240 58.350 ;
        RECT 64.475 58.150 65.240 58.290 ;
        RECT 64.475 58.105 64.765 58.150 ;
        RECT 64.920 58.090 65.240 58.150 ;
        RECT 67.680 58.290 68.000 58.350 ;
        RECT 68.690 58.290 68.830 58.785 ;
        RECT 69.060 58.770 69.380 58.830 ;
        RECT 69.520 58.770 69.840 59.030 ;
        RECT 69.980 58.770 70.300 59.030 ;
        RECT 70.455 58.785 70.745 59.015 ;
        RECT 69.610 58.630 69.750 58.770 ;
        RECT 70.530 58.630 70.670 58.785 ;
        RECT 70.900 58.770 71.220 59.030 ;
        RECT 71.360 58.770 71.680 59.030 ;
        RECT 72.280 58.770 72.600 59.030 ;
        RECT 73.215 58.970 73.505 59.015 ;
        RECT 74.580 58.970 74.900 59.030 ;
        RECT 73.215 58.830 74.900 58.970 ;
        RECT 73.215 58.785 73.505 58.830 ;
        RECT 74.580 58.770 74.900 58.830 ;
        RECT 75.040 58.770 75.360 59.030 ;
        RECT 76.970 59.015 77.110 59.510 ;
        RECT 81.060 59.510 85.020 59.650 ;
        RECT 81.060 59.465 81.350 59.510 ;
        RECT 83.160 59.465 83.450 59.510 ;
        RECT 84.730 59.465 85.020 59.510 ;
        RECT 80.100 59.310 80.420 59.370 ;
        RECT 80.575 59.310 80.865 59.355 ;
        RECT 80.100 59.170 80.865 59.310 ;
        RECT 80.100 59.110 80.420 59.170 ;
        RECT 80.575 59.125 80.865 59.170 ;
        RECT 81.455 59.310 81.745 59.355 ;
        RECT 82.645 59.310 82.935 59.355 ;
        RECT 85.165 59.310 85.455 59.355 ;
        RECT 81.455 59.170 85.455 59.310 ;
        RECT 81.455 59.125 81.745 59.170 ;
        RECT 82.645 59.125 82.935 59.170 ;
        RECT 85.165 59.125 85.455 59.170 ;
        RECT 76.895 58.785 77.185 59.015 ;
        RECT 77.340 58.970 77.660 59.030 ;
        RECT 77.815 58.970 78.105 59.015 ;
        RECT 77.340 58.830 78.105 58.970 ;
        RECT 77.340 58.770 77.660 58.830 ;
        RECT 77.815 58.785 78.105 58.830 ;
        RECT 78.720 58.770 79.040 59.030 ;
        RECT 81.940 59.015 82.260 59.030 ;
        RECT 81.910 58.970 82.260 59.015 ;
        RECT 81.745 58.830 82.260 58.970 ;
        RECT 87.550 58.970 87.690 59.805 ;
        RECT 87.920 59.790 88.240 60.050 ;
        RECT 88.855 58.970 89.145 59.015 ;
        RECT 87.550 58.830 89.145 58.970 ;
        RECT 81.910 58.785 82.260 58.830 ;
        RECT 88.855 58.785 89.145 58.830 ;
        RECT 81.940 58.770 82.260 58.785 ;
        RECT 69.610 58.490 70.670 58.630 ;
        RECT 71.820 58.630 72.140 58.690 ;
        RECT 78.275 58.630 78.565 58.675 ;
        RECT 71.820 58.490 78.565 58.630 ;
        RECT 71.820 58.430 72.140 58.490 ;
        RECT 78.275 58.445 78.565 58.490 ;
        RECT 67.680 58.150 68.830 58.290 ;
        RECT 69.075 58.290 69.365 58.335 ;
        RECT 69.520 58.290 69.840 58.350 ;
        RECT 69.075 58.150 69.840 58.290 ;
        RECT 67.680 58.090 68.000 58.150 ;
        RECT 69.075 58.105 69.365 58.150 ;
        RECT 69.520 58.090 69.840 58.150 ;
        RECT 69.980 58.290 70.300 58.350 ;
        RECT 74.580 58.290 74.900 58.350 ;
        RECT 69.980 58.150 74.900 58.290 ;
        RECT 69.980 58.090 70.300 58.150 ;
        RECT 74.580 58.090 74.900 58.150 ;
        RECT 11.950 57.470 90.610 57.950 ;
        RECT 14.795 57.270 15.085 57.315 ;
        RECT 16.620 57.270 16.940 57.330 ;
        RECT 14.795 57.130 16.940 57.270 ;
        RECT 14.795 57.085 15.085 57.130 ;
        RECT 16.620 57.070 16.940 57.130 ;
        RECT 20.300 57.270 20.620 57.330 ;
        RECT 24.915 57.270 25.205 57.315 ;
        RECT 35.480 57.270 35.800 57.330 ;
        RECT 20.300 57.130 24.670 57.270 ;
        RECT 20.300 57.070 20.620 57.130 ;
        RECT 19.380 56.930 19.700 56.990 ;
        RECT 16.710 56.790 19.700 56.930 ;
        RECT 24.530 56.930 24.670 57.130 ;
        RECT 24.915 57.130 35.800 57.270 ;
        RECT 24.915 57.085 25.205 57.130 ;
        RECT 35.480 57.070 35.800 57.130 ;
        RECT 37.780 57.270 38.100 57.330 ;
        RECT 38.255 57.270 38.545 57.315 ;
        RECT 37.780 57.130 38.545 57.270 ;
        RECT 37.780 57.070 38.100 57.130 ;
        RECT 38.255 57.085 38.545 57.130 ;
        RECT 45.600 57.270 45.920 57.330 ;
        RECT 46.075 57.270 46.365 57.315 ;
        RECT 45.600 57.130 46.365 57.270 ;
        RECT 45.600 57.070 45.920 57.130 ;
        RECT 46.075 57.085 46.365 57.130 ;
        RECT 67.220 57.070 67.540 57.330 ;
        RECT 70.900 57.270 71.220 57.330 ;
        RECT 68.230 57.130 68.830 57.270 ;
        RECT 25.820 56.930 26.140 56.990 ;
        RECT 27.660 56.930 27.980 56.990 ;
        RECT 24.530 56.790 27.980 56.930 ;
        RECT 16.710 56.635 16.850 56.790 ;
        RECT 19.380 56.730 19.700 56.790 ;
        RECT 25.820 56.730 26.140 56.790 ;
        RECT 16.175 56.405 16.465 56.635 ;
        RECT 16.635 56.405 16.925 56.635 ;
        RECT 16.250 55.910 16.390 56.405 ;
        RECT 17.080 56.390 17.400 56.650 ;
        RECT 17.540 56.590 17.860 56.650 ;
        RECT 18.015 56.590 18.305 56.635 ;
        RECT 17.540 56.450 18.305 56.590 ;
        RECT 17.540 56.390 17.860 56.450 ;
        RECT 18.015 56.405 18.305 56.450 ;
        RECT 18.460 56.590 18.780 56.650 ;
        RECT 18.460 56.540 19.150 56.590 ;
        RECT 19.855 56.540 20.145 56.635 ;
        RECT 18.460 56.450 20.145 56.540 ;
        RECT 18.460 56.390 18.780 56.450 ;
        RECT 19.010 56.405 20.145 56.450 ;
        RECT 19.010 56.400 20.070 56.405 ;
        RECT 20.285 56.390 20.605 56.650 ;
        RECT 20.880 56.620 21.170 56.665 ;
        RECT 20.880 56.480 21.450 56.620 ;
        RECT 20.880 56.435 21.170 56.480 ;
        RECT 21.310 55.970 21.450 56.480 ;
        RECT 21.680 56.390 22.000 56.650 ;
        RECT 22.155 56.405 22.445 56.635 ;
        RECT 22.615 56.590 22.905 56.635 ;
        RECT 23.060 56.590 23.380 56.650 ;
        RECT 22.615 56.450 23.380 56.590 ;
        RECT 22.615 56.405 22.905 56.450 ;
        RECT 16.250 55.770 19.150 55.910 ;
        RECT 19.010 55.630 19.150 55.770 ;
        RECT 21.220 55.710 21.540 55.970 ;
        RECT 22.230 55.910 22.370 56.405 ;
        RECT 23.060 56.390 23.380 56.450 ;
        RECT 23.520 56.390 23.840 56.650 ;
        RECT 23.980 56.390 24.300 56.650 ;
        RECT 24.900 56.590 25.220 56.650 ;
        RECT 26.830 56.635 26.970 56.790 ;
        RECT 27.660 56.730 27.980 56.790 ;
        RECT 28.595 56.930 28.885 56.975 ;
        RECT 30.280 56.930 30.570 56.975 ;
        RECT 28.595 56.790 30.570 56.930 ;
        RECT 28.595 56.745 28.885 56.790 ;
        RECT 30.280 56.745 30.570 56.790 ;
        RECT 34.100 56.930 34.420 56.990 ;
        RECT 53.880 56.930 54.200 56.990 ;
        RECT 68.230 56.975 68.370 57.130 ;
        RECT 34.100 56.790 47.670 56.930 ;
        RECT 34.100 56.730 34.420 56.790 ;
        RECT 25.375 56.590 25.665 56.635 ;
        RECT 24.900 56.450 25.665 56.590 ;
        RECT 24.900 56.390 25.220 56.450 ;
        RECT 25.375 56.405 25.665 56.450 ;
        RECT 26.295 56.405 26.585 56.635 ;
        RECT 26.755 56.405 27.045 56.635 ;
        RECT 23.520 55.910 23.840 55.970 ;
        RECT 22.230 55.770 23.840 55.910 ;
        RECT 23.520 55.710 23.840 55.770 ;
        RECT 18.460 55.370 18.780 55.630 ;
        RECT 18.920 55.570 19.240 55.630 ;
        RECT 22.600 55.570 22.920 55.630 ;
        RECT 18.920 55.430 22.920 55.570 ;
        RECT 26.370 55.570 26.510 56.405 ;
        RECT 27.200 56.390 27.520 56.650 ;
        RECT 29.055 56.590 29.345 56.635 ;
        RECT 29.500 56.590 29.820 56.650 ;
        RECT 29.055 56.450 29.820 56.590 ;
        RECT 29.055 56.405 29.345 56.450 ;
        RECT 29.500 56.390 29.820 56.450 ;
        RECT 40.095 56.590 40.385 56.635 ;
        RECT 42.395 56.590 42.685 56.635 ;
        RECT 40.095 56.450 42.685 56.590 ;
        RECT 40.095 56.405 40.385 56.450 ;
        RECT 42.395 56.405 42.685 56.450 ;
        RECT 42.840 56.590 43.160 56.650 ;
        RECT 45.155 56.590 45.445 56.635 ;
        RECT 42.840 56.450 45.445 56.590 ;
        RECT 42.840 56.390 43.160 56.450 ;
        RECT 45.155 56.405 45.445 56.450 ;
        RECT 46.980 56.390 47.300 56.650 ;
        RECT 47.530 56.635 47.670 56.790 ;
        RECT 53.880 56.790 64.230 56.930 ;
        RECT 53.880 56.730 54.200 56.790 ;
        RECT 47.455 56.405 47.745 56.635 ;
        RECT 48.375 56.405 48.665 56.635 ;
        RECT 29.935 56.250 30.225 56.295 ;
        RECT 31.125 56.250 31.415 56.295 ;
        RECT 33.645 56.250 33.935 56.295 ;
        RECT 29.935 56.110 33.935 56.250 ;
        RECT 29.935 56.065 30.225 56.110 ;
        RECT 31.125 56.065 31.415 56.110 ;
        RECT 33.645 56.065 33.935 56.110 ;
        RECT 40.540 56.050 40.860 56.310 ;
        RECT 41.475 56.250 41.765 56.295 ;
        RECT 47.900 56.250 48.220 56.310 ;
        RECT 41.475 56.110 48.220 56.250 ;
        RECT 48.450 56.250 48.590 56.405 ;
        RECT 48.820 56.390 49.140 56.650 ;
        RECT 64.090 56.635 64.230 56.790 ;
        RECT 68.155 56.745 68.445 56.975 ;
        RECT 52.975 56.590 53.265 56.635 ;
        RECT 55.275 56.590 55.565 56.635 ;
        RECT 52.975 56.450 55.565 56.590 ;
        RECT 52.975 56.405 53.265 56.450 ;
        RECT 55.275 56.405 55.565 56.450 ;
        RECT 64.015 56.405 64.305 56.635 ;
        RECT 67.680 56.390 68.000 56.650 ;
        RECT 68.690 56.590 68.830 57.130 ;
        RECT 69.150 57.130 71.220 57.270 ;
        RECT 69.150 56.975 69.290 57.130 ;
        RECT 70.900 57.070 71.220 57.130 ;
        RECT 76.420 57.070 76.740 57.330 ;
        RECT 69.075 56.745 69.365 56.975 ;
        RECT 69.535 56.930 69.825 56.975 ;
        RECT 69.980 56.930 70.300 56.990 ;
        RECT 72.740 56.930 73.060 56.990 ;
        RECT 75.500 56.930 75.820 56.990 ;
        RECT 78.260 56.930 78.580 56.990 ;
        RECT 69.535 56.790 70.300 56.930 ;
        RECT 69.535 56.745 69.825 56.790 ;
        RECT 69.980 56.730 70.300 56.790 ;
        RECT 70.990 56.790 73.060 56.930 ;
        RECT 70.440 56.590 70.760 56.650 ;
        RECT 70.990 56.635 71.130 56.790 ;
        RECT 72.740 56.730 73.060 56.790 ;
        RECT 73.750 56.790 78.580 56.930 ;
        RECT 68.690 56.450 70.760 56.590 ;
        RECT 70.440 56.390 70.760 56.450 ;
        RECT 70.915 56.405 71.205 56.635 ;
        RECT 71.360 56.590 71.680 56.650 ;
        RECT 72.295 56.590 72.585 56.635 ;
        RECT 71.360 56.450 72.585 56.590 ;
        RECT 71.360 56.390 71.680 56.450 ;
        RECT 72.295 56.405 72.585 56.450 ;
        RECT 52.040 56.250 52.360 56.310 ;
        RECT 48.450 56.110 52.360 56.250 ;
        RECT 41.475 56.065 41.765 56.110 ;
        RECT 47.900 56.050 48.220 56.110 ;
        RECT 52.040 56.050 52.360 56.110 ;
        RECT 53.420 56.050 53.740 56.310 ;
        RECT 54.340 56.050 54.660 56.310 ;
        RECT 57.560 56.250 57.880 56.310 ;
        RECT 58.035 56.250 58.325 56.295 ;
        RECT 57.560 56.110 58.325 56.250 ;
        RECT 57.560 56.050 57.880 56.110 ;
        RECT 58.035 56.065 58.325 56.110 ;
        RECT 58.940 56.250 59.260 56.310 ;
        RECT 62.175 56.250 62.465 56.295 ;
        RECT 58.940 56.110 62.465 56.250 ;
        RECT 58.940 56.050 59.260 56.110 ;
        RECT 62.175 56.065 62.465 56.110 ;
        RECT 64.460 56.250 64.780 56.310 ;
        RECT 64.460 56.110 68.600 56.250 ;
        RECT 64.460 56.050 64.780 56.110 ;
        RECT 29.540 55.910 29.830 55.955 ;
        RECT 31.640 55.910 31.930 55.955 ;
        RECT 33.210 55.910 33.500 55.955 ;
        RECT 29.540 55.770 33.500 55.910 ;
        RECT 29.540 55.725 29.830 55.770 ;
        RECT 31.640 55.725 31.930 55.770 ;
        RECT 33.210 55.725 33.500 55.770 ;
        RECT 66.300 55.910 66.620 55.970 ;
        RECT 67.695 55.910 67.985 55.955 ;
        RECT 66.300 55.770 67.985 55.910 ;
        RECT 68.460 55.910 68.600 56.110 ;
        RECT 69.520 56.050 69.840 56.310 ;
        RECT 72.755 56.250 73.045 56.295 ;
        RECT 73.750 56.250 73.890 56.790 ;
        RECT 75.500 56.730 75.820 56.790 ;
        RECT 78.260 56.730 78.580 56.790 ;
        RECT 74.135 56.405 74.425 56.635 ;
        RECT 74.595 56.590 74.885 56.635 ;
        RECT 75.040 56.590 75.360 56.650 ;
        RECT 75.975 56.590 76.265 56.635 ;
        RECT 74.595 56.450 75.360 56.590 ;
        RECT 74.595 56.405 74.885 56.450 ;
        RECT 72.755 56.110 73.890 56.250 ;
        RECT 72.755 56.065 73.045 56.110 ;
        RECT 74.210 55.910 74.350 56.405 ;
        RECT 75.040 56.390 75.360 56.450 ;
        RECT 75.590 56.450 76.265 56.590 ;
        RECT 75.590 55.955 75.730 56.450 ;
        RECT 75.975 56.405 76.265 56.450 ;
        RECT 79.195 56.590 79.485 56.635 ;
        RECT 79.640 56.590 79.960 56.650 ;
        RECT 80.560 56.635 80.880 56.650 ;
        RECT 79.195 56.450 79.960 56.590 ;
        RECT 79.195 56.405 79.485 56.450 ;
        RECT 79.640 56.390 79.960 56.450 ;
        RECT 80.530 56.405 80.880 56.635 ;
        RECT 80.560 56.390 80.880 56.405 ;
        RECT 82.400 56.590 82.720 56.650 ;
        RECT 87.475 56.590 87.765 56.635 ;
        RECT 82.400 56.450 87.765 56.590 ;
        RECT 82.400 56.390 82.720 56.450 ;
        RECT 87.475 56.405 87.765 56.450 ;
        RECT 78.275 56.250 78.565 56.295 ;
        RECT 78.720 56.250 79.040 56.310 ;
        RECT 78.275 56.110 79.040 56.250 ;
        RECT 78.275 56.065 78.565 56.110 ;
        RECT 78.720 56.050 79.040 56.110 ;
        RECT 80.075 56.250 80.365 56.295 ;
        RECT 81.265 56.250 81.555 56.295 ;
        RECT 83.785 56.250 84.075 56.295 ;
        RECT 80.075 56.110 84.075 56.250 ;
        RECT 80.075 56.065 80.365 56.110 ;
        RECT 81.265 56.065 81.555 56.110 ;
        RECT 83.785 56.065 84.075 56.110 ;
        RECT 68.460 55.770 74.350 55.910 ;
        RECT 66.300 55.710 66.620 55.770 ;
        RECT 67.695 55.725 67.985 55.770 ;
        RECT 75.515 55.725 75.805 55.955 ;
        RECT 79.680 55.910 79.970 55.955 ;
        RECT 81.780 55.910 82.070 55.955 ;
        RECT 83.350 55.910 83.640 55.955 ;
        RECT 79.680 55.770 83.640 55.910 ;
        RECT 79.680 55.725 79.970 55.770 ;
        RECT 81.780 55.725 82.070 55.770 ;
        RECT 83.350 55.725 83.640 55.770 ;
        RECT 29.960 55.570 30.280 55.630 ;
        RECT 26.370 55.430 30.280 55.570 ;
        RECT 18.920 55.370 19.240 55.430 ;
        RECT 22.600 55.370 22.920 55.430 ;
        RECT 29.960 55.370 30.280 55.430 ;
        RECT 33.640 55.570 33.960 55.630 ;
        RECT 35.955 55.570 36.245 55.615 ;
        RECT 33.640 55.430 36.245 55.570 ;
        RECT 33.640 55.370 33.960 55.430 ;
        RECT 35.955 55.385 36.245 55.430 ;
        RECT 51.120 55.370 51.440 55.630 ;
        RECT 59.400 55.370 59.720 55.630 ;
        RECT 68.600 55.570 68.920 55.630 ;
        RECT 70.455 55.570 70.745 55.615 ;
        RECT 74.120 55.570 74.440 55.630 ;
        RECT 68.600 55.430 74.440 55.570 ;
        RECT 68.600 55.370 68.920 55.430 ;
        RECT 70.455 55.385 70.745 55.430 ;
        RECT 74.120 55.370 74.440 55.430 ;
        RECT 77.355 55.570 77.645 55.615 ;
        RECT 83.780 55.570 84.100 55.630 ;
        RECT 77.355 55.430 84.100 55.570 ;
        RECT 77.355 55.385 77.645 55.430 ;
        RECT 83.780 55.370 84.100 55.430 ;
        RECT 86.080 55.370 86.400 55.630 ;
        RECT 88.380 55.370 88.700 55.630 ;
        RECT 11.950 54.750 90.610 55.230 ;
        RECT 15.255 54.550 15.545 54.595 ;
        RECT 21.220 54.550 21.540 54.610 ;
        RECT 33.195 54.550 33.485 54.595 ;
        RECT 40.540 54.550 40.860 54.610 ;
        RECT 15.255 54.410 21.540 54.550 ;
        RECT 15.255 54.365 15.545 54.410 ;
        RECT 21.220 54.350 21.540 54.410 ;
        RECT 30.510 54.410 32.950 54.550 ;
        RECT 16.200 54.210 16.490 54.255 ;
        RECT 18.300 54.210 18.590 54.255 ;
        RECT 19.870 54.210 20.160 54.255 ;
        RECT 16.200 54.070 20.160 54.210 ;
        RECT 16.200 54.025 16.490 54.070 ;
        RECT 18.300 54.025 18.590 54.070 ;
        RECT 19.870 54.025 20.160 54.070 ;
        RECT 15.240 53.870 15.560 53.930 ;
        RECT 15.715 53.870 16.005 53.915 ;
        RECT 15.240 53.730 16.005 53.870 ;
        RECT 15.240 53.670 15.560 53.730 ;
        RECT 15.715 53.685 16.005 53.730 ;
        RECT 16.595 53.870 16.885 53.915 ;
        RECT 17.785 53.870 18.075 53.915 ;
        RECT 20.305 53.870 20.595 53.915 ;
        RECT 16.595 53.730 20.595 53.870 ;
        RECT 16.595 53.685 16.885 53.730 ;
        RECT 17.785 53.685 18.075 53.730 ;
        RECT 20.305 53.685 20.595 53.730 ;
        RECT 15.790 53.530 15.930 53.685 ;
        RECT 23.980 53.530 24.300 53.590 ;
        RECT 30.510 53.575 30.650 54.410 ;
        RECT 32.810 53.870 32.950 54.410 ;
        RECT 33.195 54.410 40.860 54.550 ;
        RECT 33.195 54.365 33.485 54.410 ;
        RECT 40.540 54.350 40.860 54.410 ;
        RECT 47.455 54.550 47.745 54.595 ;
        RECT 53.420 54.550 53.740 54.610 ;
        RECT 47.455 54.410 53.740 54.550 ;
        RECT 47.455 54.365 47.745 54.410 ;
        RECT 53.420 54.350 53.740 54.410 ;
        RECT 53.880 54.550 54.200 54.610 ;
        RECT 53.880 54.410 56.870 54.550 ;
        RECT 53.880 54.350 54.200 54.410 ;
        RECT 52.540 54.210 52.830 54.255 ;
        RECT 54.640 54.210 54.930 54.255 ;
        RECT 56.210 54.210 56.500 54.255 ;
        RECT 52.540 54.070 56.500 54.210 ;
        RECT 56.730 54.210 56.870 54.410 ;
        RECT 58.940 54.350 59.260 54.610 ;
        RECT 63.080 54.550 63.400 54.610 ;
        RECT 66.775 54.550 67.065 54.595 ;
        RECT 80.560 54.550 80.880 54.610 ;
        RECT 81.035 54.550 81.325 54.595 ;
        RECT 63.080 54.410 80.330 54.550 ;
        RECT 63.080 54.350 63.400 54.410 ;
        RECT 66.775 54.365 67.065 54.410 ;
        RECT 59.415 54.210 59.705 54.255 ;
        RECT 56.730 54.070 59.705 54.210 ;
        RECT 52.540 54.025 52.830 54.070 ;
        RECT 54.640 54.025 54.930 54.070 ;
        RECT 56.210 54.025 56.500 54.070 ;
        RECT 59.415 54.025 59.705 54.070 ;
        RECT 62.160 54.210 62.450 54.255 ;
        RECT 63.730 54.210 64.020 54.255 ;
        RECT 65.830 54.210 66.120 54.255 ;
        RECT 62.160 54.070 66.120 54.210 ;
        RECT 62.160 54.025 62.450 54.070 ;
        RECT 63.730 54.025 64.020 54.070 ;
        RECT 65.830 54.025 66.120 54.070 ;
        RECT 69.520 54.210 69.810 54.255 ;
        RECT 71.090 54.210 71.380 54.255 ;
        RECT 73.190 54.210 73.480 54.255 ;
        RECT 69.520 54.070 73.480 54.210 ;
        RECT 69.520 54.025 69.810 54.070 ;
        RECT 71.090 54.025 71.380 54.070 ;
        RECT 73.190 54.025 73.480 54.070 ;
        RECT 74.580 54.010 74.900 54.270 ;
        RECT 79.640 54.010 79.960 54.270 ;
        RECT 52.935 53.870 53.225 53.915 ;
        RECT 54.125 53.870 54.415 53.915 ;
        RECT 56.645 53.870 56.935 53.915 ;
        RECT 31.430 53.730 32.490 53.870 ;
        RECT 32.810 53.730 52.730 53.870 ;
        RECT 15.790 53.390 20.300 53.530 ;
        RECT 13.400 52.990 13.720 53.250 ;
        RECT 14.335 53.005 14.625 53.235 ;
        RECT 17.050 53.190 17.340 53.235 ;
        RECT 18.460 53.190 18.780 53.250 ;
        RECT 17.050 53.050 18.780 53.190 ;
        RECT 20.160 53.190 20.300 53.390 ;
        RECT 23.980 53.390 30.190 53.530 ;
        RECT 23.980 53.330 24.300 53.390 ;
        RECT 25.375 53.190 25.665 53.235 ;
        RECT 27.200 53.190 27.520 53.250 ;
        RECT 20.160 53.050 27.520 53.190 ;
        RECT 30.050 53.190 30.190 53.390 ;
        RECT 30.435 53.345 30.725 53.575 ;
        RECT 30.880 53.330 31.200 53.590 ;
        RECT 31.430 53.190 31.570 53.730 ;
        RECT 32.350 53.575 32.490 53.730 ;
        RECT 31.815 53.345 32.105 53.575 ;
        RECT 32.275 53.530 32.565 53.575 ;
        RECT 46.980 53.530 47.300 53.590 ;
        RECT 48.360 53.530 48.680 53.590 ;
        RECT 32.275 53.390 48.680 53.530 ;
        RECT 32.275 53.345 32.565 53.390 ;
        RECT 30.050 53.050 31.570 53.190 ;
        RECT 17.050 53.005 17.340 53.050 ;
        RECT 14.410 52.850 14.550 53.005 ;
        RECT 18.460 52.990 18.780 53.050 ;
        RECT 25.375 53.005 25.665 53.050 ;
        RECT 27.200 52.990 27.520 53.050 ;
        RECT 14.780 52.850 15.100 52.910 ;
        RECT 22.615 52.850 22.905 52.895 ;
        RECT 31.890 52.850 32.030 53.345 ;
        RECT 46.980 53.330 47.300 53.390 ;
        RECT 48.360 53.330 48.680 53.390 ;
        RECT 48.835 53.345 49.125 53.575 ;
        RECT 49.755 53.345 50.045 53.575 ;
        RECT 33.180 53.190 33.500 53.250 ;
        RECT 48.910 53.190 49.050 53.345 ;
        RECT 33.180 53.050 49.050 53.190 ;
        RECT 33.180 52.990 33.500 53.050 ;
        RECT 14.410 52.710 32.030 52.850 ;
        RECT 49.830 52.850 49.970 53.345 ;
        RECT 50.200 53.330 50.520 53.590 ;
        RECT 52.055 53.345 52.345 53.575 ;
        RECT 52.590 53.530 52.730 53.730 ;
        RECT 52.935 53.730 56.935 53.870 ;
        RECT 52.935 53.685 53.225 53.730 ;
        RECT 54.125 53.685 54.415 53.730 ;
        RECT 56.645 53.685 56.935 53.730 ;
        RECT 61.725 53.870 62.015 53.915 ;
        RECT 64.245 53.870 64.535 53.915 ;
        RECT 65.435 53.870 65.725 53.915 ;
        RECT 61.725 53.730 65.725 53.870 ;
        RECT 61.725 53.685 62.015 53.730 ;
        RECT 64.245 53.685 64.535 53.730 ;
        RECT 65.435 53.685 65.725 53.730 ;
        RECT 69.085 53.870 69.375 53.915 ;
        RECT 71.605 53.870 71.895 53.915 ;
        RECT 72.795 53.870 73.085 53.915 ;
        RECT 69.085 53.730 73.085 53.870 ;
        RECT 69.085 53.685 69.375 53.730 ;
        RECT 71.605 53.685 71.895 53.730 ;
        RECT 72.795 53.685 73.085 53.730 ;
        RECT 73.675 53.870 73.965 53.915 ;
        RECT 79.730 53.870 79.870 54.010 ;
        RECT 80.190 53.915 80.330 54.410 ;
        RECT 80.560 54.410 81.325 54.550 ;
        RECT 80.560 54.350 80.880 54.410 ;
        RECT 81.035 54.365 81.325 54.410 ;
        RECT 73.675 53.730 79.870 53.870 ;
        RECT 73.675 53.685 73.965 53.730 ;
        RECT 80.115 53.685 80.405 53.915 ;
        RECT 59.860 53.530 60.180 53.590 ;
        RECT 52.590 53.390 60.180 53.530 ;
        RECT 52.130 53.190 52.270 53.345 ;
        RECT 59.860 53.330 60.180 53.390 ;
        RECT 64.920 53.575 65.240 53.590 ;
        RECT 64.920 53.530 65.270 53.575 ;
        RECT 66.315 53.530 66.605 53.575 ;
        RECT 73.750 53.530 73.890 53.685 ;
        RECT 83.320 53.670 83.640 53.930 ;
        RECT 83.780 53.670 84.100 53.930 ;
        RECT 86.080 53.870 86.400 53.930 ;
        RECT 87.935 53.870 88.225 53.915 ;
        RECT 88.840 53.870 89.160 53.930 ;
        RECT 86.080 53.730 89.160 53.870 ;
        RECT 86.080 53.670 86.400 53.730 ;
        RECT 87.935 53.685 88.225 53.730 ;
        RECT 88.840 53.670 89.160 53.730 ;
        RECT 64.920 53.390 65.435 53.530 ;
        RECT 66.315 53.390 73.890 53.530 ;
        RECT 64.920 53.345 65.270 53.390 ;
        RECT 66.315 53.345 66.605 53.390 ;
        RECT 64.920 53.330 65.240 53.345 ;
        RECT 74.120 53.330 74.440 53.590 ;
        RECT 75.055 53.530 75.345 53.575 ;
        RECT 75.500 53.530 75.820 53.590 ;
        RECT 75.055 53.390 75.820 53.530 ;
        RECT 75.055 53.345 75.345 53.390 ;
        RECT 75.500 53.330 75.820 53.390 ;
        RECT 52.500 53.190 52.820 53.250 ;
        RECT 52.130 53.050 52.820 53.190 ;
        RECT 52.500 52.990 52.820 53.050 ;
        RECT 53.390 53.190 53.680 53.235 ;
        RECT 57.100 53.190 57.420 53.250 ;
        RECT 53.390 53.050 57.420 53.190 ;
        RECT 53.390 53.005 53.680 53.050 ;
        RECT 57.100 52.990 57.420 53.050 ;
        RECT 69.980 53.190 70.300 53.250 ;
        RECT 72.340 53.190 72.630 53.235 ;
        RECT 69.980 53.050 72.630 53.190 ;
        RECT 69.980 52.990 70.300 53.050 ;
        RECT 72.340 53.005 72.630 53.050 ;
        RECT 60.780 52.850 61.100 52.910 ;
        RECT 49.830 52.710 61.100 52.850 ;
        RECT 14.780 52.650 15.100 52.710 ;
        RECT 22.615 52.665 22.905 52.710 ;
        RECT 60.780 52.650 61.100 52.710 ;
        RECT 76.880 52.650 77.200 52.910 ;
        RECT 82.875 52.850 83.165 52.895 ;
        RECT 85.175 52.850 85.465 52.895 ;
        RECT 82.875 52.710 85.465 52.850 ;
        RECT 82.875 52.665 83.165 52.710 ;
        RECT 85.175 52.665 85.465 52.710 ;
        RECT 11.950 52.030 90.610 52.510 ;
        RECT 26.740 51.830 27.060 51.890 ;
        RECT 31.800 51.830 32.120 51.890 ;
        RECT 26.740 51.690 32.120 51.830 ;
        RECT 26.740 51.630 27.060 51.690 ;
        RECT 31.800 51.630 32.120 51.690 ;
        RECT 32.260 51.830 32.580 51.890 ;
        RECT 34.560 51.830 34.880 51.890 ;
        RECT 32.260 51.690 34.880 51.830 ;
        RECT 32.260 51.630 32.580 51.690 ;
        RECT 34.560 51.630 34.880 51.690 ;
        RECT 57.100 51.630 57.420 51.890 ;
        RECT 58.955 51.830 59.245 51.875 ;
        RECT 59.400 51.830 59.720 51.890 ;
        RECT 58.955 51.690 59.720 51.830 ;
        RECT 58.955 51.645 59.245 51.690 ;
        RECT 59.400 51.630 59.720 51.690 ;
        RECT 59.860 51.830 60.180 51.890 ;
        RECT 76.420 51.830 76.740 51.890 ;
        RECT 59.860 51.690 76.740 51.830 ;
        RECT 59.860 51.630 60.180 51.690 ;
        RECT 76.420 51.630 76.740 51.690 ;
        RECT 23.075 51.490 23.365 51.535 ;
        RECT 25.360 51.490 25.680 51.550 ;
        RECT 23.075 51.350 25.680 51.490 ;
        RECT 23.075 51.305 23.365 51.350 ;
        RECT 25.360 51.290 25.680 51.350 ;
        RECT 29.975 51.490 30.265 51.535 ;
        RECT 38.240 51.490 38.560 51.550 ;
        RECT 51.120 51.535 51.440 51.550 ;
        RECT 51.090 51.490 51.440 51.535 ;
        RECT 29.975 51.350 38.560 51.490 ;
        RECT 50.925 51.350 51.440 51.490 ;
        RECT 29.975 51.305 30.265 51.350 ;
        RECT 38.240 51.290 38.560 51.350 ;
        RECT 51.090 51.305 51.440 51.350 ;
        RECT 51.120 51.290 51.440 51.305 ;
        RECT 75.960 51.490 76.280 51.550 ;
        RECT 77.355 51.490 77.645 51.535 ;
        RECT 75.960 51.350 77.645 51.490 ;
        RECT 75.960 51.290 76.280 51.350 ;
        RECT 77.355 51.305 77.645 51.350 ;
        RECT 14.780 50.950 15.100 51.210 ;
        RECT 16.635 51.150 16.925 51.195 ;
        RECT 18.920 51.150 19.240 51.210 ;
        RECT 16.635 51.010 19.240 51.150 ;
        RECT 16.635 50.965 16.925 51.010 ;
        RECT 18.920 50.950 19.240 51.010 ;
        RECT 23.995 50.965 24.285 51.195 ;
        RECT 25.450 51.150 25.590 51.290 ;
        RECT 30.435 51.150 30.725 51.195 ;
        RECT 25.450 51.010 30.725 51.150 ;
        RECT 30.435 50.965 30.725 51.010 ;
        RECT 31.355 51.150 31.645 51.195 ;
        RECT 33.180 51.150 33.500 51.210 ;
        RECT 31.355 51.010 33.500 51.150 ;
        RECT 31.355 50.965 31.645 51.010 ;
        RECT 11.560 50.470 11.880 50.530 ;
        RECT 15.715 50.470 16.005 50.515 ;
        RECT 24.070 50.470 24.210 50.965 ;
        RECT 33.180 50.950 33.500 51.010 ;
        RECT 36.875 50.965 37.165 51.195 ;
        RECT 26.295 50.810 26.585 50.855 ;
        RECT 27.200 50.810 27.520 50.870 ;
        RECT 29.500 50.810 29.820 50.870 ;
        RECT 26.295 50.670 29.820 50.810 ;
        RECT 26.295 50.625 26.585 50.670 ;
        RECT 27.200 50.610 27.520 50.670 ;
        RECT 29.500 50.610 29.820 50.670 ;
        RECT 29.960 50.810 30.280 50.870 ;
        RECT 32.275 50.810 32.565 50.855 ;
        RECT 29.960 50.670 32.565 50.810 ;
        RECT 36.950 50.810 37.090 50.965 ;
        RECT 39.620 50.950 39.940 51.210 ;
        RECT 40.080 50.950 40.400 51.210 ;
        RECT 41.000 50.950 41.320 51.210 ;
        RECT 41.475 51.150 41.765 51.195 ;
        RECT 42.840 51.150 43.160 51.210 ;
        RECT 43.760 51.195 44.080 51.210 ;
        RECT 41.475 51.010 43.160 51.150 ;
        RECT 41.475 50.965 41.765 51.010 ;
        RECT 42.840 50.950 43.160 51.010 ;
        RECT 43.730 50.965 44.080 51.195 ;
        RECT 49.755 51.150 50.045 51.195 ;
        RECT 52.500 51.150 52.820 51.210 ;
        RECT 49.755 51.010 52.820 51.150 ;
        RECT 49.755 50.965 50.045 51.010 ;
        RECT 43.760 50.950 44.080 50.965 ;
        RECT 52.500 50.950 52.820 51.010 ;
        RECT 76.880 50.950 77.200 51.210 ;
        RECT 88.840 50.950 89.160 51.210 ;
        RECT 36.950 50.670 41.230 50.810 ;
        RECT 29.960 50.610 30.280 50.670 ;
        RECT 32.275 50.625 32.565 50.670 ;
        RECT 41.090 50.530 41.230 50.670 ;
        RECT 42.395 50.625 42.685 50.855 ;
        RECT 43.275 50.810 43.565 50.855 ;
        RECT 44.465 50.810 44.755 50.855 ;
        RECT 46.985 50.810 47.275 50.855 ;
        RECT 43.275 50.670 47.275 50.810 ;
        RECT 43.275 50.625 43.565 50.670 ;
        RECT 44.465 50.625 44.755 50.670 ;
        RECT 46.985 50.625 47.275 50.670 ;
        RECT 50.635 50.810 50.925 50.855 ;
        RECT 51.825 50.810 52.115 50.855 ;
        RECT 54.345 50.810 54.635 50.855 ;
        RECT 50.635 50.670 54.635 50.810 ;
        RECT 50.635 50.625 50.925 50.670 ;
        RECT 51.825 50.625 52.115 50.670 ;
        RECT 54.345 50.625 54.635 50.670 ;
        RECT 40.080 50.470 40.400 50.530 ;
        RECT 11.560 50.330 16.005 50.470 ;
        RECT 11.560 50.270 11.880 50.330 ;
        RECT 15.715 50.285 16.005 50.330 ;
        RECT 20.160 50.330 40.400 50.470 ;
        RECT 12.940 50.130 13.260 50.190 ;
        RECT 13.875 50.130 14.165 50.175 ;
        RECT 12.940 49.990 14.165 50.130 ;
        RECT 12.940 49.930 13.260 49.990 ;
        RECT 13.875 49.945 14.165 49.990 ;
        RECT 14.780 50.130 15.100 50.190 ;
        RECT 20.160 50.130 20.300 50.330 ;
        RECT 40.080 50.270 40.400 50.330 ;
        RECT 41.000 50.470 41.320 50.530 ;
        RECT 42.470 50.470 42.610 50.625 ;
        RECT 59.400 50.610 59.720 50.870 ;
        RECT 59.875 50.625 60.165 50.855 ;
        RECT 41.000 50.330 42.610 50.470 ;
        RECT 42.880 50.470 43.170 50.515 ;
        RECT 44.980 50.470 45.270 50.515 ;
        RECT 46.550 50.470 46.840 50.515 ;
        RECT 42.880 50.330 46.840 50.470 ;
        RECT 41.000 50.270 41.320 50.330 ;
        RECT 42.880 50.285 43.170 50.330 ;
        RECT 44.980 50.285 45.270 50.330 ;
        RECT 46.550 50.285 46.840 50.330 ;
        RECT 49.280 50.270 49.600 50.530 ;
        RECT 50.240 50.470 50.530 50.515 ;
        RECT 52.340 50.470 52.630 50.515 ;
        RECT 53.910 50.470 54.200 50.515 ;
        RECT 50.240 50.330 54.200 50.470 ;
        RECT 50.240 50.285 50.530 50.330 ;
        RECT 52.340 50.285 52.630 50.330 ;
        RECT 53.910 50.285 54.200 50.330 ;
        RECT 56.655 50.470 56.945 50.515 ;
        RECT 57.560 50.470 57.880 50.530 ;
        RECT 56.655 50.330 57.880 50.470 ;
        RECT 56.655 50.285 56.945 50.330 ;
        RECT 57.560 50.270 57.880 50.330 ;
        RECT 14.780 49.990 20.300 50.130 ;
        RECT 24.915 50.130 25.205 50.175 ;
        RECT 26.740 50.130 27.060 50.190 ;
        RECT 24.915 49.990 27.060 50.130 ;
        RECT 14.780 49.930 15.100 49.990 ;
        RECT 24.915 49.945 25.205 49.990 ;
        RECT 26.740 49.930 27.060 49.990 ;
        RECT 38.715 50.130 39.005 50.175 ;
        RECT 46.060 50.130 46.380 50.190 ;
        RECT 38.715 49.990 46.380 50.130 ;
        RECT 38.715 49.945 39.005 49.990 ;
        RECT 46.060 49.930 46.380 49.990 ;
        RECT 47.900 50.130 48.220 50.190 ;
        RECT 54.340 50.130 54.660 50.190 ;
        RECT 59.950 50.130 60.090 50.625 ;
        RECT 87.460 50.470 87.780 50.530 ;
        RECT 87.935 50.470 88.225 50.515 ;
        RECT 87.460 50.330 88.225 50.470 ;
        RECT 87.460 50.270 87.780 50.330 ;
        RECT 87.935 50.285 88.225 50.330 ;
        RECT 47.900 49.990 60.090 50.130 ;
        RECT 47.900 49.930 48.220 49.990 ;
        RECT 54.340 49.930 54.660 49.990 ;
        RECT 11.950 49.310 90.610 49.790 ;
        RECT 28.580 49.110 28.900 49.170 ;
        RECT 35.940 49.110 36.260 49.170 ;
        RECT 28.580 48.970 36.260 49.110 ;
        RECT 28.580 48.910 28.900 48.970 ;
        RECT 35.940 48.910 36.260 48.970 ;
        RECT 36.415 49.110 36.705 49.155 ;
        RECT 40.080 49.110 40.400 49.170 ;
        RECT 36.415 48.970 40.400 49.110 ;
        RECT 36.415 48.925 36.705 48.970 ;
        RECT 40.080 48.910 40.400 48.970 ;
        RECT 43.760 49.110 44.080 49.170 ;
        RECT 44.235 49.110 44.525 49.155 ;
        RECT 43.760 48.970 44.525 49.110 ;
        RECT 43.760 48.910 44.080 48.970 ;
        RECT 44.235 48.925 44.525 48.970 ;
        RECT 51.580 49.110 51.900 49.170 ;
        RECT 55.735 49.110 56.025 49.155 ;
        RECT 51.580 48.970 56.025 49.110 ;
        RECT 51.580 48.910 51.900 48.970 ;
        RECT 55.735 48.925 56.025 48.970 ;
        RECT 60.780 48.910 61.100 49.170 ;
        RECT 61.700 49.110 62.020 49.170 ;
        RECT 70.440 49.110 70.760 49.170 ;
        RECT 61.700 48.970 70.760 49.110 ;
        RECT 61.700 48.910 62.020 48.970 ;
        RECT 70.440 48.910 70.760 48.970 ;
        RECT 10.640 48.770 10.960 48.830 ;
        RECT 13.875 48.770 14.165 48.815 ;
        RECT 20.300 48.770 20.620 48.830 ;
        RECT 23.980 48.770 24.300 48.830 ;
        RECT 10.640 48.630 14.165 48.770 ;
        RECT 10.640 48.570 10.960 48.630 ;
        RECT 13.875 48.585 14.165 48.630 ;
        RECT 16.250 48.630 24.300 48.770 ;
        RECT 14.780 47.890 15.100 48.150 ;
        RECT 16.250 48.135 16.390 48.630 ;
        RECT 20.300 48.570 20.620 48.630 ;
        RECT 23.980 48.570 24.300 48.630 ;
        RECT 30.000 48.770 30.290 48.815 ;
        RECT 32.100 48.770 32.390 48.815 ;
        RECT 33.670 48.770 33.960 48.815 ;
        RECT 30.000 48.630 33.960 48.770 ;
        RECT 30.000 48.585 30.290 48.630 ;
        RECT 32.100 48.585 32.390 48.630 ;
        RECT 33.670 48.585 33.960 48.630 ;
        RECT 37.360 48.770 37.650 48.815 ;
        RECT 39.460 48.770 39.750 48.815 ;
        RECT 41.030 48.770 41.320 48.815 ;
        RECT 37.360 48.630 41.320 48.770 ;
        RECT 37.360 48.585 37.650 48.630 ;
        RECT 39.460 48.585 39.750 48.630 ;
        RECT 41.030 48.585 41.320 48.630 ;
        RECT 42.840 48.770 43.160 48.830 ;
        RECT 71.375 48.770 71.665 48.815 ;
        RECT 42.840 48.630 71.665 48.770 ;
        RECT 42.840 48.570 43.160 48.630 ;
        RECT 71.375 48.585 71.665 48.630 ;
        RECT 19.380 48.430 19.700 48.490 ;
        RECT 28.120 48.430 28.440 48.490 ;
        RECT 17.630 48.290 28.440 48.430 ;
        RECT 16.175 47.905 16.465 48.135 ;
        RECT 16.620 48.090 16.940 48.150 ;
        RECT 17.630 48.135 17.770 48.290 ;
        RECT 19.380 48.230 19.700 48.290 ;
        RECT 17.095 48.090 17.385 48.135 ;
        RECT 16.620 47.950 17.385 48.090 ;
        RECT 16.620 47.890 16.940 47.950 ;
        RECT 17.095 47.905 17.385 47.950 ;
        RECT 17.555 47.905 17.845 48.135 ;
        RECT 18.000 47.890 18.320 48.150 ;
        RECT 21.220 47.890 21.540 48.150 ;
        RECT 24.900 48.090 25.220 48.150 ;
        RECT 25.835 48.090 26.125 48.135 ;
        RECT 24.900 47.950 26.125 48.090 ;
        RECT 24.900 47.890 25.220 47.950 ;
        RECT 25.835 47.905 26.125 47.950 ;
        RECT 19.380 47.210 19.700 47.470 ;
        RECT 20.300 47.210 20.620 47.470 ;
        RECT 25.910 47.410 26.050 47.905 ;
        RECT 26.740 47.890 27.060 48.150 ;
        RECT 27.290 48.135 27.430 48.290 ;
        RECT 28.120 48.230 28.440 48.290 ;
        RECT 29.500 48.230 29.820 48.490 ;
        RECT 30.395 48.430 30.685 48.475 ;
        RECT 31.585 48.430 31.875 48.475 ;
        RECT 34.105 48.430 34.395 48.475 ;
        RECT 30.395 48.290 34.395 48.430 ;
        RECT 30.395 48.245 30.685 48.290 ;
        RECT 31.585 48.245 31.875 48.290 ;
        RECT 34.105 48.245 34.395 48.290 ;
        RECT 37.755 48.430 38.045 48.475 ;
        RECT 38.945 48.430 39.235 48.475 ;
        RECT 41.465 48.430 41.755 48.475 ;
        RECT 37.755 48.290 41.755 48.430 ;
        RECT 37.755 48.245 38.045 48.290 ;
        RECT 38.945 48.245 39.235 48.290 ;
        RECT 41.465 48.245 41.755 48.290 ;
        RECT 46.060 48.430 46.380 48.490 ;
        RECT 46.535 48.430 46.825 48.475 ;
        RECT 46.060 48.290 46.825 48.430 ;
        RECT 46.060 48.230 46.380 48.290 ;
        RECT 46.535 48.245 46.825 48.290 ;
        RECT 47.455 48.430 47.745 48.475 ;
        RECT 47.900 48.430 48.220 48.490 ;
        RECT 47.455 48.290 48.220 48.430 ;
        RECT 47.455 48.245 47.745 48.290 ;
        RECT 47.900 48.230 48.220 48.290 ;
        RECT 49.280 48.430 49.600 48.490 ;
        RECT 53.895 48.430 54.185 48.475 ;
        RECT 49.280 48.290 54.185 48.430 ;
        RECT 49.280 48.230 49.600 48.290 ;
        RECT 53.895 48.245 54.185 48.290 ;
        RECT 54.340 48.430 54.660 48.490 ;
        RECT 72.740 48.430 73.060 48.490 ;
        RECT 54.340 48.290 56.870 48.430 ;
        RECT 54.340 48.230 54.660 48.290 ;
        RECT 27.215 47.905 27.505 48.135 ;
        RECT 27.675 48.090 27.965 48.135 ;
        RECT 29.960 48.090 30.280 48.150 ;
        RECT 33.640 48.090 33.960 48.150 ;
        RECT 27.675 47.950 33.960 48.090 ;
        RECT 27.675 47.905 27.965 47.950 ;
        RECT 29.960 47.890 30.280 47.950 ;
        RECT 33.640 47.890 33.960 47.950 ;
        RECT 36.875 48.090 37.165 48.135 ;
        RECT 41.000 48.090 41.320 48.150 ;
        RECT 36.875 47.950 41.320 48.090 ;
        RECT 36.875 47.905 37.165 47.950 ;
        RECT 41.000 47.890 41.320 47.950 ;
        RECT 41.550 47.950 56.410 48.090 ;
        RECT 29.055 47.750 29.345 47.795 ;
        RECT 30.740 47.750 31.030 47.795 ;
        RECT 29.055 47.610 31.030 47.750 ;
        RECT 29.055 47.565 29.345 47.610 ;
        RECT 30.740 47.565 31.030 47.610 ;
        RECT 31.800 47.750 32.120 47.810 ;
        RECT 33.180 47.750 33.500 47.810 ;
        RECT 31.800 47.610 33.500 47.750 ;
        RECT 31.800 47.550 32.120 47.610 ;
        RECT 33.180 47.550 33.500 47.610 ;
        RECT 38.210 47.750 38.500 47.795 ;
        RECT 38.700 47.750 39.020 47.810 ;
        RECT 41.550 47.750 41.690 47.950 ;
        RECT 38.210 47.610 39.020 47.750 ;
        RECT 38.210 47.565 38.500 47.610 ;
        RECT 38.700 47.550 39.020 47.610 ;
        RECT 39.250 47.610 41.690 47.750 ;
        RECT 46.075 47.750 46.365 47.795 ;
        RECT 51.135 47.750 51.425 47.795 ;
        RECT 46.075 47.610 51.425 47.750 ;
        RECT 39.250 47.410 39.390 47.610 ;
        RECT 46.075 47.565 46.365 47.610 ;
        RECT 51.135 47.565 51.425 47.610 ;
        RECT 54.800 47.550 55.120 47.810 ;
        RECT 25.910 47.270 39.390 47.410 ;
        RECT 39.620 47.410 39.940 47.470 ;
        RECT 43.760 47.410 44.080 47.470 ;
        RECT 39.620 47.270 44.080 47.410 ;
        RECT 39.620 47.210 39.940 47.270 ;
        RECT 43.760 47.210 44.080 47.270 ;
        RECT 55.720 47.210 56.040 47.470 ;
        RECT 56.270 47.410 56.410 47.950 ;
        RECT 56.730 47.750 56.870 48.290 ;
        RECT 62.250 48.290 73.060 48.430 ;
        RECT 57.115 48.090 57.405 48.135 ;
        RECT 61.700 48.090 62.020 48.150 ;
        RECT 62.250 48.135 62.390 48.290 ;
        RECT 72.740 48.230 73.060 48.290 ;
        RECT 57.115 47.950 62.020 48.090 ;
        RECT 57.115 47.905 57.405 47.950 ;
        RECT 61.700 47.890 62.020 47.950 ;
        RECT 62.175 47.905 62.465 48.135 ;
        RECT 63.540 47.890 63.860 48.150 ;
        RECT 64.015 48.090 64.305 48.135 ;
        RECT 65.395 48.090 65.685 48.135 ;
        RECT 67.220 48.090 67.540 48.150 ;
        RECT 64.015 47.950 64.690 48.090 ;
        RECT 64.015 47.905 64.305 47.950 ;
        RECT 58.035 47.750 58.325 47.795 ;
        RECT 56.730 47.610 58.325 47.750 ;
        RECT 58.035 47.565 58.325 47.610 ;
        RECT 58.955 47.750 59.245 47.795 ;
        RECT 61.240 47.750 61.560 47.810 ;
        RECT 62.635 47.750 62.925 47.795 ;
        RECT 58.955 47.610 62.925 47.750 ;
        RECT 58.955 47.565 59.245 47.610 ;
        RECT 61.240 47.550 61.560 47.610 ;
        RECT 62.635 47.565 62.925 47.610 ;
        RECT 64.550 47.410 64.690 47.950 ;
        RECT 65.395 47.950 67.540 48.090 ;
        RECT 65.395 47.905 65.685 47.950 ;
        RECT 67.220 47.890 67.540 47.950 ;
        RECT 68.615 48.090 68.905 48.135 ;
        RECT 69.060 48.090 69.380 48.150 ;
        RECT 68.615 47.950 69.380 48.090 ;
        RECT 68.615 47.905 68.905 47.950 ;
        RECT 69.060 47.890 69.380 47.950 ;
        RECT 70.440 47.890 70.760 48.150 ;
        RECT 76.895 48.090 77.185 48.135 ;
        RECT 71.910 47.950 77.185 48.090 ;
        RECT 64.920 47.750 65.240 47.810 ;
        RECT 69.535 47.750 69.825 47.795 ;
        RECT 64.920 47.610 69.825 47.750 ;
        RECT 64.920 47.550 65.240 47.610 ;
        RECT 69.535 47.565 69.825 47.610 ;
        RECT 69.995 47.750 70.285 47.795 ;
        RECT 70.900 47.750 71.220 47.810 ;
        RECT 71.910 47.750 72.050 47.950 ;
        RECT 76.895 47.905 77.185 47.950 ;
        RECT 69.995 47.610 71.220 47.750 ;
        RECT 69.995 47.565 70.285 47.610 ;
        RECT 70.900 47.550 71.220 47.610 ;
        RECT 71.450 47.610 72.050 47.750 ;
        RECT 56.270 47.270 64.690 47.410 ;
        RECT 67.220 47.410 67.540 47.470 ;
        RECT 71.450 47.410 71.590 47.610 ;
        RECT 72.740 47.550 73.060 47.810 ;
        RECT 73.660 47.550 73.980 47.810 ;
        RECT 76.970 47.750 77.110 47.905 ;
        RECT 77.800 47.890 78.120 48.150 ;
        RECT 78.260 47.890 78.580 48.150 ;
        RECT 78.720 47.890 79.040 48.150 ;
        RECT 83.320 47.750 83.640 47.810 ;
        RECT 76.970 47.610 83.640 47.750 ;
        RECT 83.320 47.550 83.640 47.610 ;
        RECT 67.220 47.270 71.590 47.410 ;
        RECT 67.220 47.210 67.540 47.270 ;
        RECT 71.820 47.210 72.140 47.470 ;
        RECT 80.100 47.210 80.420 47.470 ;
        RECT 11.950 46.590 90.610 47.070 ;
        RECT 16.620 46.190 16.940 46.450 ;
        RECT 22.140 46.390 22.460 46.450 ;
        RECT 23.995 46.390 24.285 46.435 ;
        RECT 37.320 46.390 37.640 46.450 ;
        RECT 18.090 46.250 24.285 46.390 ;
        RECT 13.400 46.050 13.720 46.110 ;
        RECT 14.795 46.050 15.085 46.095 ;
        RECT 13.400 45.910 15.085 46.050 ;
        RECT 13.400 45.850 13.720 45.910 ;
        RECT 14.795 45.865 15.085 45.910 ;
        RECT 15.715 46.050 16.005 46.095 ;
        RECT 18.090 46.050 18.230 46.250 ;
        RECT 22.140 46.190 22.460 46.250 ;
        RECT 23.995 46.205 24.285 46.250 ;
        RECT 25.910 46.250 37.640 46.390 ;
        RECT 15.715 45.910 18.230 46.050 ;
        RECT 18.430 46.050 18.720 46.095 ;
        RECT 19.380 46.050 19.700 46.110 ;
        RECT 18.430 45.910 19.700 46.050 ;
        RECT 15.715 45.865 16.005 45.910 ;
        RECT 18.430 45.865 18.720 45.910 ;
        RECT 14.870 45.710 15.010 45.865 ;
        RECT 19.380 45.850 19.700 45.910 ;
        RECT 21.220 46.050 21.540 46.110 ;
        RECT 25.415 46.050 25.705 46.095 ;
        RECT 25.910 46.050 26.050 46.250 ;
        RECT 37.320 46.190 37.640 46.250 ;
        RECT 72.740 46.390 73.060 46.450 ;
        RECT 79.655 46.390 79.945 46.435 ;
        RECT 82.400 46.390 82.720 46.450 ;
        RECT 72.740 46.250 82.720 46.390 ;
        RECT 72.740 46.190 73.060 46.250 ;
        RECT 79.655 46.205 79.945 46.250 ;
        RECT 82.400 46.190 82.720 46.250 ;
        RECT 21.220 45.910 26.050 46.050 ;
        RECT 26.295 46.050 26.585 46.095 ;
        RECT 26.295 45.910 27.890 46.050 ;
        RECT 21.220 45.850 21.540 45.910 ;
        RECT 25.415 45.865 25.705 45.910 ;
        RECT 26.295 45.865 26.585 45.910 ;
        RECT 24.455 45.710 24.745 45.755 ;
        RECT 25.820 45.710 26.140 45.770 ;
        RECT 27.750 45.755 27.890 45.910 ;
        RECT 30.510 45.910 32.490 46.050 ;
        RECT 14.870 45.570 26.140 45.710 ;
        RECT 24.455 45.525 24.745 45.570 ;
        RECT 25.820 45.510 26.140 45.570 ;
        RECT 26.755 45.525 27.045 45.755 ;
        RECT 27.675 45.525 27.965 45.755 ;
        RECT 15.240 45.370 15.560 45.430 ;
        RECT 17.095 45.370 17.385 45.415 ;
        RECT 15.240 45.230 17.385 45.370 ;
        RECT 15.240 45.170 15.560 45.230 ;
        RECT 17.095 45.185 17.385 45.230 ;
        RECT 17.975 45.370 18.265 45.415 ;
        RECT 19.165 45.370 19.455 45.415 ;
        RECT 21.685 45.370 21.975 45.415 ;
        RECT 17.975 45.230 21.975 45.370 ;
        RECT 17.975 45.185 18.265 45.230 ;
        RECT 19.165 45.185 19.455 45.230 ;
        RECT 21.685 45.185 21.975 45.230 ;
        RECT 23.980 45.370 24.300 45.430 ;
        RECT 25.360 45.370 25.680 45.430 ;
        RECT 26.830 45.370 26.970 45.525 ;
        RECT 28.120 45.510 28.440 45.770 ;
        RECT 28.580 45.510 28.900 45.770 ;
        RECT 30.510 45.755 30.650 45.910 ;
        RECT 30.435 45.525 30.725 45.755 ;
        RECT 31.715 45.710 32.005 45.755 ;
        RECT 30.970 45.570 32.005 45.710 ;
        RECT 32.350 45.710 32.490 45.910 ;
        RECT 38.240 45.850 38.560 46.110 ;
        RECT 40.080 46.050 40.400 46.110 ;
        RECT 43.315 46.050 43.605 46.095 ;
        RECT 52.975 46.050 53.265 46.095 ;
        RECT 54.340 46.050 54.660 46.110 ;
        RECT 40.080 45.910 43.605 46.050 ;
        RECT 40.080 45.850 40.400 45.910 ;
        RECT 43.315 45.865 43.605 45.910 ;
        RECT 47.990 45.910 54.660 46.050 ;
        RECT 41.000 45.710 41.320 45.770 ;
        RECT 43.760 45.710 44.080 45.770 ;
        RECT 46.075 45.710 46.365 45.755 ;
        RECT 47.455 45.710 47.745 45.755 ;
        RECT 32.350 45.570 42.150 45.710 ;
        RECT 23.980 45.230 26.970 45.370 ;
        RECT 28.210 45.370 28.350 45.510 ;
        RECT 29.500 45.370 29.820 45.430 ;
        RECT 28.210 45.230 29.820 45.370 ;
        RECT 23.980 45.170 24.300 45.230 ;
        RECT 25.360 45.170 25.680 45.230 ;
        RECT 29.500 45.170 29.820 45.230 ;
        RECT 29.975 45.370 30.265 45.415 ;
        RECT 30.970 45.370 31.110 45.570 ;
        RECT 31.715 45.525 32.005 45.570 ;
        RECT 41.000 45.510 41.320 45.570 ;
        RECT 42.010 45.415 42.150 45.570 ;
        RECT 43.760 45.570 47.745 45.710 ;
        RECT 43.760 45.510 44.080 45.570 ;
        RECT 46.075 45.525 46.365 45.570 ;
        RECT 47.455 45.525 47.745 45.570 ;
        RECT 29.975 45.230 31.110 45.370 ;
        RECT 31.315 45.370 31.605 45.415 ;
        RECT 32.505 45.370 32.795 45.415 ;
        RECT 35.025 45.370 35.315 45.415 ;
        RECT 31.315 45.230 35.315 45.370 ;
        RECT 29.975 45.185 30.265 45.230 ;
        RECT 31.315 45.185 31.605 45.230 ;
        RECT 32.505 45.185 32.795 45.230 ;
        RECT 35.025 45.185 35.315 45.230 ;
        RECT 41.935 45.370 42.225 45.415 ;
        RECT 43.300 45.370 43.620 45.430 ;
        RECT 41.935 45.230 43.620 45.370 ;
        RECT 41.935 45.185 42.225 45.230 ;
        RECT 43.300 45.170 43.620 45.230 ;
        RECT 17.580 45.030 17.870 45.075 ;
        RECT 19.680 45.030 19.970 45.075 ;
        RECT 21.250 45.030 21.540 45.075 ;
        RECT 17.580 44.890 21.540 45.030 ;
        RECT 17.580 44.845 17.870 44.890 ;
        RECT 19.680 44.845 19.970 44.890 ;
        RECT 21.250 44.845 21.540 44.890 ;
        RECT 30.920 45.030 31.210 45.075 ;
        RECT 33.020 45.030 33.310 45.075 ;
        RECT 34.590 45.030 34.880 45.075 ;
        RECT 30.920 44.890 34.880 45.030 ;
        RECT 30.920 44.845 31.210 44.890 ;
        RECT 33.020 44.845 33.310 44.890 ;
        RECT 34.590 44.845 34.880 44.890 ;
        RECT 37.320 44.830 37.640 45.090 ;
        RECT 21.680 44.690 22.000 44.750 ;
        RECT 47.990 44.690 48.130 45.910 ;
        RECT 52.975 45.865 53.265 45.910 ;
        RECT 54.340 45.850 54.660 45.910 ;
        RECT 65.840 46.050 66.160 46.110 ;
        RECT 71.835 46.050 72.125 46.095 ;
        RECT 76.880 46.050 77.200 46.110 ;
        RECT 65.840 45.910 67.910 46.050 ;
        RECT 65.840 45.850 66.160 45.910 ;
        RECT 67.770 45.770 67.910 45.910 ;
        RECT 71.835 45.910 77.200 46.050 ;
        RECT 71.835 45.865 72.125 45.910 ;
        RECT 48.360 45.710 48.680 45.770 ;
        RECT 49.295 45.710 49.585 45.755 ;
        RECT 50.215 45.710 50.505 45.755 ;
        RECT 50.660 45.710 50.980 45.770 ;
        RECT 48.360 45.570 50.980 45.710 ;
        RECT 48.360 45.510 48.680 45.570 ;
        RECT 49.295 45.525 49.585 45.570 ;
        RECT 50.215 45.525 50.505 45.570 ;
        RECT 50.660 45.510 50.980 45.570 ;
        RECT 51.580 45.510 51.900 45.770 ;
        RECT 52.500 45.710 52.820 45.770 ;
        RECT 55.260 45.710 55.580 45.770 ;
        RECT 52.500 45.570 55.580 45.710 ;
        RECT 52.500 45.510 52.820 45.570 ;
        RECT 55.260 45.510 55.580 45.570 ;
        RECT 59.860 45.510 60.180 45.770 ;
        RECT 60.795 45.710 61.085 45.755 ;
        RECT 61.240 45.710 61.560 45.770 ;
        RECT 64.920 45.710 65.240 45.770 ;
        RECT 60.795 45.570 65.240 45.710 ;
        RECT 60.795 45.525 61.085 45.570 ;
        RECT 61.240 45.510 61.560 45.570 ;
        RECT 64.920 45.510 65.240 45.570 ;
        RECT 67.235 45.525 67.525 45.755 ;
        RECT 52.055 45.185 52.345 45.415 ;
        RECT 52.130 45.030 52.270 45.185 ;
        RECT 58.940 45.170 59.260 45.430 ;
        RECT 65.840 45.370 66.160 45.430 ;
        RECT 67.310 45.370 67.450 45.525 ;
        RECT 67.680 45.510 68.000 45.770 ;
        RECT 71.910 45.370 72.050 45.865 ;
        RECT 76.880 45.850 77.200 45.910 ;
        RECT 72.280 45.710 72.600 45.770 ;
        RECT 74.035 45.710 74.325 45.755 ;
        RECT 72.280 45.570 74.325 45.710 ;
        RECT 72.280 45.510 72.600 45.570 ;
        RECT 74.035 45.525 74.325 45.570 ;
        RECT 87.460 45.510 87.780 45.770 ;
        RECT 72.755 45.370 73.045 45.415 ;
        RECT 65.840 45.230 73.045 45.370 ;
        RECT 65.840 45.170 66.160 45.230 ;
        RECT 72.755 45.185 73.045 45.230 ;
        RECT 73.635 45.370 73.925 45.415 ;
        RECT 74.825 45.370 75.115 45.415 ;
        RECT 77.345 45.370 77.635 45.415 ;
        RECT 73.635 45.230 77.635 45.370 ;
        RECT 73.635 45.185 73.925 45.230 ;
        RECT 74.825 45.185 75.115 45.230 ;
        RECT 77.345 45.185 77.635 45.230 ;
        RECT 55.720 45.030 56.040 45.090 ;
        RECT 52.130 44.890 56.040 45.030 ;
        RECT 55.720 44.830 56.040 44.890 ;
        RECT 73.240 45.030 73.530 45.075 ;
        RECT 75.340 45.030 75.630 45.075 ;
        RECT 76.910 45.030 77.200 45.075 ;
        RECT 73.240 44.890 77.200 45.030 ;
        RECT 73.240 44.845 73.530 44.890 ;
        RECT 75.340 44.845 75.630 44.890 ;
        RECT 76.910 44.845 77.200 44.890 ;
        RECT 88.395 45.030 88.685 45.075 ;
        RECT 89.300 45.030 89.620 45.090 ;
        RECT 88.395 44.890 89.620 45.030 ;
        RECT 88.395 44.845 88.685 44.890 ;
        RECT 89.300 44.830 89.620 44.890 ;
        RECT 21.680 44.550 48.130 44.690 ;
        RECT 21.680 44.490 22.000 44.550 ;
        RECT 11.950 43.870 90.610 44.350 ;
        RECT 15.240 43.670 15.560 43.730 ;
        RECT 13.490 43.530 15.560 43.670 ;
        RECT 13.490 43.035 13.630 43.530 ;
        RECT 15.240 43.470 15.560 43.530 ;
        RECT 18.920 43.670 19.240 43.730 ;
        RECT 20.315 43.670 20.605 43.715 ;
        RECT 18.920 43.530 20.605 43.670 ;
        RECT 18.920 43.470 19.240 43.530 ;
        RECT 20.315 43.485 20.605 43.530 ;
        RECT 29.055 43.670 29.345 43.715 ;
        RECT 29.500 43.670 29.820 43.730 ;
        RECT 29.055 43.530 29.820 43.670 ;
        RECT 29.055 43.485 29.345 43.530 ;
        RECT 29.500 43.470 29.820 43.530 ;
        RECT 38.255 43.670 38.545 43.715 ;
        RECT 38.700 43.670 39.020 43.730 ;
        RECT 50.215 43.670 50.505 43.715 ;
        RECT 51.580 43.670 51.900 43.730 ;
        RECT 59.860 43.670 60.180 43.730 ;
        RECT 70.900 43.670 71.220 43.730 ;
        RECT 38.255 43.530 39.020 43.670 ;
        RECT 38.255 43.485 38.545 43.530 ;
        RECT 38.700 43.470 39.020 43.530 ;
        RECT 39.250 43.530 48.130 43.670 ;
        RECT 13.900 43.330 14.190 43.375 ;
        RECT 16.000 43.330 16.290 43.375 ;
        RECT 17.570 43.330 17.860 43.375 ;
        RECT 13.900 43.190 17.860 43.330 ;
        RECT 13.900 43.145 14.190 43.190 ;
        RECT 16.000 43.145 16.290 43.190 ;
        RECT 17.570 43.145 17.860 43.190 ;
        RECT 24.440 43.330 24.760 43.390 ;
        RECT 28.135 43.330 28.425 43.375 ;
        RECT 36.860 43.330 37.180 43.390 ;
        RECT 24.440 43.190 27.430 43.330 ;
        RECT 24.440 43.130 24.760 43.190 ;
        RECT 13.415 42.805 13.705 43.035 ;
        RECT 14.295 42.990 14.585 43.035 ;
        RECT 15.485 42.990 15.775 43.035 ;
        RECT 18.005 42.990 18.295 43.035 ;
        RECT 27.290 42.990 27.430 43.190 ;
        RECT 28.135 43.190 37.180 43.330 ;
        RECT 28.135 43.145 28.425 43.190 ;
        RECT 36.860 43.130 37.180 43.190 ;
        RECT 29.040 42.990 29.360 43.050 ;
        RECT 14.295 42.850 18.295 42.990 ;
        RECT 14.295 42.805 14.585 42.850 ;
        RECT 15.485 42.805 15.775 42.850 ;
        RECT 18.005 42.805 18.295 42.850 ;
        RECT 22.230 42.850 26.970 42.990 ;
        RECT 22.230 42.710 22.370 42.850 ;
        RECT 22.140 42.450 22.460 42.710 ;
        RECT 23.520 42.650 23.840 42.710 ;
        RECT 25.375 42.650 25.665 42.695 ;
        RECT 23.520 42.510 25.665 42.650 ;
        RECT 23.520 42.450 23.840 42.510 ;
        RECT 25.375 42.465 25.665 42.510 ;
        RECT 25.835 42.650 26.125 42.695 ;
        RECT 26.280 42.650 26.600 42.710 ;
        RECT 26.830 42.695 26.970 42.850 ;
        RECT 27.290 42.850 29.360 42.990 ;
        RECT 27.290 42.695 27.430 42.850 ;
        RECT 29.040 42.790 29.360 42.850 ;
        RECT 31.355 42.990 31.645 43.035 ;
        RECT 33.180 42.990 33.500 43.050 ;
        RECT 39.250 42.990 39.390 43.530 ;
        RECT 43.800 43.330 44.090 43.375 ;
        RECT 45.900 43.330 46.190 43.375 ;
        RECT 47.470 43.330 47.760 43.375 ;
        RECT 43.800 43.190 47.760 43.330 ;
        RECT 47.990 43.330 48.130 43.530 ;
        RECT 50.215 43.530 51.900 43.670 ;
        RECT 50.215 43.485 50.505 43.530 ;
        RECT 51.580 43.470 51.900 43.530 ;
        RECT 52.130 43.530 71.220 43.670 ;
        RECT 52.130 43.330 52.270 43.530 ;
        RECT 59.860 43.470 60.180 43.530 ;
        RECT 70.900 43.470 71.220 43.530 ;
        RECT 72.280 43.470 72.600 43.730 ;
        RECT 74.595 43.670 74.885 43.715 ;
        RECT 77.800 43.670 78.120 43.730 ;
        RECT 74.595 43.530 78.120 43.670 ;
        RECT 74.595 43.485 74.885 43.530 ;
        RECT 77.800 43.470 78.120 43.530 ;
        RECT 47.990 43.190 52.270 43.330 ;
        RECT 53.000 43.330 53.290 43.375 ;
        RECT 55.100 43.330 55.390 43.375 ;
        RECT 56.670 43.330 56.960 43.375 ;
        RECT 53.000 43.190 56.960 43.330 ;
        RECT 43.800 43.145 44.090 43.190 ;
        RECT 45.900 43.145 46.190 43.190 ;
        RECT 47.470 43.145 47.760 43.190 ;
        RECT 53.000 43.145 53.290 43.190 ;
        RECT 55.100 43.145 55.390 43.190 ;
        RECT 56.670 43.145 56.960 43.190 ;
        RECT 61.280 43.330 61.570 43.375 ;
        RECT 63.380 43.330 63.670 43.375 ;
        RECT 64.950 43.330 65.240 43.375 ;
        RECT 61.280 43.190 65.240 43.330 ;
        RECT 61.280 43.145 61.570 43.190 ;
        RECT 63.380 43.145 63.670 43.190 ;
        RECT 64.950 43.145 65.240 43.190 ;
        RECT 77.380 43.330 77.670 43.375 ;
        RECT 79.480 43.330 79.770 43.375 ;
        RECT 81.050 43.330 81.340 43.375 ;
        RECT 77.380 43.190 81.340 43.330 ;
        RECT 77.380 43.145 77.670 43.190 ;
        RECT 79.480 43.145 79.770 43.190 ;
        RECT 81.050 43.145 81.340 43.190 ;
        RECT 40.555 42.990 40.845 43.035 ;
        RECT 31.355 42.850 39.390 42.990 ;
        RECT 39.710 42.850 40.845 42.990 ;
        RECT 31.355 42.805 31.645 42.850 ;
        RECT 33.180 42.790 33.500 42.850 ;
        RECT 25.835 42.510 26.600 42.650 ;
        RECT 25.835 42.465 26.125 42.510 ;
        RECT 26.280 42.450 26.600 42.510 ;
        RECT 26.755 42.465 27.045 42.695 ;
        RECT 27.215 42.465 27.505 42.695 ;
        RECT 27.660 42.650 27.980 42.710 ;
        RECT 30.435 42.650 30.725 42.695 ;
        RECT 30.895 42.650 31.185 42.695 ;
        RECT 32.720 42.650 33.040 42.710 ;
        RECT 27.660 42.510 33.040 42.650 ;
        RECT 27.660 42.450 27.980 42.510 ;
        RECT 30.435 42.465 30.725 42.510 ;
        RECT 30.895 42.465 31.185 42.510 ;
        RECT 32.720 42.450 33.040 42.510 ;
        RECT 36.400 42.650 36.720 42.710 ;
        RECT 39.710 42.650 39.850 42.850 ;
        RECT 40.555 42.805 40.845 42.850 ;
        RECT 41.475 42.990 41.765 43.035 ;
        RECT 44.195 42.990 44.485 43.035 ;
        RECT 45.385 42.990 45.675 43.035 ;
        RECT 47.905 42.990 48.195 43.035 ;
        RECT 41.475 42.850 43.990 42.990 ;
        RECT 41.475 42.805 41.765 42.850 ;
        RECT 36.400 42.510 39.850 42.650 ;
        RECT 36.400 42.450 36.720 42.510 ;
        RECT 40.080 42.450 40.400 42.710 ;
        RECT 43.300 42.450 43.620 42.710 ;
        RECT 43.850 42.650 43.990 42.850 ;
        RECT 44.195 42.850 48.195 42.990 ;
        RECT 44.195 42.805 44.485 42.850 ;
        RECT 45.385 42.805 45.675 42.850 ;
        RECT 47.905 42.805 48.195 42.850 ;
        RECT 53.395 42.990 53.685 43.035 ;
        RECT 54.585 42.990 54.875 43.035 ;
        RECT 57.105 42.990 57.395 43.035 ;
        RECT 53.395 42.850 57.395 42.990 ;
        RECT 53.395 42.805 53.685 42.850 ;
        RECT 54.585 42.805 54.875 42.850 ;
        RECT 57.105 42.805 57.395 42.850 ;
        RECT 61.675 42.990 61.965 43.035 ;
        RECT 62.865 42.990 63.155 43.035 ;
        RECT 65.385 42.990 65.675 43.035 ;
        RECT 71.820 42.990 72.140 43.050 ;
        RECT 61.675 42.850 65.675 42.990 ;
        RECT 61.675 42.805 61.965 42.850 ;
        RECT 62.865 42.805 63.155 42.850 ;
        RECT 65.385 42.805 65.675 42.850 ;
        RECT 70.070 42.850 72.140 42.990 ;
        RECT 50.660 42.650 50.980 42.710 ;
        RECT 51.135 42.650 51.425 42.695 ;
        RECT 43.850 42.510 48.130 42.650 ;
        RECT 47.990 42.370 48.130 42.510 ;
        RECT 50.660 42.510 51.425 42.650 ;
        RECT 50.660 42.450 50.980 42.510 ;
        RECT 51.135 42.465 51.425 42.510 ;
        RECT 52.515 42.650 52.805 42.695 ;
        RECT 55.260 42.650 55.580 42.710 ;
        RECT 60.795 42.650 61.085 42.695 ;
        RECT 65.840 42.650 66.160 42.710 ;
        RECT 52.515 42.510 57.330 42.650 ;
        RECT 52.515 42.465 52.805 42.510 ;
        RECT 55.260 42.450 55.580 42.510 ;
        RECT 57.190 42.370 57.330 42.510 ;
        RECT 60.795 42.510 66.160 42.650 ;
        RECT 60.795 42.465 61.085 42.510 ;
        RECT 65.840 42.450 66.160 42.510 ;
        RECT 67.220 42.650 67.540 42.710 ;
        RECT 70.070 42.695 70.210 42.850 ;
        RECT 71.820 42.790 72.140 42.850 ;
        RECT 77.775 42.990 78.065 43.035 ;
        RECT 78.965 42.990 79.255 43.035 ;
        RECT 81.485 42.990 81.775 43.035 ;
        RECT 77.775 42.850 81.775 42.990 ;
        RECT 77.775 42.805 78.065 42.850 ;
        RECT 78.965 42.805 79.255 42.850 ;
        RECT 81.485 42.805 81.775 42.850 ;
        RECT 69.075 42.650 69.365 42.695 ;
        RECT 67.220 42.510 69.365 42.650 ;
        RECT 67.220 42.450 67.540 42.510 ;
        RECT 69.075 42.465 69.365 42.510 ;
        RECT 69.995 42.465 70.285 42.695 ;
        RECT 70.440 42.450 70.760 42.710 ;
        RECT 70.915 42.465 71.205 42.695 ;
        RECT 71.360 42.650 71.680 42.710 ;
        RECT 73.675 42.650 73.965 42.695 ;
        RECT 71.360 42.510 73.965 42.650 ;
        RECT 14.780 42.355 15.100 42.370 ;
        RECT 14.750 42.125 15.100 42.355 ;
        RECT 14.780 42.110 15.100 42.125 ;
        RECT 29.500 42.310 29.820 42.370 ;
        RECT 44.650 42.310 44.940 42.355 ;
        RECT 46.520 42.310 46.840 42.370 ;
        RECT 29.500 42.170 43.530 42.310 ;
        RECT 29.500 42.110 29.820 42.170 ;
        RECT 21.220 41.770 21.540 42.030 ;
        RECT 43.390 41.970 43.530 42.170 ;
        RECT 44.650 42.170 46.840 42.310 ;
        RECT 44.650 42.125 44.940 42.170 ;
        RECT 46.520 42.110 46.840 42.170 ;
        RECT 47.900 42.310 48.220 42.370 ;
        RECT 49.740 42.310 50.060 42.370 ;
        RECT 53.880 42.355 54.200 42.370 ;
        RECT 47.900 42.170 50.060 42.310 ;
        RECT 47.900 42.110 48.220 42.170 ;
        RECT 49.740 42.110 50.060 42.170 ;
        RECT 53.850 42.125 54.200 42.355 ;
        RECT 53.880 42.110 54.200 42.125 ;
        RECT 57.100 42.110 57.420 42.370 ;
        RECT 62.130 42.310 62.420 42.355 ;
        RECT 64.000 42.310 64.320 42.370 ;
        RECT 62.130 42.170 64.320 42.310 ;
        RECT 62.130 42.125 62.420 42.170 ;
        RECT 64.000 42.110 64.320 42.170 ;
        RECT 68.600 42.310 68.920 42.370 ;
        RECT 70.990 42.310 71.130 42.465 ;
        RECT 71.360 42.450 71.680 42.510 ;
        RECT 73.675 42.465 73.965 42.510 ;
        RECT 76.880 42.650 77.200 42.710 ;
        RECT 81.940 42.650 82.260 42.710 ;
        RECT 76.880 42.510 82.260 42.650 ;
        RECT 68.600 42.170 71.130 42.310 ;
        RECT 72.755 42.310 73.045 42.355 ;
        RECT 72.755 42.170 73.430 42.310 ;
        RECT 68.600 42.110 68.920 42.170 ;
        RECT 72.755 42.125 73.045 42.170 ;
        RECT 73.290 42.030 73.430 42.170 ;
        RECT 51.595 41.970 51.885 42.015 ;
        RECT 52.960 41.970 53.280 42.030 ;
        RECT 54.800 41.970 55.120 42.030 ;
        RECT 43.390 41.830 55.120 41.970 ;
        RECT 51.595 41.785 51.885 41.830 ;
        RECT 52.960 41.770 53.280 41.830 ;
        RECT 54.800 41.770 55.120 41.830 ;
        RECT 59.415 41.970 59.705 42.015 ;
        RECT 60.780 41.970 61.100 42.030 ;
        RECT 59.415 41.830 61.100 41.970 ;
        RECT 59.415 41.785 59.705 41.830 ;
        RECT 60.780 41.770 61.100 41.830 ;
        RECT 67.695 41.970 67.985 42.015 ;
        RECT 69.520 41.970 69.840 42.030 ;
        RECT 67.695 41.830 69.840 41.970 ;
        RECT 67.695 41.785 67.985 41.830 ;
        RECT 69.520 41.770 69.840 41.830 ;
        RECT 70.440 41.970 70.760 42.030 ;
        RECT 71.820 41.970 72.140 42.030 ;
        RECT 70.440 41.830 72.140 41.970 ;
        RECT 70.440 41.770 70.760 41.830 ;
        RECT 71.820 41.770 72.140 41.830 ;
        RECT 73.200 41.770 73.520 42.030 ;
        RECT 73.750 41.970 73.890 42.465 ;
        RECT 76.880 42.450 77.200 42.510 ;
        RECT 81.940 42.450 82.260 42.510 ;
        RECT 78.230 42.310 78.520 42.355 ;
        RECT 80.100 42.310 80.420 42.370 ;
        RECT 78.230 42.170 80.420 42.310 ;
        RECT 78.230 42.125 78.520 42.170 ;
        RECT 80.100 42.110 80.420 42.170 ;
        RECT 83.795 41.970 84.085 42.015 ;
        RECT 87.460 41.970 87.780 42.030 ;
        RECT 73.750 41.830 87.780 41.970 ;
        RECT 83.795 41.785 84.085 41.830 ;
        RECT 87.460 41.770 87.780 41.830 ;
        RECT 11.950 41.150 90.610 41.630 ;
        RECT 14.335 40.950 14.625 40.995 ;
        RECT 14.780 40.950 15.100 41.010 ;
        RECT 14.335 40.810 15.100 40.950 ;
        RECT 14.335 40.765 14.625 40.810 ;
        RECT 14.780 40.750 15.100 40.810 ;
        RECT 23.075 40.950 23.365 40.995 ;
        RECT 30.420 40.950 30.740 41.010 ;
        RECT 23.075 40.810 30.740 40.950 ;
        RECT 23.075 40.765 23.365 40.810 ;
        RECT 30.420 40.750 30.740 40.810 ;
        RECT 46.520 40.750 46.840 41.010 ;
        RECT 48.375 40.950 48.665 40.995 ;
        RECT 51.580 40.950 51.900 41.010 ;
        RECT 48.375 40.810 51.900 40.950 ;
        RECT 48.375 40.765 48.665 40.810 ;
        RECT 51.580 40.750 51.900 40.810 ;
        RECT 52.055 40.950 52.345 40.995 ;
        RECT 53.420 40.950 53.740 41.010 ;
        RECT 54.355 40.950 54.645 40.995 ;
        RECT 63.080 40.950 63.400 41.010 ;
        RECT 52.055 40.810 54.645 40.950 ;
        RECT 52.055 40.765 52.345 40.810 ;
        RECT 53.420 40.750 53.740 40.810 ;
        RECT 54.355 40.765 54.645 40.810 ;
        RECT 59.490 40.810 63.400 40.950 ;
        RECT 18.015 40.610 18.305 40.655 ;
        RECT 16.710 40.470 18.305 40.610 ;
        RECT 15.715 40.085 16.005 40.315 ;
        RECT 15.790 39.250 15.930 40.085 ;
        RECT 16.160 40.070 16.480 40.330 ;
        RECT 16.710 40.315 16.850 40.470 ;
        RECT 18.015 40.425 18.305 40.470 ;
        RECT 18.920 40.610 19.240 40.670 ;
        RECT 20.760 40.610 21.080 40.670 ;
        RECT 21.695 40.610 21.985 40.655 ;
        RECT 27.200 40.610 27.520 40.670 ;
        RECT 28.135 40.610 28.425 40.655 ;
        RECT 18.920 40.470 20.530 40.610 ;
        RECT 18.920 40.410 19.240 40.470 ;
        RECT 16.635 40.085 16.925 40.315 ;
        RECT 17.555 40.085 17.845 40.315 ;
        RECT 19.380 40.270 19.700 40.330 ;
        RECT 20.390 40.315 20.530 40.470 ;
        RECT 20.760 40.470 21.985 40.610 ;
        RECT 20.760 40.410 21.080 40.470 ;
        RECT 21.695 40.425 21.985 40.470 ;
        RECT 22.230 40.470 25.590 40.610 ;
        RECT 19.855 40.270 20.145 40.315 ;
        RECT 19.380 40.130 20.145 40.270 ;
        RECT 16.250 39.590 16.390 40.070 ;
        RECT 17.630 39.930 17.770 40.085 ;
        RECT 19.380 40.070 19.700 40.130 ;
        RECT 19.855 40.085 20.145 40.130 ;
        RECT 20.315 40.085 20.605 40.315 ;
        RECT 21.220 40.070 21.540 40.330 ;
        RECT 22.230 40.315 22.370 40.470 ;
        RECT 22.230 40.130 22.565 40.315 ;
        RECT 25.450 40.270 25.590 40.470 ;
        RECT 27.200 40.470 28.425 40.610 ;
        RECT 27.200 40.410 27.520 40.470 ;
        RECT 28.135 40.425 28.425 40.470 ;
        RECT 29.040 40.610 29.360 40.670 ;
        RECT 37.320 40.610 37.640 40.670 ;
        RECT 29.040 40.470 33.870 40.610 ;
        RECT 29.040 40.410 29.360 40.470 ;
        RECT 25.450 40.130 27.430 40.270 ;
        RECT 22.275 40.085 22.565 40.130 ;
        RECT 24.900 39.930 25.220 39.990 ;
        RECT 17.630 39.790 25.220 39.930 ;
        RECT 27.290 39.930 27.430 40.130 ;
        RECT 27.660 40.070 27.980 40.330 ;
        RECT 28.595 40.270 28.885 40.315 ;
        RECT 29.500 40.270 29.820 40.330 ;
        RECT 28.595 40.130 29.820 40.270 ;
        RECT 28.595 40.085 28.885 40.130 ;
        RECT 29.500 40.070 29.820 40.130 ;
        RECT 31.355 40.085 31.645 40.315 ;
        RECT 32.275 40.270 32.565 40.315 ;
        RECT 33.180 40.270 33.500 40.330 ;
        RECT 32.275 40.130 33.500 40.270 ;
        RECT 33.730 40.270 33.870 40.470 ;
        RECT 37.320 40.470 41.690 40.610 ;
        RECT 37.320 40.410 37.640 40.470 ;
        RECT 41.550 40.315 41.690 40.470 ;
        RECT 52.960 40.410 53.280 40.670 ;
        RECT 59.490 40.610 59.630 40.810 ;
        RECT 63.080 40.750 63.400 40.810 ;
        RECT 64.000 40.750 64.320 41.010 ;
        RECT 82.415 40.765 82.705 40.995 ;
        RECT 54.430 40.470 59.630 40.610 ;
        RECT 59.875 40.610 60.165 40.655 ;
        RECT 67.680 40.610 68.000 40.670 ;
        RECT 59.875 40.470 68.000 40.610 ;
        RECT 41.015 40.270 41.305 40.315 ;
        RECT 33.730 40.130 41.305 40.270 ;
        RECT 32.275 40.085 32.565 40.130 ;
        RECT 31.430 39.930 31.570 40.085 ;
        RECT 33.180 40.070 33.500 40.130 ;
        RECT 41.015 40.085 41.305 40.130 ;
        RECT 41.475 40.085 41.765 40.315 ;
        RECT 42.380 40.070 42.700 40.330 ;
        RECT 42.855 40.270 43.145 40.315 ;
        RECT 54.430 40.270 54.570 40.470 ;
        RECT 59.875 40.425 60.165 40.470 ;
        RECT 67.680 40.410 68.000 40.470 ;
        RECT 69.980 40.610 70.300 40.670 ;
        RECT 82.490 40.610 82.630 40.765 ;
        RECT 69.980 40.470 73.890 40.610 ;
        RECT 69.980 40.410 70.300 40.470 ;
        RECT 42.855 40.130 54.570 40.270 ;
        RECT 54.815 40.270 55.105 40.315 ;
        RECT 55.720 40.270 56.040 40.330 ;
        RECT 60.780 40.270 61.100 40.330 ;
        RECT 54.815 40.130 61.100 40.270 ;
        RECT 42.855 40.085 43.145 40.130 ;
        RECT 54.815 40.085 55.105 40.130 ;
        RECT 55.720 40.070 56.040 40.130 ;
        RECT 60.780 40.070 61.100 40.130 ;
        RECT 61.240 40.070 61.560 40.330 ;
        RECT 65.380 40.070 65.700 40.330 ;
        RECT 65.855 40.085 66.145 40.315 ;
        RECT 66.315 40.085 66.605 40.315 ;
        RECT 33.640 39.930 33.960 39.990 ;
        RECT 27.290 39.790 33.960 39.930 ;
        RECT 24.900 39.730 25.220 39.790 ;
        RECT 33.640 39.730 33.960 39.790 ;
        RECT 48.360 39.930 48.680 39.990 ;
        RECT 48.835 39.930 49.125 39.975 ;
        RECT 48.360 39.790 49.125 39.930 ;
        RECT 48.360 39.730 48.680 39.790 ;
        RECT 48.835 39.745 49.125 39.790 ;
        RECT 49.740 39.730 50.060 39.990 ;
        RECT 56.195 39.930 56.485 39.975 ;
        RECT 57.100 39.930 57.420 39.990 ;
        RECT 56.195 39.790 57.420 39.930 ;
        RECT 56.195 39.745 56.485 39.790 ;
        RECT 57.100 39.730 57.420 39.790 ;
        RECT 59.860 39.930 60.180 39.990 ;
        RECT 60.335 39.930 60.625 39.975 ;
        RECT 65.930 39.930 66.070 40.085 ;
        RECT 59.860 39.790 60.625 39.930 ;
        RECT 59.860 39.730 60.180 39.790 ;
        RECT 60.335 39.745 60.625 39.790 ;
        RECT 60.870 39.790 66.070 39.930 ;
        RECT 66.390 39.930 66.530 40.085 ;
        RECT 67.220 40.070 67.540 40.330 ;
        RECT 68.140 40.070 68.460 40.330 ;
        RECT 69.075 40.270 69.365 40.315 ;
        RECT 69.520 40.270 69.840 40.330 ;
        RECT 70.530 40.315 70.670 40.470 ;
        RECT 69.075 40.130 69.840 40.270 ;
        RECT 69.075 40.085 69.365 40.130 ;
        RECT 69.520 40.070 69.840 40.130 ;
        RECT 70.455 40.085 70.745 40.315 ;
        RECT 70.900 40.270 71.220 40.330 ;
        RECT 73.750 40.315 73.890 40.470 ;
        RECT 78.810 40.470 82.630 40.610 ;
        RECT 71.375 40.270 71.665 40.315 ;
        RECT 72.755 40.270 73.045 40.315 ;
        RECT 70.900 40.130 73.045 40.270 ;
        RECT 70.900 40.070 71.220 40.130 ;
        RECT 71.375 40.085 71.665 40.130 ;
        RECT 72.755 40.085 73.045 40.130 ;
        RECT 73.675 40.270 73.965 40.315 ;
        RECT 74.120 40.270 74.440 40.330 ;
        RECT 73.675 40.130 74.440 40.270 ;
        RECT 73.675 40.085 73.965 40.130 ;
        RECT 74.120 40.070 74.440 40.130 ;
        RECT 77.800 40.270 78.120 40.330 ;
        RECT 78.810 40.315 78.950 40.470 ;
        RECT 78.735 40.270 79.025 40.315 ;
        RECT 77.800 40.130 79.025 40.270 ;
        RECT 77.800 40.070 78.120 40.130 ;
        RECT 78.735 40.085 79.025 40.130 ;
        RECT 79.640 40.070 79.960 40.330 ;
        RECT 80.115 40.085 80.405 40.315 ;
        RECT 80.575 40.270 80.865 40.315 ;
        RECT 81.020 40.270 81.340 40.330 ;
        RECT 80.575 40.130 81.340 40.270 ;
        RECT 80.575 40.085 80.865 40.130 ;
        RECT 69.995 39.930 70.285 39.975 ;
        RECT 66.390 39.790 70.285 39.930 ;
        RECT 40.095 39.590 40.385 39.635 ;
        RECT 59.400 39.590 59.720 39.650 ;
        RECT 16.250 39.450 39.850 39.590 ;
        RECT 19.840 39.250 20.160 39.310 ;
        RECT 21.220 39.250 21.540 39.310 ;
        RECT 15.790 39.110 21.540 39.250 ;
        RECT 19.840 39.050 20.160 39.110 ;
        RECT 21.220 39.050 21.540 39.110 ;
        RECT 29.500 39.250 29.820 39.310 ;
        RECT 30.435 39.250 30.725 39.295 ;
        RECT 29.500 39.110 30.725 39.250 ;
        RECT 39.710 39.250 39.850 39.450 ;
        RECT 40.095 39.450 59.720 39.590 ;
        RECT 40.095 39.405 40.385 39.450 ;
        RECT 59.400 39.390 59.720 39.450 ;
        RECT 49.280 39.250 49.600 39.310 ;
        RECT 39.710 39.110 49.600 39.250 ;
        RECT 29.500 39.050 29.820 39.110 ;
        RECT 30.435 39.065 30.725 39.110 ;
        RECT 49.280 39.050 49.600 39.110 ;
        RECT 51.120 39.050 51.440 39.310 ;
        RECT 51.580 39.250 51.900 39.310 ;
        RECT 52.055 39.250 52.345 39.295 ;
        RECT 51.580 39.110 52.345 39.250 ;
        RECT 51.580 39.050 51.900 39.110 ;
        RECT 52.055 39.065 52.345 39.110 ;
        RECT 58.940 39.250 59.260 39.310 ;
        RECT 60.870 39.250 61.010 39.790 ;
        RECT 69.995 39.745 70.285 39.790 ;
        RECT 71.820 39.930 72.140 39.990 ;
        RECT 78.260 39.930 78.580 39.990 ;
        RECT 80.190 39.930 80.330 40.085 ;
        RECT 81.020 40.070 81.340 40.130 ;
        RECT 83.320 40.070 83.640 40.330 ;
        RECT 71.820 39.790 80.330 39.930 ;
        RECT 71.820 39.730 72.140 39.790 ;
        RECT 78.260 39.730 78.580 39.790 ;
        RECT 68.140 39.590 68.460 39.650 ;
        RECT 78.720 39.590 79.040 39.650 ;
        RECT 62.250 39.450 68.460 39.590 ;
        RECT 58.940 39.110 61.010 39.250 ;
        RECT 61.700 39.250 62.020 39.310 ;
        RECT 62.250 39.295 62.390 39.450 ;
        RECT 68.140 39.390 68.460 39.450 ;
        RECT 70.530 39.450 79.040 39.590 ;
        RECT 62.175 39.250 62.465 39.295 ;
        RECT 61.700 39.110 62.465 39.250 ;
        RECT 58.940 39.050 59.260 39.110 ;
        RECT 61.700 39.050 62.020 39.110 ;
        RECT 62.175 39.065 62.465 39.110 ;
        RECT 65.380 39.250 65.700 39.310 ;
        RECT 70.530 39.250 70.670 39.450 ;
        RECT 78.720 39.390 79.040 39.450 ;
        RECT 81.955 39.590 82.245 39.635 ;
        RECT 83.320 39.590 83.640 39.650 ;
        RECT 81.955 39.450 83.640 39.590 ;
        RECT 81.955 39.405 82.245 39.450 ;
        RECT 83.320 39.390 83.640 39.450 ;
        RECT 65.380 39.110 70.670 39.250 ;
        RECT 65.380 39.050 65.700 39.110 ;
        RECT 70.900 39.050 71.220 39.310 ;
        RECT 73.660 39.250 73.980 39.310 ;
        RECT 74.595 39.250 74.885 39.295 ;
        RECT 73.660 39.110 74.885 39.250 ;
        RECT 73.660 39.050 73.980 39.110 ;
        RECT 74.595 39.065 74.885 39.110 ;
        RECT 11.950 38.430 90.610 38.910 ;
        RECT 20.300 38.230 20.620 38.290 ;
        RECT 21.680 38.230 22.000 38.290 ;
        RECT 33.655 38.230 33.945 38.275 ;
        RECT 20.300 38.090 22.000 38.230 ;
        RECT 20.300 38.030 20.620 38.090 ;
        RECT 21.680 38.030 22.000 38.090 ;
        RECT 29.590 38.090 33.945 38.230 ;
        RECT 17.120 37.890 17.410 37.935 ;
        RECT 19.220 37.890 19.510 37.935 ;
        RECT 20.790 37.890 21.080 37.935 ;
        RECT 17.120 37.750 21.080 37.890 ;
        RECT 17.120 37.705 17.410 37.750 ;
        RECT 19.220 37.705 19.510 37.750 ;
        RECT 20.790 37.705 21.080 37.750 ;
        RECT 15.240 37.550 15.560 37.610 ;
        RECT 16.620 37.550 16.940 37.610 ;
        RECT 15.240 37.410 16.940 37.550 ;
        RECT 15.240 37.350 15.560 37.410 ;
        RECT 16.620 37.350 16.940 37.410 ;
        RECT 17.515 37.550 17.805 37.595 ;
        RECT 18.705 37.550 18.995 37.595 ;
        RECT 21.225 37.550 21.515 37.595 ;
        RECT 17.515 37.410 21.515 37.550 ;
        RECT 29.590 37.550 29.730 38.090 ;
        RECT 29.590 37.410 30.190 37.550 ;
        RECT 17.515 37.365 17.805 37.410 ;
        RECT 18.705 37.365 18.995 37.410 ;
        RECT 21.225 37.365 21.515 37.410 ;
        RECT 25.360 37.210 25.680 37.270 ;
        RECT 28.580 37.210 28.900 37.270 ;
        RECT 25.360 37.070 28.900 37.210 ;
        RECT 25.360 37.010 25.680 37.070 ;
        RECT 28.580 37.010 28.900 37.070 ;
        RECT 29.040 37.210 29.360 37.270 ;
        RECT 30.050 37.255 30.190 37.410 ;
        RECT 33.270 37.270 33.410 38.090 ;
        RECT 33.655 38.045 33.945 38.090 ;
        RECT 53.880 38.030 54.200 38.290 ;
        RECT 75.975 38.230 76.265 38.275 ;
        RECT 79.640 38.230 79.960 38.290 ;
        RECT 75.975 38.090 79.960 38.230 ;
        RECT 75.975 38.045 76.265 38.090 ;
        RECT 79.640 38.030 79.960 38.090 ;
        RECT 39.160 37.890 39.450 37.935 ;
        RECT 40.730 37.890 41.020 37.935 ;
        RECT 42.830 37.890 43.120 37.935 ;
        RECT 39.160 37.750 43.120 37.890 ;
        RECT 39.160 37.705 39.450 37.750 ;
        RECT 40.730 37.705 41.020 37.750 ;
        RECT 42.830 37.705 43.120 37.750 ;
        RECT 48.360 37.890 48.680 37.950 ;
        RECT 73.200 37.890 73.520 37.950 ;
        RECT 48.360 37.750 73.520 37.890 ;
        RECT 48.360 37.690 48.680 37.750 ;
        RECT 73.200 37.690 73.520 37.750 ;
        RECT 81.980 37.890 82.270 37.935 ;
        RECT 84.080 37.890 84.370 37.935 ;
        RECT 85.650 37.890 85.940 37.935 ;
        RECT 81.980 37.750 85.940 37.890 ;
        RECT 81.980 37.705 82.270 37.750 ;
        RECT 84.080 37.705 84.370 37.750 ;
        RECT 85.650 37.705 85.940 37.750 ;
        RECT 38.725 37.550 39.015 37.595 ;
        RECT 41.245 37.550 41.535 37.595 ;
        RECT 42.435 37.550 42.725 37.595 ;
        RECT 38.725 37.410 42.725 37.550 ;
        RECT 38.725 37.365 39.015 37.410 ;
        RECT 41.245 37.365 41.535 37.410 ;
        RECT 42.435 37.365 42.725 37.410 ;
        RECT 49.740 37.550 50.060 37.610 ;
        RECT 56.655 37.550 56.945 37.595 ;
        RECT 49.740 37.410 56.945 37.550 ;
        RECT 49.740 37.350 50.060 37.410 ;
        RECT 56.655 37.365 56.945 37.410 ;
        RECT 60.780 37.350 61.100 37.610 ;
        RECT 81.020 37.550 81.340 37.610 ;
        RECT 79.730 37.410 81.340 37.550 ;
        RECT 29.515 37.210 29.805 37.255 ;
        RECT 29.040 37.070 29.805 37.210 ;
        RECT 29.040 37.010 29.360 37.070 ;
        RECT 29.515 37.025 29.805 37.070 ;
        RECT 29.975 37.025 30.265 37.255 ;
        RECT 30.420 37.010 30.740 37.270 ;
        RECT 32.720 37.010 33.040 37.270 ;
        RECT 33.180 37.010 33.500 37.270 ;
        RECT 33.640 37.210 33.960 37.270 ;
        RECT 34.115 37.210 34.405 37.255 ;
        RECT 39.160 37.210 39.480 37.270 ;
        RECT 43.300 37.210 43.620 37.270 ;
        RECT 33.640 37.070 39.480 37.210 ;
        RECT 33.640 37.010 33.960 37.070 ;
        RECT 34.115 37.025 34.405 37.070 ;
        RECT 39.160 37.010 39.480 37.070 ;
        RECT 41.090 37.070 43.620 37.210 ;
        RECT 17.970 36.870 18.260 36.915 ;
        RECT 19.840 36.870 20.160 36.930 ;
        RECT 26.295 36.870 26.585 36.915 ;
        RECT 17.970 36.730 20.160 36.870 ;
        RECT 17.970 36.685 18.260 36.730 ;
        RECT 19.840 36.670 20.160 36.730 ;
        RECT 23.610 36.730 26.585 36.870 ;
        RECT 20.760 36.530 21.080 36.590 ;
        RECT 23.610 36.575 23.750 36.730 ;
        RECT 26.295 36.685 26.585 36.730 ;
        RECT 27.200 36.670 27.520 36.930 ;
        RECT 30.510 36.870 30.650 37.010 ;
        RECT 41.090 36.930 41.230 37.070 ;
        RECT 43.300 37.010 43.620 37.070 ;
        RECT 45.155 37.025 45.445 37.255 ;
        RECT 30.510 36.730 37.090 36.870 ;
        RECT 23.535 36.530 23.825 36.575 ;
        RECT 20.760 36.390 23.825 36.530 ;
        RECT 20.760 36.330 21.080 36.390 ;
        RECT 23.535 36.345 23.825 36.390 ;
        RECT 25.360 36.330 25.680 36.590 ;
        RECT 27.290 36.530 27.430 36.670 ;
        RECT 29.500 36.530 29.820 36.590 ;
        RECT 27.290 36.390 29.820 36.530 ;
        RECT 29.500 36.330 29.820 36.390 ;
        RECT 29.960 36.530 30.280 36.590 ;
        RECT 31.815 36.530 32.105 36.575 ;
        RECT 29.960 36.390 32.105 36.530 ;
        RECT 29.960 36.330 30.280 36.390 ;
        RECT 31.815 36.345 32.105 36.390 ;
        RECT 36.400 36.330 36.720 36.590 ;
        RECT 36.950 36.530 37.090 36.730 ;
        RECT 41.000 36.670 41.320 36.930 ;
        RECT 42.090 36.870 42.380 36.915 ;
        RECT 43.775 36.870 44.065 36.915 ;
        RECT 42.090 36.730 44.065 36.870 ;
        RECT 42.090 36.685 42.380 36.730 ;
        RECT 43.775 36.685 44.065 36.730 ;
        RECT 45.230 36.870 45.370 37.025 ;
        RECT 45.600 37.010 45.920 37.270 ;
        RECT 46.060 37.010 46.380 37.270 ;
        RECT 46.520 37.210 46.840 37.270 ;
        RECT 46.995 37.210 47.285 37.255 ;
        RECT 65.380 37.210 65.700 37.270 ;
        RECT 46.520 37.070 47.285 37.210 ;
        RECT 46.520 37.010 46.840 37.070 ;
        RECT 46.995 37.025 47.285 37.070 ;
        RECT 55.350 37.070 65.700 37.210 ;
        RECT 55.350 36.870 55.490 37.070 ;
        RECT 65.380 37.010 65.700 37.070 ;
        RECT 77.800 37.010 78.120 37.270 ;
        RECT 78.720 37.010 79.040 37.270 ;
        RECT 79.730 37.255 79.870 37.410 ;
        RECT 81.020 37.350 81.340 37.410 ;
        RECT 82.375 37.550 82.665 37.595 ;
        RECT 83.565 37.550 83.855 37.595 ;
        RECT 86.085 37.550 86.375 37.595 ;
        RECT 82.375 37.410 86.375 37.550 ;
        RECT 82.375 37.365 82.665 37.410 ;
        RECT 83.565 37.365 83.855 37.410 ;
        RECT 86.085 37.365 86.375 37.410 ;
        RECT 79.195 37.025 79.485 37.255 ;
        RECT 79.655 37.025 79.945 37.255 ;
        RECT 81.495 37.210 81.785 37.255 ;
        RECT 81.940 37.210 82.260 37.270 ;
        RECT 81.495 37.070 82.260 37.210 ;
        RECT 81.495 37.025 81.785 37.070 ;
        RECT 45.230 36.730 55.490 36.870 ;
        RECT 55.735 36.870 56.025 36.915 ;
        RECT 58.035 36.870 58.325 36.915 ;
        RECT 55.735 36.730 58.325 36.870 ;
        RECT 45.230 36.530 45.370 36.730 ;
        RECT 55.735 36.685 56.025 36.730 ;
        RECT 58.035 36.685 58.325 36.730 ;
        RECT 62.160 36.670 62.480 36.930 ;
        RECT 73.660 36.870 73.980 36.930 ;
        RECT 74.135 36.870 74.425 36.915 ;
        RECT 73.660 36.730 74.425 36.870 ;
        RECT 73.660 36.670 73.980 36.730 ;
        RECT 74.135 36.685 74.425 36.730 ;
        RECT 75.055 36.870 75.345 36.915 ;
        RECT 78.260 36.870 78.580 36.930 ;
        RECT 75.055 36.730 78.580 36.870 ;
        RECT 75.055 36.685 75.345 36.730 ;
        RECT 78.260 36.670 78.580 36.730 ;
        RECT 36.950 36.390 45.370 36.530 ;
        RECT 56.195 36.530 56.485 36.575 ;
        RECT 56.640 36.530 56.960 36.590 ;
        RECT 56.195 36.390 56.960 36.530 ;
        RECT 56.195 36.345 56.485 36.390 ;
        RECT 56.640 36.330 56.960 36.390 ;
        RECT 62.620 36.330 62.940 36.590 ;
        RECT 72.740 36.530 73.060 36.590 ;
        RECT 79.270 36.530 79.410 37.025 ;
        RECT 81.940 37.010 82.260 37.070 ;
        RECT 81.035 36.870 81.325 36.915 ;
        RECT 82.720 36.870 83.010 36.915 ;
        RECT 81.035 36.730 83.010 36.870 ;
        RECT 81.035 36.685 81.325 36.730 ;
        RECT 82.720 36.685 83.010 36.730 ;
        RECT 72.740 36.390 79.410 36.530 ;
        RECT 85.620 36.530 85.940 36.590 ;
        RECT 88.395 36.530 88.685 36.575 ;
        RECT 85.620 36.390 88.685 36.530 ;
        RECT 72.740 36.330 73.060 36.390 ;
        RECT 85.620 36.330 85.940 36.390 ;
        RECT 88.395 36.345 88.685 36.390 ;
        RECT 11.950 35.710 90.610 36.190 ;
        RECT 19.840 35.310 20.160 35.570 ;
        RECT 29.040 35.310 29.360 35.570 ;
        RECT 29.500 35.510 29.820 35.570 ;
        RECT 32.720 35.510 33.040 35.570 ;
        RECT 29.500 35.370 33.040 35.510 ;
        RECT 29.500 35.310 29.820 35.370 ;
        RECT 32.720 35.310 33.040 35.370 ;
        RECT 41.015 35.510 41.305 35.555 ;
        RECT 41.460 35.510 41.780 35.570 ;
        RECT 41.015 35.370 41.780 35.510 ;
        RECT 41.015 35.325 41.305 35.370 ;
        RECT 41.460 35.310 41.780 35.370 ;
        RECT 43.315 35.510 43.605 35.555 ;
        RECT 46.060 35.510 46.380 35.570 ;
        RECT 43.315 35.370 46.380 35.510 ;
        RECT 43.315 35.325 43.605 35.370 ;
        RECT 46.060 35.310 46.380 35.370 ;
        RECT 49.740 35.510 50.060 35.570 ;
        RECT 51.595 35.510 51.885 35.555 ;
        RECT 62.160 35.510 62.480 35.570 ;
        RECT 49.740 35.370 62.480 35.510 ;
        RECT 49.740 35.310 50.060 35.370 ;
        RECT 51.595 35.325 51.885 35.370 ;
        RECT 62.160 35.310 62.480 35.370 ;
        RECT 65.840 35.510 66.160 35.570 ;
        RECT 77.355 35.510 77.645 35.555 ;
        RECT 78.720 35.510 79.040 35.570 ;
        RECT 87.460 35.510 87.780 35.570 ;
        RECT 88.855 35.510 89.145 35.555 ;
        RECT 65.840 35.370 74.350 35.510 ;
        RECT 65.840 35.310 66.160 35.370 ;
        RECT 74.210 35.230 74.350 35.370 ;
        RECT 77.355 35.370 79.040 35.510 ;
        RECT 77.355 35.325 77.645 35.370 ;
        RECT 78.720 35.310 79.040 35.370 ;
        RECT 79.270 35.370 89.145 35.510 ;
        RECT 25.360 35.170 25.680 35.230 ;
        RECT 28.580 35.170 28.900 35.230 ;
        RECT 33.640 35.170 33.960 35.230 ;
        RECT 22.230 35.030 25.680 35.170 ;
        RECT 21.220 34.630 21.540 34.890 ;
        RECT 21.680 34.630 22.000 34.890 ;
        RECT 22.230 34.875 22.370 35.030 ;
        RECT 25.360 34.970 25.680 35.030 ;
        RECT 25.910 35.030 28.900 35.170 ;
        RECT 22.155 34.645 22.445 34.875 ;
        RECT 23.075 34.645 23.365 34.875 ;
        RECT 23.535 34.830 23.825 34.875 ;
        RECT 25.910 34.830 26.050 35.030 ;
        RECT 28.580 34.970 28.900 35.030 ;
        RECT 29.590 35.030 33.960 35.170 ;
        RECT 23.535 34.690 26.050 34.830 ;
        RECT 23.535 34.645 23.825 34.690 ;
        RECT 23.150 34.490 23.290 34.645 ;
        RECT 27.200 34.630 27.520 34.890 ;
        RECT 29.590 34.875 29.730 35.030 ;
        RECT 33.640 34.970 33.960 35.030 ;
        RECT 36.400 35.170 36.720 35.230 ;
        RECT 39.635 35.170 39.925 35.215 ;
        RECT 42.395 35.170 42.685 35.215 ;
        RECT 36.400 35.030 42.685 35.170 ;
        RECT 36.400 34.970 36.720 35.030 ;
        RECT 39.635 34.985 39.925 35.030 ;
        RECT 42.395 34.985 42.685 35.030 ;
        RECT 54.340 35.170 54.660 35.230 ;
        RECT 68.140 35.170 68.460 35.230 ;
        RECT 54.340 35.030 68.460 35.170 ;
        RECT 54.340 34.970 54.660 35.030 ;
        RECT 68.140 34.970 68.460 35.030 ;
        RECT 74.120 35.170 74.440 35.230 ;
        RECT 78.260 35.170 78.580 35.230 ;
        RECT 79.270 35.215 79.410 35.370 ;
        RECT 87.460 35.310 87.780 35.370 ;
        RECT 88.855 35.325 89.145 35.370 ;
        RECT 83.320 35.215 83.640 35.230 ;
        RECT 79.195 35.170 79.485 35.215 ;
        RECT 83.290 35.170 83.640 35.215 ;
        RECT 74.120 35.030 77.110 35.170 ;
        RECT 74.120 34.970 74.440 35.030 ;
        RECT 28.135 34.830 28.425 34.875 ;
        RECT 28.135 34.690 29.270 34.830 ;
        RECT 28.135 34.645 28.425 34.690 ;
        RECT 23.150 34.350 24.670 34.490 ;
        RECT 24.530 33.855 24.670 34.350 ;
        RECT 24.455 33.810 24.745 33.855 ;
        RECT 25.820 33.810 26.140 33.870 ;
        RECT 24.455 33.670 26.140 33.810 ;
        RECT 29.130 33.810 29.270 34.690 ;
        RECT 29.515 34.645 29.805 34.875 ;
        RECT 29.960 34.830 30.280 34.890 ;
        RECT 30.795 34.830 31.085 34.875 ;
        RECT 38.255 34.830 38.545 34.875 ;
        RECT 29.960 34.690 31.085 34.830 ;
        RECT 29.960 34.630 30.280 34.690 ;
        RECT 30.795 34.645 31.085 34.690 ;
        RECT 36.490 34.690 38.545 34.830 ;
        RECT 30.395 34.490 30.685 34.535 ;
        RECT 31.585 34.490 31.875 34.535 ;
        RECT 34.105 34.490 34.395 34.535 ;
        RECT 30.395 34.350 34.395 34.490 ;
        RECT 30.395 34.305 30.685 34.350 ;
        RECT 31.585 34.305 31.875 34.350 ;
        RECT 34.105 34.305 34.395 34.350 ;
        RECT 30.000 34.150 30.290 34.195 ;
        RECT 32.100 34.150 32.390 34.195 ;
        RECT 33.670 34.150 33.960 34.195 ;
        RECT 30.000 34.010 33.960 34.150 ;
        RECT 30.000 33.965 30.290 34.010 ;
        RECT 32.100 33.965 32.390 34.010 ;
        RECT 33.670 33.965 33.960 34.010 ;
        RECT 30.420 33.810 30.740 33.870 ;
        RECT 36.490 33.855 36.630 34.690 ;
        RECT 38.255 34.645 38.545 34.690 ;
        RECT 39.160 34.630 39.480 34.890 ;
        RECT 40.095 34.645 40.385 34.875 ;
        RECT 39.250 34.150 39.390 34.630 ;
        RECT 40.170 34.490 40.310 34.645 ;
        RECT 41.460 34.630 41.780 34.890 ;
        RECT 50.660 34.830 50.980 34.890 ;
        RECT 51.135 34.830 51.425 34.875 ;
        RECT 50.660 34.690 51.425 34.830 ;
        RECT 50.660 34.630 50.980 34.690 ;
        RECT 51.135 34.645 51.425 34.690 ;
        RECT 51.580 34.830 51.900 34.890 ;
        RECT 52.515 34.830 52.805 34.875 ;
        RECT 51.580 34.690 52.805 34.830 ;
        RECT 51.580 34.630 51.900 34.690 ;
        RECT 52.515 34.645 52.805 34.690 ;
        RECT 53.420 34.630 53.740 34.890 ;
        RECT 55.720 34.830 56.040 34.890 ;
        RECT 57.475 34.830 57.765 34.875 ;
        RECT 55.720 34.690 57.765 34.830 ;
        RECT 55.720 34.630 56.040 34.690 ;
        RECT 57.475 34.645 57.765 34.690 ;
        RECT 62.620 34.830 62.940 34.890 ;
        RECT 69.535 34.830 69.825 34.875 ;
        RECT 70.915 34.830 71.205 34.875 ;
        RECT 62.620 34.690 71.205 34.830 ;
        RECT 62.620 34.630 62.940 34.690 ;
        RECT 41.920 34.490 42.240 34.550 ;
        RECT 40.170 34.350 42.240 34.490 ;
        RECT 41.920 34.290 42.240 34.350 ;
        RECT 56.195 34.305 56.485 34.535 ;
        RECT 57.075 34.490 57.365 34.535 ;
        RECT 58.265 34.490 58.555 34.535 ;
        RECT 60.785 34.490 61.075 34.535 ;
        RECT 57.075 34.350 61.075 34.490 ;
        RECT 57.075 34.305 57.365 34.350 ;
        RECT 58.265 34.305 58.555 34.350 ;
        RECT 60.785 34.305 61.075 34.350 ;
        RECT 51.120 34.150 51.440 34.210 ;
        RECT 39.250 34.010 51.440 34.150 ;
        RECT 51.120 33.950 51.440 34.010 ;
        RECT 36.415 33.810 36.705 33.855 ;
        RECT 29.130 33.670 36.705 33.810 ;
        RECT 56.270 33.810 56.410 34.305 ;
        RECT 56.680 34.150 56.970 34.195 ;
        RECT 58.780 34.150 59.070 34.195 ;
        RECT 60.350 34.150 60.640 34.195 ;
        RECT 56.680 34.010 60.640 34.150 ;
        RECT 56.680 33.965 56.970 34.010 ;
        RECT 58.780 33.965 59.070 34.010 ;
        RECT 60.350 33.965 60.640 34.010 ;
        RECT 57.100 33.810 57.420 33.870 ;
        RECT 56.270 33.670 57.420 33.810 ;
        RECT 24.455 33.625 24.745 33.670 ;
        RECT 25.820 33.610 26.140 33.670 ;
        RECT 30.420 33.610 30.740 33.670 ;
        RECT 36.415 33.625 36.705 33.670 ;
        RECT 57.100 33.610 57.420 33.670 ;
        RECT 57.560 33.810 57.880 33.870 ;
        RECT 63.095 33.810 63.385 33.855 ;
        RECT 63.540 33.810 63.860 33.870 ;
        RECT 57.560 33.670 63.860 33.810 ;
        RECT 68.230 33.810 68.370 34.690 ;
        RECT 69.535 34.645 69.825 34.690 ;
        RECT 70.915 34.645 71.205 34.690 ;
        RECT 71.835 34.645 72.125 34.875 ;
        RECT 75.515 34.645 75.805 34.875 ;
        RECT 75.960 34.830 76.280 34.890 ;
        RECT 76.435 34.830 76.725 34.875 ;
        RECT 75.960 34.690 76.725 34.830 ;
        RECT 76.970 34.830 77.110 35.030 ;
        RECT 78.260 35.030 79.485 35.170 ;
        RECT 83.125 35.030 83.640 35.170 ;
        RECT 78.260 34.970 78.580 35.030 ;
        RECT 79.195 34.985 79.485 35.030 ;
        RECT 83.290 34.985 83.640 35.030 ;
        RECT 83.320 34.970 83.640 34.985 ;
        RECT 78.720 34.830 79.040 34.890 ;
        RECT 76.970 34.690 79.040 34.830 ;
        RECT 70.440 34.490 70.760 34.550 ;
        RECT 71.910 34.490 72.050 34.645 ;
        RECT 70.440 34.350 72.050 34.490 ;
        RECT 70.440 34.290 70.760 34.350 ;
        RECT 72.740 34.290 73.060 34.550 ;
        RECT 75.590 34.210 75.730 34.645 ;
        RECT 75.960 34.630 76.280 34.690 ;
        RECT 76.435 34.645 76.725 34.690 ;
        RECT 78.720 34.630 79.040 34.690 ;
        RECT 79.640 34.630 79.960 34.890 ;
        RECT 80.560 34.830 80.880 34.890 ;
        RECT 85.620 34.830 85.940 34.890 ;
        RECT 80.560 34.690 85.940 34.830 ;
        RECT 80.560 34.630 80.880 34.690 ;
        RECT 85.620 34.630 85.940 34.690 ;
        RECT 81.940 34.290 82.260 34.550 ;
        RECT 82.835 34.490 83.125 34.535 ;
        RECT 84.025 34.490 84.315 34.535 ;
        RECT 86.545 34.490 86.835 34.535 ;
        RECT 82.835 34.350 86.835 34.490 ;
        RECT 82.835 34.305 83.125 34.350 ;
        RECT 84.025 34.305 84.315 34.350 ;
        RECT 86.545 34.305 86.835 34.350 ;
        RECT 68.615 34.150 68.905 34.195 ;
        RECT 75.500 34.150 75.820 34.210 ;
        RECT 68.615 34.010 75.820 34.150 ;
        RECT 68.615 33.965 68.905 34.010 ;
        RECT 75.500 33.950 75.820 34.010 ;
        RECT 76.420 34.150 76.740 34.210 ;
        RECT 77.815 34.150 78.105 34.195 ;
        RECT 76.420 34.010 78.105 34.150 ;
        RECT 76.420 33.950 76.740 34.010 ;
        RECT 77.815 33.965 78.105 34.010 ;
        RECT 78.720 34.150 79.040 34.210 ;
        RECT 81.020 34.150 81.340 34.210 ;
        RECT 78.720 34.010 81.340 34.150 ;
        RECT 78.720 33.950 79.040 34.010 ;
        RECT 81.020 33.950 81.340 34.010 ;
        RECT 82.440 34.150 82.730 34.195 ;
        RECT 84.540 34.150 84.830 34.195 ;
        RECT 86.110 34.150 86.400 34.195 ;
        RECT 82.440 34.010 86.400 34.150 ;
        RECT 82.440 33.965 82.730 34.010 ;
        RECT 84.540 33.965 84.830 34.010 ;
        RECT 86.110 33.965 86.400 34.010 ;
        RECT 79.640 33.810 79.960 33.870 ;
        RECT 68.230 33.670 79.960 33.810 ;
        RECT 57.560 33.610 57.880 33.670 ;
        RECT 63.095 33.625 63.385 33.670 ;
        RECT 63.540 33.610 63.860 33.670 ;
        RECT 79.640 33.610 79.960 33.670 ;
        RECT 11.950 32.990 90.610 33.470 ;
        RECT 20.160 32.650 49.970 32.790 ;
        RECT 17.540 32.450 17.860 32.510 ;
        RECT 19.380 32.450 19.700 32.510 ;
        RECT 20.160 32.450 20.300 32.650 ;
        RECT 17.540 32.310 20.300 32.450 ;
        RECT 21.680 32.450 22.000 32.510 ;
        RECT 21.680 32.310 22.370 32.450 ;
        RECT 17.540 32.250 17.860 32.310 ;
        RECT 19.380 32.250 19.700 32.310 ;
        RECT 21.680 32.250 22.000 32.310 ;
        RECT 20.760 32.110 21.080 32.170 ;
        RECT 14.870 31.970 21.080 32.110 ;
        RECT 14.870 31.815 15.010 31.970 ;
        RECT 20.760 31.910 21.080 31.970 ;
        RECT 22.230 32.110 22.370 32.310 ;
        RECT 41.460 32.250 41.780 32.510 ;
        RECT 49.830 32.450 49.970 32.650 ;
        RECT 50.200 32.590 50.520 32.850 ;
        RECT 55.720 32.590 56.040 32.850 ;
        RECT 67.310 32.650 75.270 32.790 ;
        RECT 58.980 32.450 59.270 32.495 ;
        RECT 61.080 32.450 61.370 32.495 ;
        RECT 62.650 32.450 62.940 32.495 ;
        RECT 49.830 32.310 56.870 32.450 ;
        RECT 33.180 32.110 33.500 32.170 ;
        RECT 41.550 32.110 41.690 32.250 ;
        RECT 48.360 32.110 48.680 32.170 ;
        RECT 50.660 32.110 50.980 32.170 ;
        RECT 56.195 32.110 56.485 32.155 ;
        RECT 22.230 31.970 33.500 32.110 ;
        RECT 14.795 31.585 15.085 31.815 ;
        RECT 15.240 31.770 15.560 31.830 ;
        RECT 17.540 31.770 17.860 31.830 ;
        RECT 15.240 31.630 17.860 31.770 ;
        RECT 15.240 31.570 15.560 31.630 ;
        RECT 17.540 31.570 17.860 31.630 ;
        RECT 18.000 31.770 18.320 31.830 ;
        RECT 22.230 31.815 22.370 31.970 ;
        RECT 33.180 31.910 33.500 31.970 ;
        RECT 41.090 31.970 48.680 32.110 ;
        RECT 21.695 31.770 21.985 31.815 ;
        RECT 18.000 31.630 21.985 31.770 ;
        RECT 18.000 31.570 18.320 31.630 ;
        RECT 21.695 31.585 21.985 31.630 ;
        RECT 22.155 31.585 22.445 31.815 ;
        RECT 22.600 31.570 22.920 31.830 ;
        RECT 23.535 31.770 23.825 31.815 ;
        RECT 23.980 31.770 24.300 31.830 ;
        RECT 25.820 31.770 26.140 31.830 ;
        RECT 23.535 31.630 26.140 31.770 ;
        RECT 23.535 31.585 23.825 31.630 ;
        RECT 23.980 31.570 24.300 31.630 ;
        RECT 25.820 31.570 26.140 31.630 ;
        RECT 16.635 31.430 16.925 31.475 ;
        RECT 17.080 31.430 17.400 31.490 ;
        RECT 16.635 31.290 17.400 31.430 ;
        RECT 41.090 31.430 41.230 31.970 ;
        RECT 48.360 31.910 48.680 31.970 ;
        RECT 48.910 31.970 50.980 32.110 ;
        RECT 41.460 31.770 41.780 31.830 ;
        RECT 47.455 31.770 47.745 31.815 ;
        RECT 41.460 31.630 47.745 31.770 ;
        RECT 41.460 31.570 41.780 31.630 ;
        RECT 47.455 31.585 47.745 31.630 ;
        RECT 42.855 31.430 43.145 31.475 ;
        RECT 41.090 31.290 43.145 31.430 ;
        RECT 16.635 31.245 16.925 31.290 ;
        RECT 17.080 31.230 17.400 31.290 ;
        RECT 42.855 31.245 43.145 31.290 ;
        RECT 43.775 31.430 44.065 31.475 ;
        RECT 44.220 31.430 44.540 31.490 ;
        RECT 48.910 31.475 49.050 31.970 ;
        RECT 50.660 31.910 50.980 31.970 ;
        RECT 53.510 31.970 56.485 32.110 ;
        RECT 49.295 31.770 49.585 31.815 ;
        RECT 50.200 31.770 50.520 31.830 ;
        RECT 49.295 31.630 50.520 31.770 ;
        RECT 49.295 31.585 49.585 31.630 ;
        RECT 50.200 31.570 50.520 31.630 ;
        RECT 52.500 31.570 52.820 31.830 ;
        RECT 53.510 31.815 53.650 31.970 ;
        RECT 56.195 31.925 56.485 31.970 ;
        RECT 53.435 31.585 53.725 31.815 ;
        RECT 53.895 31.585 54.185 31.815 ;
        RECT 43.775 31.290 44.540 31.430 ;
        RECT 43.775 31.245 44.065 31.290 ;
        RECT 44.220 31.230 44.540 31.290 ;
        RECT 48.375 31.245 48.665 31.475 ;
        RECT 48.835 31.245 49.125 31.475 ;
        RECT 49.740 31.430 50.060 31.490 ;
        RECT 53.970 31.430 54.110 31.585 ;
        RECT 54.340 31.570 54.660 31.830 ;
        RECT 56.730 31.770 56.870 32.310 ;
        RECT 58.980 32.310 62.940 32.450 ;
        RECT 58.980 32.265 59.270 32.310 ;
        RECT 61.080 32.265 61.370 32.310 ;
        RECT 62.650 32.265 62.940 32.310 ;
        RECT 57.100 32.110 57.420 32.170 ;
        RECT 58.495 32.110 58.785 32.155 ;
        RECT 57.100 31.970 58.785 32.110 ;
        RECT 57.100 31.910 57.420 31.970 ;
        RECT 58.495 31.925 58.785 31.970 ;
        RECT 59.375 32.110 59.665 32.155 ;
        RECT 60.565 32.110 60.855 32.155 ;
        RECT 63.085 32.110 63.375 32.155 ;
        RECT 59.375 31.970 63.375 32.110 ;
        RECT 59.375 31.925 59.665 31.970 ;
        RECT 60.565 31.925 60.855 31.970 ;
        RECT 63.085 31.925 63.375 31.970 ;
        RECT 58.035 31.770 58.325 31.815 ;
        RECT 61.700 31.770 62.020 31.830 ;
        RECT 62.620 31.770 62.940 31.830 ;
        RECT 56.730 31.630 62.940 31.770 ;
        RECT 58.035 31.585 58.325 31.630 ;
        RECT 61.700 31.570 62.020 31.630 ;
        RECT 62.620 31.570 62.940 31.630 ;
        RECT 66.300 31.770 66.620 31.830 ;
        RECT 66.775 31.770 67.065 31.815 ;
        RECT 67.310 31.770 67.450 32.650 ;
        RECT 75.130 32.495 75.270 32.650 ;
        RECT 68.640 32.450 68.930 32.495 ;
        RECT 70.740 32.450 71.030 32.495 ;
        RECT 72.310 32.450 72.600 32.495 ;
        RECT 68.640 32.310 72.600 32.450 ;
        RECT 68.640 32.265 68.930 32.310 ;
        RECT 70.740 32.265 71.030 32.310 ;
        RECT 72.310 32.265 72.600 32.310 ;
        RECT 75.055 32.450 75.345 32.495 ;
        RECT 82.400 32.450 82.720 32.510 ;
        RECT 75.055 32.310 82.720 32.450 ;
        RECT 75.055 32.265 75.345 32.310 ;
        RECT 82.400 32.250 82.720 32.310 ;
        RECT 69.035 32.110 69.325 32.155 ;
        RECT 70.225 32.110 70.515 32.155 ;
        RECT 72.745 32.110 73.035 32.155 ;
        RECT 69.035 31.970 73.035 32.110 ;
        RECT 69.035 31.925 69.325 31.970 ;
        RECT 70.225 31.925 70.515 31.970 ;
        RECT 72.745 31.925 73.035 31.970 ;
        RECT 66.300 31.630 67.450 31.770 ;
        RECT 68.155 31.770 68.445 31.815 ;
        RECT 71.820 31.770 72.140 31.830 ;
        RECT 68.155 31.630 72.140 31.770 ;
        RECT 66.300 31.570 66.620 31.630 ;
        RECT 66.775 31.585 67.065 31.630 ;
        RECT 68.155 31.585 68.445 31.630 ;
        RECT 71.820 31.570 72.140 31.630 ;
        RECT 87.460 31.570 87.780 31.830 ;
        RECT 49.740 31.290 54.110 31.430 ;
        RECT 13.875 31.090 14.165 31.135 ;
        RECT 14.320 31.090 14.640 31.150 ;
        RECT 13.875 30.950 14.640 31.090 ;
        RECT 13.875 30.905 14.165 30.950 ;
        RECT 14.320 30.890 14.640 30.950 ;
        RECT 15.715 31.090 16.005 31.135 ;
        RECT 16.160 31.090 16.480 31.150 ;
        RECT 15.715 30.950 16.480 31.090 ;
        RECT 15.715 30.905 16.005 30.950 ;
        RECT 16.160 30.890 16.480 30.950 ;
        RECT 20.300 30.890 20.620 31.150 ;
        RECT 44.680 30.890 45.000 31.150 ;
        RECT 48.450 31.090 48.590 31.245 ;
        RECT 49.740 31.230 50.060 31.290 ;
        RECT 51.120 31.090 51.440 31.150 ;
        RECT 48.450 30.950 51.440 31.090 ;
        RECT 53.970 31.090 54.110 31.290 ;
        RECT 56.180 31.430 56.500 31.490 ;
        RECT 57.115 31.430 57.405 31.475 ;
        RECT 57.560 31.430 57.880 31.490 ;
        RECT 56.180 31.290 57.880 31.430 ;
        RECT 56.180 31.230 56.500 31.290 ;
        RECT 57.115 31.245 57.405 31.290 ;
        RECT 57.560 31.230 57.880 31.290 ;
        RECT 58.480 31.430 58.800 31.490 ;
        RECT 59.720 31.430 60.010 31.475 ;
        RECT 58.480 31.290 60.010 31.430 ;
        RECT 58.480 31.230 58.800 31.290 ;
        RECT 59.720 31.245 60.010 31.290 ;
        RECT 67.695 31.430 67.985 31.475 ;
        RECT 69.490 31.430 69.780 31.475 ;
        RECT 71.360 31.430 71.680 31.490 ;
        RECT 67.695 31.290 69.290 31.430 ;
        RECT 67.695 31.245 67.985 31.290 ;
        RECT 58.940 31.090 59.260 31.150 ;
        RECT 53.970 30.950 59.260 31.090 ;
        RECT 51.120 30.890 51.440 30.950 ;
        RECT 58.940 30.890 59.260 30.950 ;
        RECT 61.700 31.090 62.020 31.150 ;
        RECT 65.395 31.090 65.685 31.135 ;
        RECT 61.700 30.950 65.685 31.090 ;
        RECT 61.700 30.890 62.020 30.950 ;
        RECT 65.395 30.905 65.685 30.950 ;
        RECT 65.855 31.090 66.145 31.135 ;
        RECT 68.600 31.090 68.920 31.150 ;
        RECT 65.855 30.950 68.920 31.090 ;
        RECT 69.150 31.090 69.290 31.290 ;
        RECT 69.490 31.290 71.680 31.430 ;
        RECT 69.490 31.245 69.780 31.290 ;
        RECT 71.360 31.230 71.680 31.290 ;
        RECT 73.660 31.430 73.980 31.490 ;
        RECT 77.355 31.430 77.645 31.475 ;
        RECT 73.660 31.290 77.645 31.430 ;
        RECT 73.660 31.230 73.980 31.290 ;
        RECT 77.355 31.245 77.645 31.290 ;
        RECT 78.260 31.230 78.580 31.490 ;
        RECT 73.750 31.090 73.890 31.230 ;
        RECT 69.150 30.950 73.890 31.090 ;
        RECT 65.855 30.905 66.145 30.950 ;
        RECT 68.600 30.890 68.920 30.950 ;
        RECT 79.180 30.890 79.500 31.150 ;
        RECT 88.395 31.090 88.685 31.135 ;
        RECT 89.300 31.090 89.620 31.150 ;
        RECT 88.395 30.950 89.620 31.090 ;
        RECT 88.395 30.905 88.685 30.950 ;
        RECT 89.300 30.890 89.620 30.950 ;
        RECT 11.950 30.270 90.610 30.750 ;
        RECT 18.000 30.070 18.320 30.130 ;
        RECT 15.790 29.930 18.320 30.070 ;
        RECT 15.790 29.730 15.930 29.930 ;
        RECT 18.000 29.870 18.320 29.930 ;
        RECT 22.600 30.070 22.920 30.130 ;
        RECT 24.915 30.070 25.205 30.115 ;
        RECT 22.600 29.930 25.205 30.070 ;
        RECT 22.600 29.870 22.920 29.930 ;
        RECT 24.915 29.885 25.205 29.930 ;
        RECT 25.820 30.070 26.140 30.130 ;
        RECT 46.520 30.070 46.840 30.130 ;
        RECT 63.080 30.070 63.400 30.130 ;
        RECT 64.935 30.070 65.225 30.115 ;
        RECT 68.140 30.070 68.460 30.130 ;
        RECT 25.820 29.930 46.840 30.070 ;
        RECT 25.820 29.870 26.140 29.930 ;
        RECT 15.330 29.590 15.930 29.730 ;
        RECT 18.890 29.730 19.180 29.775 ;
        RECT 20.300 29.730 20.620 29.790 ;
        RECT 18.890 29.590 20.620 29.730 ;
        RECT 15.330 29.435 15.470 29.590 ;
        RECT 18.890 29.545 19.180 29.590 ;
        RECT 20.300 29.530 20.620 29.590 ;
        RECT 15.255 29.205 15.545 29.435 ;
        RECT 15.700 29.190 16.020 29.450 ;
        RECT 16.160 29.190 16.480 29.450 ;
        RECT 17.095 29.390 17.385 29.435 ;
        RECT 18.550 29.390 19.150 29.405 ;
        RECT 23.980 29.390 24.300 29.450 ;
        RECT 25.835 29.390 26.125 29.435 ;
        RECT 17.095 29.265 24.300 29.390 ;
        RECT 17.095 29.250 18.690 29.265 ;
        RECT 19.010 29.250 24.300 29.265 ;
        RECT 17.095 29.205 17.385 29.250 ;
        RECT 23.980 29.190 24.300 29.250 ;
        RECT 24.530 29.250 26.125 29.390 ;
        RECT 16.620 29.050 16.940 29.110 ;
        RECT 17.555 29.050 17.845 29.095 ;
        RECT 16.620 28.910 17.845 29.050 ;
        RECT 16.620 28.850 16.940 28.910 ;
        RECT 17.555 28.865 17.845 28.910 ;
        RECT 18.435 29.050 18.725 29.095 ;
        RECT 19.625 29.050 19.915 29.095 ;
        RECT 22.145 29.050 22.435 29.095 ;
        RECT 18.435 28.910 22.435 29.050 ;
        RECT 18.435 28.865 18.725 28.910 ;
        RECT 19.625 28.865 19.915 28.910 ;
        RECT 22.145 28.865 22.435 28.910 ;
        RECT 18.040 28.710 18.330 28.755 ;
        RECT 20.140 28.710 20.430 28.755 ;
        RECT 21.710 28.710 22.000 28.755 ;
        RECT 18.040 28.570 22.000 28.710 ;
        RECT 18.040 28.525 18.330 28.570 ;
        RECT 20.140 28.525 20.430 28.570 ;
        RECT 21.710 28.525 22.000 28.570 ;
        RECT 13.860 28.170 14.180 28.430 ;
        RECT 21.220 28.370 21.540 28.430 ;
        RECT 24.530 28.415 24.670 29.250 ;
        RECT 25.835 29.205 26.125 29.250 ;
        RECT 26.740 29.190 27.060 29.450 ;
        RECT 29.055 29.205 29.345 29.435 ;
        RECT 29.515 29.205 29.805 29.435 ;
        RECT 29.130 28.710 29.270 29.205 ;
        RECT 29.590 29.050 29.730 29.205 ;
        RECT 29.960 29.190 30.280 29.450 ;
        RECT 30.970 29.435 31.110 29.930 ;
        RECT 46.520 29.870 46.840 29.930 ;
        RECT 49.370 29.930 62.850 30.070 ;
        RECT 37.335 29.730 37.625 29.775 ;
        RECT 32.810 29.590 37.625 29.730 ;
        RECT 30.895 29.205 31.185 29.435 ;
        RECT 31.815 29.390 32.105 29.435 ;
        RECT 32.260 29.390 32.580 29.450 ;
        RECT 32.810 29.435 32.950 29.590 ;
        RECT 37.335 29.545 37.625 29.590 ;
        RECT 40.540 29.730 40.860 29.790 ;
        RECT 49.370 29.730 49.510 29.930 ;
        RECT 57.100 29.730 57.420 29.790 ;
        RECT 40.540 29.590 49.510 29.730 ;
        RECT 49.830 29.590 57.420 29.730 ;
        RECT 40.540 29.530 40.860 29.590 ;
        RECT 31.815 29.250 32.580 29.390 ;
        RECT 31.815 29.205 32.105 29.250 ;
        RECT 32.260 29.190 32.580 29.250 ;
        RECT 32.735 29.205 33.025 29.435 ;
        RECT 33.180 29.190 33.500 29.450 ;
        RECT 33.655 29.390 33.945 29.435 ;
        RECT 34.100 29.390 34.420 29.450 ;
        RECT 33.655 29.250 34.420 29.390 ;
        RECT 33.655 29.205 33.945 29.250 ;
        RECT 34.100 29.190 34.420 29.250 ;
        RECT 35.480 29.190 35.800 29.450 ;
        RECT 36.415 29.390 36.705 29.435 ;
        RECT 41.460 29.390 41.780 29.450 ;
        RECT 42.380 29.435 42.700 29.450 ;
        RECT 49.830 29.435 49.970 29.590 ;
        RECT 57.100 29.530 57.420 29.590 ;
        RECT 51.120 29.435 51.440 29.450 ;
        RECT 36.415 29.250 41.780 29.390 ;
        RECT 36.415 29.205 36.705 29.250 ;
        RECT 41.460 29.190 41.780 29.250 ;
        RECT 42.350 29.205 42.700 29.435 ;
        RECT 49.755 29.205 50.045 29.435 ;
        RECT 51.090 29.205 51.440 29.435 ;
        RECT 42.380 29.190 42.700 29.205 ;
        RECT 51.120 29.190 51.440 29.205 ;
        RECT 52.500 29.390 52.820 29.450 ;
        RECT 59.030 29.435 59.170 29.930 ;
        RECT 61.255 29.730 61.545 29.775 ;
        RECT 59.950 29.590 61.545 29.730 ;
        RECT 62.710 29.730 62.850 29.930 ;
        RECT 63.080 29.930 65.225 30.070 ;
        RECT 63.080 29.870 63.400 29.930 ;
        RECT 64.935 29.885 65.225 29.930 ;
        RECT 65.930 29.930 68.460 30.070 ;
        RECT 65.930 29.730 66.070 29.930 ;
        RECT 68.140 29.870 68.460 29.930 ;
        RECT 71.360 29.870 71.680 30.130 ;
        RECT 78.260 30.070 78.580 30.130 ;
        RECT 81.035 30.070 81.325 30.115 ;
        RECT 78.260 29.930 83.090 30.070 ;
        RECT 78.260 29.870 78.580 29.930 ;
        RECT 81.035 29.885 81.325 29.930 ;
        RECT 62.710 29.590 66.070 29.730 ;
        RECT 52.500 29.250 55.030 29.390 ;
        RECT 52.500 29.190 52.820 29.250 ;
        RECT 33.270 29.050 33.410 29.190 ;
        RECT 54.890 29.110 55.030 29.250 ;
        RECT 58.955 29.205 59.245 29.435 ;
        RECT 59.400 29.190 59.720 29.450 ;
        RECT 59.950 29.435 60.090 29.590 ;
        RECT 61.255 29.545 61.545 29.590 ;
        RECT 66.300 29.530 66.620 29.790 ;
        RECT 70.440 29.730 70.760 29.790 ;
        RECT 69.610 29.590 70.760 29.730 ;
        RECT 59.875 29.205 60.165 29.435 ;
        RECT 60.795 29.205 61.085 29.435 ;
        RECT 61.700 29.390 62.020 29.450 ;
        RECT 62.175 29.390 62.465 29.435 ;
        RECT 61.700 29.250 62.465 29.390 ;
        RECT 41.000 29.050 41.320 29.110 ;
        RECT 29.590 28.910 33.410 29.050 ;
        RECT 34.190 28.910 41.320 29.050 ;
        RECT 34.190 28.770 34.330 28.910 ;
        RECT 41.000 28.850 41.320 28.910 ;
        RECT 41.895 29.050 42.185 29.095 ;
        RECT 43.085 29.050 43.375 29.095 ;
        RECT 45.605 29.050 45.895 29.095 ;
        RECT 41.895 28.910 45.895 29.050 ;
        RECT 41.895 28.865 42.185 28.910 ;
        RECT 43.085 28.865 43.375 28.910 ;
        RECT 45.605 28.865 45.895 28.910 ;
        RECT 50.635 29.050 50.925 29.095 ;
        RECT 51.825 29.050 52.115 29.095 ;
        RECT 54.345 29.050 54.635 29.095 ;
        RECT 50.635 28.910 54.635 29.050 ;
        RECT 50.635 28.865 50.925 28.910 ;
        RECT 51.825 28.865 52.115 28.910 ;
        RECT 54.345 28.865 54.635 28.910 ;
        RECT 54.800 29.050 55.120 29.110 ;
        RECT 60.870 29.050 61.010 29.205 ;
        RECT 61.700 29.190 62.020 29.250 ;
        RECT 62.175 29.205 62.465 29.250 ;
        RECT 62.620 29.390 62.940 29.450 ;
        RECT 63.095 29.390 63.385 29.435 ;
        RECT 62.620 29.250 63.385 29.390 ;
        RECT 54.800 28.910 61.010 29.050 ;
        RECT 62.250 29.050 62.390 29.205 ;
        RECT 62.620 29.190 62.940 29.250 ;
        RECT 63.095 29.205 63.385 29.250 ;
        RECT 65.840 29.190 66.160 29.450 ;
        RECT 66.760 29.190 67.080 29.450 ;
        RECT 67.695 29.390 67.985 29.435 ;
        RECT 67.310 29.250 67.985 29.390 ;
        RECT 67.310 29.050 67.450 29.250 ;
        RECT 67.695 29.205 67.985 29.250 ;
        RECT 68.155 29.205 68.445 29.435 ;
        RECT 68.600 29.390 68.920 29.450 ;
        RECT 69.610 29.435 69.750 29.590 ;
        RECT 70.440 29.530 70.760 29.590 ;
        RECT 71.820 29.730 72.140 29.790 ;
        RECT 81.940 29.730 82.260 29.790 ;
        RECT 82.950 29.775 83.090 29.930 ;
        RECT 71.820 29.590 82.260 29.730 ;
        RECT 71.820 29.530 72.140 29.590 ;
        RECT 74.210 29.435 74.350 29.590 ;
        RECT 81.940 29.530 82.260 29.590 ;
        RECT 82.875 29.730 83.165 29.775 ;
        RECT 84.700 29.730 85.020 29.790 ;
        RECT 82.875 29.590 85.020 29.730 ;
        RECT 82.875 29.545 83.165 29.590 ;
        RECT 84.700 29.530 85.020 29.590 ;
        RECT 69.075 29.390 69.365 29.435 ;
        RECT 68.600 29.250 69.365 29.390 ;
        RECT 68.230 29.050 68.370 29.205 ;
        RECT 68.600 29.190 68.920 29.250 ;
        RECT 69.075 29.205 69.365 29.250 ;
        RECT 69.535 29.205 69.825 29.435 ;
        RECT 69.995 29.205 70.285 29.435 ;
        RECT 74.135 29.205 74.425 29.435 ;
        RECT 75.470 29.390 75.760 29.435 ;
        RECT 76.880 29.390 77.200 29.450 ;
        RECT 75.470 29.250 77.200 29.390 ;
        RECT 75.470 29.205 75.760 29.250 ;
        RECT 62.250 28.910 67.450 29.050 ;
        RECT 67.770 28.910 68.370 29.050 ;
        RECT 54.800 28.850 55.120 28.910 ;
        RECT 29.130 28.570 30.190 28.710 ;
        RECT 24.455 28.370 24.745 28.415 ;
        RECT 21.220 28.230 24.745 28.370 ;
        RECT 21.220 28.170 21.540 28.230 ;
        RECT 24.455 28.185 24.745 28.230 ;
        RECT 27.675 28.370 27.965 28.415 ;
        RECT 29.500 28.370 29.820 28.430 ;
        RECT 27.675 28.230 29.820 28.370 ;
        RECT 30.050 28.370 30.190 28.570 ;
        RECT 34.100 28.510 34.420 28.770 ;
        RECT 35.940 28.710 36.260 28.770 ;
        RECT 34.650 28.570 36.260 28.710 ;
        RECT 34.650 28.370 34.790 28.570 ;
        RECT 35.940 28.510 36.260 28.570 ;
        RECT 41.500 28.710 41.790 28.755 ;
        RECT 43.600 28.710 43.890 28.755 ;
        RECT 45.170 28.710 45.460 28.755 ;
        RECT 41.500 28.570 45.460 28.710 ;
        RECT 41.500 28.525 41.790 28.570 ;
        RECT 43.600 28.525 43.890 28.570 ;
        RECT 45.170 28.525 45.460 28.570 ;
        RECT 50.240 28.710 50.530 28.755 ;
        RECT 52.340 28.710 52.630 28.755 ;
        RECT 53.910 28.710 54.200 28.755 ;
        RECT 50.240 28.570 54.200 28.710 ;
        RECT 50.240 28.525 50.530 28.570 ;
        RECT 52.340 28.525 52.630 28.570 ;
        RECT 53.910 28.525 54.200 28.570 ;
        RECT 57.575 28.710 57.865 28.755 ;
        RECT 58.480 28.710 58.800 28.770 ;
        RECT 57.575 28.570 58.800 28.710 ;
        RECT 57.575 28.525 57.865 28.570 ;
        RECT 58.480 28.510 58.800 28.570 ;
        RECT 30.050 28.230 34.790 28.370 ;
        RECT 27.675 28.185 27.965 28.230 ;
        RECT 29.500 28.170 29.820 28.230 ;
        RECT 35.020 28.170 35.340 28.430 ;
        RECT 44.220 28.370 44.540 28.430 ;
        RECT 47.915 28.370 48.205 28.415 ;
        RECT 44.220 28.230 48.205 28.370 ;
        RECT 44.220 28.170 44.540 28.230 ;
        RECT 47.915 28.185 48.205 28.230 ;
        RECT 54.340 28.370 54.660 28.430 ;
        RECT 56.655 28.370 56.945 28.415 ;
        RECT 54.340 28.230 56.945 28.370 ;
        RECT 60.870 28.370 61.010 28.910 ;
        RECT 61.240 28.710 61.560 28.770 ;
        RECT 65.840 28.710 66.160 28.770 ;
        RECT 61.240 28.570 66.160 28.710 ;
        RECT 61.240 28.510 61.560 28.570 ;
        RECT 65.840 28.510 66.160 28.570 ;
        RECT 67.770 28.370 67.910 28.910 ;
        RECT 68.140 28.710 68.460 28.770 ;
        RECT 70.070 28.710 70.210 29.205 ;
        RECT 76.880 29.190 77.200 29.250 ;
        RECT 77.340 29.390 77.660 29.450 ;
        RECT 81.020 29.390 81.340 29.450 ;
        RECT 82.415 29.390 82.705 29.435 ;
        RECT 77.340 29.250 79.870 29.390 ;
        RECT 77.340 29.190 77.660 29.250 ;
        RECT 79.730 29.110 79.870 29.250 ;
        RECT 81.020 29.250 82.705 29.390 ;
        RECT 81.020 29.190 81.340 29.250 ;
        RECT 82.415 29.205 82.705 29.250 ;
        RECT 83.335 29.205 83.625 29.435 ;
        RECT 75.015 29.050 75.305 29.095 ;
        RECT 76.205 29.050 76.495 29.095 ;
        RECT 78.725 29.050 79.015 29.095 ;
        RECT 75.015 28.910 79.015 29.050 ;
        RECT 75.015 28.865 75.305 28.910 ;
        RECT 76.205 28.865 76.495 28.910 ;
        RECT 78.725 28.865 79.015 28.910 ;
        RECT 79.640 29.050 79.960 29.110 ;
        RECT 83.410 29.050 83.550 29.205 ;
        RECT 84.240 29.190 84.560 29.450 ;
        RECT 79.640 28.910 83.550 29.050 ;
        RECT 79.640 28.850 79.960 28.910 ;
        RECT 68.140 28.570 70.210 28.710 ;
        RECT 74.620 28.710 74.910 28.755 ;
        RECT 76.720 28.710 77.010 28.755 ;
        RECT 78.290 28.710 78.580 28.755 ;
        RECT 74.620 28.570 78.580 28.710 ;
        RECT 68.140 28.510 68.460 28.570 ;
        RECT 74.620 28.525 74.910 28.570 ;
        RECT 76.720 28.525 77.010 28.570 ;
        RECT 78.290 28.525 78.580 28.570 ;
        RECT 80.100 28.370 80.420 28.430 ;
        RECT 60.870 28.230 80.420 28.370 ;
        RECT 54.340 28.170 54.660 28.230 ;
        RECT 56.655 28.185 56.945 28.230 ;
        RECT 80.100 28.170 80.420 28.230 ;
        RECT 81.480 28.170 81.800 28.430 ;
        RECT 11.950 27.550 90.610 28.030 ;
        RECT 17.080 27.350 17.400 27.410 ;
        RECT 20.315 27.350 20.605 27.395 ;
        RECT 17.080 27.210 20.605 27.350 ;
        RECT 17.080 27.150 17.400 27.210 ;
        RECT 20.315 27.165 20.605 27.210 ;
        RECT 13.900 27.010 14.190 27.055 ;
        RECT 16.000 27.010 16.290 27.055 ;
        RECT 17.570 27.010 17.860 27.055 ;
        RECT 13.900 26.870 17.860 27.010 ;
        RECT 13.900 26.825 14.190 26.870 ;
        RECT 16.000 26.825 16.290 26.870 ;
        RECT 17.570 26.825 17.860 26.870 ;
        RECT 14.295 26.670 14.585 26.715 ;
        RECT 15.485 26.670 15.775 26.715 ;
        RECT 18.005 26.670 18.295 26.715 ;
        RECT 14.295 26.530 18.295 26.670 ;
        RECT 14.295 26.485 14.585 26.530 ;
        RECT 15.485 26.485 15.775 26.530 ;
        RECT 18.005 26.485 18.295 26.530 ;
        RECT 13.415 26.330 13.705 26.375 ;
        RECT 16.620 26.330 16.940 26.390 ;
        RECT 13.415 26.190 16.940 26.330 ;
        RECT 20.390 26.330 20.530 27.165 ;
        RECT 23.520 27.150 23.840 27.410 ;
        RECT 26.280 27.350 26.600 27.410 ;
        RECT 41.015 27.350 41.305 27.395 ;
        RECT 41.460 27.350 41.780 27.410 ;
        RECT 26.280 27.210 40.770 27.350 ;
        RECT 26.280 27.150 26.600 27.210 ;
        RECT 27.240 27.010 27.530 27.055 ;
        RECT 29.340 27.010 29.630 27.055 ;
        RECT 30.910 27.010 31.200 27.055 ;
        RECT 27.240 26.870 31.200 27.010 ;
        RECT 27.240 26.825 27.530 26.870 ;
        RECT 29.340 26.825 29.630 26.870 ;
        RECT 30.910 26.825 31.200 26.870 ;
        RECT 34.600 27.010 34.890 27.055 ;
        RECT 36.700 27.010 36.990 27.055 ;
        RECT 38.270 27.010 38.560 27.055 ;
        RECT 34.600 26.870 38.560 27.010 ;
        RECT 40.630 27.010 40.770 27.210 ;
        RECT 41.015 27.210 41.780 27.350 ;
        RECT 41.015 27.165 41.305 27.210 ;
        RECT 41.460 27.150 41.780 27.210 ;
        RECT 42.380 27.150 42.700 27.410 ;
        RECT 45.230 27.210 68.600 27.350 ;
        RECT 45.230 27.010 45.370 27.210 ;
        RECT 40.630 26.870 45.370 27.010 ;
        RECT 34.600 26.825 34.890 26.870 ;
        RECT 36.700 26.825 36.990 26.870 ;
        RECT 38.270 26.825 38.560 26.870 ;
        RECT 45.600 26.810 45.920 27.070 ;
        RECT 51.120 26.810 51.440 27.070 ;
        RECT 68.460 27.010 68.600 27.210 ;
        RECT 76.880 27.150 77.200 27.410 ;
        RECT 81.480 27.010 81.800 27.070 ;
        RECT 68.460 26.870 81.800 27.010 ;
        RECT 81.480 26.810 81.800 26.870 ;
        RECT 82.440 27.010 82.730 27.055 ;
        RECT 84.540 27.010 84.830 27.055 ;
        RECT 86.110 27.010 86.400 27.055 ;
        RECT 82.440 26.870 86.400 27.010 ;
        RECT 82.440 26.825 82.730 26.870 ;
        RECT 84.540 26.825 84.830 26.870 ;
        RECT 86.110 26.825 86.400 26.870 ;
        RECT 27.635 26.670 27.925 26.715 ;
        RECT 28.825 26.670 29.115 26.715 ;
        RECT 31.345 26.670 31.635 26.715 ;
        RECT 27.635 26.530 31.635 26.670 ;
        RECT 27.635 26.485 27.925 26.530 ;
        RECT 28.825 26.485 29.115 26.530 ;
        RECT 31.345 26.485 31.635 26.530 ;
        RECT 34.995 26.670 35.285 26.715 ;
        RECT 36.185 26.670 36.475 26.715 ;
        RECT 38.705 26.670 38.995 26.715 ;
        RECT 45.690 26.670 45.830 26.810 ;
        RECT 47.440 26.670 47.760 26.730 ;
        RECT 72.740 26.670 73.060 26.730 ;
        RECT 76.880 26.670 77.200 26.730 ;
        RECT 79.640 26.670 79.960 26.730 ;
        RECT 81.940 26.670 82.260 26.730 ;
        RECT 34.995 26.530 38.995 26.670 ;
        RECT 34.995 26.485 35.285 26.530 ;
        RECT 36.185 26.485 36.475 26.530 ;
        RECT 38.705 26.485 38.995 26.530 ;
        RECT 44.310 26.530 76.650 26.670 ;
        RECT 20.775 26.330 21.065 26.375 ;
        RECT 20.390 26.190 21.065 26.330 ;
        RECT 13.415 26.145 13.705 26.190 ;
        RECT 16.620 26.130 16.940 26.190 ;
        RECT 20.775 26.145 21.065 26.190 ;
        RECT 21.220 26.330 21.540 26.390 ;
        RECT 22.155 26.330 22.445 26.375 ;
        RECT 21.220 26.190 22.445 26.330 ;
        RECT 21.220 26.130 21.540 26.190 ;
        RECT 22.155 26.145 22.445 26.190 ;
        RECT 22.615 26.330 22.905 26.375 ;
        RECT 23.980 26.330 24.300 26.390 ;
        RECT 22.615 26.190 24.300 26.330 ;
        RECT 22.615 26.145 22.905 26.190 ;
        RECT 23.980 26.130 24.300 26.190 ;
        RECT 26.740 26.130 27.060 26.390 ;
        RECT 28.090 26.330 28.380 26.375 ;
        RECT 29.500 26.330 29.820 26.390 ;
        RECT 28.090 26.190 29.820 26.330 ;
        RECT 28.090 26.145 28.380 26.190 ;
        RECT 29.500 26.130 29.820 26.190 ;
        RECT 34.100 26.130 34.420 26.390 ;
        RECT 44.310 26.375 44.450 26.530 ;
        RECT 47.440 26.470 47.760 26.530 ;
        RECT 35.450 26.145 35.740 26.375 ;
        RECT 43.775 26.145 44.065 26.375 ;
        RECT 44.235 26.145 44.525 26.375 ;
        RECT 13.860 25.990 14.180 26.050 ;
        RECT 14.640 25.990 14.930 26.035 ;
        RECT 21.695 25.990 21.985 26.035 ;
        RECT 13.860 25.850 14.930 25.990 ;
        RECT 13.860 25.790 14.180 25.850 ;
        RECT 14.640 25.805 14.930 25.850 ;
        RECT 20.850 25.850 21.985 25.990 ;
        RECT 20.850 25.710 20.990 25.850 ;
        RECT 21.695 25.805 21.985 25.850 ;
        RECT 35.020 25.990 35.340 26.050 ;
        RECT 35.570 25.990 35.710 26.145 ;
        RECT 35.020 25.850 35.710 25.990 ;
        RECT 35.940 25.990 36.260 26.050 ;
        RECT 40.540 25.990 40.860 26.050 ;
        RECT 43.850 25.990 43.990 26.145 ;
        RECT 44.680 26.130 45.000 26.390 ;
        RECT 45.615 26.330 45.905 26.375 ;
        RECT 46.520 26.330 46.840 26.390 ;
        RECT 52.500 26.330 52.820 26.390 ;
        RECT 53.050 26.375 53.190 26.530 ;
        RECT 72.740 26.470 73.060 26.530 ;
        RECT 45.615 26.190 46.840 26.330 ;
        RECT 45.615 26.145 45.905 26.190 ;
        RECT 46.520 26.130 46.840 26.190 ;
        RECT 48.910 26.190 52.820 26.330 ;
        RECT 35.940 25.850 43.990 25.990 ;
        RECT 35.020 25.790 35.340 25.850 ;
        RECT 35.940 25.790 36.260 25.850 ;
        RECT 40.540 25.790 40.860 25.850 ;
        RECT 48.360 25.790 48.680 26.050 ;
        RECT 20.760 25.450 21.080 25.710 ;
        RECT 29.500 25.650 29.820 25.710 ;
        RECT 33.655 25.650 33.945 25.695 ;
        RECT 29.500 25.510 33.945 25.650 ;
        RECT 29.500 25.450 29.820 25.510 ;
        RECT 33.655 25.465 33.945 25.510 ;
        RECT 34.560 25.650 34.880 25.710 ;
        RECT 48.910 25.650 49.050 26.190 ;
        RECT 52.500 26.130 52.820 26.190 ;
        RECT 52.975 26.145 53.265 26.375 ;
        RECT 53.435 26.145 53.725 26.375 ;
        RECT 54.355 26.145 54.645 26.375 ;
        RECT 58.035 26.330 58.325 26.375 ;
        RECT 67.220 26.330 67.540 26.390 ;
        RECT 74.135 26.330 74.425 26.375 ;
        RECT 75.960 26.330 76.280 26.390 ;
        RECT 58.035 26.190 67.540 26.330 ;
        RECT 58.035 26.145 58.325 26.190 ;
        RECT 49.295 25.805 49.585 26.035 ;
        RECT 50.215 25.990 50.505 26.035 ;
        RECT 53.510 25.990 53.650 26.145 ;
        RECT 50.215 25.850 53.650 25.990 ;
        RECT 50.215 25.805 50.505 25.850 ;
        RECT 34.560 25.510 49.050 25.650 ;
        RECT 49.370 25.650 49.510 25.805 ;
        RECT 54.430 25.710 54.570 26.145 ;
        RECT 67.220 26.130 67.540 26.190 ;
        RECT 68.460 26.190 76.280 26.330 ;
        RECT 76.510 26.330 76.650 26.530 ;
        RECT 76.880 26.530 78.950 26.670 ;
        RECT 76.880 26.470 77.200 26.530 ;
        RECT 77.800 26.330 78.120 26.390 ;
        RECT 76.510 26.190 78.120 26.330 ;
        RECT 54.800 25.990 55.120 26.050 ;
        RECT 68.460 25.990 68.600 26.190 ;
        RECT 74.135 26.145 74.425 26.190 ;
        RECT 75.960 26.130 76.280 26.190 ;
        RECT 77.800 26.130 78.120 26.190 ;
        RECT 78.260 26.130 78.580 26.390 ;
        RECT 78.810 26.375 78.950 26.530 ;
        RECT 79.640 26.530 82.260 26.670 ;
        RECT 79.640 26.470 79.960 26.530 ;
        RECT 81.940 26.470 82.260 26.530 ;
        RECT 82.835 26.670 83.125 26.715 ;
        RECT 84.025 26.670 84.315 26.715 ;
        RECT 86.545 26.670 86.835 26.715 ;
        RECT 82.835 26.530 86.835 26.670 ;
        RECT 82.835 26.485 83.125 26.530 ;
        RECT 84.025 26.485 84.315 26.530 ;
        RECT 86.545 26.485 86.835 26.530 ;
        RECT 78.735 26.145 79.025 26.375 ;
        RECT 79.180 26.130 79.500 26.390 ;
        RECT 80.100 26.130 80.420 26.390 ;
        RECT 54.800 25.850 68.600 25.990 ;
        RECT 75.055 25.990 75.345 26.035 ;
        RECT 81.940 25.990 82.260 26.050 ;
        RECT 83.180 25.990 83.470 26.035 ;
        RECT 75.055 25.850 81.710 25.990 ;
        RECT 54.800 25.790 55.120 25.850 ;
        RECT 75.055 25.805 75.345 25.850 ;
        RECT 50.660 25.650 50.980 25.710 ;
        RECT 53.880 25.650 54.200 25.710 ;
        RECT 49.370 25.510 54.200 25.650 ;
        RECT 34.560 25.450 34.880 25.510 ;
        RECT 50.660 25.450 50.980 25.510 ;
        RECT 53.880 25.450 54.200 25.510 ;
        RECT 54.340 25.650 54.660 25.710 ;
        RECT 57.115 25.650 57.405 25.695 ;
        RECT 54.340 25.510 57.405 25.650 ;
        RECT 54.340 25.450 54.660 25.510 ;
        RECT 57.115 25.465 57.405 25.510 ;
        RECT 75.975 25.650 76.265 25.695 ;
        RECT 79.180 25.650 79.500 25.710 ;
        RECT 75.975 25.510 79.500 25.650 ;
        RECT 81.570 25.650 81.710 25.850 ;
        RECT 81.940 25.850 83.470 25.990 ;
        RECT 81.940 25.790 82.260 25.850 ;
        RECT 83.180 25.805 83.470 25.850 ;
        RECT 84.240 25.650 84.560 25.710 ;
        RECT 88.840 25.650 89.160 25.710 ;
        RECT 81.570 25.510 89.160 25.650 ;
        RECT 75.975 25.465 76.265 25.510 ;
        RECT 79.180 25.450 79.500 25.510 ;
        RECT 84.240 25.450 84.560 25.510 ;
        RECT 88.840 25.450 89.160 25.510 ;
        RECT 11.950 24.830 90.610 25.310 ;
        RECT 29.055 24.630 29.345 24.675 ;
        RECT 29.960 24.630 30.280 24.690 ;
        RECT 29.055 24.490 30.280 24.630 ;
        RECT 29.055 24.445 29.345 24.490 ;
        RECT 29.960 24.430 30.280 24.490 ;
        RECT 42.380 24.630 42.700 24.690 ;
        RECT 48.360 24.630 48.680 24.690 ;
        RECT 54.800 24.630 55.120 24.690 ;
        RECT 42.380 24.490 46.290 24.630 ;
        RECT 42.380 24.430 42.700 24.490 ;
        RECT 20.760 24.290 21.080 24.350 ;
        RECT 22.155 24.290 22.445 24.335 ;
        RECT 20.760 24.150 22.445 24.290 ;
        RECT 20.760 24.090 21.080 24.150 ;
        RECT 22.155 24.105 22.445 24.150 ;
        RECT 26.280 24.290 26.600 24.350 ;
        RECT 27.215 24.290 27.505 24.335 ;
        RECT 26.280 24.150 27.505 24.290 ;
        RECT 26.280 24.090 26.600 24.150 ;
        RECT 27.215 24.105 27.505 24.150 ;
        RECT 28.135 24.290 28.425 24.335 ;
        RECT 29.500 24.290 29.820 24.350 ;
        RECT 28.135 24.150 29.820 24.290 ;
        RECT 28.135 24.105 28.425 24.150 ;
        RECT 29.500 24.090 29.820 24.150 ;
        RECT 39.160 24.290 39.480 24.350 ;
        RECT 41.015 24.290 41.305 24.335 ;
        RECT 44.220 24.290 44.540 24.350 ;
        RECT 39.160 24.150 41.305 24.290 ;
        RECT 39.160 24.090 39.480 24.150 ;
        RECT 41.015 24.105 41.305 24.150 ;
        RECT 41.550 24.150 44.540 24.290 ;
        RECT 14.795 23.765 15.085 23.995 ;
        RECT 17.080 23.950 17.400 24.010 ;
        RECT 18.015 23.950 18.305 23.995 ;
        RECT 17.080 23.810 18.305 23.950 ;
        RECT 14.870 23.270 15.010 23.765 ;
        RECT 17.080 23.750 17.400 23.810 ;
        RECT 18.015 23.765 18.305 23.810 ;
        RECT 19.855 23.950 20.145 23.995 ;
        RECT 20.300 23.950 20.620 24.010 ;
        RECT 21.235 23.950 21.525 23.995 ;
        RECT 19.855 23.810 21.525 23.950 ;
        RECT 19.855 23.765 20.145 23.810 ;
        RECT 20.300 23.750 20.620 23.810 ;
        RECT 21.235 23.765 21.525 23.810 ;
        RECT 22.615 23.765 22.905 23.995 ;
        RECT 23.075 23.950 23.365 23.995 ;
        RECT 23.980 23.950 24.300 24.010 ;
        RECT 23.075 23.810 24.300 23.950 ;
        RECT 23.075 23.765 23.365 23.810 ;
        RECT 22.690 23.610 22.830 23.765 ;
        RECT 23.980 23.750 24.300 23.810 ;
        RECT 24.455 23.950 24.745 23.995 ;
        RECT 24.900 23.950 25.220 24.010 ;
        RECT 24.455 23.810 25.220 23.950 ;
        RECT 29.590 23.950 29.730 24.090 ;
        RECT 41.550 23.995 41.690 24.150 ;
        RECT 44.220 24.090 44.540 24.150 ;
        RECT 45.600 24.090 45.920 24.350 ;
        RECT 46.150 24.290 46.290 24.490 ;
        RECT 48.360 24.490 55.120 24.630 ;
        RECT 48.360 24.430 48.680 24.490 ;
        RECT 54.800 24.430 55.120 24.490 ;
        RECT 64.460 24.630 64.780 24.690 ;
        RECT 70.440 24.630 70.760 24.690 ;
        RECT 76.880 24.630 77.200 24.690 ;
        RECT 64.460 24.490 66.990 24.630 ;
        RECT 64.460 24.430 64.780 24.490 ;
        RECT 50.200 24.290 50.520 24.350 ;
        RECT 46.150 24.150 50.520 24.290 ;
        RECT 40.095 23.950 40.385 23.995 ;
        RECT 29.590 23.810 40.385 23.950 ;
        RECT 24.455 23.765 24.745 23.810 ;
        RECT 24.530 23.610 24.670 23.765 ;
        RECT 24.900 23.750 25.220 23.810 ;
        RECT 40.095 23.765 40.385 23.810 ;
        RECT 41.475 23.765 41.765 23.995 ;
        RECT 41.935 23.950 42.225 23.995 ;
        RECT 42.380 23.950 42.700 24.010 ;
        RECT 46.610 23.995 46.750 24.150 ;
        RECT 50.200 24.090 50.520 24.150 ;
        RECT 54.340 24.290 54.660 24.350 ;
        RECT 62.175 24.290 62.465 24.335 ;
        RECT 66.850 24.290 66.990 24.490 ;
        RECT 69.150 24.490 77.200 24.630 ;
        RECT 54.340 24.150 61.010 24.290 ;
        RECT 54.340 24.090 54.660 24.150 ;
        RECT 41.935 23.810 42.700 23.950 ;
        RECT 41.935 23.765 42.225 23.810 ;
        RECT 42.380 23.750 42.700 23.810 ;
        RECT 44.695 23.765 44.985 23.995 ;
        RECT 46.075 23.765 46.365 23.995 ;
        RECT 46.535 23.765 46.825 23.995 ;
        RECT 56.640 23.950 56.960 24.010 ;
        RECT 58.955 23.950 59.245 23.995 ;
        RECT 56.640 23.810 59.245 23.950 ;
        RECT 22.690 23.470 24.670 23.610 ;
        RECT 40.540 23.610 40.860 23.670 ;
        RECT 44.770 23.610 44.910 23.765 ;
        RECT 40.540 23.470 44.910 23.610 ;
        RECT 46.150 23.610 46.290 23.765 ;
        RECT 56.640 23.750 56.960 23.810 ;
        RECT 58.955 23.765 59.245 23.810 ;
        RECT 59.400 23.750 59.720 24.010 ;
        RECT 60.870 23.995 61.010 24.150 ;
        RECT 62.175 24.150 66.530 24.290 ;
        RECT 66.850 24.150 67.450 24.290 ;
        RECT 62.175 24.105 62.465 24.150 ;
        RECT 66.390 24.010 66.530 24.150 ;
        RECT 59.875 23.765 60.165 23.995 ;
        RECT 60.795 23.765 61.085 23.995 ;
        RECT 62.620 23.950 62.940 24.010 ;
        RECT 63.095 23.950 63.385 23.995 ;
        RECT 62.620 23.810 63.385 23.950 ;
        RECT 47.900 23.610 48.220 23.670 ;
        RECT 46.150 23.470 48.220 23.610 ;
        RECT 40.540 23.410 40.860 23.470 ;
        RECT 47.900 23.410 48.220 23.470 ;
        RECT 55.260 23.610 55.580 23.670 ;
        RECT 59.490 23.610 59.630 23.750 ;
        RECT 55.260 23.470 59.630 23.610 ;
        RECT 59.950 23.610 60.090 23.765 ;
        RECT 62.620 23.750 62.940 23.810 ;
        RECT 63.095 23.765 63.385 23.810 ;
        RECT 64.920 23.750 65.240 24.010 ;
        RECT 65.395 23.765 65.685 23.995 ;
        RECT 61.255 23.610 61.545 23.655 ;
        RECT 64.460 23.610 64.780 23.670 ;
        RECT 59.950 23.470 61.545 23.610 ;
        RECT 55.260 23.410 55.580 23.470 ;
        RECT 61.255 23.425 61.545 23.470 ;
        RECT 61.790 23.470 64.780 23.610 ;
        RECT 65.470 23.610 65.610 23.765 ;
        RECT 65.840 23.750 66.160 24.010 ;
        RECT 66.300 23.950 66.620 24.010 ;
        RECT 66.775 23.950 67.065 23.995 ;
        RECT 66.300 23.810 67.065 23.950 ;
        RECT 67.310 23.950 67.450 24.150 ;
        RECT 69.150 23.995 69.290 24.490 ;
        RECT 70.440 24.430 70.760 24.490 ;
        RECT 76.880 24.430 77.200 24.490 ;
        RECT 77.800 24.430 78.120 24.690 ;
        RECT 78.260 24.630 78.580 24.690 ;
        RECT 78.260 24.490 80.790 24.630 ;
        RECT 78.260 24.430 78.580 24.490 ;
        RECT 72.755 24.290 73.045 24.335 ;
        RECT 73.660 24.290 73.980 24.350 ;
        RECT 72.755 24.150 73.980 24.290 ;
        RECT 72.755 24.105 73.045 24.150 ;
        RECT 73.660 24.090 73.980 24.150 ;
        RECT 74.120 24.290 74.440 24.350 ;
        RECT 77.890 24.290 78.030 24.430 ;
        RECT 80.650 24.290 80.790 24.490 ;
        RECT 81.020 24.290 81.340 24.350 ;
        RECT 74.120 24.150 76.650 24.290 ;
        RECT 77.890 24.150 80.330 24.290 ;
        RECT 74.120 24.090 74.440 24.150 ;
        RECT 68.615 23.950 68.905 23.995 ;
        RECT 67.310 23.810 68.905 23.950 ;
        RECT 66.300 23.750 66.620 23.810 ;
        RECT 66.775 23.765 67.065 23.810 ;
        RECT 68.615 23.765 68.905 23.810 ;
        RECT 69.075 23.765 69.365 23.995 ;
        RECT 69.535 23.765 69.825 23.995 ;
        RECT 70.455 23.950 70.745 23.995 ;
        RECT 70.455 23.810 71.590 23.950 ;
        RECT 70.455 23.765 70.745 23.810 ;
        RECT 67.680 23.610 68.000 23.670 ;
        RECT 65.470 23.470 68.000 23.610 ;
        RECT 69.610 23.610 69.750 23.765 ;
        RECT 70.915 23.610 71.205 23.655 ;
        RECT 69.610 23.470 71.205 23.610 ;
        RECT 71.450 23.610 71.590 23.810 ;
        RECT 71.820 23.750 72.140 24.010 ;
        RECT 75.500 23.950 75.820 24.010 ;
        RECT 76.510 23.995 76.650 24.150 ;
        RECT 72.370 23.810 75.820 23.950 ;
        RECT 72.370 23.610 72.510 23.810 ;
        RECT 75.500 23.750 75.820 23.810 ;
        RECT 76.435 23.765 76.725 23.995 ;
        RECT 76.895 23.765 77.185 23.995 ;
        RECT 71.450 23.470 72.510 23.610 ;
        RECT 76.970 23.610 77.110 23.765 ;
        RECT 77.340 23.750 77.660 24.010 ;
        RECT 77.800 23.950 78.120 24.010 ;
        RECT 78.275 23.950 78.565 23.995 ;
        RECT 77.800 23.810 78.565 23.950 ;
        RECT 77.800 23.750 78.120 23.810 ;
        RECT 78.275 23.765 78.565 23.810 ;
        RECT 78.720 23.750 79.040 24.010 ;
        RECT 79.180 23.950 79.500 24.010 ;
        RECT 80.190 23.995 80.330 24.150 ;
        RECT 80.650 24.150 81.340 24.290 ;
        RECT 80.650 23.995 80.790 24.150 ;
        RECT 81.020 24.090 81.340 24.150 ;
        RECT 79.655 23.950 79.945 23.995 ;
        RECT 79.180 23.810 79.945 23.950 ;
        RECT 79.180 23.750 79.500 23.810 ;
        RECT 79.655 23.765 79.945 23.810 ;
        RECT 80.115 23.765 80.405 23.995 ;
        RECT 80.575 23.765 80.865 23.995 ;
        RECT 83.795 23.950 84.085 23.995 ;
        RECT 84.240 23.950 84.560 24.010 ;
        RECT 81.065 23.810 84.560 23.950 ;
        RECT 81.065 23.610 81.205 23.810 ;
        RECT 83.795 23.765 84.085 23.810 ;
        RECT 84.240 23.750 84.560 23.810 ;
        RECT 85.620 23.750 85.940 24.010 ;
        RECT 88.840 23.750 89.160 24.010 ;
        RECT 76.970 23.470 81.205 23.610 ;
        RECT 22.140 23.270 22.460 23.330 ;
        RECT 14.870 23.130 22.460 23.270 ;
        RECT 22.140 23.070 22.460 23.130 ;
        RECT 23.060 23.270 23.380 23.330 ;
        RECT 25.375 23.270 25.665 23.315 ;
        RECT 23.060 23.130 25.665 23.270 ;
        RECT 23.060 23.070 23.380 23.130 ;
        RECT 25.375 23.085 25.665 23.130 ;
        RECT 42.840 23.070 43.160 23.330 ;
        RECT 47.455 23.270 47.745 23.315 ;
        RECT 48.820 23.270 49.140 23.330 ;
        RECT 47.455 23.130 49.140 23.270 ;
        RECT 47.455 23.085 47.745 23.130 ;
        RECT 48.820 23.070 49.140 23.130 ;
        RECT 54.800 23.270 55.120 23.330 ;
        RECT 61.790 23.270 61.930 23.470 ;
        RECT 64.460 23.410 64.780 23.470 ;
        RECT 67.680 23.410 68.000 23.470 ;
        RECT 70.915 23.425 71.205 23.470 ;
        RECT 81.940 23.410 82.260 23.670 ;
        RECT 93.440 23.610 93.760 23.670 ;
        RECT 84.790 23.470 93.760 23.610 ;
        RECT 54.800 23.130 61.930 23.270 ;
        RECT 54.800 23.070 55.120 23.130 ;
        RECT 64.000 23.070 64.320 23.330 ;
        RECT 69.060 23.270 69.380 23.330 ;
        RECT 84.790 23.315 84.930 23.470 ;
        RECT 93.440 23.410 93.760 23.470 ;
        RECT 75.515 23.270 75.805 23.315 ;
        RECT 69.060 23.130 75.805 23.270 ;
        RECT 69.060 23.070 69.380 23.130 ;
        RECT 75.515 23.085 75.805 23.130 ;
        RECT 84.715 23.085 85.005 23.315 ;
        RECT 86.555 23.270 86.845 23.315 ;
        RECT 90.220 23.270 90.540 23.330 ;
        RECT 86.555 23.130 90.540 23.270 ;
        RECT 86.555 23.085 86.845 23.130 ;
        RECT 90.220 23.070 90.540 23.130 ;
        RECT 13.400 22.930 13.720 22.990 ;
        RECT 13.875 22.930 14.165 22.975 ;
        RECT 13.400 22.790 14.165 22.930 ;
        RECT 13.400 22.730 13.720 22.790 ;
        RECT 13.875 22.745 14.165 22.790 ;
        RECT 17.080 22.730 17.400 22.990 ;
        RECT 18.000 22.930 18.320 22.990 ;
        RECT 18.935 22.930 19.225 22.975 ;
        RECT 18.000 22.790 19.225 22.930 ;
        RECT 18.000 22.730 18.320 22.790 ;
        RECT 18.935 22.745 19.225 22.790 ;
        RECT 23.520 22.930 23.840 22.990 ;
        RECT 23.995 22.930 24.285 22.975 ;
        RECT 23.520 22.790 24.285 22.930 ;
        RECT 23.520 22.730 23.840 22.790 ;
        RECT 23.995 22.745 24.285 22.790 ;
        RECT 57.560 22.730 57.880 22.990 ;
        RECT 65.840 22.930 66.160 22.990 ;
        RECT 67.235 22.930 67.525 22.975 ;
        RECT 65.840 22.790 67.525 22.930 ;
        RECT 65.840 22.730 66.160 22.790 ;
        RECT 67.235 22.745 67.525 22.790 ;
        RECT 76.880 22.930 77.200 22.990 ;
        RECT 78.720 22.930 79.040 22.990 ;
        RECT 76.880 22.790 79.040 22.930 ;
        RECT 76.880 22.730 77.200 22.790 ;
        RECT 78.720 22.730 79.040 22.790 ;
        RECT 87.000 22.930 87.320 22.990 ;
        RECT 87.935 22.930 88.225 22.975 ;
        RECT 87.000 22.790 88.225 22.930 ;
        RECT 87.000 22.730 87.320 22.790 ;
        RECT 87.935 22.745 88.225 22.790 ;
        RECT 11.950 22.110 90.610 22.590 ;
        RECT 24.440 21.910 24.760 21.970 ;
        RECT 40.095 21.910 40.385 21.955 ;
        RECT 40.540 21.910 40.860 21.970 ;
        RECT 24.440 21.770 39.850 21.910 ;
        RECT 24.440 21.710 24.760 21.770 ;
        RECT 21.680 21.570 22.000 21.630 ;
        RECT 33.680 21.570 33.970 21.615 ;
        RECT 35.780 21.570 36.070 21.615 ;
        RECT 37.350 21.570 37.640 21.615 ;
        RECT 21.680 21.430 22.370 21.570 ;
        RECT 21.680 21.370 22.000 21.430 ;
        RECT 18.460 21.230 18.780 21.290 ;
        RECT 22.230 21.230 22.370 21.430 ;
        RECT 33.680 21.430 37.640 21.570 ;
        RECT 33.680 21.385 33.970 21.430 ;
        RECT 35.780 21.385 36.070 21.430 ;
        RECT 37.350 21.385 37.640 21.430 ;
        RECT 34.075 21.230 34.365 21.275 ;
        RECT 35.265 21.230 35.555 21.275 ;
        RECT 37.785 21.230 38.075 21.275 ;
        RECT 15.330 21.090 21.910 21.230 ;
        RECT 15.330 20.935 15.470 21.090 ;
        RECT 18.460 21.030 18.780 21.090 ;
        RECT 15.255 20.705 15.545 20.935 ;
        RECT 15.700 20.690 16.020 20.950 ;
        RECT 16.160 20.690 16.480 20.950 ;
        RECT 17.095 20.705 17.385 20.935 ;
        RECT 19.855 20.890 20.145 20.935 ;
        RECT 21.220 20.890 21.540 20.950 ;
        RECT 21.770 20.935 21.910 21.090 ;
        RECT 22.230 21.090 31.110 21.230 ;
        RECT 22.230 20.935 22.370 21.090 ;
        RECT 19.855 20.750 21.540 20.890 ;
        RECT 19.855 20.705 20.145 20.750 ;
        RECT 17.170 20.550 17.310 20.705 ;
        RECT 21.220 20.690 21.540 20.750 ;
        RECT 21.695 20.705 21.985 20.935 ;
        RECT 22.155 20.705 22.445 20.935 ;
        RECT 22.600 20.690 22.920 20.950 ;
        RECT 23.535 20.890 23.825 20.935 ;
        RECT 25.820 20.890 26.140 20.950 ;
        RECT 27.290 20.935 27.430 21.090 ;
        RECT 23.535 20.750 26.140 20.890 ;
        RECT 23.535 20.705 23.825 20.750 ;
        RECT 23.610 20.550 23.750 20.705 ;
        RECT 25.820 20.690 26.140 20.750 ;
        RECT 26.755 20.705 27.045 20.935 ;
        RECT 27.215 20.705 27.505 20.935 ;
        RECT 17.170 20.410 23.750 20.550 ;
        RECT 13.860 20.010 14.180 20.270 ;
        RECT 18.920 20.010 19.240 20.270 ;
        RECT 19.380 20.210 19.700 20.270 ;
        RECT 20.315 20.210 20.605 20.255 ;
        RECT 19.380 20.070 20.605 20.210 ;
        RECT 26.830 20.210 26.970 20.705 ;
        RECT 27.660 20.690 27.980 20.950 ;
        RECT 29.515 20.705 29.805 20.935 ;
        RECT 29.590 20.550 29.730 20.705 ;
        RECT 30.420 20.690 30.740 20.950 ;
        RECT 30.970 20.935 31.110 21.090 ;
        RECT 34.075 21.090 38.075 21.230 ;
        RECT 39.710 21.230 39.850 21.770 ;
        RECT 40.095 21.770 40.860 21.910 ;
        RECT 40.095 21.725 40.385 21.770 ;
        RECT 40.540 21.710 40.860 21.770 ;
        RECT 42.840 21.910 43.160 21.970 ;
        RECT 56.640 21.910 56.960 21.970 ;
        RECT 68.140 21.910 68.460 21.970 ;
        RECT 42.840 21.770 56.960 21.910 ;
        RECT 42.840 21.710 43.160 21.770 ;
        RECT 56.640 21.710 56.960 21.770 ;
        RECT 57.190 21.770 68.460 21.910 ;
        RECT 57.190 21.570 57.330 21.770 ;
        RECT 68.140 21.710 68.460 21.770 ;
        RECT 71.375 21.910 71.665 21.955 ;
        RECT 71.820 21.910 72.140 21.970 ;
        RECT 71.375 21.770 72.140 21.910 ;
        RECT 71.375 21.725 71.665 21.770 ;
        RECT 71.820 21.710 72.140 21.770 ;
        RECT 73.200 21.910 73.520 21.970 ;
        RECT 73.200 21.770 82.630 21.910 ;
        RECT 73.200 21.710 73.520 21.770 ;
        RECT 42.930 21.430 57.330 21.570 ;
        RECT 57.600 21.570 57.890 21.615 ;
        RECT 59.700 21.570 59.990 21.615 ;
        RECT 61.270 21.570 61.560 21.615 ;
        RECT 57.600 21.430 61.560 21.570 ;
        RECT 42.930 21.230 43.070 21.430 ;
        RECT 57.600 21.385 57.890 21.430 ;
        RECT 59.700 21.385 59.990 21.430 ;
        RECT 61.270 21.385 61.560 21.430 ;
        RECT 64.960 21.570 65.250 21.615 ;
        RECT 67.060 21.570 67.350 21.615 ;
        RECT 68.630 21.570 68.920 21.615 ;
        RECT 64.960 21.430 68.920 21.570 ;
        RECT 64.960 21.385 65.250 21.430 ;
        RECT 67.060 21.385 67.350 21.430 ;
        RECT 68.630 21.385 68.920 21.430 ;
        RECT 78.260 21.370 78.580 21.630 ;
        RECT 82.490 21.570 82.630 21.770 ;
        RECT 83.780 21.570 84.100 21.630 ;
        RECT 87.475 21.570 87.765 21.615 ;
        RECT 82.490 21.430 83.090 21.570 ;
        RECT 47.440 21.230 47.760 21.290 ;
        RECT 57.995 21.230 58.285 21.275 ;
        RECT 59.185 21.230 59.475 21.275 ;
        RECT 61.705 21.230 61.995 21.275 ;
        RECT 39.710 21.090 43.070 21.230 ;
        RECT 43.390 21.090 49.050 21.230 ;
        RECT 34.075 21.045 34.365 21.090 ;
        RECT 35.265 21.045 35.555 21.090 ;
        RECT 37.785 21.045 38.075 21.090 ;
        RECT 30.895 20.705 31.185 20.935 ;
        RECT 31.340 20.690 31.660 20.950 ;
        RECT 33.195 20.890 33.485 20.935 ;
        RECT 33.640 20.890 33.960 20.950 ;
        RECT 33.195 20.750 33.960 20.890 ;
        RECT 33.195 20.705 33.485 20.750 ;
        RECT 33.640 20.690 33.960 20.750 ;
        RECT 42.840 20.690 43.160 20.950 ;
        RECT 43.390 20.935 43.530 21.090 ;
        RECT 47.440 21.030 47.760 21.090 ;
        RECT 43.315 20.705 43.605 20.935 ;
        RECT 43.760 20.690 44.080 20.950 ;
        RECT 44.695 20.890 44.985 20.935 ;
        RECT 46.520 20.890 46.840 20.950 ;
        RECT 48.910 20.935 49.050 21.090 ;
        RECT 49.830 21.090 55.030 21.230 ;
        RECT 44.695 20.750 46.840 20.890 ;
        RECT 44.695 20.705 44.985 20.750 ;
        RECT 46.520 20.690 46.840 20.750 ;
        RECT 48.375 20.705 48.665 20.935 ;
        RECT 48.835 20.705 49.125 20.935 ;
        RECT 32.260 20.550 32.580 20.610 ;
        RECT 29.590 20.410 32.580 20.550 ;
        RECT 32.260 20.350 32.580 20.410 ;
        RECT 32.735 20.550 33.025 20.595 ;
        RECT 34.420 20.550 34.710 20.595 ;
        RECT 48.450 20.550 48.590 20.705 ;
        RECT 49.280 20.690 49.600 20.950 ;
        RECT 49.830 20.550 49.970 21.090 ;
        RECT 54.890 20.950 55.030 21.090 ;
        RECT 57.995 21.090 61.995 21.230 ;
        RECT 57.995 21.045 58.285 21.090 ;
        RECT 59.185 21.045 59.475 21.090 ;
        RECT 61.705 21.045 61.995 21.090 ;
        RECT 65.355 21.230 65.645 21.275 ;
        RECT 66.545 21.230 66.835 21.275 ;
        RECT 69.065 21.230 69.355 21.275 ;
        RECT 65.355 21.090 69.355 21.230 ;
        RECT 65.355 21.045 65.645 21.090 ;
        RECT 66.545 21.045 66.835 21.090 ;
        RECT 69.065 21.045 69.355 21.090 ;
        RECT 72.740 21.230 73.060 21.290 ;
        RECT 75.500 21.230 75.820 21.290 ;
        RECT 78.350 21.230 78.490 21.370 ;
        RECT 72.740 21.090 73.890 21.230 ;
        RECT 72.740 21.030 73.060 21.090 ;
        RECT 50.215 20.705 50.505 20.935 ;
        RECT 32.735 20.410 34.710 20.550 ;
        RECT 32.735 20.365 33.025 20.410 ;
        RECT 34.420 20.365 34.710 20.410 ;
        RECT 35.110 20.410 49.970 20.550 ;
        RECT 50.290 20.550 50.430 20.705 ;
        RECT 54.340 20.690 54.660 20.950 ;
        RECT 54.800 20.690 55.120 20.950 ;
        RECT 55.260 20.690 55.580 20.950 ;
        RECT 55.720 20.690 56.040 20.950 ;
        RECT 56.655 20.705 56.945 20.935 ;
        RECT 54.430 20.550 54.570 20.690 ;
        RECT 56.730 20.550 56.870 20.705 ;
        RECT 57.100 20.690 57.420 20.950 ;
        RECT 57.560 20.890 57.880 20.950 ;
        RECT 58.395 20.890 58.685 20.935 ;
        RECT 57.560 20.750 58.685 20.890 ;
        RECT 57.560 20.690 57.880 20.750 ;
        RECT 58.395 20.705 58.685 20.750 ;
        RECT 64.475 20.890 64.765 20.935 ;
        RECT 68.600 20.890 68.920 20.950 ;
        RECT 64.475 20.750 68.920 20.890 ;
        RECT 64.475 20.705 64.765 20.750 ;
        RECT 68.600 20.690 68.920 20.750 ;
        RECT 73.200 20.690 73.520 20.950 ;
        RECT 73.750 20.935 73.890 21.090 ;
        RECT 75.130 21.090 78.490 21.230 ;
        RECT 78.825 21.090 82.630 21.230 ;
        RECT 73.675 20.705 73.965 20.935 ;
        RECT 74.120 20.690 74.440 20.950 ;
        RECT 75.130 20.935 75.270 21.090 ;
        RECT 75.500 21.030 75.820 21.090 ;
        RECT 78.825 20.950 78.965 21.090 ;
        RECT 75.055 20.705 75.345 20.935 ;
        RECT 77.340 20.690 77.660 20.950 ;
        RECT 78.260 20.690 78.580 20.950 ;
        RECT 78.720 20.690 79.040 20.950 ;
        RECT 79.180 20.690 79.500 20.950 ;
        RECT 80.100 20.890 80.420 20.950 ;
        RECT 82.490 20.935 82.630 21.090 ;
        RECT 82.950 20.935 83.090 21.430 ;
        RECT 83.780 21.430 87.765 21.570 ;
        RECT 83.780 21.370 84.100 21.430 ;
        RECT 87.475 21.385 87.765 21.430 ;
        RECT 81.035 20.890 81.325 20.935 ;
        RECT 80.100 20.750 81.325 20.890 ;
        RECT 80.100 20.690 80.420 20.750 ;
        RECT 81.035 20.705 81.325 20.750 ;
        RECT 81.955 20.690 82.245 20.920 ;
        RECT 82.415 20.705 82.705 20.935 ;
        RECT 82.875 20.705 83.165 20.935 ;
        RECT 84.700 20.690 85.020 20.950 ;
        RECT 86.540 20.690 86.860 20.950 ;
        RECT 65.840 20.595 66.160 20.610 ;
        RECT 65.810 20.550 66.160 20.595 ;
        RECT 50.290 20.410 56.870 20.550 ;
        RECT 65.645 20.410 66.160 20.550 ;
        RECT 27.200 20.210 27.520 20.270 ;
        RECT 26.830 20.070 27.520 20.210 ;
        RECT 19.380 20.010 19.700 20.070 ;
        RECT 20.315 20.025 20.605 20.070 ;
        RECT 27.200 20.010 27.520 20.070 ;
        RECT 29.040 20.010 29.360 20.270 ;
        RECT 31.340 20.210 31.660 20.270 ;
        RECT 35.110 20.210 35.250 20.410 ;
        RECT 65.810 20.365 66.160 20.410 ;
        RECT 65.840 20.350 66.160 20.365 ;
        RECT 82.030 20.270 82.170 20.690 ;
        RECT 31.340 20.070 35.250 20.210 ;
        RECT 31.340 20.010 31.660 20.070 ;
        RECT 41.460 20.010 41.780 20.270 ;
        RECT 46.980 20.010 47.300 20.270 ;
        RECT 53.435 20.210 53.725 20.255 ;
        RECT 54.340 20.210 54.660 20.270 ;
        RECT 53.435 20.070 54.660 20.210 ;
        RECT 53.435 20.025 53.725 20.070 ;
        RECT 54.340 20.010 54.660 20.070 ;
        RECT 56.640 20.210 56.960 20.270 ;
        RECT 61.240 20.210 61.560 20.270 ;
        RECT 56.640 20.070 61.560 20.210 ;
        RECT 56.640 20.010 56.960 20.070 ;
        RECT 61.240 20.010 61.560 20.070 ;
        RECT 64.015 20.210 64.305 20.255 ;
        RECT 66.300 20.210 66.620 20.270 ;
        RECT 64.015 20.070 66.620 20.210 ;
        RECT 64.015 20.025 64.305 20.070 ;
        RECT 66.300 20.010 66.620 20.070 ;
        RECT 71.820 20.010 72.140 20.270 ;
        RECT 77.340 20.210 77.660 20.270 ;
        RECT 80.100 20.210 80.420 20.270 ;
        RECT 77.340 20.070 80.420 20.210 ;
        RECT 77.340 20.010 77.660 20.070 ;
        RECT 80.100 20.010 80.420 20.070 ;
        RECT 80.575 20.210 80.865 20.255 ;
        RECT 81.020 20.210 81.340 20.270 ;
        RECT 80.575 20.070 81.340 20.210 ;
        RECT 80.575 20.025 80.865 20.070 ;
        RECT 81.020 20.010 81.340 20.070 ;
        RECT 81.940 20.010 82.260 20.270 ;
        RECT 83.320 20.210 83.640 20.270 ;
        RECT 84.255 20.210 84.545 20.255 ;
        RECT 83.320 20.070 84.545 20.210 ;
        RECT 83.320 20.010 83.640 20.070 ;
        RECT 84.255 20.025 84.545 20.070 ;
        RECT 85.620 20.010 85.940 20.270 ;
        RECT 11.950 19.390 90.610 19.870 ;
        RECT 16.160 18.990 16.480 19.250 ;
        RECT 20.300 19.190 20.620 19.250 ;
        RECT 16.710 19.050 20.620 19.190 ;
        RECT 14.335 18.850 14.625 18.895 ;
        RECT 14.780 18.850 15.100 18.910 ;
        RECT 14.335 18.710 15.100 18.850 ;
        RECT 14.335 18.665 14.625 18.710 ;
        RECT 14.780 18.650 15.100 18.710 ;
        RECT 15.255 18.850 15.545 18.895 ;
        RECT 16.710 18.850 16.850 19.050 ;
        RECT 20.300 18.990 20.620 19.050 ;
        RECT 27.200 18.990 27.520 19.250 ;
        RECT 30.420 19.190 30.740 19.250 ;
        RECT 35.035 19.190 35.325 19.235 ;
        RECT 30.420 19.050 35.325 19.190 ;
        RECT 30.420 18.990 30.740 19.050 ;
        RECT 35.035 19.005 35.325 19.050 ;
        RECT 47.900 19.190 48.220 19.250 ;
        RECT 53.435 19.190 53.725 19.235 ;
        RECT 47.900 19.050 53.725 19.190 ;
        RECT 47.900 18.990 48.220 19.050 ;
        RECT 53.435 19.005 53.725 19.050 ;
        RECT 55.720 19.190 56.040 19.250 ;
        RECT 61.255 19.190 61.545 19.235 ;
        RECT 71.360 19.190 71.680 19.250 ;
        RECT 55.720 19.050 61.545 19.190 ;
        RECT 55.720 18.990 56.040 19.050 ;
        RECT 61.255 19.005 61.545 19.050 ;
        RECT 65.470 19.050 71.680 19.190 ;
        RECT 29.040 18.895 29.360 18.910 ;
        RECT 29.010 18.850 29.360 18.895 ;
        RECT 15.255 18.710 16.850 18.850 ;
        RECT 17.170 18.710 26.970 18.850 ;
        RECT 28.845 18.710 29.360 18.850 ;
        RECT 15.255 18.665 15.545 18.710 ;
        RECT 16.620 18.510 16.940 18.570 ;
        RECT 17.170 18.510 17.310 18.710 ;
        RECT 26.830 18.570 26.970 18.710 ;
        RECT 29.010 18.665 29.360 18.710 ;
        RECT 29.040 18.650 29.360 18.665 ;
        RECT 33.640 18.850 33.960 18.910 ;
        RECT 35.955 18.850 36.245 18.895 ;
        RECT 40.540 18.850 40.860 18.910 ;
        RECT 33.640 18.710 40.860 18.850 ;
        RECT 33.640 18.650 33.960 18.710 ;
        RECT 35.955 18.665 36.245 18.710 ;
        RECT 40.540 18.650 40.860 18.710 ;
        RECT 41.460 18.850 41.780 18.910 ;
        RECT 44.280 18.850 44.570 18.895 ;
        RECT 57.100 18.850 57.420 18.910 ;
        RECT 41.460 18.710 44.570 18.850 ;
        RECT 41.460 18.650 41.780 18.710 ;
        RECT 44.280 18.665 44.570 18.710 ;
        RECT 46.610 18.710 57.420 18.850 ;
        RECT 17.540 18.510 17.860 18.570 ;
        RECT 19.380 18.555 19.700 18.570 ;
        RECT 18.015 18.510 18.305 18.555 ;
        RECT 19.350 18.510 19.700 18.555 ;
        RECT 16.620 18.370 18.305 18.510 ;
        RECT 19.185 18.370 19.700 18.510 ;
        RECT 16.620 18.310 16.940 18.370 ;
        RECT 17.540 18.310 17.860 18.370 ;
        RECT 18.015 18.325 18.305 18.370 ;
        RECT 19.350 18.325 19.700 18.370 ;
        RECT 19.380 18.310 19.700 18.325 ;
        RECT 22.140 18.510 22.460 18.570 ;
        RECT 25.375 18.510 25.665 18.555 ;
        RECT 25.820 18.510 26.140 18.570 ;
        RECT 22.140 18.370 25.130 18.510 ;
        RECT 22.140 18.310 22.460 18.370 ;
        RECT 18.895 18.170 19.185 18.215 ;
        RECT 20.085 18.170 20.375 18.215 ;
        RECT 22.605 18.170 22.895 18.215 ;
        RECT 18.895 18.030 22.895 18.170 ;
        RECT 24.990 18.170 25.130 18.370 ;
        RECT 25.375 18.370 26.140 18.510 ;
        RECT 25.375 18.325 25.665 18.370 ;
        RECT 25.820 18.310 26.140 18.370 ;
        RECT 26.295 18.325 26.585 18.555 ;
        RECT 26.740 18.510 27.060 18.570 ;
        RECT 46.610 18.555 46.750 18.710 ;
        RECT 27.675 18.510 27.965 18.555 ;
        RECT 26.740 18.370 27.965 18.510 ;
        RECT 26.370 18.170 26.510 18.325 ;
        RECT 26.740 18.310 27.060 18.370 ;
        RECT 27.675 18.325 27.965 18.370 ;
        RECT 28.210 18.370 34.330 18.510 ;
        RECT 28.210 18.170 28.350 18.370 ;
        RECT 24.990 18.030 26.510 18.170 ;
        RECT 18.895 17.985 19.185 18.030 ;
        RECT 20.085 17.985 20.375 18.030 ;
        RECT 22.605 17.985 22.895 18.030 ;
        RECT 18.500 17.830 18.790 17.875 ;
        RECT 20.600 17.830 20.890 17.875 ;
        RECT 22.170 17.830 22.460 17.875 ;
        RECT 18.500 17.690 22.460 17.830 ;
        RECT 18.500 17.645 18.790 17.690 ;
        RECT 20.600 17.645 20.890 17.690 ;
        RECT 22.170 17.645 22.460 17.690 ;
        RECT 24.900 17.290 25.220 17.550 ;
        RECT 26.370 17.490 26.510 18.030 ;
        RECT 26.830 18.030 28.350 18.170 ;
        RECT 28.555 18.170 28.845 18.215 ;
        RECT 29.745 18.170 30.035 18.215 ;
        RECT 32.265 18.170 32.555 18.215 ;
        RECT 28.555 18.030 32.555 18.170 ;
        RECT 34.190 18.170 34.330 18.370 ;
        RECT 36.875 18.325 37.165 18.555 ;
        RECT 45.615 18.510 45.905 18.555 ;
        RECT 46.535 18.510 46.825 18.555 ;
        RECT 45.615 18.370 46.825 18.510 ;
        RECT 45.615 18.325 45.905 18.370 ;
        RECT 46.535 18.325 46.825 18.370 ;
        RECT 46.980 18.510 47.300 18.570 ;
        RECT 53.970 18.555 54.110 18.710 ;
        RECT 57.100 18.650 57.420 18.710 ;
        RECT 62.620 18.850 62.940 18.910 ;
        RECT 65.470 18.895 65.610 19.050 ;
        RECT 71.360 18.990 71.680 19.050 ;
        RECT 74.120 19.190 74.440 19.250 ;
        RECT 77.815 19.190 78.105 19.235 ;
        RECT 74.120 19.050 78.105 19.190 ;
        RECT 74.120 18.990 74.440 19.050 ;
        RECT 77.815 19.005 78.105 19.050 ;
        RECT 78.720 19.190 79.040 19.250 ;
        RECT 86.540 19.190 86.860 19.250 ;
        RECT 78.720 19.050 86.860 19.190 ;
        RECT 78.720 18.990 79.040 19.050 ;
        RECT 86.540 18.990 86.860 19.050 ;
        RECT 63.095 18.850 63.385 18.895 ;
        RECT 62.620 18.710 63.385 18.850 ;
        RECT 62.620 18.650 62.940 18.710 ;
        RECT 63.095 18.665 63.385 18.710 ;
        RECT 65.395 18.665 65.685 18.895 ;
        RECT 65.840 18.650 66.160 18.910 ;
        RECT 79.640 18.850 79.960 18.910 ;
        RECT 69.610 18.710 79.960 18.850 ;
        RECT 47.815 18.510 48.105 18.555 ;
        RECT 46.980 18.370 48.105 18.510 ;
        RECT 35.480 18.170 35.800 18.230 ;
        RECT 36.950 18.170 37.090 18.325 ;
        RECT 46.980 18.310 47.300 18.370 ;
        RECT 47.815 18.325 48.105 18.370 ;
        RECT 53.895 18.325 54.185 18.555 ;
        RECT 54.340 18.510 54.660 18.570 ;
        RECT 55.175 18.510 55.465 18.555 ;
        RECT 54.340 18.370 55.465 18.510 ;
        RECT 54.340 18.310 54.660 18.370 ;
        RECT 55.175 18.325 55.465 18.370 ;
        RECT 62.175 18.325 62.465 18.555 ;
        RECT 34.190 18.030 37.090 18.170 ;
        RECT 41.025 18.170 41.315 18.215 ;
        RECT 43.545 18.170 43.835 18.215 ;
        RECT 44.735 18.170 45.025 18.215 ;
        RECT 41.025 18.030 45.025 18.170 ;
        RECT 26.830 17.890 26.970 18.030 ;
        RECT 28.555 17.985 28.845 18.030 ;
        RECT 29.745 17.985 30.035 18.030 ;
        RECT 32.265 17.985 32.555 18.030 ;
        RECT 35.480 17.970 35.800 18.030 ;
        RECT 41.025 17.985 41.315 18.030 ;
        RECT 43.545 17.985 43.835 18.030 ;
        RECT 44.735 17.985 45.025 18.030 ;
        RECT 47.415 18.170 47.705 18.215 ;
        RECT 48.605 18.170 48.895 18.215 ;
        RECT 51.125 18.170 51.415 18.215 ;
        RECT 47.415 18.030 51.415 18.170 ;
        RECT 47.415 17.985 47.705 18.030 ;
        RECT 48.605 17.985 48.895 18.030 ;
        RECT 51.125 17.985 51.415 18.030 ;
        RECT 54.775 18.170 55.065 18.215 ;
        RECT 55.965 18.170 56.255 18.215 ;
        RECT 58.485 18.170 58.775 18.215 ;
        RECT 62.250 18.170 62.390 18.325 ;
        RECT 64.920 18.310 65.240 18.570 ;
        RECT 66.775 18.325 67.065 18.555 ;
        RECT 69.610 18.510 69.750 18.710 ;
        RECT 79.640 18.650 79.960 18.710 ;
        RECT 69.150 18.370 69.750 18.510 ;
        RECT 69.950 18.510 70.240 18.555 ;
        RECT 71.820 18.510 72.140 18.570 ;
        RECT 69.950 18.370 72.140 18.510 ;
        RECT 63.540 18.170 63.860 18.230 ;
        RECT 66.850 18.170 66.990 18.325 ;
        RECT 54.775 18.030 58.775 18.170 ;
        RECT 54.775 17.985 55.065 18.030 ;
        RECT 55.965 17.985 56.255 18.030 ;
        RECT 58.485 17.985 58.775 18.030 ;
        RECT 60.870 18.030 66.990 18.170 ;
        RECT 68.600 18.170 68.920 18.230 ;
        RECT 69.150 18.170 69.290 18.370 ;
        RECT 69.950 18.325 70.240 18.370 ;
        RECT 71.820 18.310 72.140 18.370 ;
        RECT 75.960 18.310 76.280 18.570 ;
        RECT 76.895 18.510 77.185 18.555 ;
        RECT 77.800 18.510 78.120 18.570 ;
        RECT 81.020 18.555 81.340 18.570 ;
        RECT 80.990 18.510 81.340 18.555 ;
        RECT 76.895 18.370 78.120 18.510 ;
        RECT 80.825 18.370 81.340 18.510 ;
        RECT 76.895 18.325 77.185 18.370 ;
        RECT 68.600 18.030 69.290 18.170 ;
        RECT 69.495 18.170 69.785 18.215 ;
        RECT 70.685 18.170 70.975 18.215 ;
        RECT 73.205 18.170 73.495 18.215 ;
        RECT 69.495 18.030 73.495 18.170 ;
        RECT 26.740 17.630 27.060 17.890 ;
        RECT 28.160 17.830 28.450 17.875 ;
        RECT 30.260 17.830 30.550 17.875 ;
        RECT 31.830 17.830 32.120 17.875 ;
        RECT 39.160 17.830 39.480 17.890 ;
        RECT 60.870 17.875 61.010 18.030 ;
        RECT 63.540 17.970 63.860 18.030 ;
        RECT 68.600 17.970 68.920 18.030 ;
        RECT 69.495 17.985 69.785 18.030 ;
        RECT 70.685 17.985 70.975 18.030 ;
        RECT 73.205 17.985 73.495 18.030 ;
        RECT 28.160 17.690 32.120 17.830 ;
        RECT 28.160 17.645 28.450 17.690 ;
        RECT 30.260 17.645 30.550 17.690 ;
        RECT 31.830 17.645 32.120 17.690 ;
        RECT 34.650 17.690 39.480 17.830 ;
        RECT 34.650 17.535 34.790 17.690 ;
        RECT 39.160 17.630 39.480 17.690 ;
        RECT 41.460 17.830 41.750 17.875 ;
        RECT 43.030 17.830 43.320 17.875 ;
        RECT 45.130 17.830 45.420 17.875 ;
        RECT 41.460 17.690 45.420 17.830 ;
        RECT 41.460 17.645 41.750 17.690 ;
        RECT 43.030 17.645 43.320 17.690 ;
        RECT 45.130 17.645 45.420 17.690 ;
        RECT 47.020 17.830 47.310 17.875 ;
        RECT 49.120 17.830 49.410 17.875 ;
        RECT 50.690 17.830 50.980 17.875 ;
        RECT 47.020 17.690 50.980 17.830 ;
        RECT 47.020 17.645 47.310 17.690 ;
        RECT 49.120 17.645 49.410 17.690 ;
        RECT 50.690 17.645 50.980 17.690 ;
        RECT 54.380 17.830 54.670 17.875 ;
        RECT 56.480 17.830 56.770 17.875 ;
        RECT 58.050 17.830 58.340 17.875 ;
        RECT 54.380 17.690 58.340 17.830 ;
        RECT 54.380 17.645 54.670 17.690 ;
        RECT 56.480 17.645 56.770 17.690 ;
        RECT 58.050 17.645 58.340 17.690 ;
        RECT 60.795 17.645 61.085 17.875 ;
        RECT 61.240 17.830 61.560 17.890 ;
        RECT 69.100 17.830 69.390 17.875 ;
        RECT 71.200 17.830 71.490 17.875 ;
        RECT 72.770 17.830 73.060 17.875 ;
        RECT 61.240 17.690 68.600 17.830 ;
        RECT 61.240 17.630 61.560 17.690 ;
        RECT 34.575 17.490 34.865 17.535 ;
        RECT 26.370 17.350 34.865 17.490 ;
        RECT 34.575 17.305 34.865 17.350 ;
        RECT 37.320 17.490 37.640 17.550 ;
        RECT 38.715 17.490 39.005 17.535 ;
        RECT 37.320 17.350 39.005 17.490 ;
        RECT 37.320 17.290 37.640 17.350 ;
        RECT 38.715 17.305 39.005 17.350 ;
        RECT 52.040 17.490 52.360 17.550 ;
        RECT 64.015 17.490 64.305 17.535 ;
        RECT 52.040 17.350 64.305 17.490 ;
        RECT 68.460 17.490 68.600 17.690 ;
        RECT 69.100 17.690 73.060 17.830 ;
        RECT 69.100 17.645 69.390 17.690 ;
        RECT 71.200 17.645 71.490 17.690 ;
        RECT 72.770 17.645 73.060 17.690 ;
        RECT 75.515 17.830 75.805 17.875 ;
        RECT 75.960 17.830 76.280 17.890 ;
        RECT 76.970 17.830 77.110 18.325 ;
        RECT 77.800 18.310 78.120 18.370 ;
        RECT 80.990 18.325 81.340 18.370 ;
        RECT 81.020 18.310 81.340 18.325 ;
        RECT 82.400 18.510 82.720 18.570 ;
        RECT 87.015 18.510 87.305 18.555 ;
        RECT 82.400 18.370 87.305 18.510 ;
        RECT 82.400 18.310 82.720 18.370 ;
        RECT 87.015 18.325 87.305 18.370 ;
        RECT 79.640 17.970 79.960 18.230 ;
        RECT 80.535 18.170 80.825 18.215 ;
        RECT 81.725 18.170 82.015 18.215 ;
        RECT 84.245 18.170 84.535 18.215 ;
        RECT 80.535 18.030 84.535 18.170 ;
        RECT 80.535 17.985 80.825 18.030 ;
        RECT 81.725 17.985 82.015 18.030 ;
        RECT 84.245 17.985 84.535 18.030 ;
        RECT 75.515 17.690 77.110 17.830 ;
        RECT 80.140 17.830 80.430 17.875 ;
        RECT 82.240 17.830 82.530 17.875 ;
        RECT 83.810 17.830 84.100 17.875 ;
        RECT 80.140 17.690 84.100 17.830 ;
        RECT 75.515 17.645 75.805 17.690 ;
        RECT 75.960 17.630 76.280 17.690 ;
        RECT 80.140 17.645 80.430 17.690 ;
        RECT 82.240 17.645 82.530 17.690 ;
        RECT 83.810 17.645 84.100 17.690 ;
        RECT 79.180 17.490 79.500 17.550 ;
        RECT 68.460 17.350 79.500 17.490 ;
        RECT 52.040 17.290 52.360 17.350 ;
        RECT 64.015 17.305 64.305 17.350 ;
        RECT 79.180 17.290 79.500 17.350 ;
        RECT 87.920 17.290 88.240 17.550 ;
        RECT 11.950 16.670 90.610 17.150 ;
        RECT 20.300 16.270 20.620 16.530 ;
        RECT 21.695 16.470 21.985 16.515 ;
        RECT 22.600 16.470 22.920 16.530 ;
        RECT 41.000 16.470 41.320 16.530 ;
        RECT 21.695 16.330 22.920 16.470 ;
        RECT 21.695 16.285 21.985 16.330 ;
        RECT 22.600 16.270 22.920 16.330 ;
        RECT 31.890 16.330 41.320 16.470 ;
        RECT 13.900 16.130 14.190 16.175 ;
        RECT 16.000 16.130 16.290 16.175 ;
        RECT 17.570 16.130 17.860 16.175 ;
        RECT 13.900 15.990 17.860 16.130 ;
        RECT 13.900 15.945 14.190 15.990 ;
        RECT 16.000 15.945 16.290 15.990 ;
        RECT 17.570 15.945 17.860 15.990 ;
        RECT 14.295 15.790 14.585 15.835 ;
        RECT 15.485 15.790 15.775 15.835 ;
        RECT 18.005 15.790 18.295 15.835 ;
        RECT 14.295 15.650 18.295 15.790 ;
        RECT 14.295 15.605 14.585 15.650 ;
        RECT 15.485 15.605 15.775 15.650 ;
        RECT 18.005 15.605 18.295 15.650 ;
        RECT 13.415 15.450 13.705 15.495 ;
        RECT 17.540 15.450 17.860 15.510 ;
        RECT 13.415 15.310 17.860 15.450 ;
        RECT 13.415 15.265 13.705 15.310 ;
        RECT 17.540 15.250 17.860 15.310 ;
        RECT 22.615 15.450 22.905 15.495 ;
        RECT 24.900 15.450 25.220 15.510 ;
        RECT 22.615 15.310 25.220 15.450 ;
        RECT 22.615 15.265 22.905 15.310 ;
        RECT 24.900 15.250 25.220 15.310 ;
        RECT 27.675 15.450 27.965 15.495 ;
        RECT 29.500 15.450 29.820 15.510 ;
        RECT 27.675 15.310 29.820 15.450 ;
        RECT 27.675 15.265 27.965 15.310 ;
        RECT 29.500 15.250 29.820 15.310 ;
        RECT 29.960 15.250 30.280 15.510 ;
        RECT 31.890 15.495 32.030 16.330 ;
        RECT 41.000 16.270 41.320 16.330 ;
        RECT 43.760 16.470 44.080 16.530 ;
        RECT 44.235 16.470 44.525 16.515 ;
        RECT 43.760 16.330 44.525 16.470 ;
        RECT 43.760 16.270 44.080 16.330 ;
        RECT 44.235 16.285 44.525 16.330 ;
        RECT 49.280 16.470 49.600 16.530 ;
        RECT 50.215 16.470 50.505 16.515 ;
        RECT 49.280 16.330 50.505 16.470 ;
        RECT 49.280 16.270 49.600 16.330 ;
        RECT 50.215 16.285 50.505 16.330 ;
        RECT 78.260 16.470 78.580 16.530 ;
        RECT 78.735 16.470 79.025 16.515 ;
        RECT 78.260 16.330 79.025 16.470 ;
        RECT 78.260 16.270 78.580 16.330 ;
        RECT 78.735 16.285 79.025 16.330 ;
        RECT 81.035 16.470 81.325 16.515 ;
        RECT 81.940 16.470 82.260 16.530 ;
        RECT 81.035 16.330 82.260 16.470 ;
        RECT 81.035 16.285 81.325 16.330 ;
        RECT 81.940 16.270 82.260 16.330 ;
        RECT 32.735 16.130 33.025 16.175 ;
        RECT 35.480 16.130 35.800 16.190 ;
        RECT 32.735 15.990 35.800 16.130 ;
        RECT 32.735 15.945 33.025 15.990 ;
        RECT 35.480 15.930 35.800 15.990 ;
        RECT 41.935 16.130 42.225 16.175 ;
        RECT 46.520 16.130 46.840 16.190 ;
        RECT 41.935 15.990 46.840 16.130 ;
        RECT 41.935 15.945 42.225 15.990 ;
        RECT 46.520 15.930 46.840 15.990 ;
        RECT 82.440 16.130 82.730 16.175 ;
        RECT 84.540 16.130 84.830 16.175 ;
        RECT 86.110 16.130 86.400 16.175 ;
        RECT 82.440 15.990 86.400 16.130 ;
        RECT 82.440 15.945 82.730 15.990 ;
        RECT 84.540 15.945 84.830 15.990 ;
        RECT 86.110 15.945 86.400 15.990 ;
        RECT 53.880 15.790 54.200 15.850 ;
        RECT 67.680 15.790 68.000 15.850 ;
        RECT 78.720 15.790 79.040 15.850 ;
        RECT 37.410 15.650 43.530 15.790 ;
        RECT 37.410 15.510 37.550 15.650 ;
        RECT 31.815 15.265 32.105 15.495 ;
        RECT 33.640 15.250 33.960 15.510 ;
        RECT 35.495 15.450 35.785 15.495 ;
        RECT 36.400 15.450 36.720 15.510 ;
        RECT 35.495 15.310 36.720 15.450 ;
        RECT 35.495 15.265 35.785 15.310 ;
        RECT 36.400 15.250 36.720 15.310 ;
        RECT 37.320 15.250 37.640 15.510 ;
        RECT 39.160 15.250 39.480 15.510 ;
        RECT 39.620 15.450 39.940 15.510 ;
        RECT 40.630 15.495 40.770 15.650 ;
        RECT 40.095 15.450 40.385 15.495 ;
        RECT 39.620 15.310 40.385 15.450 ;
        RECT 39.620 15.250 39.940 15.310 ;
        RECT 40.095 15.265 40.385 15.310 ;
        RECT 40.555 15.265 40.845 15.495 ;
        RECT 41.015 15.450 41.305 15.495 ;
        RECT 42.840 15.450 43.160 15.510 ;
        RECT 43.390 15.495 43.530 15.650 ;
        RECT 53.880 15.650 58.710 15.790 ;
        RECT 53.880 15.590 54.200 15.650 ;
        RECT 41.015 15.310 43.160 15.450 ;
        RECT 41.015 15.265 41.305 15.310 ;
        RECT 42.840 15.250 43.160 15.310 ;
        RECT 43.315 15.265 43.605 15.495 ;
        RECT 44.220 15.450 44.540 15.510 ;
        RECT 46.075 15.450 46.365 15.495 ;
        RECT 44.220 15.310 46.365 15.450 ;
        RECT 44.220 15.250 44.540 15.310 ;
        RECT 46.075 15.265 46.365 15.310 ;
        RECT 46.535 15.450 46.825 15.495 ;
        RECT 47.900 15.450 48.220 15.510 ;
        RECT 49.295 15.450 49.585 15.495 ;
        RECT 46.535 15.310 49.585 15.450 ;
        RECT 46.535 15.265 46.825 15.310 ;
        RECT 47.900 15.250 48.220 15.310 ;
        RECT 49.295 15.265 49.585 15.310 ;
        RECT 53.435 15.450 53.725 15.495 ;
        RECT 56.180 15.450 56.500 15.510 ;
        RECT 58.570 15.495 58.710 15.650 ;
        RECT 67.680 15.650 79.040 15.790 ;
        RECT 67.680 15.590 68.000 15.650 ;
        RECT 53.435 15.310 56.500 15.450 ;
        RECT 53.435 15.265 53.725 15.310 ;
        RECT 56.180 15.250 56.500 15.310 ;
        RECT 56.655 15.265 56.945 15.495 ;
        RECT 58.495 15.265 58.785 15.495 ;
        RECT 63.095 15.450 63.385 15.495 ;
        RECT 63.540 15.450 63.860 15.510 ;
        RECT 63.095 15.310 63.860 15.450 ;
        RECT 63.095 15.265 63.385 15.310 ;
        RECT 13.860 15.110 14.180 15.170 ;
        RECT 14.640 15.110 14.930 15.155 ;
        RECT 13.860 14.970 14.930 15.110 ;
        RECT 13.860 14.910 14.180 14.970 ;
        RECT 14.640 14.925 14.930 14.970 ;
        RECT 23.535 15.110 23.825 15.155 ;
        RECT 25.360 15.110 25.680 15.170 ;
        RECT 38.700 15.110 39.020 15.170 ;
        RECT 23.535 14.970 25.680 15.110 ;
        RECT 23.535 14.925 23.825 14.970 ;
        RECT 25.360 14.910 25.680 14.970 ;
        RECT 34.650 14.970 39.020 15.110 ;
        RECT 25.820 14.770 26.140 14.830 ;
        RECT 26.755 14.770 27.045 14.815 ;
        RECT 25.820 14.630 27.045 14.770 ;
        RECT 25.820 14.570 26.140 14.630 ;
        RECT 26.755 14.585 27.045 14.630 ;
        RECT 29.040 14.570 29.360 14.830 ;
        RECT 30.895 14.770 31.185 14.815 ;
        RECT 32.260 14.770 32.580 14.830 ;
        RECT 34.650 14.815 34.790 14.970 ;
        RECT 38.700 14.910 39.020 14.970 ;
        RECT 42.395 15.110 42.685 15.155 ;
        RECT 48.360 15.110 48.680 15.170 ;
        RECT 42.395 14.970 48.680 15.110 ;
        RECT 56.730 15.110 56.870 15.265 ;
        RECT 63.540 15.250 63.860 15.310 ;
        RECT 66.300 15.250 66.620 15.510 ;
        RECT 69.520 15.250 69.840 15.510 ;
        RECT 71.360 15.250 71.680 15.510 ;
        RECT 75.960 15.250 76.280 15.510 ;
        RECT 77.890 15.495 78.030 15.650 ;
        RECT 78.720 15.590 79.040 15.650 ;
        RECT 79.640 15.790 79.960 15.850 ;
        RECT 81.955 15.790 82.245 15.835 ;
        RECT 79.640 15.650 82.245 15.790 ;
        RECT 79.640 15.590 79.960 15.650 ;
        RECT 81.955 15.605 82.245 15.650 ;
        RECT 82.835 15.790 83.125 15.835 ;
        RECT 84.025 15.790 84.315 15.835 ;
        RECT 86.545 15.790 86.835 15.835 ;
        RECT 82.835 15.650 86.835 15.790 ;
        RECT 82.835 15.605 83.125 15.650 ;
        RECT 84.025 15.605 84.315 15.650 ;
        RECT 86.545 15.605 86.835 15.650 ;
        RECT 83.320 15.495 83.640 15.510 ;
        RECT 77.815 15.265 78.105 15.495 ;
        RECT 83.290 15.450 83.640 15.495 ;
        RECT 83.125 15.310 83.640 15.450 ;
        RECT 83.290 15.265 83.640 15.310 ;
        RECT 83.320 15.250 83.640 15.265 ;
        RECT 61.700 15.110 62.020 15.170 ;
        RECT 56.730 14.970 62.020 15.110 ;
        RECT 42.395 14.925 42.685 14.970 ;
        RECT 48.360 14.910 48.680 14.970 ;
        RECT 61.700 14.910 62.020 14.970 ;
        RECT 72.740 15.110 73.060 15.170 ;
        RECT 76.895 15.110 77.185 15.155 ;
        RECT 79.195 15.110 79.485 15.155 ;
        RECT 72.740 14.970 79.485 15.110 ;
        RECT 72.740 14.910 73.060 14.970 ;
        RECT 76.895 14.925 77.185 14.970 ;
        RECT 79.195 14.925 79.485 14.970 ;
        RECT 80.115 15.110 80.405 15.155 ;
        RECT 84.240 15.110 84.560 15.170 ;
        RECT 80.115 14.970 89.070 15.110 ;
        RECT 80.115 14.925 80.405 14.970 ;
        RECT 84.240 14.910 84.560 14.970 ;
        RECT 30.895 14.630 32.580 14.770 ;
        RECT 30.895 14.585 31.185 14.630 ;
        RECT 32.260 14.570 32.580 14.630 ;
        RECT 34.575 14.585 34.865 14.815 ;
        RECT 36.415 14.770 36.705 14.815 ;
        RECT 41.460 14.770 41.780 14.830 ;
        RECT 36.415 14.630 41.780 14.770 ;
        RECT 36.415 14.585 36.705 14.630 ;
        RECT 41.460 14.570 41.780 14.630 ;
        RECT 45.140 14.570 45.460 14.830 ;
        RECT 47.455 14.770 47.745 14.815 ;
        RECT 47.900 14.770 48.220 14.830 ;
        RECT 47.455 14.630 48.220 14.770 ;
        RECT 47.455 14.585 47.745 14.630 ;
        RECT 47.900 14.570 48.220 14.630 ;
        RECT 51.580 14.770 51.900 14.830 ;
        RECT 52.515 14.770 52.805 14.815 ;
        RECT 51.580 14.630 52.805 14.770 ;
        RECT 51.580 14.570 51.900 14.630 ;
        RECT 52.515 14.585 52.805 14.630 ;
        RECT 54.800 14.770 55.120 14.830 ;
        RECT 55.735 14.770 56.025 14.815 ;
        RECT 54.800 14.630 56.025 14.770 ;
        RECT 54.800 14.570 55.120 14.630 ;
        RECT 55.735 14.585 56.025 14.630 ;
        RECT 58.020 14.770 58.340 14.830 ;
        RECT 59.415 14.770 59.705 14.815 ;
        RECT 58.020 14.630 59.705 14.770 ;
        RECT 58.020 14.570 58.340 14.630 ;
        RECT 59.415 14.585 59.705 14.630 ;
        RECT 61.240 14.770 61.560 14.830 ;
        RECT 62.175 14.770 62.465 14.815 ;
        RECT 61.240 14.630 62.465 14.770 ;
        RECT 61.240 14.570 61.560 14.630 ;
        RECT 62.175 14.585 62.465 14.630 ;
        RECT 64.460 14.770 64.780 14.830 ;
        RECT 65.395 14.770 65.685 14.815 ;
        RECT 64.460 14.630 65.685 14.770 ;
        RECT 64.460 14.570 64.780 14.630 ;
        RECT 65.395 14.585 65.685 14.630 ;
        RECT 67.680 14.770 68.000 14.830 ;
        RECT 68.615 14.770 68.905 14.815 ;
        RECT 67.680 14.630 68.905 14.770 ;
        RECT 67.680 14.570 68.000 14.630 ;
        RECT 68.615 14.585 68.905 14.630 ;
        RECT 70.900 14.770 71.220 14.830 ;
        RECT 72.295 14.770 72.585 14.815 ;
        RECT 70.900 14.630 72.585 14.770 ;
        RECT 70.900 14.570 71.220 14.630 ;
        RECT 72.295 14.585 72.585 14.630 ;
        RECT 74.120 14.770 74.440 14.830 ;
        RECT 88.930 14.815 89.070 14.970 ;
        RECT 75.055 14.770 75.345 14.815 ;
        RECT 74.120 14.630 75.345 14.770 ;
        RECT 74.120 14.570 74.440 14.630 ;
        RECT 75.055 14.585 75.345 14.630 ;
        RECT 88.855 14.585 89.145 14.815 ;
        RECT 11.950 13.950 90.610 14.430 ;
        RECT 6.500 10.010 6.820 10.070 ;
        RECT 14.320 10.010 14.640 10.070 ;
        RECT 6.500 9.870 14.640 10.010 ;
        RECT 6.500 9.810 6.820 9.870 ;
        RECT 14.320 9.810 14.640 9.870 ;
        RECT 77.340 10.010 77.660 10.070 ;
        RECT 87.920 10.010 88.240 10.070 ;
        RECT 77.340 9.870 88.240 10.010 ;
        RECT 77.340 9.810 77.660 9.870 ;
        RECT 87.920 9.810 88.240 9.870 ;
        RECT 9.720 9.670 10.040 9.730 ;
        RECT 18.000 9.670 18.320 9.730 ;
        RECT 9.720 9.530 18.320 9.670 ;
        RECT 9.720 9.470 10.040 9.530 ;
        RECT 18.000 9.470 18.320 9.530 ;
        RECT 80.560 8.990 80.880 9.050 ;
        RECT 85.620 8.990 85.940 9.050 ;
        RECT 80.560 8.850 85.940 8.990 ;
        RECT 80.560 8.790 80.880 8.850 ;
        RECT 85.620 8.790 85.940 8.850 ;
      LAYER met2 ;
        RECT 69.205 222.560 69.595 222.640 ;
        RECT 69.205 222.420 127.660 222.560 ;
        RECT 69.205 222.340 69.595 222.420 ;
        RECT 72.120 222.090 72.420 222.215 ;
        RECT 72.120 221.950 126.920 222.090 ;
        RECT 72.120 221.825 72.420 221.950 ;
        RECT 74.770 221.725 75.160 221.785 ;
        RECT 125.240 221.770 125.770 221.780 ;
        RECT 125.240 221.725 125.805 221.770 ;
        RECT 74.770 221.540 125.805 221.725 ;
        RECT 74.770 221.485 75.160 221.540 ;
        RECT 125.240 221.490 125.805 221.540 ;
        RECT 126.780 221.620 126.920 221.950 ;
        RECT 127.520 222.060 127.660 222.420 ;
        RECT 149.680 222.060 150.000 222.120 ;
        RECT 127.520 221.920 150.000 222.060 ;
        RECT 149.680 221.860 150.000 221.920 ;
        RECT 125.240 221.480 125.770 221.490 ;
        RECT 126.780 221.480 140.200 221.620 ;
        RECT 138.880 221.310 139.370 221.320 ;
        RECT 80.275 221.240 80.665 221.305 ;
        RECT 82.770 221.240 83.840 221.280 ;
        RECT 80.275 221.160 117.550 221.240 ;
        RECT 138.880 221.160 139.405 221.310 ;
        RECT 80.275 221.120 139.405 221.160 ;
        RECT 80.275 221.070 82.940 221.120 ;
        RECT 83.620 221.070 139.405 221.120 ;
        RECT 80.275 221.005 80.665 221.070 ;
        RECT 117.055 221.030 139.405 221.070 ;
        RECT 117.055 221.020 139.370 221.030 ;
        RECT 83.085 220.900 83.475 220.980 ;
        RECT 117.055 220.965 139.130 221.020 ;
        RECT 140.060 221.000 140.200 221.480 ;
        RECT 149.120 221.000 149.440 221.060 ;
        RECT 83.085 220.800 116.760 220.900 ;
        RECT 140.060 220.860 149.440 221.000 ;
        RECT 149.120 220.800 149.440 220.860 ;
        RECT 83.085 220.760 133.370 220.800 ;
        RECT 83.085 220.680 83.475 220.760 ;
        RECT 116.620 220.660 133.370 220.760 ;
        RECT 85.785 220.525 86.175 220.595 ;
        RECT 115.915 220.580 116.285 220.585 ;
        RECT 115.570 220.525 116.285 220.580 ;
        RECT 85.785 220.365 116.285 220.525 ;
        RECT 85.785 220.295 86.175 220.365 ;
        RECT 115.570 220.310 116.285 220.365 ;
        RECT 115.915 220.305 116.285 220.310 ;
        RECT 91.280 220.140 91.670 220.220 ;
        RECT 132.220 220.210 132.610 220.480 ;
        RECT 93.670 220.140 94.650 220.160 ;
        RECT 116.845 220.140 132.610 220.210 ;
        RECT 91.280 220.040 132.610 220.140 ;
        RECT 133.230 220.250 133.370 220.660 ;
        RECT 148.660 220.250 148.920 220.340 ;
        RECT 133.230 220.110 148.920 220.250 ;
        RECT 91.280 220.035 132.510 220.040 ;
        RECT 91.280 220.020 117.005 220.035 ;
        RECT 148.660 220.020 148.920 220.110 ;
        RECT 91.280 219.995 93.810 220.020 ;
        RECT 94.490 220.000 117.005 220.020 ;
        RECT 94.490 219.995 116.860 220.000 ;
        RECT 91.280 219.920 91.670 219.995 ;
        RECT 93.955 219.800 94.345 219.880 ;
        RECT 148.110 219.800 148.430 219.860 ;
        RECT 93.955 219.660 148.430 219.800 ;
        RECT 88.600 219.490 88.900 219.615 ;
        RECT 93.955 219.580 94.345 219.660 ;
        RECT 148.110 219.600 148.430 219.660 ;
        RECT 88.600 219.440 93.810 219.490 ;
        RECT 94.490 219.440 111.950 219.490 ;
        RECT 88.600 219.350 111.950 219.440 ;
        RECT 88.600 219.225 88.900 219.350 ;
        RECT 93.560 219.310 94.730 219.350 ;
        RECT 93.670 219.290 94.610 219.310 ;
        RECT 77.535 219.090 77.925 219.170 ;
        RECT 96.090 219.090 111.560 219.180 ;
        RECT 77.535 219.080 88.440 219.090 ;
        RECT 89.070 219.080 111.560 219.090 ;
        RECT 77.535 219.040 111.560 219.080 ;
        RECT 77.535 218.950 96.230 219.040 ;
        RECT 77.535 218.870 77.925 218.950 ;
        RECT 88.330 218.940 89.190 218.950 ;
        RECT 66.485 218.730 66.875 218.810 ;
        RECT 96.750 218.730 111.150 218.830 ;
        RECT 66.485 218.690 111.150 218.730 ;
        RECT 66.485 218.590 96.890 218.690 ;
        RECT 66.485 218.510 66.875 218.590 ;
        RECT 63.655 218.200 64.045 218.280 ;
        RECT 63.655 218.060 110.150 218.200 ;
        RECT 63.655 217.980 64.045 218.060 ;
        RECT 61.260 209.310 61.540 213.310 ;
        RECT 70.920 209.310 71.200 213.310 ;
        RECT 27.500 201.685 29.040 202.055 ;
        RECT 49.770 201.200 50.030 201.520 ;
        RECT 47.470 199.840 47.730 200.160 ;
        RECT 6.980 198.625 7.260 198.995 ;
        RECT 30.800 198.965 32.340 199.335 ;
        RECT 7.050 113.120 7.190 198.625 ;
        RECT 41.490 198.140 41.750 198.460 ;
        RECT 43.330 198.140 43.590 198.460 ;
        RECT 41.030 197.800 41.290 198.120 ;
        RECT 36.890 197.460 37.150 197.780 ;
        RECT 27.500 196.245 29.040 196.615 ;
        RECT 36.950 195.400 37.090 197.460 ;
        RECT 36.890 195.080 37.150 195.400 ;
        RECT 30.800 193.525 32.340 193.895 ;
        RECT 27.500 190.805 29.040 191.175 ;
        RECT 30.800 188.085 32.340 188.455 ;
        RECT 21.250 187.260 21.510 187.580 ;
        RECT 16.650 186.580 16.910 186.900 ;
        RECT 16.710 185.200 16.850 186.580 ;
        RECT 20.330 185.900 20.590 186.220 ;
        RECT 16.650 184.880 16.910 185.200 ;
        RECT 20.390 184.180 20.530 185.900 ;
        RECT 17.110 183.860 17.370 184.180 ;
        RECT 20.330 183.860 20.590 184.180 ;
        RECT 17.170 181.800 17.310 183.860 ;
        RECT 21.310 182.480 21.450 187.260 ;
        RECT 36.950 187.240 37.090 195.080 ;
        RECT 39.650 194.400 39.910 194.720 ;
        RECT 39.710 193.360 39.850 194.400 ;
        RECT 39.650 193.040 39.910 193.360 ;
        RECT 41.090 191.660 41.230 197.800 ;
        RECT 41.550 193.020 41.690 198.140 ;
        RECT 41.950 198.030 42.210 198.120 ;
        RECT 41.950 197.890 42.610 198.030 ;
        RECT 41.950 197.800 42.210 197.890 ;
        RECT 41.950 196.780 42.210 197.100 ;
        RECT 42.010 193.360 42.150 196.780 ;
        RECT 42.470 193.360 42.610 197.890 ;
        RECT 43.390 195.740 43.530 198.140 ;
        RECT 47.530 198.120 47.670 199.840 ;
        RECT 47.470 197.800 47.730 198.120 ;
        RECT 46.090 196.780 46.350 197.100 ;
        RECT 46.150 196.080 46.290 196.780 ;
        RECT 45.170 195.760 45.430 196.080 ;
        RECT 46.090 195.760 46.350 196.080 ;
        RECT 43.330 195.420 43.590 195.740 ;
        RECT 44.250 194.060 44.510 194.380 ;
        RECT 44.710 194.060 44.970 194.380 ;
        RECT 41.950 193.040 42.210 193.360 ;
        RECT 42.410 193.040 42.670 193.360 ;
        RECT 41.490 192.700 41.750 193.020 ;
        RECT 40.570 191.340 40.830 191.660 ;
        RECT 41.030 191.340 41.290 191.660 ;
        RECT 40.630 190.640 40.770 191.340 ;
        RECT 40.570 190.320 40.830 190.640 ;
        RECT 40.110 188.620 40.370 188.940 ;
        RECT 40.170 187.580 40.310 188.620 ;
        RECT 40.110 187.260 40.370 187.580 ;
        RECT 26.770 186.920 27.030 187.240 ;
        RECT 36.890 186.920 37.150 187.240 ;
        RECT 24.470 186.580 24.730 186.900 ;
        RECT 24.530 184.180 24.670 186.580 ;
        RECT 26.310 185.900 26.570 186.220 ;
        RECT 26.370 184.600 26.510 185.900 ;
        RECT 26.830 185.200 26.970 186.920 ;
        RECT 33.210 185.900 33.470 186.220 ;
        RECT 27.500 185.365 29.040 185.735 ;
        RECT 26.770 184.880 27.030 185.200 ;
        RECT 27.230 184.880 27.490 185.200 ;
        RECT 27.290 184.600 27.430 184.880 ;
        RECT 26.370 184.460 27.430 184.600 ;
        RECT 24.470 183.860 24.730 184.180 ;
        RECT 22.630 183.180 22.890 183.500 ;
        RECT 21.250 182.160 21.510 182.480 ;
        RECT 22.690 182.140 22.830 183.180 ;
        RECT 22.630 181.820 22.890 182.140 ;
        RECT 17.110 181.480 17.370 181.800 ;
        RECT 17.170 179.760 17.310 181.480 ;
        RECT 17.110 179.440 17.370 179.760 ;
        RECT 17.170 176.700 17.310 179.440 ;
        RECT 24.530 178.740 24.670 183.860 ;
        RECT 27.290 181.200 27.430 184.460 ;
        RECT 29.990 184.200 30.250 184.520 ;
        RECT 30.510 184.460 31.570 184.600 ;
        RECT 29.070 183.860 29.330 184.180 ;
        RECT 29.130 182.140 29.270 183.860 ;
        RECT 29.530 183.180 29.790 183.500 ;
        RECT 29.070 181.820 29.330 182.140 ;
        RECT 26.370 181.060 27.430 181.200 ;
        RECT 24.470 178.420 24.730 178.740 ;
        RECT 26.370 178.480 26.510 181.060 ;
        RECT 27.230 180.690 27.490 180.780 ;
        RECT 26.830 180.550 27.490 180.690 ;
        RECT 26.830 179.420 26.970 180.550 ;
        RECT 27.230 180.460 27.490 180.550 ;
        RECT 27.500 179.925 29.040 180.295 ;
        RECT 29.590 179.760 29.730 183.180 ;
        RECT 30.050 181.710 30.190 184.200 ;
        RECT 30.510 184.180 30.650 184.460 ;
        RECT 30.450 183.860 30.710 184.180 ;
        RECT 30.910 183.860 31.170 184.180 ;
        RECT 30.970 183.410 31.110 183.860 ;
        RECT 31.430 183.500 31.570 184.460 ;
        RECT 33.270 184.180 33.410 185.900 ;
        RECT 33.210 183.860 33.470 184.180 ;
        RECT 34.590 183.860 34.850 184.180 ;
        RECT 35.970 183.860 36.230 184.180 ;
        RECT 32.290 183.750 32.550 183.840 ;
        RECT 32.290 183.610 32.950 183.750 ;
        RECT 32.290 183.520 32.550 183.610 ;
        RECT 30.510 183.270 31.110 183.410 ;
        RECT 30.510 182.480 30.650 183.270 ;
        RECT 31.370 183.180 31.630 183.500 ;
        RECT 30.800 182.645 32.340 183.015 ;
        RECT 32.810 182.480 32.950 183.610 ;
        RECT 33.210 183.180 33.470 183.500 ;
        RECT 30.450 182.160 30.710 182.480 ;
        RECT 32.750 182.160 33.010 182.480 ;
        RECT 30.450 181.710 30.710 181.800 ;
        RECT 30.050 181.570 30.710 181.710 ;
        RECT 30.450 181.480 30.710 181.570 ;
        RECT 33.270 181.460 33.410 183.180 ;
        RECT 34.130 182.160 34.390 182.480 ;
        RECT 34.190 181.800 34.330 182.160 ;
        RECT 34.650 181.800 34.790 183.860 ;
        RECT 34.130 181.480 34.390 181.800 ;
        RECT 34.590 181.480 34.850 181.800 ;
        RECT 35.050 181.480 35.310 181.800 ;
        RECT 33.210 181.140 33.470 181.460 ;
        RECT 29.990 180.460 30.250 180.780 ;
        RECT 33.210 180.460 33.470 180.780 ;
        RECT 29.530 179.440 29.790 179.760 ;
        RECT 26.770 179.100 27.030 179.420 ;
        RECT 21.710 178.080 21.970 178.400 ;
        RECT 21.770 177.040 21.910 178.080 ;
        RECT 21.710 176.720 21.970 177.040 ;
        RECT 17.110 176.380 17.370 176.700 ;
        RECT 20.790 175.360 21.050 175.680 ;
        RECT 20.850 162.330 20.990 175.360 ;
        RECT 24.530 171.260 24.670 178.420 ;
        RECT 26.370 178.340 27.430 178.480 ;
        RECT 27.290 178.060 27.430 178.340 ;
        RECT 27.230 177.740 27.490 178.060 ;
        RECT 27.290 175.680 27.430 177.740 ;
        RECT 27.230 175.360 27.490 175.680 ;
        RECT 27.500 174.485 29.040 174.855 ;
        RECT 29.070 174.000 29.330 174.320 ;
        RECT 27.230 173.660 27.490 173.980 ;
        RECT 26.310 172.640 26.570 172.960 ;
        RECT 24.470 170.940 24.730 171.260 ;
        RECT 21.250 170.600 21.510 170.920 ;
        RECT 21.310 168.880 21.450 170.600 ;
        RECT 25.850 169.580 26.110 169.900 ;
        RECT 21.250 168.560 21.510 168.880 ;
        RECT 25.910 167.860 26.050 169.580 ;
        RECT 25.850 167.540 26.110 167.860 ;
        RECT 26.370 167.180 26.510 172.640 ;
        RECT 27.290 169.810 27.430 173.660 ;
        RECT 28.610 173.320 28.870 173.640 ;
        RECT 28.150 172.980 28.410 173.300 ;
        RECT 28.210 170.920 28.350 172.980 ;
        RECT 28.670 170.920 28.810 173.320 ;
        RECT 29.130 171.600 29.270 174.000 ;
        RECT 30.050 173.300 30.190 180.460 ;
        RECT 30.800 177.205 32.340 177.575 ;
        RECT 29.990 172.980 30.250 173.300 ;
        RECT 29.530 172.300 29.790 172.620 ;
        RECT 30.450 172.300 30.710 172.620 ;
        RECT 29.590 171.680 29.730 172.300 ;
        RECT 29.070 171.280 29.330 171.600 ;
        RECT 29.590 171.540 30.190 171.680 ;
        RECT 29.530 170.940 29.790 171.260 ;
        RECT 28.150 170.600 28.410 170.920 ;
        RECT 28.610 170.600 28.870 170.920 ;
        RECT 28.210 169.900 28.350 170.600 ;
        RECT 26.830 169.670 27.430 169.810 ;
        RECT 26.830 168.540 26.970 169.670 ;
        RECT 28.150 169.580 28.410 169.900 ;
        RECT 27.500 169.045 29.040 169.415 ;
        RECT 26.770 168.280 27.030 168.540 ;
        RECT 26.770 168.220 27.430 168.280 ;
        RECT 26.830 168.140 27.430 168.220 ;
        RECT 24.010 166.860 24.270 167.180 ;
        RECT 26.310 166.860 26.570 167.180 ;
        RECT 26.770 166.860 27.030 167.180 ;
        RECT 21.250 162.330 21.510 162.420 ;
        RECT 20.850 162.190 21.510 162.330 ;
        RECT 21.250 162.100 21.510 162.190 ;
        RECT 21.310 154.940 21.450 162.100 ;
        RECT 22.170 155.980 22.430 156.300 ;
        RECT 21.250 154.620 21.510 154.940 ;
        RECT 17.570 151.220 17.830 151.540 ;
        RECT 17.630 141.000 17.770 151.220 ;
        RECT 18.950 150.880 19.210 151.200 ;
        RECT 19.010 149.840 19.150 150.880 ;
        RECT 21.310 149.840 21.450 154.620 ;
        RECT 22.230 153.580 22.370 155.980 ;
        RECT 22.170 153.260 22.430 153.580 ;
        RECT 18.950 149.520 19.210 149.840 ;
        RECT 21.250 149.520 21.510 149.840 ;
        RECT 17.570 140.680 17.830 141.000 ;
        RECT 19.870 140.000 20.130 140.320 ;
        RECT 19.930 138.960 20.070 140.000 ;
        RECT 21.310 139.980 21.450 149.520 ;
        RECT 22.630 148.160 22.890 148.480 ;
        RECT 22.690 143.720 22.830 148.160 ;
        RECT 22.630 143.400 22.890 143.720 ;
        RECT 21.710 140.340 21.970 140.660 ;
        RECT 21.250 139.660 21.510 139.980 ;
        RECT 21.310 138.960 21.450 139.660 ;
        RECT 19.870 138.640 20.130 138.960 ;
        RECT 21.250 138.640 21.510 138.960 ;
        RECT 10.670 137.115 10.930 137.260 ;
        RECT 10.660 136.745 10.940 137.115 ;
        RECT 21.770 121.960 21.910 140.340 ;
        RECT 24.070 140.320 24.210 166.860 ;
        RECT 26.830 165.560 26.970 166.860 ;
        RECT 27.290 165.820 27.430 168.140 ;
        RECT 29.590 167.860 29.730 170.940 ;
        RECT 27.690 167.540 27.950 167.860 ;
        RECT 29.530 167.540 29.790 167.860 ;
        RECT 27.750 166.160 27.890 167.540 ;
        RECT 28.150 167.200 28.410 167.520 ;
        RECT 27.690 165.840 27.950 166.160 ;
        RECT 26.370 165.480 26.970 165.560 ;
        RECT 27.230 165.500 27.490 165.820 ;
        RECT 28.210 165.480 28.350 167.200 ;
        RECT 26.310 165.420 26.970 165.480 ;
        RECT 26.310 165.160 26.570 165.420 ;
        RECT 28.150 165.160 28.410 165.480 ;
        RECT 29.590 165.140 29.730 167.540 ;
        RECT 29.530 164.820 29.790 165.140 ;
        RECT 24.470 164.140 24.730 164.460 ;
        RECT 24.930 164.140 25.190 164.460 ;
        RECT 24.530 163.440 24.670 164.140 ;
        RECT 24.470 163.120 24.730 163.440 ;
        RECT 24.990 163.100 25.130 164.140 ;
        RECT 27.500 163.605 29.040 163.975 ;
        RECT 24.930 162.780 25.190 163.100 ;
        RECT 24.990 157.320 25.130 162.780 ;
        RECT 28.150 161.420 28.410 161.740 ;
        RECT 28.210 160.380 28.350 161.420 ;
        RECT 28.150 160.060 28.410 160.380 ;
        RECT 29.590 160.120 29.730 164.820 ;
        RECT 30.050 163.440 30.190 171.540 ;
        RECT 30.510 170.830 30.650 172.300 ;
        RECT 30.800 171.765 32.340 172.135 ;
        RECT 30.910 170.830 31.170 170.920 ;
        RECT 30.510 170.690 31.170 170.830 ;
        RECT 30.910 170.600 31.170 170.690 ;
        RECT 30.450 169.580 30.710 169.900 ;
        RECT 30.510 168.200 30.650 169.580 ;
        RECT 30.450 167.880 30.710 168.200 ;
        RECT 30.510 165.560 30.650 167.880 ;
        RECT 30.800 166.325 32.340 166.695 ;
        RECT 32.290 165.840 32.550 166.160 ;
        RECT 30.510 165.420 31.110 165.560 ;
        RECT 30.450 164.480 30.710 164.800 ;
        RECT 29.990 163.120 30.250 163.440 ;
        RECT 30.510 162.840 30.650 164.480 ;
        RECT 30.050 162.700 30.650 162.840 ;
        RECT 30.050 160.720 30.190 162.700 ;
        RECT 30.970 162.420 31.110 165.420 ;
        RECT 31.370 164.140 31.630 164.460 ;
        RECT 31.430 162.420 31.570 164.140 ;
        RECT 32.350 163.100 32.490 165.840 ;
        RECT 32.750 165.160 33.010 165.480 ;
        RECT 32.290 162.780 32.550 163.100 ;
        RECT 30.910 162.100 31.170 162.420 ;
        RECT 31.370 162.100 31.630 162.420 ;
        RECT 30.450 161.760 30.710 162.080 ;
        RECT 30.510 160.720 30.650 161.760 ;
        RECT 30.800 160.885 32.340 161.255 ;
        RECT 29.990 160.400 30.250 160.720 ;
        RECT 30.450 160.400 30.710 160.720 ;
        RECT 29.590 159.980 30.190 160.120 ;
        RECT 30.050 159.700 30.190 159.980 ;
        RECT 32.290 159.720 32.550 160.040 ;
        RECT 29.990 159.380 30.250 159.700 ;
        RECT 27.500 158.165 29.040 158.535 ;
        RECT 24.930 157.000 25.190 157.320 ;
        RECT 24.990 154.940 25.130 157.000 ;
        RECT 25.850 156.660 26.110 156.980 ;
        RECT 25.910 155.280 26.050 156.660 ;
        RECT 25.850 154.960 26.110 155.280 ;
        RECT 24.930 154.620 25.190 154.940 ;
        RECT 24.990 151.880 25.130 154.620 ;
        RECT 24.930 151.560 25.190 151.880 ;
        RECT 24.470 150.540 24.730 150.860 ;
        RECT 24.530 149.500 24.670 150.540 ;
        RECT 24.990 149.840 25.130 151.560 ;
        RECT 25.910 150.860 26.050 154.960 ;
        RECT 30.050 154.940 30.190 159.380 ;
        RECT 32.350 157.320 32.490 159.720 ;
        RECT 32.290 157.000 32.550 157.320 ;
        RECT 30.450 155.980 30.710 156.300 ;
        RECT 29.990 154.620 30.250 154.940 ;
        RECT 27.500 152.725 29.040 153.095 ;
        RECT 29.990 151.560 30.250 151.880 ;
        RECT 25.390 150.540 25.650 150.860 ;
        RECT 25.850 150.540 26.110 150.860 ;
        RECT 24.930 149.520 25.190 149.840 ;
        RECT 24.470 149.180 24.730 149.500 ;
        RECT 25.450 148.480 25.590 150.540 ;
        RECT 25.390 148.160 25.650 148.480 ;
        RECT 25.910 148.140 26.050 150.540 ;
        RECT 30.050 149.840 30.190 151.560 ;
        RECT 29.990 149.520 30.250 149.840 ;
        RECT 30.510 149.750 30.650 155.980 ;
        RECT 30.800 155.445 32.340 155.815 ;
        RECT 30.800 150.005 32.340 150.375 ;
        RECT 30.510 149.610 31.110 149.750 ;
        RECT 25.850 147.820 26.110 148.140 ;
        RECT 27.500 147.285 29.040 147.655 ;
        RECT 27.690 146.460 27.950 146.780 ;
        RECT 26.310 146.120 26.570 146.440 ;
        RECT 24.930 145.100 25.190 145.420 ;
        RECT 24.470 144.080 24.730 144.400 ;
        RECT 24.010 140.000 24.270 140.320 ;
        RECT 24.070 133.520 24.210 140.000 ;
        RECT 24.530 138.620 24.670 144.080 ;
        RECT 24.990 143.040 25.130 145.100 ;
        RECT 26.370 143.800 26.510 146.120 ;
        RECT 27.750 146.100 27.890 146.460 ;
        RECT 30.050 146.100 30.190 149.520 ;
        RECT 30.970 149.160 31.110 149.610 ;
        RECT 30.450 148.840 30.710 149.160 ;
        RECT 30.910 148.840 31.170 149.160 ;
        RECT 30.510 147.120 30.650 148.840 ;
        RECT 30.450 146.800 30.710 147.120 ;
        RECT 26.770 145.780 27.030 146.100 ;
        RECT 27.690 145.780 27.950 146.100 ;
        RECT 28.150 145.780 28.410 146.100 ;
        RECT 29.990 145.780 30.250 146.100 ;
        RECT 26.830 144.400 26.970 145.780 ;
        RECT 26.770 144.080 27.030 144.400 ;
        RECT 27.750 144.060 27.890 145.780 ;
        RECT 25.910 143.720 26.510 143.800 ;
        RECT 27.690 143.740 27.950 144.060 ;
        RECT 28.210 143.720 28.350 145.780 ;
        RECT 30.450 145.100 30.710 145.420 ;
        RECT 25.850 143.660 26.510 143.720 ;
        RECT 25.850 143.400 26.110 143.660 ;
        RECT 25.390 143.060 25.650 143.380 ;
        RECT 24.930 142.720 25.190 143.040 ;
        RECT 24.470 138.300 24.730 138.620 ;
        RECT 24.990 137.600 25.130 142.720 ;
        RECT 25.450 138.280 25.590 143.060 ;
        RECT 26.370 142.700 26.510 143.660 ;
        RECT 28.150 143.400 28.410 143.720 ;
        RECT 29.530 143.060 29.790 143.380 ;
        RECT 25.850 142.380 26.110 142.700 ;
        RECT 26.310 142.380 26.570 142.700 ;
        RECT 25.390 137.960 25.650 138.280 ;
        RECT 24.930 137.280 25.190 137.600 ;
        RECT 25.910 137.260 26.050 142.380 ;
        RECT 26.370 141.680 26.510 142.380 ;
        RECT 27.500 141.845 29.040 142.215 ;
        RECT 26.310 141.360 26.570 141.680 ;
        RECT 26.770 141.020 27.030 141.340 ;
        RECT 26.830 139.980 26.970 141.020 ;
        RECT 29.590 140.660 29.730 143.060 ;
        RECT 29.990 142.380 30.250 142.700 ;
        RECT 29.530 140.340 29.790 140.660 ;
        RECT 26.770 139.660 27.030 139.980 ;
        RECT 26.830 138.620 26.970 139.660 ;
        RECT 26.770 138.300 27.030 138.620 ;
        RECT 29.590 138.280 29.730 140.340 ;
        RECT 29.530 137.960 29.790 138.280 ;
        RECT 26.770 137.620 27.030 137.940 ;
        RECT 25.850 136.940 26.110 137.260 ;
        RECT 26.830 135.640 26.970 137.620 ;
        RECT 27.500 136.405 29.040 136.775 ;
        RECT 26.830 135.500 27.430 135.640 ;
        RECT 24.010 133.200 24.270 133.520 ;
        RECT 27.290 132.240 27.430 135.500 ;
        RECT 29.590 135.220 29.730 137.960 ;
        RECT 29.530 134.900 29.790 135.220 ;
        RECT 30.050 134.960 30.190 142.380 ;
        RECT 30.510 139.980 30.650 145.100 ;
        RECT 30.800 144.565 32.340 144.935 ;
        RECT 32.810 144.060 32.950 165.160 ;
        RECT 33.270 162.760 33.410 180.460 ;
        RECT 35.110 179.760 35.250 181.480 ;
        RECT 35.050 179.440 35.310 179.760 ;
        RECT 36.030 179.420 36.170 183.860 ;
        RECT 36.430 181.140 36.690 181.460 ;
        RECT 36.490 179.760 36.630 181.140 ;
        RECT 36.430 179.440 36.690 179.760 ;
        RECT 35.970 179.100 36.230 179.420 ;
        RECT 36.950 178.740 37.090 186.920 ;
        RECT 41.090 184.520 41.230 191.340 ;
        RECT 41.550 189.620 41.690 192.700 ;
        RECT 44.310 192.680 44.450 194.060 ;
        RECT 44.770 193.360 44.910 194.060 ;
        RECT 44.710 193.040 44.970 193.360 ;
        RECT 44.700 192.760 44.980 192.875 ;
        RECT 45.230 192.760 45.370 195.760 ;
        RECT 47.010 194.740 47.270 195.060 ;
        RECT 45.630 194.060 45.890 194.380 ;
        RECT 45.690 193.020 45.830 194.060 ;
        RECT 47.070 193.360 47.210 194.740 ;
        RECT 47.530 194.720 47.670 197.800 ;
        RECT 47.930 196.780 48.190 197.100 ;
        RECT 47.470 194.400 47.730 194.720 ;
        RECT 47.010 193.040 47.270 193.360 ;
        RECT 44.250 192.360 44.510 192.680 ;
        RECT 44.700 192.620 45.370 192.760 ;
        RECT 45.630 192.700 45.890 193.020 ;
        RECT 44.700 192.505 44.980 192.620 ;
        RECT 44.710 192.360 44.970 192.505 ;
        RECT 41.490 189.300 41.750 189.620 ;
        RECT 41.490 188.620 41.750 188.940 ;
        RECT 41.550 185.200 41.690 188.620 ;
        RECT 42.870 185.960 43.130 186.220 ;
        RECT 42.470 185.900 43.130 185.960 ;
        RECT 42.470 185.820 43.070 185.900 ;
        RECT 41.490 184.880 41.750 185.200 ;
        RECT 41.030 184.200 41.290 184.520 ;
        RECT 40.110 181.480 40.370 181.800 ;
        RECT 36.890 178.420 37.150 178.740 ;
        RECT 34.130 178.080 34.390 178.400 ;
        RECT 33.670 172.640 33.930 172.960 ;
        RECT 33.730 165.140 33.870 172.640 ;
        RECT 34.190 167.860 34.330 178.080 ;
        RECT 35.970 174.000 36.230 174.320 ;
        RECT 36.030 169.900 36.170 174.000 ;
        RECT 36.950 173.640 37.090 178.420 ;
        RECT 40.170 178.400 40.310 181.480 ;
        RECT 40.570 179.100 40.830 179.420 ;
        RECT 40.110 178.080 40.370 178.400 ;
        RECT 36.890 173.320 37.150 173.640 ;
        RECT 36.950 171.260 37.090 173.320 ;
        RECT 36.890 170.940 37.150 171.260 ;
        RECT 35.970 169.580 36.230 169.900 ;
        RECT 34.130 167.540 34.390 167.860 ;
        RECT 33.670 164.820 33.930 165.140 ;
        RECT 33.670 162.780 33.930 163.100 ;
        RECT 33.210 162.440 33.470 162.760 ;
        RECT 33.210 161.760 33.470 162.080 ;
        RECT 33.270 156.980 33.410 161.760 ;
        RECT 33.210 156.660 33.470 156.980 ;
        RECT 33.210 154.960 33.470 155.280 ;
        RECT 33.270 150.860 33.410 154.960 ;
        RECT 33.210 150.540 33.470 150.860 ;
        RECT 33.210 148.840 33.470 149.160 ;
        RECT 33.270 146.780 33.410 148.840 ;
        RECT 33.730 148.820 33.870 162.780 ;
        RECT 34.190 162.080 34.330 167.540 ;
        RECT 35.510 166.920 35.770 167.180 ;
        RECT 36.030 166.920 36.170 169.580 ;
        RECT 36.950 167.860 37.090 170.940 ;
        RECT 40.630 170.920 40.770 179.100 ;
        RECT 41.090 173.210 41.230 184.200 ;
        RECT 42.470 184.180 42.610 185.820 ;
        RECT 42.410 183.860 42.670 184.180 ;
        RECT 41.950 183.520 42.210 183.840 ;
        RECT 41.490 173.210 41.750 173.300 ;
        RECT 41.090 173.070 41.750 173.210 ;
        RECT 41.490 172.980 41.750 173.070 ;
        RECT 41.030 172.300 41.290 172.620 ;
        RECT 42.010 172.360 42.150 183.520 ;
        RECT 42.470 181.800 42.610 183.860 ;
        RECT 43.790 183.180 44.050 183.500 ;
        RECT 43.850 181.800 43.990 183.180 ;
        RECT 42.410 181.480 42.670 181.800 ;
        RECT 43.790 181.480 44.050 181.800 ;
        RECT 44.310 178.740 44.450 192.360 ;
        RECT 47.530 186.560 47.670 194.400 ;
        RECT 47.990 194.380 48.130 196.780 ;
        RECT 49.830 196.080 49.970 201.200 ;
        RECT 61.330 200.500 61.470 209.310 ;
        RECT 70.990 200.500 71.130 209.310 ;
        RECT 110.010 206.150 110.150 218.060 ;
        RECT 111.010 206.600 111.150 218.690 ;
        RECT 110.920 206.340 111.240 206.600 ;
        RECT 109.920 205.890 110.240 206.150 ;
        RECT 111.420 206.120 111.560 219.040 ;
        RECT 111.330 205.860 111.650 206.120 ;
        RECT 101.480 205.335 105.480 205.405 ;
        RECT 111.810 205.335 111.950 219.350 ;
        RECT 121.210 218.215 121.530 218.275 ;
        RECT 125.435 218.215 125.805 218.285 ;
        RECT 121.210 218.075 125.805 218.215 ;
        RECT 121.210 218.015 121.530 218.075 ;
        RECT 125.435 218.005 125.805 218.075 ;
        RECT 128.010 218.215 128.330 218.275 ;
        RECT 132.235 218.215 132.605 218.285 ;
        RECT 139.035 218.275 139.405 218.285 ;
        RECT 128.010 218.075 132.605 218.215 ;
        RECT 128.010 218.015 128.330 218.075 ;
        RECT 132.235 218.005 132.605 218.075 ;
        RECT 138.890 218.015 139.405 218.275 ;
        RECT 139.035 218.005 139.405 218.015 ;
        RECT 116.450 217.755 116.770 217.815 ;
        RECT 119.850 217.755 120.170 217.815 ;
        RECT 121.550 217.755 121.870 217.815 ;
        RECT 116.450 217.615 121.870 217.755 ;
        RECT 116.450 217.555 116.770 217.615 ;
        RECT 119.850 217.555 120.170 217.615 ;
        RECT 121.550 217.555 121.870 217.615 ;
        RECT 124.610 217.755 124.930 217.815 ;
        RECT 126.650 217.755 126.970 217.815 ;
        RECT 124.610 217.615 126.970 217.755 ;
        RECT 124.610 217.555 124.930 217.615 ;
        RECT 126.650 217.555 126.970 217.615 ;
        RECT 127.330 217.755 127.650 217.815 ;
        RECT 130.050 217.755 130.370 217.815 ;
        RECT 131.750 217.755 132.070 217.815 ;
        RECT 127.330 217.615 132.070 217.755 ;
        RECT 127.330 217.555 127.650 217.615 ;
        RECT 130.050 217.555 130.370 217.615 ;
        RECT 131.750 217.555 132.070 217.615 ;
        RECT 133.110 217.755 133.430 217.815 ;
        RECT 134.470 217.755 134.790 217.815 ;
        RECT 133.110 217.615 134.790 217.755 ;
        RECT 133.110 217.555 133.430 217.615 ;
        RECT 134.470 217.555 134.790 217.615 ;
        RECT 138.890 215.915 139.210 215.975 ;
        RECT 140.250 215.915 140.570 215.975 ;
        RECT 138.890 215.775 140.570 215.915 ;
        RECT 138.890 215.715 139.210 215.775 ;
        RECT 140.250 215.715 140.570 215.775 ;
        RECT 123.930 215.455 124.250 215.515 ;
        RECT 126.310 215.455 126.630 215.515 ;
        RECT 123.930 215.315 126.630 215.455 ;
        RECT 123.930 215.255 124.250 215.315 ;
        RECT 126.310 215.255 126.630 215.315 ;
        RECT 135.490 215.455 135.810 215.515 ;
        RECT 137.530 215.455 137.850 215.515 ;
        RECT 135.490 215.315 137.850 215.455 ;
        RECT 135.490 215.255 135.810 215.315 ;
        RECT 137.530 215.255 137.850 215.315 ;
        RECT 117.130 214.995 117.450 215.055 ;
        RECT 118.490 214.995 118.810 215.055 ;
        RECT 117.130 214.855 118.810 214.995 ;
        RECT 117.130 214.795 117.450 214.855 ;
        RECT 118.490 214.795 118.810 214.855 ;
        RECT 144.330 213.615 144.650 213.675 ;
        RECT 146.030 213.615 146.350 213.675 ;
        RECT 144.330 213.475 146.350 213.615 ;
        RECT 144.330 213.415 144.650 213.475 ;
        RECT 146.030 213.415 146.350 213.475 ;
        RECT 117.130 213.155 117.450 213.215 ;
        RECT 120.870 213.155 121.190 213.215 ;
        RECT 117.130 213.015 121.190 213.155 ;
        RECT 117.130 212.955 117.450 213.015 ;
        RECT 120.870 212.955 121.190 213.015 ;
        RECT 130.730 213.155 131.050 213.215 ;
        RECT 134.470 213.155 134.790 213.215 ;
        RECT 130.730 213.015 134.790 213.155 ;
        RECT 130.730 212.955 131.050 213.015 ;
        RECT 134.470 212.955 134.790 213.015 ;
        RECT 117.130 212.695 117.450 212.755 ;
        RECT 121.210 212.695 121.530 212.755 ;
        RECT 126.990 212.695 127.310 212.755 ;
        RECT 117.130 212.555 127.310 212.695 ;
        RECT 117.130 212.495 117.450 212.555 ;
        RECT 121.210 212.495 121.530 212.555 ;
        RECT 126.990 212.495 127.310 212.555 ;
        RECT 128.010 212.695 128.330 212.755 ;
        RECT 129.030 212.695 129.350 212.755 ;
        RECT 128.010 212.555 129.350 212.695 ;
        RECT 128.010 212.495 128.330 212.555 ;
        RECT 129.030 212.495 129.350 212.555 ;
        RECT 126.990 212.235 127.310 212.295 ;
        RECT 134.810 212.235 135.130 212.295 ;
        RECT 137.870 212.235 138.190 212.295 ;
        RECT 126.990 212.095 138.190 212.235 ;
        RECT 126.990 212.035 127.310 212.095 ;
        RECT 134.810 212.035 135.130 212.095 ;
        RECT 137.870 212.035 138.190 212.095 ;
        RECT 119.170 210.855 119.490 210.915 ;
        RECT 124.270 210.855 124.590 210.915 ;
        RECT 119.170 210.715 124.590 210.855 ;
        RECT 119.170 210.655 119.490 210.715 ;
        RECT 124.270 210.655 124.590 210.715 ;
        RECT 132.770 210.855 133.090 210.915 ;
        RECT 135.150 210.855 135.470 210.915 ;
        RECT 132.770 210.715 135.470 210.855 ;
        RECT 132.770 210.655 133.090 210.715 ;
        RECT 135.150 210.655 135.470 210.715 ;
        RECT 138.210 210.855 138.530 210.915 ;
        RECT 139.910 210.855 140.230 210.915 ;
        RECT 138.210 210.715 140.230 210.855 ;
        RECT 138.210 210.655 138.530 210.715 ;
        RECT 139.910 210.655 140.230 210.715 ;
        RECT 117.130 210.395 117.450 210.455 ;
        RECT 121.550 210.395 121.870 210.455 ;
        RECT 117.130 210.255 121.870 210.395 ;
        RECT 117.130 210.195 117.450 210.255 ;
        RECT 121.550 210.195 121.870 210.255 ;
        RECT 138.890 210.395 139.210 210.455 ;
        RECT 139.910 210.395 140.230 210.455 ;
        RECT 138.890 210.255 140.230 210.395 ;
        RECT 138.890 210.195 139.210 210.255 ;
        RECT 139.910 210.195 140.230 210.255 ;
        RECT 121.890 209.935 122.210 209.995 ;
        RECT 125.290 209.935 125.610 209.995 ;
        RECT 129.710 209.935 130.030 209.995 ;
        RECT 121.890 209.795 130.030 209.935 ;
        RECT 121.890 209.735 122.210 209.795 ;
        RECT 125.290 209.735 125.610 209.795 ;
        RECT 129.710 209.735 130.030 209.795 ;
        RECT 144.330 209.015 144.650 209.075 ;
        RECT 146.030 209.015 146.350 209.075 ;
        RECT 144.330 208.875 146.350 209.015 ;
        RECT 144.330 208.815 144.650 208.875 ;
        RECT 146.030 208.815 146.350 208.875 ;
        RECT 143.795 208.555 144.165 208.625 ;
        RECT 146.030 208.555 146.350 208.615 ;
        RECT 143.795 208.415 146.350 208.555 ;
        RECT 143.795 208.345 144.165 208.415 ;
        RECT 146.030 208.355 146.350 208.415 ;
        RECT 113.390 208.095 113.710 208.155 ;
        RECT 117.130 208.095 117.450 208.155 ;
        RECT 113.390 207.955 117.450 208.095 ;
        RECT 113.390 207.895 113.710 207.955 ;
        RECT 117.130 207.895 117.450 207.955 ;
        RECT 135.150 208.095 135.470 208.155 ;
        RECT 138.890 208.095 139.210 208.155 ;
        RECT 140.590 208.095 140.910 208.155 ;
        RECT 142.630 208.095 142.950 208.155 ;
        RECT 135.150 207.955 142.950 208.095 ;
        RECT 135.150 207.895 135.470 207.955 ;
        RECT 138.890 207.895 139.210 207.955 ;
        RECT 140.590 207.895 140.910 207.955 ;
        RECT 142.630 207.895 142.950 207.955 ;
        RECT 133.110 207.175 133.430 207.235 ;
        RECT 142.435 207.175 142.805 207.245 ;
        RECT 133.110 207.035 142.805 207.175 ;
        RECT 133.110 206.975 133.430 207.035 ;
        RECT 142.435 206.965 142.805 207.035 ;
        RECT 143.990 206.715 144.310 206.775 ;
        RECT 145.350 206.715 145.670 206.775 ;
        RECT 143.990 206.575 145.670 206.715 ;
        RECT 143.990 206.515 144.310 206.575 ;
        RECT 145.350 206.515 145.670 206.575 ;
        RECT 116.110 206.255 116.430 206.315 ;
        RECT 121.550 206.255 121.870 206.315 ;
        RECT 127.670 206.255 127.990 206.315 ;
        RECT 116.110 206.115 127.990 206.255 ;
        RECT 116.110 206.055 116.430 206.115 ;
        RECT 121.550 206.055 121.870 206.115 ;
        RECT 127.670 206.055 127.990 206.115 ;
        RECT 135.490 205.795 135.810 205.855 ;
        RECT 138.890 205.795 139.210 205.855 ;
        RECT 135.490 205.655 139.210 205.795 ;
        RECT 135.490 205.595 135.810 205.655 ;
        RECT 138.890 205.595 139.210 205.655 ;
        RECT 141.610 205.795 141.930 205.855 ;
        RECT 143.650 205.795 143.970 205.855 ;
        RECT 141.610 205.655 143.970 205.795 ;
        RECT 141.610 205.595 141.930 205.655 ;
        RECT 143.650 205.595 143.970 205.655 ;
        RECT 112.710 205.335 113.030 205.395 ;
        RECT 101.480 205.195 113.030 205.335 ;
        RECT 101.480 205.125 105.480 205.195 ;
        RECT 112.710 205.135 113.030 205.195 ;
        RECT 147.050 205.335 147.370 205.395 ;
        RECT 149.680 205.335 150.000 205.430 ;
        RECT 155.245 205.335 159.245 205.405 ;
        RECT 147.050 205.195 159.245 205.335 ;
        RECT 147.050 205.135 147.370 205.195 ;
        RECT 149.680 205.100 150.000 205.195 ;
        RECT 155.245 205.125 159.245 205.195 ;
        RECT 123.930 204.875 124.250 204.935 ;
        RECT 126.650 204.875 126.970 204.935 ;
        RECT 123.930 204.735 126.970 204.875 ;
        RECT 123.930 204.675 124.250 204.735 ;
        RECT 126.650 204.675 126.970 204.735 ;
        RECT 127.670 204.875 127.990 204.935 ;
        RECT 130.730 204.875 131.050 204.935 ;
        RECT 136.170 204.875 136.490 204.935 ;
        RECT 138.890 204.875 139.210 204.935 ;
        RECT 127.670 204.735 139.210 204.875 ;
        RECT 127.670 204.675 127.990 204.735 ;
        RECT 130.730 204.675 131.050 204.735 ;
        RECT 136.170 204.675 136.490 204.735 ;
        RECT 138.890 204.675 139.210 204.735 ;
        RECT 128.010 204.415 128.330 204.475 ;
        RECT 129.710 204.415 130.030 204.475 ;
        RECT 128.010 204.275 130.030 204.415 ;
        RECT 128.010 204.215 128.330 204.275 ;
        RECT 129.710 204.215 130.030 204.275 ;
        RECT 130.730 204.415 131.050 204.475 ;
        RECT 143.795 204.415 144.165 204.485 ;
        RECT 130.730 204.275 144.165 204.415 ;
        RECT 130.730 204.215 131.050 204.275 ;
        RECT 143.795 204.205 144.165 204.275 ;
        RECT 113.390 202.835 113.710 203.095 ;
        RECT 111.360 202.575 111.620 202.665 ;
        RECT 112.710 202.575 113.030 202.635 ;
        RECT 107.190 202.435 113.030 202.575 ;
        RECT 101.480 202.115 105.480 202.185 ;
        RECT 107.190 202.115 107.330 202.435 ;
        RECT 111.360 202.345 111.620 202.435 ;
        RECT 112.710 202.375 113.030 202.435 ;
        RECT 101.480 201.975 107.330 202.115 ;
        RECT 101.480 201.905 105.480 201.975 ;
        RECT 113.480 201.655 113.620 202.835 ;
        RECT 114.895 202.205 115.265 203.745 ;
        RECT 120.335 202.205 120.705 203.745 ;
        RECT 125.775 202.205 126.145 203.745 ;
        RECT 131.215 202.205 131.585 203.745 ;
        RECT 136.655 202.205 137.025 203.745 ;
        RECT 142.095 202.205 142.465 203.745 ;
        RECT 147.535 202.205 147.905 203.745 ;
        RECT 155.245 202.115 159.245 202.185 ;
        RECT 148.670 201.975 159.245 202.115 ;
        RECT 117.130 201.655 117.450 201.715 ;
        RECT 120.870 201.655 121.190 201.715 ;
        RECT 113.480 201.515 116.850 201.655 ;
        RECT 116.710 200.795 116.850 201.515 ;
        RECT 117.130 201.515 121.190 201.655 ;
        RECT 117.130 201.455 117.450 201.515 ;
        RECT 120.870 201.455 121.190 201.515 ;
        RECT 129.710 201.655 130.030 201.715 ;
        RECT 139.910 201.655 140.230 201.715 ;
        RECT 129.710 201.515 140.230 201.655 ;
        RECT 129.710 201.455 130.030 201.515 ;
        RECT 139.910 201.455 140.230 201.515 ;
        RECT 140.590 201.655 140.910 201.715 ;
        RECT 145.350 201.655 145.670 201.715 ;
        RECT 140.590 201.515 145.670 201.655 ;
        RECT 140.590 201.455 140.910 201.515 ;
        RECT 145.350 201.455 145.670 201.515 ;
        RECT 118.830 201.195 119.150 201.255 ;
        RECT 131.750 201.195 132.070 201.255 ;
        RECT 138.210 201.195 138.530 201.255 ;
        RECT 118.830 201.055 138.530 201.195 ;
        RECT 118.830 200.995 119.150 201.055 ;
        RECT 131.750 200.995 132.070 201.055 ;
        RECT 138.210 200.995 138.530 201.055 ;
        RECT 138.890 201.195 139.210 201.255 ;
        RECT 140.590 201.195 140.910 201.255 ;
        RECT 138.890 201.055 140.910 201.195 ;
        RECT 138.890 200.995 139.210 201.055 ;
        RECT 140.590 200.995 140.910 201.055 ;
        RECT 142.970 201.195 143.290 201.255 ;
        RECT 148.110 201.195 148.440 201.290 ;
        RECT 148.670 201.195 148.810 201.975 ;
        RECT 155.245 201.905 159.245 201.975 ;
        RECT 142.970 201.055 148.810 201.195 ;
        RECT 142.970 200.995 143.290 201.055 ;
        RECT 148.110 200.960 148.440 201.055 ;
        RECT 113.050 200.735 113.370 200.795 ;
        RECT 115.430 200.735 115.750 200.795 ;
        RECT 113.050 200.595 115.750 200.735 ;
        RECT 116.710 200.735 117.110 200.795 ;
        RECT 119.850 200.735 120.170 200.795 ;
        RECT 121.890 200.735 122.210 200.795 ;
        RECT 123.590 200.735 123.910 200.795 ;
        RECT 116.710 200.595 123.910 200.735 ;
        RECT 113.050 200.535 113.370 200.595 ;
        RECT 115.430 200.535 115.750 200.595 ;
        RECT 116.790 200.535 117.110 200.595 ;
        RECT 119.850 200.535 120.170 200.595 ;
        RECT 121.890 200.535 122.210 200.595 ;
        RECT 123.590 200.535 123.910 200.595 ;
        RECT 129.710 200.735 130.030 200.795 ;
        RECT 132.430 200.735 132.750 200.795 ;
        RECT 137.190 200.735 137.510 200.795 ;
        RECT 129.710 200.595 132.750 200.735 ;
        RECT 129.710 200.535 130.030 200.595 ;
        RECT 132.430 200.535 132.750 200.595 ;
        RECT 133.030 200.595 137.510 200.735 ;
        RECT 61.270 200.180 61.530 200.500 ;
        RECT 70.930 200.180 71.190 200.500 ;
        RECT 56.670 199.500 56.930 199.820 ;
        RECT 60.350 199.500 60.610 199.820 ;
        RECT 63.110 199.500 63.370 199.820 ;
        RECT 69.550 199.500 69.810 199.820 ;
        RECT 56.730 198.800 56.870 199.500 ;
        RECT 56.670 198.480 56.930 198.800 ;
        RECT 55.290 197.460 55.550 197.780 ;
        RECT 49.770 195.760 50.030 196.080 ;
        RECT 48.850 194.740 49.110 195.060 ;
        RECT 47.930 194.060 48.190 194.380 ;
        RECT 47.990 192.000 48.130 194.060 ;
        RECT 47.930 191.680 48.190 192.000 ;
        RECT 46.090 186.240 46.350 186.560 ;
        RECT 47.470 186.240 47.730 186.560 ;
        RECT 45.630 180.800 45.890 181.120 ;
        RECT 45.690 178.740 45.830 180.800 ;
        RECT 44.250 178.420 44.510 178.740 ;
        RECT 45.630 178.420 45.890 178.740 ;
        RECT 43.790 176.040 44.050 176.360 ;
        RECT 42.870 175.360 43.130 175.680 ;
        RECT 42.410 175.020 42.670 175.340 ;
        RECT 42.470 172.960 42.610 175.020 ;
        RECT 42.930 174.320 43.070 175.360 ;
        RECT 42.870 174.000 43.130 174.320 ;
        RECT 43.330 173.660 43.590 173.980 ;
        RECT 43.390 172.960 43.530 173.660 ;
        RECT 42.410 172.640 42.670 172.960 ;
        RECT 43.330 172.640 43.590 172.960 ;
        RECT 40.570 170.600 40.830 170.920 ;
        RECT 40.630 168.880 40.770 170.600 ;
        RECT 40.570 168.560 40.830 168.880 ;
        RECT 41.090 167.860 41.230 172.300 ;
        RECT 41.550 172.220 42.150 172.360 ;
        RECT 36.890 167.540 37.150 167.860 ;
        RECT 38.730 167.540 38.990 167.860 ;
        RECT 41.030 167.540 41.290 167.860 ;
        RECT 35.510 166.860 36.170 166.920 ;
        RECT 37.810 166.860 38.070 167.180 ;
        RECT 35.570 166.780 36.170 166.860 ;
        RECT 36.030 165.480 36.170 166.780 ;
        RECT 37.870 165.820 38.010 166.860 ;
        RECT 37.810 165.500 38.070 165.820 ;
        RECT 35.970 165.160 36.230 165.480 ;
        RECT 36.030 163.440 36.170 165.160 ;
        RECT 36.430 164.820 36.690 165.140 ;
        RECT 35.970 163.120 36.230 163.440 ;
        RECT 36.030 162.760 36.170 163.120 ;
        RECT 35.970 162.440 36.230 162.760 ;
        RECT 36.490 162.420 36.630 164.820 ;
        RECT 37.350 162.780 37.610 163.100 ;
        RECT 36.430 162.100 36.690 162.420 ;
        RECT 34.190 161.940 34.790 162.080 ;
        RECT 34.650 159.700 34.790 161.940 ;
        RECT 37.410 160.040 37.550 162.780 ;
        RECT 37.870 162.420 38.010 165.500 ;
        RECT 37.810 162.100 38.070 162.420 ;
        RECT 37.350 159.720 37.610 160.040 ;
        RECT 34.590 159.380 34.850 159.700 ;
        RECT 34.130 158.700 34.390 159.020 ;
        RECT 34.190 155.280 34.330 158.700 ;
        RECT 34.130 154.960 34.390 155.280 ;
        RECT 34.650 153.920 34.790 159.380 ;
        RECT 37.870 156.720 38.010 162.100 ;
        RECT 38.790 160.040 38.930 167.540 ;
        RECT 41.550 167.520 41.690 172.220 ;
        RECT 43.390 167.860 43.530 172.640 ;
        RECT 43.850 172.620 43.990 176.040 ;
        RECT 45.690 174.320 45.830 178.420 ;
        RECT 45.630 174.000 45.890 174.320 ;
        RECT 45.690 173.210 45.830 174.000 ;
        RECT 46.150 173.980 46.290 186.240 ;
        RECT 47.470 183.180 47.730 183.500 ;
        RECT 46.550 181.140 46.810 181.460 ;
        RECT 46.610 179.760 46.750 181.140 ;
        RECT 47.530 180.780 47.670 183.180 ;
        RECT 47.010 180.460 47.270 180.780 ;
        RECT 47.470 180.460 47.730 180.780 ;
        RECT 46.550 179.440 46.810 179.760 ;
        RECT 47.070 179.080 47.210 180.460 ;
        RECT 47.010 178.760 47.270 179.080 ;
        RECT 46.090 173.660 46.350 173.980 ;
        RECT 46.550 173.210 46.810 173.300 ;
        RECT 45.690 173.070 46.810 173.210 ;
        RECT 46.550 172.980 46.810 173.070 ;
        RECT 43.790 172.300 44.050 172.620 ;
        RECT 43.330 167.540 43.590 167.860 ;
        RECT 43.850 167.520 43.990 172.300 ;
        RECT 44.710 169.920 44.970 170.240 ;
        RECT 41.490 167.200 41.750 167.520 ;
        RECT 43.790 167.200 44.050 167.520 ;
        RECT 41.550 163.440 41.690 167.200 ;
        RECT 44.770 166.160 44.910 169.920 ;
        RECT 46.610 168.880 46.750 172.980 ;
        RECT 47.070 172.620 47.210 178.760 ;
        RECT 47.990 178.400 48.130 191.680 ;
        RECT 48.390 179.440 48.650 179.760 ;
        RECT 47.930 178.080 48.190 178.400 ;
        RECT 48.450 177.040 48.590 179.440 ;
        RECT 48.390 176.720 48.650 177.040 ;
        RECT 47.470 176.040 47.730 176.360 ;
        RECT 47.530 174.320 47.670 176.040 ;
        RECT 47.470 174.000 47.730 174.320 ;
        RECT 47.010 172.300 47.270 172.620 ;
        RECT 48.910 170.920 49.050 194.740 ;
        RECT 49.310 194.060 49.570 194.380 ;
        RECT 49.370 192.340 49.510 194.060 ;
        RECT 49.310 192.020 49.570 192.340 ;
        RECT 49.830 190.640 49.970 195.760 ;
        RECT 55.350 195.060 55.490 197.460 ;
        RECT 60.410 196.080 60.550 199.500 ;
        RECT 61.730 196.780 61.990 197.100 ;
        RECT 60.350 195.760 60.610 196.080 ;
        RECT 61.790 195.060 61.930 196.780 ;
        RECT 55.290 194.740 55.550 195.060 ;
        RECT 59.430 194.740 59.690 195.060 ;
        RECT 61.730 194.740 61.990 195.060 ;
        RECT 58.050 194.060 58.310 194.380 ;
        RECT 58.110 193.360 58.250 194.060 ;
        RECT 59.490 193.360 59.630 194.740 ;
        RECT 50.230 193.040 50.490 193.360 ;
        RECT 56.210 193.040 56.470 193.360 ;
        RECT 58.050 193.040 58.310 193.360 ;
        RECT 59.430 193.040 59.690 193.360 ;
        RECT 50.290 192.875 50.430 193.040 ;
        RECT 50.220 192.505 50.500 192.875 ;
        RECT 50.230 192.360 50.490 192.505 ;
        RECT 49.770 190.320 50.030 190.640 ;
        RECT 49.310 183.520 49.570 183.840 ;
        RECT 49.370 182.480 49.510 183.520 ;
        RECT 49.310 182.160 49.570 182.480 ;
        RECT 49.830 175.680 49.970 190.320 ;
        RECT 56.270 189.620 56.410 193.040 ;
        RECT 61.790 192.680 61.930 194.740 ;
        RECT 61.730 192.360 61.990 192.680 ;
        RECT 60.810 191.340 61.070 191.660 ;
        RECT 60.870 190.300 61.010 191.340 ;
        RECT 59.430 189.980 59.690 190.300 ;
        RECT 60.810 189.980 61.070 190.300 ;
        RECT 55.750 189.300 56.010 189.620 ;
        RECT 56.210 189.300 56.470 189.620 ;
        RECT 51.610 187.260 51.870 187.580 ;
        RECT 51.670 183.500 51.810 187.260 ;
        RECT 55.810 186.900 55.950 189.300 ;
        RECT 56.270 187.920 56.410 189.300 ;
        RECT 56.670 188.620 56.930 188.940 ;
        RECT 56.210 187.600 56.470 187.920 ;
        RECT 56.730 187.240 56.870 188.620 ;
        RECT 56.670 186.920 56.930 187.240 ;
        RECT 58.510 186.920 58.770 187.240 ;
        RECT 55.750 186.580 56.010 186.900 ;
        RECT 56.730 185.200 56.870 186.920 ;
        RECT 57.590 186.580 57.850 186.900 ;
        RECT 56.670 184.880 56.930 185.200 ;
        RECT 52.070 183.860 52.330 184.180 ;
        RECT 56.210 183.860 56.470 184.180 ;
        RECT 51.610 183.180 51.870 183.500 ;
        RECT 51.150 181.140 51.410 181.460 ;
        RECT 51.210 179.760 51.350 181.140 ;
        RECT 51.150 179.440 51.410 179.760 ;
        RECT 49.770 175.360 50.030 175.680 ;
        RECT 51.670 175.340 51.810 183.180 ;
        RECT 52.130 182.480 52.270 183.860 ;
        RECT 56.270 182.480 56.410 183.860 ;
        RECT 57.650 182.480 57.790 186.580 ;
        RECT 52.070 182.160 52.330 182.480 ;
        RECT 56.210 182.160 56.470 182.480 ;
        RECT 57.590 182.160 57.850 182.480 ;
        RECT 58.050 181.820 58.310 182.140 ;
        RECT 53.910 181.480 54.170 181.800 ;
        RECT 56.210 181.480 56.470 181.800 ;
        RECT 57.590 181.480 57.850 181.800 ;
        RECT 52.990 179.100 53.250 179.420 ;
        RECT 52.530 175.360 52.790 175.680 ;
        RECT 51.610 175.020 51.870 175.340 ;
        RECT 51.670 173.300 51.810 175.020 ;
        RECT 51.610 172.980 51.870 173.300 ;
        RECT 52.590 172.960 52.730 175.360 ;
        RECT 52.530 172.640 52.790 172.960 ;
        RECT 47.930 170.600 48.190 170.920 ;
        RECT 48.850 170.600 49.110 170.920 ;
        RECT 49.770 170.600 50.030 170.920 ;
        RECT 46.550 168.560 46.810 168.880 ;
        RECT 47.990 168.540 48.130 170.600 ;
        RECT 49.830 168.880 49.970 170.600 ;
        RECT 50.230 169.580 50.490 169.900 ;
        RECT 49.770 168.560 50.030 168.880 ;
        RECT 47.930 168.220 48.190 168.540 ;
        RECT 50.290 167.860 50.430 169.580 ;
        RECT 47.930 167.600 48.190 167.860 ;
        RECT 47.930 167.540 49.510 167.600 ;
        RECT 50.230 167.540 50.490 167.860 ;
        RECT 51.610 167.600 51.870 167.860 ;
        RECT 52.590 167.600 52.730 172.640 ;
        RECT 53.050 168.880 53.190 179.100 ;
        RECT 53.970 178.740 54.110 181.480 ;
        RECT 54.830 181.140 55.090 181.460 ;
        RECT 55.290 181.140 55.550 181.460 ;
        RECT 54.890 178.740 55.030 181.140 ;
        RECT 55.350 179.760 55.490 181.140 ;
        RECT 55.750 180.460 56.010 180.780 ;
        RECT 55.290 179.440 55.550 179.760 ;
        RECT 55.810 179.160 55.950 180.460 ;
        RECT 56.270 179.760 56.410 181.480 ;
        RECT 57.650 179.760 57.790 181.480 ;
        RECT 56.210 179.440 56.470 179.760 ;
        RECT 57.590 179.440 57.850 179.760 ;
        RECT 55.810 179.080 56.410 179.160 ;
        RECT 55.810 179.020 56.470 179.080 ;
        RECT 53.910 178.420 54.170 178.740 ;
        RECT 54.830 178.420 55.090 178.740 ;
        RECT 53.970 169.900 54.110 178.420 ;
        RECT 55.810 173.300 55.950 179.020 ;
        RECT 56.210 178.760 56.470 179.020 ;
        RECT 58.110 178.400 58.250 181.820 ;
        RECT 58.570 179.420 58.710 186.920 ;
        RECT 58.970 185.900 59.230 186.220 ;
        RECT 59.030 181.800 59.170 185.900 ;
        RECT 59.490 184.180 59.630 189.980 ;
        RECT 60.350 189.530 60.610 189.620 ;
        RECT 60.870 189.530 61.010 189.980 ;
        RECT 61.790 189.620 61.930 192.360 ;
        RECT 62.650 192.020 62.910 192.340 ;
        RECT 62.190 191.340 62.450 191.660 ;
        RECT 60.350 189.390 61.010 189.530 ;
        RECT 60.350 189.300 60.610 189.390 ;
        RECT 60.350 185.900 60.610 186.220 ;
        RECT 60.410 184.860 60.550 185.900 ;
        RECT 60.350 184.540 60.610 184.860 ;
        RECT 59.430 184.035 59.690 184.180 ;
        RECT 59.420 183.665 59.700 184.035 ;
        RECT 59.430 183.180 59.690 183.500 ;
        RECT 59.490 181.800 59.630 183.180 ;
        RECT 58.970 181.480 59.230 181.800 ;
        RECT 59.430 181.480 59.690 181.800 ;
        RECT 60.410 179.420 60.550 184.540 ;
        RECT 60.870 181.120 61.010 189.390 ;
        RECT 61.730 189.300 61.990 189.620 ;
        RECT 62.250 187.580 62.390 191.340 ;
        RECT 62.710 189.620 62.850 192.020 ;
        RECT 62.650 189.300 62.910 189.620 ;
        RECT 62.710 188.940 62.850 189.300 ;
        RECT 62.650 188.620 62.910 188.940 ;
        RECT 62.190 187.260 62.450 187.580 ;
        RECT 62.710 187.240 62.850 188.620 ;
        RECT 62.650 186.920 62.910 187.240 ;
        RECT 63.170 184.600 63.310 199.500 ;
        RECT 66.790 196.780 67.050 197.100 ;
        RECT 64.030 194.740 64.290 195.060 ;
        RECT 64.090 190.640 64.230 194.740 ;
        RECT 65.870 194.400 66.130 194.720 ;
        RECT 64.950 191.680 65.210 192.000 ;
        RECT 65.010 190.640 65.150 191.680 ;
        RECT 65.930 191.660 66.070 194.400 ;
        RECT 66.850 192.680 66.990 196.780 ;
        RECT 67.250 195.990 67.510 196.080 ;
        RECT 67.250 195.850 67.910 195.990 ;
        RECT 67.250 195.760 67.510 195.850 ;
        RECT 67.250 194.740 67.510 195.060 ;
        RECT 66.790 192.360 67.050 192.680 ;
        RECT 65.870 191.340 66.130 191.660 ;
        RECT 64.030 190.320 64.290 190.640 ;
        RECT 64.950 190.320 65.210 190.640 ;
        RECT 65.010 189.960 65.150 190.320 ;
        RECT 64.950 189.640 65.210 189.960 ;
        RECT 65.010 186.900 65.150 189.640 ;
        RECT 66.850 189.280 66.990 192.360 ;
        RECT 67.310 192.000 67.450 194.740 ;
        RECT 67.770 193.360 67.910 195.850 ;
        RECT 68.170 194.060 68.430 194.380 ;
        RECT 67.710 193.040 67.970 193.360 ;
        RECT 67.250 191.680 67.510 192.000 ;
        RECT 66.790 188.960 67.050 189.280 ;
        RECT 64.950 186.580 65.210 186.900 ;
        RECT 67.250 186.240 67.510 186.560 ;
        RECT 67.310 185.200 67.450 186.240 ;
        RECT 63.570 184.880 63.830 185.200 ;
        RECT 67.250 184.880 67.510 185.200 ;
        RECT 62.710 184.460 63.310 184.600 ;
        RECT 63.630 184.520 63.770 184.880 ;
        RECT 66.790 184.540 67.050 184.860 ;
        RECT 62.190 184.035 62.450 184.180 ;
        RECT 62.180 183.665 62.460 184.035 ;
        RECT 61.730 183.180 61.990 183.500 ;
        RECT 61.790 182.140 61.930 183.180 ;
        RECT 61.730 181.820 61.990 182.140 ;
        RECT 61.270 181.370 61.530 181.460 ;
        RECT 62.710 181.370 62.850 184.460 ;
        RECT 63.570 184.200 63.830 184.520 ;
        RECT 64.030 183.860 64.290 184.180 ;
        RECT 63.110 183.520 63.370 183.840 ;
        RECT 61.270 181.230 62.850 181.370 ;
        RECT 61.270 181.140 61.530 181.230 ;
        RECT 60.810 180.800 61.070 181.120 ;
        RECT 58.510 179.100 58.770 179.420 ;
        RECT 60.350 179.100 60.610 179.420 ;
        RECT 58.970 178.420 59.230 178.740 ;
        RECT 60.870 178.480 61.010 180.800 ;
        RECT 57.590 178.080 57.850 178.400 ;
        RECT 58.050 178.080 58.310 178.400 ;
        RECT 58.510 178.080 58.770 178.400 ;
        RECT 56.670 173.320 56.930 173.640 ;
        RECT 55.750 172.980 56.010 173.300 ;
        RECT 56.210 172.980 56.470 173.300 ;
        RECT 56.270 171.600 56.410 172.980 ;
        RECT 56.210 171.280 56.470 171.600 ;
        RECT 56.210 170.600 56.470 170.920 ;
        RECT 53.910 169.580 54.170 169.900 ;
        RECT 52.990 168.560 53.250 168.880 ;
        RECT 55.750 168.560 56.010 168.880 ;
        RECT 53.450 168.220 53.710 168.540 ;
        RECT 51.610 167.540 52.730 167.600 ;
        RECT 47.990 167.520 49.510 167.540 ;
        RECT 47.990 167.460 49.570 167.520 ;
        RECT 51.670 167.460 52.730 167.540 ;
        RECT 49.310 167.200 49.570 167.460 ;
        RECT 52.590 167.180 52.730 167.460 ;
        RECT 52.070 166.860 52.330 167.180 ;
        RECT 52.530 166.860 52.790 167.180 ;
        RECT 44.710 165.840 44.970 166.160 ;
        RECT 41.490 163.120 41.750 163.440 ;
        RECT 41.490 162.440 41.750 162.760 ;
        RECT 41.030 162.100 41.290 162.420 ;
        RECT 40.570 161.760 40.830 162.080 ;
        RECT 39.190 161.420 39.450 161.740 ;
        RECT 38.270 159.720 38.530 160.040 ;
        RECT 38.730 159.720 38.990 160.040 ;
        RECT 37.410 156.580 38.010 156.720 ;
        RECT 34.590 153.600 34.850 153.920 ;
        RECT 35.510 151.560 35.770 151.880 ;
        RECT 34.130 150.540 34.390 150.860 ;
        RECT 34.190 149.500 34.330 150.540 ;
        RECT 34.130 149.180 34.390 149.500 ;
        RECT 33.670 148.500 33.930 148.820 ;
        RECT 35.570 147.120 35.710 151.560 ;
        RECT 37.410 151.540 37.550 156.580 ;
        RECT 38.330 154.940 38.470 159.720 ;
        RECT 39.250 157.320 39.390 161.420 ;
        RECT 40.630 160.380 40.770 161.760 ;
        RECT 41.090 160.380 41.230 162.100 ;
        RECT 41.550 160.720 41.690 162.440 ;
        RECT 48.850 162.100 49.110 162.420 ;
        RECT 46.090 161.420 46.350 161.740 ;
        RECT 47.010 161.420 47.270 161.740 ;
        RECT 41.490 160.400 41.750 160.720 ;
        RECT 40.570 160.060 40.830 160.380 ;
        RECT 41.030 160.060 41.290 160.380 ;
        RECT 40.110 159.720 40.370 160.040 ;
        RECT 40.170 158.000 40.310 159.720 ;
        RECT 40.110 157.680 40.370 158.000 ;
        RECT 39.190 157.000 39.450 157.320 ;
        RECT 38.270 154.620 38.530 154.940 ;
        RECT 37.810 153.600 38.070 153.920 ;
        RECT 37.870 151.540 38.010 153.600 ;
        RECT 38.330 151.540 38.470 154.620 ;
        RECT 40.630 151.540 40.770 160.060 ;
        RECT 46.150 156.300 46.290 161.420 ;
        RECT 46.550 156.890 46.810 156.980 ;
        RECT 47.070 156.890 47.210 161.420 ;
        RECT 48.910 160.720 49.050 162.100 ;
        RECT 52.130 162.080 52.270 166.860 ;
        RECT 52.990 162.100 53.250 162.420 ;
        RECT 52.130 161.940 52.730 162.080 ;
        RECT 52.070 161.420 52.330 161.740 ;
        RECT 48.850 160.400 49.110 160.720 ;
        RECT 47.470 159.720 47.730 160.040 ;
        RECT 47.530 158.000 47.670 159.720 ;
        RECT 47.470 157.680 47.730 158.000 ;
        RECT 46.550 156.750 47.210 156.890 ;
        RECT 46.550 156.660 46.810 156.750 ;
        RECT 48.390 156.320 48.650 156.640 ;
        RECT 41.490 155.980 41.750 156.300 ;
        RECT 46.090 155.980 46.350 156.300 ;
        RECT 41.550 152.640 41.690 155.980 ;
        RECT 47.930 154.280 48.190 154.600 ;
        RECT 41.090 152.500 41.690 152.640 ;
        RECT 37.350 151.220 37.610 151.540 ;
        RECT 37.810 151.220 38.070 151.540 ;
        RECT 38.270 151.220 38.530 151.540 ;
        RECT 40.570 151.220 40.830 151.540 ;
        RECT 38.330 149.840 38.470 151.220 ;
        RECT 38.270 149.520 38.530 149.840 ;
        RECT 40.110 148.160 40.370 148.480 ;
        RECT 35.510 146.800 35.770 147.120 ;
        RECT 33.210 146.460 33.470 146.780 ;
        RECT 37.810 145.100 38.070 145.420 ;
        RECT 37.870 144.060 38.010 145.100 ;
        RECT 32.750 143.800 33.010 144.060 ;
        RECT 32.750 143.740 34.330 143.800 ;
        RECT 37.810 143.740 38.070 144.060 ;
        RECT 32.810 143.660 34.330 143.740 ;
        RECT 40.170 143.720 40.310 148.160 ;
        RECT 41.090 146.440 41.230 152.500 ;
        RECT 41.490 151.560 41.750 151.880 ;
        RECT 41.550 146.440 41.690 151.560 ;
        RECT 43.330 151.220 43.590 151.540 ;
        RECT 42.410 148.840 42.670 149.160 ;
        RECT 42.470 147.120 42.610 148.840 ;
        RECT 42.410 146.800 42.670 147.120 ;
        RECT 41.030 146.120 41.290 146.440 ;
        RECT 41.490 146.120 41.750 146.440 ;
        RECT 43.390 143.720 43.530 151.220 ;
        RECT 47.990 149.160 48.130 154.280 ;
        RECT 47.930 148.840 48.190 149.160 ;
        RECT 45.170 148.500 45.430 148.820 ;
        RECT 45.230 144.060 45.370 148.500 ;
        RECT 45.630 146.460 45.890 146.780 ;
        RECT 45.170 143.740 45.430 144.060 ;
        RECT 30.450 139.660 30.710 139.980 ;
        RECT 30.800 139.125 32.340 139.495 ;
        RECT 34.190 138.620 34.330 143.660 ;
        RECT 38.270 143.400 38.530 143.720 ;
        RECT 40.110 143.400 40.370 143.720 ;
        RECT 43.330 143.400 43.590 143.720 ;
        RECT 35.050 143.060 35.310 143.380 ;
        RECT 35.110 141.680 35.250 143.060 ;
        RECT 37.810 142.380 38.070 142.700 ;
        RECT 35.050 141.360 35.310 141.680 ;
        RECT 37.870 140.660 38.010 142.380 ;
        RECT 38.330 141.000 38.470 143.400 ;
        RECT 41.030 142.380 41.290 142.700 ;
        RECT 44.250 142.380 44.510 142.700 ;
        RECT 38.270 140.680 38.530 141.000 ;
        RECT 35.510 140.340 35.770 140.660 ;
        RECT 37.810 140.340 38.070 140.660 ;
        RECT 34.130 138.300 34.390 138.620 ;
        RECT 35.570 137.940 35.710 140.340 ;
        RECT 35.510 137.620 35.770 137.940 ;
        RECT 32.750 135.580 33.010 135.900 ;
        RECT 30.450 134.960 30.710 135.220 ;
        RECT 30.050 134.900 30.710 134.960 ;
        RECT 30.050 134.820 30.650 134.900 ;
        RECT 27.690 134.220 27.950 134.540 ;
        RECT 26.830 132.100 27.430 132.240 ;
        RECT 26.830 130.370 26.970 132.100 ;
        RECT 27.750 131.820 27.890 134.220 ;
        RECT 30.050 133.520 30.190 134.820 ;
        RECT 30.800 133.685 32.340 134.055 ;
        RECT 29.990 133.200 30.250 133.520 ;
        RECT 29.530 132.180 29.790 132.500 ;
        RECT 27.690 131.500 27.950 131.820 ;
        RECT 27.500 130.965 29.040 131.335 ;
        RECT 26.830 130.230 27.430 130.370 ;
        RECT 27.290 129.440 27.430 130.230 ;
        RECT 27.230 129.120 27.490 129.440 ;
        RECT 25.390 128.780 25.650 129.100 ;
        RECT 25.450 124.680 25.590 128.780 ;
        RECT 27.290 128.080 27.430 129.120 ;
        RECT 27.230 127.760 27.490 128.080 ;
        RECT 27.500 125.525 29.040 125.895 ;
        RECT 25.390 124.360 25.650 124.680 ;
        RECT 29.590 122.640 29.730 132.180 ;
        RECT 29.990 131.500 30.250 131.820 ;
        RECT 29.530 122.320 29.790 122.640 ;
        RECT 21.710 121.640 21.970 121.960 ;
        RECT 22.170 121.640 22.430 121.960 ;
        RECT 21.770 119.240 21.910 121.640 ;
        RECT 22.230 119.920 22.370 121.640 ;
        RECT 27.500 120.085 29.040 120.455 ;
        RECT 30.050 119.920 30.190 131.500 ;
        RECT 32.810 130.120 32.950 135.580 ;
        RECT 35.570 135.220 35.710 137.620 ;
        RECT 41.090 135.220 41.230 142.380 ;
        RECT 43.790 140.000 44.050 140.320 ;
        RECT 43.850 138.960 43.990 140.000 ;
        RECT 43.790 138.640 44.050 138.960 ;
        RECT 44.310 138.280 44.450 142.380 ;
        RECT 45.690 138.960 45.830 146.460 ;
        RECT 47.470 145.780 47.730 146.100 ;
        RECT 46.090 145.440 46.350 145.760 ;
        RECT 46.150 142.700 46.290 145.440 ;
        RECT 46.090 142.380 46.350 142.700 ;
        RECT 46.150 138.960 46.290 142.380 ;
        RECT 47.530 139.980 47.670 145.780 ;
        RECT 48.450 145.760 48.590 156.320 ;
        RECT 48.910 155.280 49.050 160.400 ;
        RECT 52.130 160.040 52.270 161.420 ;
        RECT 52.070 159.720 52.330 160.040 ;
        RECT 51.150 159.040 51.410 159.360 ;
        RECT 51.210 157.660 51.350 159.040 ;
        RECT 51.150 157.340 51.410 157.660 ;
        RECT 48.850 155.190 49.110 155.280 ;
        RECT 48.850 155.050 49.510 155.190 ;
        RECT 48.850 154.960 49.110 155.050 ;
        RECT 48.850 153.260 49.110 153.580 ;
        RECT 48.910 152.560 49.050 153.260 ;
        RECT 48.850 152.240 49.110 152.560 ;
        RECT 49.370 151.540 49.510 155.050 ;
        RECT 52.130 154.600 52.270 159.720 ;
        RECT 52.070 154.280 52.330 154.600 ;
        RECT 50.230 153.260 50.490 153.580 ;
        RECT 50.290 151.880 50.430 153.260 ;
        RECT 50.230 151.560 50.490 151.880 ;
        RECT 49.310 151.220 49.570 151.540 ;
        RECT 49.770 150.880 50.030 151.200 ;
        RECT 48.850 148.840 49.110 149.160 ;
        RECT 48.390 145.440 48.650 145.760 ;
        RECT 48.910 144.060 49.050 148.840 ;
        RECT 49.830 144.400 49.970 150.880 ;
        RECT 49.770 144.080 50.030 144.400 ;
        RECT 48.850 143.740 49.110 144.060 ;
        RECT 47.930 143.400 48.190 143.720 ;
        RECT 47.990 141.340 48.130 143.400 ;
        RECT 48.390 142.720 48.650 143.040 ;
        RECT 47.930 141.020 48.190 141.340 ;
        RECT 47.470 139.660 47.730 139.980 ;
        RECT 45.630 138.640 45.890 138.960 ;
        RECT 46.090 138.640 46.350 138.960 ;
        RECT 44.250 137.960 44.510 138.280 ;
        RECT 45.690 136.240 45.830 138.640 ;
        RECT 47.530 137.940 47.670 139.660 ;
        RECT 48.450 138.960 48.590 142.720 ;
        RECT 48.910 141.680 49.050 143.740 ;
        RECT 48.850 141.360 49.110 141.680 ;
        RECT 48.910 138.960 49.050 141.360 ;
        RECT 49.830 141.000 49.970 144.080 ;
        RECT 52.070 142.380 52.330 142.700 ;
        RECT 51.150 141.020 51.410 141.340 ;
        RECT 49.770 140.680 50.030 141.000 ;
        RECT 49.310 140.000 49.570 140.320 ;
        RECT 48.390 138.640 48.650 138.960 ;
        RECT 48.850 138.640 49.110 138.960 ;
        RECT 49.370 138.360 49.510 140.000 ;
        RECT 48.910 138.280 49.510 138.360 ;
        RECT 49.830 138.280 49.970 140.680 ;
        RECT 51.210 138.280 51.350 141.020 ;
        RECT 52.130 140.660 52.270 142.380 ;
        RECT 52.070 140.340 52.330 140.660 ;
        RECT 51.610 140.000 51.870 140.320 ;
        RECT 51.670 138.960 51.810 140.000 ;
        RECT 51.610 138.640 51.870 138.960 ;
        RECT 52.130 138.360 52.270 140.340 ;
        RECT 48.850 138.220 49.510 138.280 ;
        RECT 48.850 137.960 49.110 138.220 ;
        RECT 49.770 137.960 50.030 138.280 ;
        RECT 51.150 137.960 51.410 138.280 ;
        RECT 51.670 138.220 52.270 138.360 ;
        RECT 47.470 137.620 47.730 137.940 ;
        RECT 41.490 135.920 41.750 136.240 ;
        RECT 45.630 135.920 45.890 136.240 ;
        RECT 35.510 134.900 35.770 135.220 ;
        RECT 41.030 134.900 41.290 135.220 ;
        RECT 33.210 134.560 33.470 134.880 ;
        RECT 33.270 131.820 33.410 134.560 ;
        RECT 34.590 132.180 34.850 132.500 ;
        RECT 33.210 131.500 33.470 131.820 ;
        RECT 32.750 129.800 33.010 130.120 ;
        RECT 30.800 128.245 32.340 128.615 ;
        RECT 34.650 128.080 34.790 132.180 ;
        RECT 35.570 129.780 35.710 134.900 ;
        RECT 38.270 134.560 38.530 134.880 ;
        RECT 38.330 132.160 38.470 134.560 ;
        RECT 41.550 132.840 41.690 135.920 ;
        RECT 47.530 135.560 47.670 137.620 ;
        RECT 48.390 136.940 48.650 137.260 ;
        RECT 47.470 135.240 47.730 135.560 ;
        RECT 46.090 134.220 46.350 134.540 ;
        RECT 46.150 132.840 46.290 134.220 ;
        RECT 47.530 133.180 47.670 135.240 ;
        RECT 47.470 132.860 47.730 133.180 ;
        RECT 41.490 132.520 41.750 132.840 ;
        RECT 45.630 132.520 45.890 132.840 ;
        RECT 46.090 132.520 46.350 132.840 ;
        RECT 38.270 131.840 38.530 132.160 ;
        RECT 36.430 131.500 36.690 131.820 ;
        RECT 41.490 131.500 41.750 131.820 ;
        RECT 44.250 131.500 44.510 131.820 ;
        RECT 36.490 129.780 36.630 131.500 ;
        RECT 41.030 130.140 41.290 130.460 ;
        RECT 35.510 129.460 35.770 129.780 ;
        RECT 36.430 129.460 36.690 129.780 ;
        RECT 39.190 129.520 39.450 129.780 ;
        RECT 39.190 129.460 39.850 129.520 ;
        RECT 34.590 127.760 34.850 128.080 ;
        RECT 33.670 127.080 33.930 127.400 ;
        RECT 33.730 125.360 33.870 127.080 ;
        RECT 35.570 126.720 35.710 129.460 ;
        RECT 39.250 129.380 39.850 129.460 ;
        RECT 39.190 128.780 39.450 129.100 ;
        RECT 35.970 126.740 36.230 127.060 ;
        RECT 38.730 126.740 38.990 127.060 ;
        RECT 35.510 126.400 35.770 126.720 ;
        RECT 36.030 125.440 36.170 126.740 ;
        RECT 38.270 126.060 38.530 126.380 ;
        RECT 33.670 125.040 33.930 125.360 ;
        RECT 35.570 125.300 36.170 125.440 ;
        RECT 35.570 124.680 35.710 125.300 ;
        RECT 35.970 124.700 36.230 125.020 ;
        RECT 38.330 124.760 38.470 126.060 ;
        RECT 38.790 125.360 38.930 126.740 ;
        RECT 38.730 125.040 38.990 125.360 ;
        RECT 35.510 124.360 35.770 124.680 ;
        RECT 30.450 123.340 30.710 123.660 ;
        RECT 22.170 119.600 22.430 119.920 ;
        RECT 23.090 119.600 23.350 119.920 ;
        RECT 29.990 119.600 30.250 119.920 ;
        RECT 21.710 118.920 21.970 119.240 ;
        RECT 16.650 117.900 16.910 118.220 ;
        RECT 10.660 116.345 10.940 116.715 ;
        RECT 10.670 116.200 10.930 116.345 ;
        RECT 15.270 115.520 15.530 115.840 ;
        RECT 10.670 113.315 10.930 113.460 ;
        RECT 6.990 112.800 7.250 113.120 ;
        RECT 10.660 112.945 10.940 113.315 ;
        RECT 15.330 111.080 15.470 115.520 ;
        RECT 15.730 113.140 15.990 113.460 ;
        RECT 15.270 110.760 15.530 111.080 ;
        RECT 12.960 108.865 13.240 109.235 ;
        RECT 13.030 104.960 13.170 108.865 ;
        RECT 15.330 107.680 15.470 110.760 ;
        RECT 13.890 107.360 14.150 107.680 ;
        RECT 15.270 107.360 15.530 107.680 ;
        RECT 13.950 106.320 14.090 107.360 ;
        RECT 13.890 106.000 14.150 106.320 ;
        RECT 15.330 105.980 15.470 107.360 ;
        RECT 15.790 105.980 15.930 113.140 ;
        RECT 16.710 111.080 16.850 117.900 ;
        RECT 21.770 113.460 21.910 118.920 ;
        RECT 23.150 118.900 23.290 119.600 ;
        RECT 23.090 118.580 23.350 118.900 ;
        RECT 23.550 118.580 23.810 118.900 ;
        RECT 22.630 118.240 22.890 118.560 ;
        RECT 22.690 116.860 22.830 118.240 ;
        RECT 23.090 117.900 23.350 118.220 ;
        RECT 22.630 116.540 22.890 116.860 ;
        RECT 20.330 113.140 20.590 113.460 ;
        RECT 21.710 113.140 21.970 113.460 ;
        RECT 18.030 112.460 18.290 112.780 ;
        RECT 16.650 110.760 16.910 111.080 ;
        RECT 16.190 110.420 16.450 110.740 ;
        RECT 15.270 105.660 15.530 105.980 ;
        RECT 15.730 105.660 15.990 105.980 ;
        RECT 16.250 105.300 16.390 110.420 ;
        RECT 16.190 104.980 16.450 105.300 ;
        RECT 12.970 104.640 13.230 104.960 ;
        RECT 10.660 102.745 10.940 103.115 ;
        RECT 10.730 102.580 10.870 102.745 ;
        RECT 16.710 102.580 16.850 110.760 ;
        RECT 17.110 109.740 17.370 110.060 ;
        RECT 17.170 105.640 17.310 109.740 ;
        RECT 18.090 105.980 18.230 112.460 ;
        RECT 20.390 111.670 20.530 113.140 ;
        RECT 21.770 111.760 21.910 113.140 ;
        RECT 19.930 111.530 20.530 111.670 ;
        RECT 19.930 109.040 20.070 111.530 ;
        RECT 20.790 111.440 21.050 111.760 ;
        RECT 21.710 111.440 21.970 111.760 ;
        RECT 20.330 110.760 20.590 111.080 ;
        RECT 19.870 108.720 20.130 109.040 ;
        RECT 18.030 105.660 18.290 105.980 ;
        RECT 19.930 105.640 20.070 108.720 ;
        RECT 20.390 108.020 20.530 110.760 ;
        RECT 20.330 107.700 20.590 108.020 ;
        RECT 20.850 105.980 20.990 111.440 ;
        RECT 21.710 110.760 21.970 111.080 ;
        RECT 21.770 109.040 21.910 110.760 ;
        RECT 21.710 108.720 21.970 109.040 ;
        RECT 22.170 108.040 22.430 108.360 ;
        RECT 21.250 107.700 21.510 108.020 ;
        RECT 20.790 105.660 21.050 105.980 ;
        RECT 17.110 105.320 17.370 105.640 ;
        RECT 19.870 105.320 20.130 105.640 ;
        RECT 21.310 103.600 21.450 107.700 ;
        RECT 22.230 106.320 22.370 108.040 ;
        RECT 23.150 108.020 23.290 117.900 ;
        RECT 23.610 116.520 23.750 118.580 ;
        RECT 24.930 118.240 25.190 118.560 ;
        RECT 23.550 116.200 23.810 116.520 ;
        RECT 24.990 115.840 25.130 118.240 ;
        RECT 29.530 117.900 29.790 118.220 ;
        RECT 25.850 116.540 26.110 116.860 ;
        RECT 25.910 116.180 26.050 116.540 ;
        RECT 25.850 115.860 26.110 116.180 ;
        RECT 24.930 115.520 25.190 115.840 ;
        RECT 25.390 112.800 25.650 113.120 ;
        RECT 24.930 108.380 25.190 108.700 ;
        RECT 23.090 107.700 23.350 108.020 ;
        RECT 24.470 107.700 24.730 108.020 ;
        RECT 24.530 106.400 24.670 107.700 ;
        RECT 22.170 106.000 22.430 106.320 ;
        RECT 22.690 106.260 24.670 106.400 ;
        RECT 21.700 105.465 21.980 105.835 ;
        RECT 21.710 105.320 21.970 105.465 ;
        RECT 22.170 104.980 22.430 105.300 ;
        RECT 20.330 103.280 20.590 103.600 ;
        RECT 21.250 103.280 21.510 103.600 ;
        RECT 10.670 102.260 10.930 102.580 ;
        RECT 16.650 102.260 16.910 102.580 ;
        RECT 18.030 102.260 18.290 102.580 ;
        RECT 17.110 101.580 17.370 101.900 ;
        RECT 13.430 99.880 13.690 100.200 ;
        RECT 13.490 92.040 13.630 99.880 ;
        RECT 17.170 98.160 17.310 101.580 ;
        RECT 18.090 98.160 18.230 102.260 ;
        RECT 20.390 99.600 20.530 103.280 ;
        RECT 22.230 102.920 22.370 104.980 ;
        RECT 22.690 103.260 22.830 106.260 ;
        RECT 24.010 105.660 24.270 105.980 ;
        RECT 23.090 104.640 23.350 104.960 ;
        RECT 22.630 102.940 22.890 103.260 ;
        RECT 22.170 102.600 22.430 102.920 ;
        RECT 22.170 101.920 22.430 102.240 ;
        RECT 20.790 101.580 21.050 101.900 ;
        RECT 20.850 100.200 20.990 101.580 ;
        RECT 22.230 100.880 22.370 101.920 ;
        RECT 22.690 100.880 22.830 102.940 ;
        RECT 22.170 100.560 22.430 100.880 ;
        RECT 22.630 100.560 22.890 100.880 ;
        RECT 20.790 99.880 21.050 100.200 ;
        RECT 23.150 99.980 23.290 104.640 ;
        RECT 19.930 99.460 20.530 99.600 ;
        RECT 22.690 99.840 23.290 99.980 ;
        RECT 24.070 99.860 24.210 105.660 ;
        RECT 24.530 105.300 24.670 106.260 ;
        RECT 24.990 105.640 25.130 108.380 ;
        RECT 25.450 107.680 25.590 112.800 ;
        RECT 25.910 111.080 26.050 115.860 ;
        RECT 29.590 115.840 29.730 117.900 ;
        RECT 30.510 116.520 30.650 123.340 ;
        RECT 30.800 122.805 32.340 123.175 ;
        RECT 32.750 117.900 33.010 118.220 ;
        RECT 30.800 117.365 32.340 117.735 ;
        RECT 32.810 116.860 32.950 117.900 ;
        RECT 32.750 116.540 33.010 116.860 ;
        RECT 30.450 116.200 30.710 116.520 ;
        RECT 29.530 115.520 29.790 115.840 ;
        RECT 27.500 114.645 29.040 115.015 ;
        RECT 29.590 111.080 29.730 115.520 ;
        RECT 30.510 115.500 30.650 116.200 ;
        RECT 35.510 115.860 35.770 116.180 ;
        RECT 36.030 115.920 36.170 124.700 ;
        RECT 36.950 124.620 38.470 124.760 ;
        RECT 36.430 124.250 36.690 124.340 ;
        RECT 36.950 124.250 37.090 124.620 ;
        RECT 38.330 124.340 38.470 124.620 ;
        RECT 36.430 124.110 37.090 124.250 ;
        RECT 36.430 124.020 36.690 124.110 ;
        RECT 36.430 117.900 36.690 118.220 ;
        RECT 36.490 116.520 36.630 117.900 ;
        RECT 36.430 116.200 36.690 116.520 ;
        RECT 30.450 115.180 30.710 115.500 ;
        RECT 34.590 115.180 34.850 115.500 ;
        RECT 29.990 113.140 30.250 113.460 ;
        RECT 30.050 111.080 30.190 113.140 ;
        RECT 30.800 111.925 32.340 112.295 ;
        RECT 34.650 111.420 34.790 115.180 ;
        RECT 35.570 113.200 35.710 115.860 ;
        RECT 36.030 115.780 36.630 115.920 ;
        RECT 35.970 115.180 36.230 115.500 ;
        RECT 35.110 113.060 35.710 113.200 ;
        RECT 34.590 111.100 34.850 111.420 ;
        RECT 35.110 111.080 35.250 113.060 ;
        RECT 35.510 112.460 35.770 112.780 ;
        RECT 25.850 110.760 26.110 111.080 ;
        RECT 29.530 110.760 29.790 111.080 ;
        RECT 29.990 110.760 30.250 111.080 ;
        RECT 35.050 110.760 35.310 111.080 ;
        RECT 25.910 109.040 26.050 110.760 ;
        RECT 26.310 109.740 26.570 110.060 ;
        RECT 26.770 109.740 27.030 110.060 ;
        RECT 26.370 109.040 26.510 109.740 ;
        RECT 25.850 108.720 26.110 109.040 ;
        RECT 26.310 108.720 26.570 109.040 ;
        RECT 26.830 108.700 26.970 109.740 ;
        RECT 27.500 109.205 29.040 109.575 ;
        RECT 26.770 108.380 27.030 108.700 ;
        RECT 29.590 108.020 29.730 110.760 ;
        RECT 35.110 109.040 35.250 110.760 ;
        RECT 35.050 108.720 35.310 109.040 ;
        RECT 35.570 108.360 35.710 112.460 ;
        RECT 35.510 108.040 35.770 108.360 ;
        RECT 36.030 108.020 36.170 115.180 ;
        RECT 29.530 107.700 29.790 108.020 ;
        RECT 35.970 107.700 36.230 108.020 ;
        RECT 25.390 107.360 25.650 107.680 ;
        RECT 29.990 107.360 30.250 107.680 ;
        RECT 24.930 105.320 25.190 105.640 ;
        RECT 25.390 105.320 25.650 105.640 ;
        RECT 24.470 104.980 24.730 105.300 ;
        RECT 24.470 104.300 24.730 104.620 ;
        RECT 24.930 104.300 25.190 104.620 ;
        RECT 17.110 97.840 17.370 98.160 ;
        RECT 18.030 97.840 18.290 98.160 ;
        RECT 17.170 95.100 17.310 97.840 ;
        RECT 17.110 94.780 17.370 95.100 ;
        RECT 19.930 94.420 20.070 99.460 ;
        RECT 20.330 98.860 20.590 99.180 ;
        RECT 20.790 98.860 21.050 99.180 ;
        RECT 20.390 97.140 20.530 98.860 ;
        RECT 20.330 96.820 20.590 97.140 ;
        RECT 17.570 94.100 17.830 94.420 ;
        RECT 19.870 94.100 20.130 94.420 ;
        RECT 14.810 93.420 15.070 93.740 ;
        RECT 13.430 91.720 13.690 92.040 ;
        RECT 14.870 91.360 15.010 93.420 ;
        RECT 17.630 92.120 17.770 94.100 ;
        RECT 20.390 93.740 20.530 96.820 ;
        RECT 20.330 93.420 20.590 93.740 ;
        RECT 17.170 91.980 17.770 92.120 ;
        RECT 14.810 91.040 15.070 91.360 ;
        RECT 17.170 90.000 17.310 91.980 ;
        RECT 20.330 91.380 20.590 91.700 ;
        RECT 17.570 91.040 17.830 91.360 ;
        RECT 17.110 89.680 17.370 90.000 ;
        RECT 17.630 89.320 17.770 91.040 ;
        RECT 20.390 89.660 20.530 91.380 ;
        RECT 20.850 91.020 20.990 98.860 ;
        RECT 21.250 96.480 21.510 96.800 ;
        RECT 21.310 94.760 21.450 96.480 ;
        RECT 21.710 95.120 21.970 95.440 ;
        RECT 21.250 94.440 21.510 94.760 ;
        RECT 21.250 93.760 21.510 94.080 ;
        RECT 21.310 92.720 21.450 93.760 ;
        RECT 21.250 92.400 21.510 92.720 ;
        RECT 21.770 92.120 21.910 95.120 ;
        RECT 21.770 92.040 22.370 92.120 ;
        RECT 21.710 91.980 22.370 92.040 ;
        RECT 21.710 91.720 21.970 91.980 ;
        RECT 21.710 91.040 21.970 91.360 ;
        RECT 20.790 90.930 21.050 91.020 ;
        RECT 20.790 90.790 21.450 90.930 ;
        RECT 20.790 90.700 21.050 90.790 ;
        RECT 20.330 89.340 20.590 89.660 ;
        RECT 17.570 89.000 17.830 89.320 ;
        RECT 18.950 85.260 19.210 85.580 ;
        RECT 19.010 80.820 19.150 85.260 ;
        RECT 18.950 80.730 19.210 80.820 ;
        RECT 18.950 80.590 19.610 80.730 ;
        RECT 18.950 80.500 19.210 80.590 ;
        RECT 19.470 80.140 19.610 80.590 ;
        RECT 19.870 80.160 20.130 80.480 ;
        RECT 17.110 79.820 17.370 80.140 ;
        RECT 19.410 79.820 19.670 80.140 ;
        RECT 15.730 78.120 15.990 78.440 ;
        RECT 15.790 76.400 15.930 78.120 ;
        RECT 15.730 76.080 15.990 76.400 ;
        RECT 16.650 75.400 16.910 75.720 ;
        RECT 16.710 72.660 16.850 75.400 ;
        RECT 17.170 75.380 17.310 79.820 ;
        RECT 17.110 75.060 17.370 75.380 ;
        RECT 19.470 75.040 19.610 79.820 ;
        RECT 19.930 75.720 20.070 80.160 ;
        RECT 20.390 78.780 20.530 89.340 ;
        RECT 20.790 89.000 21.050 89.320 ;
        RECT 20.850 87.280 20.990 89.000 ;
        RECT 20.790 86.960 21.050 87.280 ;
        RECT 20.790 85.600 21.050 85.920 ;
        RECT 20.850 84.640 20.990 85.600 ;
        RECT 21.310 85.580 21.450 90.790 ;
        RECT 21.770 88.300 21.910 91.040 ;
        RECT 21.710 87.980 21.970 88.300 ;
        RECT 21.250 85.260 21.510 85.580 ;
        RECT 21.770 84.640 21.910 87.980 ;
        RECT 22.230 86.940 22.370 91.980 ;
        RECT 22.170 86.620 22.430 86.940 ;
        RECT 22.170 85.940 22.430 86.260 ;
        RECT 20.850 84.500 21.910 84.640 ;
        RECT 20.850 81.500 20.990 84.500 ;
        RECT 21.250 81.520 21.510 81.840 ;
        RECT 20.790 81.180 21.050 81.500 ;
        RECT 21.310 80.820 21.450 81.520 ;
        RECT 22.230 81.160 22.370 85.940 ;
        RECT 22.170 80.840 22.430 81.160 ;
        RECT 21.250 80.500 21.510 80.820 ;
        RECT 21.310 79.120 21.450 80.500 ;
        RECT 22.170 80.160 22.430 80.480 ;
        RECT 21.250 78.800 21.510 79.120 ;
        RECT 20.330 78.460 20.590 78.780 ;
        RECT 19.870 75.400 20.130 75.720 ;
        RECT 19.410 74.720 19.670 75.040 ;
        RECT 20.390 73.340 20.530 78.460 ;
        RECT 21.310 76.400 21.450 78.800 ;
        RECT 22.230 78.440 22.370 80.160 ;
        RECT 22.170 78.120 22.430 78.440 ;
        RECT 22.230 76.400 22.370 78.120 ;
        RECT 21.250 76.080 21.510 76.400 ;
        RECT 22.170 76.080 22.430 76.400 ;
        RECT 21.310 75.380 21.450 76.080 ;
        RECT 21.250 75.060 21.510 75.380 ;
        RECT 20.790 74.380 21.050 74.700 ;
        RECT 20.330 73.020 20.590 73.340 ;
        RECT 19.870 72.680 20.130 73.000 ;
        RECT 16.650 72.340 16.910 72.660 ;
        RECT 19.410 72.000 19.670 72.320 ;
        RECT 13.890 71.660 14.150 71.980 ;
        RECT 17.570 71.660 17.830 71.980 ;
        RECT 13.950 69.600 14.090 71.660 ;
        RECT 13.890 69.280 14.150 69.600 ;
        RECT 12.960 68.065 13.240 68.435 ;
        RECT 12.970 67.920 13.230 68.065 ;
        RECT 17.630 67.560 17.770 71.660 ;
        RECT 19.470 70.960 19.610 72.000 ;
        RECT 18.030 70.640 18.290 70.960 ;
        RECT 19.410 70.640 19.670 70.960 ;
        RECT 17.570 67.240 17.830 67.560 ;
        RECT 18.090 66.540 18.230 70.640 ;
        RECT 19.930 70.620 20.070 72.680 ;
        RECT 19.870 70.300 20.130 70.620 ;
        RECT 19.930 66.960 20.070 70.300 ;
        RECT 20.390 69.940 20.530 73.020 ;
        RECT 20.850 72.660 20.990 74.380 ;
        RECT 21.250 73.360 21.510 73.680 ;
        RECT 21.310 73.000 21.450 73.360 ;
        RECT 21.250 72.680 21.510 73.000 ;
        RECT 20.790 72.340 21.050 72.660 ;
        RECT 20.330 69.620 20.590 69.940 ;
        RECT 20.390 67.900 20.530 69.620 ;
        RECT 20.330 67.580 20.590 67.900 ;
        RECT 19.470 66.820 20.070 66.960 ;
        RECT 18.030 66.220 18.290 66.540 ;
        RECT 10.660 63.985 10.940 64.355 ;
        RECT 14.810 64.180 15.070 64.500 ;
        RECT 10.730 63.820 10.870 63.985 ;
        RECT 10.670 63.500 10.930 63.820 ;
        RECT 12.040 61.265 12.320 61.635 ;
        RECT 14.870 61.440 15.010 64.180 ;
        RECT 15.730 63.500 15.990 63.820 ;
        RECT 12.110 60.080 12.250 61.265 ;
        RECT 14.810 61.120 15.070 61.440 ;
        RECT 12.050 59.760 12.310 60.080 ;
        RECT 15.270 58.740 15.530 59.060 ;
        RECT 12.960 54.465 13.240 54.835 ;
        RECT 11.580 51.065 11.860 51.435 ;
        RECT 11.650 50.560 11.790 51.065 ;
        RECT 11.590 50.240 11.850 50.560 ;
        RECT 13.030 50.220 13.170 54.465 ;
        RECT 15.330 53.960 15.470 58.740 ;
        RECT 15.790 58.235 15.930 63.500 ;
        RECT 17.110 60.780 17.370 61.100 ;
        RECT 16.650 58.400 16.910 58.720 ;
        RECT 15.720 57.865 16.000 58.235 ;
        RECT 16.710 57.360 16.850 58.400 ;
        RECT 16.650 57.040 16.910 57.360 ;
        RECT 17.170 56.680 17.310 60.780 ;
        RECT 17.570 58.400 17.830 58.720 ;
        RECT 17.630 56.680 17.770 58.400 ;
        RECT 18.030 58.060 18.290 58.380 ;
        RECT 17.110 56.360 17.370 56.680 ;
        RECT 17.570 56.360 17.830 56.680 ;
        RECT 15.270 53.640 15.530 53.960 ;
        RECT 13.430 52.960 13.690 53.280 ;
        RECT 12.970 49.900 13.230 50.220 ;
        RECT 10.670 48.715 10.930 48.860 ;
        RECT 10.660 48.345 10.940 48.715 ;
        RECT 13.490 46.140 13.630 52.960 ;
        RECT 14.810 52.620 15.070 52.940 ;
        RECT 14.870 51.240 15.010 52.620 ;
        RECT 14.810 50.920 15.070 51.240 ;
        RECT 14.810 49.900 15.070 50.220 ;
        RECT 14.870 48.180 15.010 49.900 ;
        RECT 14.810 47.860 15.070 48.180 ;
        RECT 13.430 45.820 13.690 46.140 ;
        RECT 15.330 45.460 15.470 53.640 ;
        RECT 18.090 48.180 18.230 58.060 ;
        RECT 19.470 57.440 19.610 66.820 ;
        RECT 19.870 66.220 20.130 66.540 ;
        RECT 19.930 58.380 20.070 66.220 ;
        RECT 20.390 62.120 20.530 67.580 ;
        RECT 21.250 64.180 21.510 64.500 ;
        RECT 20.790 62.140 21.050 62.460 ;
        RECT 20.330 61.800 20.590 62.120 ;
        RECT 20.850 59.740 20.990 62.140 ;
        RECT 21.310 61.780 21.450 64.180 ;
        RECT 21.710 63.500 21.970 63.820 ;
        RECT 21.250 61.460 21.510 61.780 ;
        RECT 21.310 60.080 21.450 61.460 ;
        RECT 21.250 59.760 21.510 60.080 ;
        RECT 20.790 59.420 21.050 59.740 ;
        RECT 20.850 59.060 20.990 59.420 ;
        RECT 20.790 58.740 21.050 59.060 ;
        RECT 21.770 58.720 21.910 63.500 ;
        RECT 22.690 61.780 22.830 99.840 ;
        RECT 24.010 99.540 24.270 99.860 ;
        RECT 24.070 96.800 24.210 99.540 ;
        RECT 24.010 96.480 24.270 96.800 ;
        RECT 24.010 94.100 24.270 94.420 ;
        RECT 23.550 93.760 23.810 94.080 ;
        RECT 23.090 92.400 23.350 92.720 ;
        RECT 23.150 90.000 23.290 92.400 ;
        RECT 23.090 89.680 23.350 90.000 ;
        RECT 23.150 88.640 23.290 89.680 ;
        RECT 23.090 88.320 23.350 88.640 ;
        RECT 23.150 81.840 23.290 88.320 ;
        RECT 23.090 81.520 23.350 81.840 ;
        RECT 23.610 78.350 23.750 93.760 ;
        RECT 24.070 91.700 24.210 94.100 ;
        RECT 24.530 92.720 24.670 104.300 ;
        RECT 24.990 102.580 25.130 104.300 ;
        RECT 25.450 102.920 25.590 105.320 ;
        RECT 27.500 103.765 29.040 104.135 ;
        RECT 25.390 102.600 25.650 102.920 ;
        RECT 24.930 102.260 25.190 102.580 ;
        RECT 24.930 99.540 25.190 99.860 ;
        RECT 24.990 95.440 25.130 99.540 ;
        RECT 25.450 97.480 25.590 102.600 ;
        RECT 27.500 98.325 29.040 98.695 ;
        RECT 25.390 97.160 25.650 97.480 ;
        RECT 24.930 95.120 25.190 95.440 ;
        RECT 25.450 94.760 25.590 97.160 ;
        RECT 25.390 94.440 25.650 94.760 ;
        RECT 26.310 94.440 26.570 94.760 ;
        RECT 24.470 92.400 24.730 92.720 ;
        RECT 24.010 91.380 24.270 91.700 ;
        RECT 24.930 89.680 25.190 90.000 ;
        RECT 24.990 88.300 25.130 89.680 ;
        RECT 25.450 88.980 25.590 94.440 ;
        RECT 26.370 92.720 26.510 94.440 ;
        RECT 27.500 92.885 29.040 93.255 ;
        RECT 26.310 92.400 26.570 92.720 ;
        RECT 26.310 91.380 26.570 91.700 ;
        RECT 25.850 89.340 26.110 89.660 ;
        RECT 25.390 88.660 25.650 88.980 ;
        RECT 24.930 87.980 25.190 88.300 ;
        RECT 25.450 86.600 25.590 88.660 ;
        RECT 25.910 87.280 26.050 89.340 ;
        RECT 25.850 86.960 26.110 87.280 ;
        RECT 24.010 86.280 24.270 86.600 ;
        RECT 25.390 86.280 25.650 86.600 ;
        RECT 23.150 78.210 23.750 78.350 ;
        RECT 22.630 61.460 22.890 61.780 ;
        RECT 21.710 58.400 21.970 58.720 ;
        RECT 19.870 58.060 20.130 58.380 ;
        RECT 18.550 57.300 20.070 57.440 ;
        RECT 18.550 56.680 18.690 57.300 ;
        RECT 19.410 56.875 19.670 57.020 ;
        RECT 18.490 56.360 18.750 56.680 ;
        RECT 19.400 56.505 19.680 56.875 ;
        RECT 18.490 55.340 18.750 55.660 ;
        RECT 18.950 55.340 19.210 55.660 ;
        RECT 18.550 53.280 18.690 55.340 ;
        RECT 18.490 52.960 18.750 53.280 ;
        RECT 19.010 52.680 19.150 55.340 ;
        RECT 18.550 52.540 19.150 52.680 ;
        RECT 16.650 47.860 16.910 48.180 ;
        RECT 18.030 47.860 18.290 48.180 ;
        RECT 16.710 46.480 16.850 47.860 ;
        RECT 16.650 46.160 16.910 46.480 ;
        RECT 15.270 45.140 15.530 45.460 ;
        RECT 15.330 43.760 15.470 45.140 ;
        RECT 15.270 43.440 15.530 43.760 ;
        RECT 14.810 42.080 15.070 42.400 ;
        RECT 14.870 41.040 15.010 42.080 ;
        RECT 14.810 40.720 15.070 41.040 ;
        RECT 15.330 37.640 15.470 43.440 ;
        RECT 16.190 40.270 16.450 40.360 ;
        RECT 15.790 40.130 16.450 40.270 ;
        RECT 15.270 37.320 15.530 37.640 ;
        RECT 15.270 31.600 15.530 31.860 ;
        RECT 14.870 31.540 15.530 31.600 ;
        RECT 14.870 31.460 15.470 31.540 ;
        RECT 14.350 30.860 14.610 31.180 ;
        RECT 13.890 28.140 14.150 28.460 ;
        RECT 13.950 26.080 14.090 28.140 ;
        RECT 13.890 25.760 14.150 26.080 ;
        RECT 13.430 22.700 13.690 23.020 ;
        RECT 6.530 9.780 6.790 10.100 ;
        RECT 13.490 9.840 13.630 22.700 ;
        RECT 13.890 19.980 14.150 20.300 ;
        RECT 13.950 15.200 14.090 19.980 ;
        RECT 13.890 14.880 14.150 15.200 ;
        RECT 14.410 10.100 14.550 30.860 ;
        RECT 14.870 18.940 15.010 31.460 ;
        RECT 15.790 29.480 15.930 40.130 ;
        RECT 16.190 40.040 16.450 40.130 ;
        RECT 16.650 37.320 16.910 37.640 ;
        RECT 16.190 30.860 16.450 31.180 ;
        RECT 16.250 29.480 16.390 30.860 ;
        RECT 15.730 29.160 15.990 29.480 ;
        RECT 16.190 29.160 16.450 29.480 ;
        RECT 15.790 20.980 15.930 29.160 ;
        RECT 16.710 29.140 16.850 37.320 ;
        RECT 17.570 32.220 17.830 32.540 ;
        RECT 17.630 31.860 17.770 32.220 ;
        RECT 18.090 31.860 18.230 47.860 ;
        RECT 18.550 39.875 18.690 52.540 ;
        RECT 18.950 50.920 19.210 51.240 ;
        RECT 19.010 43.760 19.150 50.920 ;
        RECT 19.470 48.520 19.610 56.505 ;
        RECT 19.410 48.200 19.670 48.520 ;
        RECT 19.410 47.180 19.670 47.500 ;
        RECT 19.470 46.140 19.610 47.180 ;
        RECT 19.410 45.820 19.670 46.140 ;
        RECT 18.950 43.440 19.210 43.760 ;
        RECT 19.010 40.700 19.150 43.440 ;
        RECT 18.950 40.380 19.210 40.700 ;
        RECT 19.410 40.040 19.670 40.360 ;
        RECT 18.480 39.505 18.760 39.875 ;
        RECT 17.570 31.540 17.830 31.860 ;
        RECT 18.030 31.540 18.290 31.860 ;
        RECT 17.110 31.200 17.370 31.520 ;
        RECT 16.650 28.820 16.910 29.140 ;
        RECT 16.710 26.420 16.850 28.820 ;
        RECT 17.170 27.440 17.310 31.200 ;
        RECT 18.090 30.160 18.230 31.540 ;
        RECT 18.030 29.840 18.290 30.160 ;
        RECT 17.110 27.120 17.370 27.440 ;
        RECT 16.650 26.100 16.910 26.420 ;
        RECT 15.730 20.660 15.990 20.980 ;
        RECT 16.190 20.660 16.450 20.980 ;
        RECT 16.250 19.280 16.390 20.660 ;
        RECT 16.190 18.960 16.450 19.280 ;
        RECT 14.810 18.620 15.070 18.940 ;
        RECT 16.710 18.600 16.850 26.100 ;
        RECT 17.170 24.040 17.310 27.120 ;
        RECT 17.110 23.720 17.370 24.040 ;
        RECT 17.110 22.700 17.370 23.020 ;
        RECT 18.030 22.700 18.290 23.020 ;
        RECT 16.650 18.280 16.910 18.600 ;
        RECT 17.170 17.180 17.310 22.700 ;
        RECT 17.570 18.280 17.830 18.600 ;
        RECT 16.710 17.040 17.310 17.180 ;
        RECT 16.710 13.240 16.850 17.040 ;
        RECT 17.630 15.540 17.770 18.280 ;
        RECT 17.570 15.220 17.830 15.540 ;
        RECT 16.250 13.100 16.850 13.240 ;
        RECT 6.590 7.310 6.730 9.780 ;
        RECT 9.750 9.440 10.010 9.760 ;
        RECT 13.030 9.700 13.630 9.840 ;
        RECT 14.350 9.780 14.610 10.100 ;
        RECT 9.810 7.310 9.950 9.440 ;
        RECT 13.030 7.310 13.170 9.700 ;
        RECT 16.250 7.310 16.390 13.100 ;
        RECT 18.090 9.760 18.230 22.700 ;
        RECT 18.550 21.320 18.690 39.505 ;
        RECT 19.470 32.540 19.610 40.040 ;
        RECT 19.930 39.340 20.070 57.300 ;
        RECT 20.330 57.040 20.590 57.360 ;
        RECT 20.390 56.875 20.530 57.040 ;
        RECT 20.320 56.680 20.600 56.875 ;
        RECT 21.770 56.680 21.910 58.400 ;
        RECT 23.150 57.440 23.290 78.210 ;
        RECT 23.550 77.440 23.810 77.760 ;
        RECT 23.610 72.660 23.750 77.440 ;
        RECT 24.070 77.420 24.210 86.280 ;
        RECT 26.370 84.220 26.510 91.380 ;
        RECT 29.530 87.980 29.790 88.300 ;
        RECT 27.500 87.445 29.040 87.815 ;
        RECT 26.770 85.600 27.030 85.920 ;
        RECT 26.830 84.560 26.970 85.600 ;
        RECT 26.770 84.240 27.030 84.560 ;
        RECT 26.310 83.900 26.570 84.220 ;
        RECT 26.370 80.820 26.510 83.900 ;
        RECT 29.590 83.540 29.730 87.980 ;
        RECT 30.050 86.680 30.190 107.360 ;
        RECT 35.050 107.020 35.310 107.340 ;
        RECT 30.800 106.485 32.340 106.855 ;
        RECT 35.110 105.980 35.250 107.020 ;
        RECT 35.050 105.660 35.310 105.980 ;
        RECT 30.800 101.045 32.340 101.415 ;
        RECT 32.750 98.860 33.010 99.180 ;
        RECT 30.800 95.605 32.340 95.975 ;
        RECT 32.810 95.440 32.950 98.860 ;
        RECT 36.490 98.160 36.630 115.780 ;
        RECT 36.430 97.840 36.690 98.160 ;
        RECT 34.130 96.480 34.390 96.800 ;
        RECT 34.190 95.440 34.330 96.480 ;
        RECT 32.750 95.120 33.010 95.440 ;
        RECT 34.130 95.120 34.390 95.440 ;
        RECT 32.810 91.360 32.950 95.120 ;
        RECT 36.490 95.100 36.630 97.840 ;
        RECT 36.430 94.780 36.690 95.100 ;
        RECT 36.950 94.420 37.090 124.110 ;
        RECT 37.810 124.020 38.070 124.340 ;
        RECT 38.270 124.020 38.530 124.340 ;
        RECT 37.870 117.200 38.010 124.020 ;
        RECT 39.250 124.000 39.390 128.780 ;
        RECT 39.190 123.680 39.450 124.000 ;
        RECT 39.710 121.280 39.850 129.380 ;
        RECT 40.570 126.740 40.830 127.060 ;
        RECT 40.630 126.380 40.770 126.740 ;
        RECT 40.570 126.060 40.830 126.380 ;
        RECT 40.110 124.760 40.370 125.020 ;
        RECT 41.090 124.760 41.230 130.140 ;
        RECT 41.550 125.360 41.690 131.500 ;
        RECT 44.310 129.780 44.450 131.500 ;
        RECT 41.950 129.460 42.210 129.780 ;
        RECT 44.250 129.460 44.510 129.780 ;
        RECT 41.490 125.040 41.750 125.360 ;
        RECT 40.110 124.700 41.230 124.760 ;
        RECT 40.170 124.620 41.230 124.700 ;
        RECT 39.650 120.960 39.910 121.280 ;
        RECT 39.710 119.320 39.850 120.960 ;
        RECT 39.250 119.180 39.850 119.320 ;
        RECT 37.810 116.880 38.070 117.200 ;
        RECT 39.250 116.520 39.390 119.180 ;
        RECT 39.650 118.580 39.910 118.900 ;
        RECT 39.190 116.200 39.450 116.520 ;
        RECT 39.190 112.460 39.450 112.780 ;
        RECT 39.250 110.060 39.390 112.460 ;
        RECT 39.710 111.080 39.850 118.580 ;
        RECT 40.570 116.200 40.830 116.520 ;
        RECT 40.110 115.860 40.370 116.180 ;
        RECT 40.170 112.780 40.310 115.860 ;
        RECT 40.110 112.460 40.370 112.780 ;
        RECT 40.170 111.420 40.310 112.460 ;
        RECT 40.110 111.100 40.370 111.420 ;
        RECT 39.650 110.760 39.910 111.080 ;
        RECT 38.730 109.740 38.990 110.060 ;
        RECT 39.190 109.740 39.450 110.060 ;
        RECT 38.270 108.380 38.530 108.700 ;
        RECT 38.790 108.610 38.930 109.740 ;
        RECT 39.190 108.610 39.450 108.700 ;
        RECT 38.790 108.470 39.450 108.610 ;
        RECT 39.190 108.380 39.450 108.470 ;
        RECT 40.630 108.440 40.770 116.200 ;
        RECT 41.490 115.520 41.750 115.840 ;
        RECT 41.550 113.460 41.690 115.520 ;
        RECT 41.490 113.140 41.750 113.460 ;
        RECT 41.550 111.760 41.690 113.140 ;
        RECT 41.490 111.440 41.750 111.760 ;
        RECT 41.030 110.760 41.290 111.080 ;
        RECT 41.090 109.040 41.230 110.760 ;
        RECT 41.030 108.720 41.290 109.040 ;
        RECT 37.350 107.360 37.610 107.680 ;
        RECT 37.410 106.320 37.550 107.360 ;
        RECT 38.330 106.320 38.470 108.380 ;
        RECT 40.170 108.300 40.770 108.440 ;
        RECT 37.350 106.000 37.610 106.320 ;
        RECT 38.270 106.000 38.530 106.320 ;
        RECT 38.270 105.320 38.530 105.640 ;
        RECT 38.330 103.600 38.470 105.320 ;
        RECT 38.270 103.280 38.530 103.600 ;
        RECT 39.650 102.260 39.910 102.580 ;
        RECT 39.710 100.880 39.850 102.260 ;
        RECT 40.170 101.900 40.310 108.300 ;
        RECT 40.570 107.700 40.830 108.020 ;
        RECT 40.630 106.320 40.770 107.700 ;
        RECT 40.570 106.000 40.830 106.320 ;
        RECT 40.630 102.580 40.770 106.000 ;
        RECT 41.490 105.320 41.750 105.640 ;
        RECT 41.550 103.000 41.690 105.320 ;
        RECT 42.010 103.600 42.150 129.460 ;
        RECT 43.790 129.120 44.050 129.440 ;
        RECT 43.850 127.400 43.990 129.120 ;
        RECT 44.310 127.740 44.450 129.460 ;
        RECT 44.710 128.780 44.970 129.100 ;
        RECT 44.250 127.420 44.510 127.740 ;
        RECT 44.770 127.400 44.910 128.780 ;
        RECT 43.790 127.080 44.050 127.400 ;
        RECT 44.710 127.080 44.970 127.400 ;
        RECT 42.870 126.800 43.130 127.060 ;
        RECT 42.870 126.740 43.990 126.800 ;
        RECT 44.250 126.740 44.510 127.060 ;
        RECT 45.170 126.740 45.430 127.060 ;
        RECT 42.930 126.660 43.990 126.740 ;
        RECT 42.410 126.060 42.670 126.380 ;
        RECT 43.330 126.060 43.590 126.380 ;
        RECT 42.470 124.000 42.610 126.060 ;
        RECT 43.390 124.340 43.530 126.060 ;
        RECT 43.850 125.360 43.990 126.660 ;
        RECT 44.310 126.380 44.450 126.740 ;
        RECT 44.250 126.060 44.510 126.380 ;
        RECT 43.790 125.040 44.050 125.360 ;
        RECT 43.330 124.020 43.590 124.340 ;
        RECT 42.410 123.680 42.670 124.000 ;
        RECT 42.870 116.200 43.130 116.520 ;
        RECT 42.410 115.180 42.670 115.500 ;
        RECT 42.470 113.460 42.610 115.180 ;
        RECT 42.930 113.460 43.070 116.200 ;
        RECT 43.390 113.800 43.530 124.020 ;
        RECT 45.230 123.660 45.370 126.740 ;
        RECT 45.690 125.360 45.830 132.520 ;
        RECT 46.150 130.120 46.290 132.520 ;
        RECT 47.530 132.160 47.670 132.860 ;
        RECT 48.450 132.840 48.590 136.940 ;
        RECT 48.390 132.520 48.650 132.840 ;
        RECT 48.910 132.500 49.050 137.960 ;
        RECT 51.670 133.180 51.810 138.220 ;
        RECT 52.070 137.280 52.330 137.600 ;
        RECT 52.130 135.220 52.270 137.280 ;
        RECT 52.070 134.900 52.330 135.220 ;
        RECT 51.610 132.860 51.870 133.180 ;
        RECT 48.850 132.180 49.110 132.500 ;
        RECT 47.470 131.840 47.730 132.160 ;
        RECT 46.090 129.800 46.350 130.120 ;
        RECT 47.530 126.380 47.670 131.840 ;
        RECT 47.930 129.460 48.190 129.780 ;
        RECT 47.470 126.060 47.730 126.380 ;
        RECT 45.630 125.040 45.890 125.360 ;
        RECT 47.010 125.040 47.270 125.360 ;
        RECT 45.170 123.340 45.430 123.660 ;
        RECT 45.230 122.640 45.370 123.340 ;
        RECT 45.170 122.320 45.430 122.640 ;
        RECT 47.070 121.960 47.210 125.040 ;
        RECT 47.990 124.680 48.130 129.460 ;
        RECT 48.390 128.780 48.650 129.100 ;
        RECT 47.930 124.360 48.190 124.680 ;
        RECT 47.470 124.020 47.730 124.340 ;
        RECT 47.530 122.640 47.670 124.020 ;
        RECT 47.470 122.320 47.730 122.640 ;
        RECT 48.450 121.960 48.590 128.780 ;
        RECT 52.130 126.720 52.270 134.900 ;
        RECT 52.070 126.400 52.330 126.720 ;
        RECT 49.770 123.340 50.030 123.660 ;
        RECT 47.010 121.640 47.270 121.960 ;
        RECT 48.390 121.640 48.650 121.960 ;
        RECT 43.790 120.620 44.050 120.940 ;
        RECT 43.850 116.520 43.990 120.620 ;
        RECT 48.850 118.580 49.110 118.900 ;
        RECT 48.910 116.520 49.050 118.580 ;
        RECT 43.790 116.200 44.050 116.520 ;
        RECT 48.850 116.200 49.110 116.520 ;
        RECT 48.390 115.860 48.650 116.180 ;
        RECT 43.790 115.520 44.050 115.840 ;
        RECT 43.330 113.480 43.590 113.800 ;
        RECT 42.410 113.140 42.670 113.460 ;
        RECT 42.870 113.140 43.130 113.460 ;
        RECT 42.930 111.080 43.070 113.140 ;
        RECT 43.330 112.800 43.590 113.120 ;
        RECT 42.870 110.760 43.130 111.080 ;
        RECT 43.390 110.480 43.530 112.800 ;
        RECT 43.850 111.080 43.990 115.520 ;
        RECT 44.250 115.180 44.510 115.500 ;
        RECT 43.790 110.760 44.050 111.080 ;
        RECT 44.310 110.740 44.450 115.180 ;
        RECT 48.450 114.140 48.590 115.860 ;
        RECT 48.390 113.820 48.650 114.140 ;
        RECT 44.710 112.800 44.970 113.120 ;
        RECT 44.770 111.760 44.910 112.800 ;
        RECT 44.710 111.440 44.970 111.760 ;
        RECT 42.930 110.340 43.530 110.480 ;
        RECT 44.250 110.420 44.510 110.740 ;
        RECT 42.930 108.020 43.070 110.340 ;
        RECT 43.330 109.740 43.590 110.060 ;
        RECT 42.870 107.700 43.130 108.020 ;
        RECT 42.410 104.980 42.670 105.300 ;
        RECT 41.950 103.280 42.210 103.600 ;
        RECT 41.550 102.860 42.150 103.000 ;
        RECT 40.570 102.260 40.830 102.580 ;
        RECT 41.490 102.260 41.750 102.580 ;
        RECT 40.110 101.580 40.370 101.900 ;
        RECT 39.650 100.560 39.910 100.880 ;
        RECT 40.570 94.440 40.830 94.760 ;
        RECT 36.890 94.100 37.150 94.420 ;
        RECT 32.750 91.040 33.010 91.360 ;
        RECT 30.800 90.165 32.340 90.535 ;
        RECT 30.050 86.540 30.650 86.680 ;
        RECT 29.990 83.560 30.250 83.880 ;
        RECT 29.530 83.220 29.790 83.540 ;
        RECT 27.500 82.005 29.040 82.375 ;
        RECT 26.310 80.500 26.570 80.820 ;
        RECT 24.010 77.100 24.270 77.420 ;
        RECT 24.070 75.380 24.210 77.100 ;
        RECT 24.010 75.060 24.270 75.380 ;
        RECT 24.470 74.380 24.730 74.700 ;
        RECT 23.550 72.340 23.810 72.660 ;
        RECT 23.550 70.300 23.810 70.620 ;
        RECT 23.610 67.900 23.750 70.300 ;
        RECT 23.550 67.580 23.810 67.900 ;
        RECT 24.530 67.220 24.670 74.380 ;
        RECT 26.370 73.680 26.510 80.500 ;
        RECT 27.690 79.820 27.950 80.140 ;
        RECT 27.750 78.440 27.890 79.820 ;
        RECT 27.690 78.120 27.950 78.440 ;
        RECT 27.500 76.565 29.040 76.935 ;
        RECT 26.770 74.720 27.030 75.040 ;
        RECT 26.830 73.680 26.970 74.720 ;
        RECT 26.310 73.360 26.570 73.680 ;
        RECT 26.770 73.360 27.030 73.680 ;
        RECT 25.390 73.020 25.650 73.340 ;
        RECT 25.450 70.280 25.590 73.020 ;
        RECT 25.390 69.960 25.650 70.280 ;
        RECT 26.370 68.240 26.510 73.360 ;
        RECT 27.500 71.125 29.040 71.495 ;
        RECT 27.690 69.280 27.950 69.600 ;
        RECT 27.750 68.240 27.890 69.280 ;
        RECT 26.310 67.920 26.570 68.240 ;
        RECT 27.690 67.920 27.950 68.240 ;
        RECT 30.050 67.640 30.190 83.560 ;
        RECT 29.590 67.500 30.190 67.640 ;
        RECT 24.470 66.900 24.730 67.220 ;
        RECT 26.770 66.900 27.030 67.220 ;
        RECT 26.830 65.520 26.970 66.900 ;
        RECT 27.500 65.685 29.040 66.055 ;
        RECT 26.770 65.480 27.030 65.520 ;
        RECT 25.910 65.340 27.030 65.480 ;
        RECT 25.910 64.840 26.050 65.340 ;
        RECT 26.770 65.200 27.030 65.340 ;
        RECT 25.850 64.520 26.110 64.840 ;
        RECT 28.610 64.180 28.870 64.500 ;
        RECT 25.850 63.840 26.110 64.160 ;
        RECT 24.470 63.500 24.730 63.820 ;
        RECT 24.530 62.120 24.670 63.500 ;
        RECT 25.390 62.480 25.650 62.800 ;
        RECT 24.470 61.800 24.730 62.120 ;
        RECT 24.930 59.760 25.190 60.080 ;
        RECT 23.550 59.420 23.810 59.740 ;
        RECT 22.690 57.300 23.290 57.440 ;
        RECT 20.315 56.505 20.600 56.680 ;
        RECT 20.315 56.360 20.575 56.505 ;
        RECT 21.710 56.360 21.970 56.680 ;
        RECT 21.250 55.680 21.510 56.000 ;
        RECT 21.310 54.640 21.450 55.680 ;
        RECT 21.250 54.320 21.510 54.640 ;
        RECT 21.770 51.680 21.910 56.360 ;
        RECT 22.690 55.660 22.830 57.300 ;
        RECT 23.610 56.680 23.750 59.420 ;
        RECT 24.990 56.680 25.130 59.760 ;
        RECT 25.450 59.060 25.590 62.480 ;
        RECT 25.390 58.740 25.650 59.060 ;
        RECT 23.090 56.360 23.350 56.680 ;
        RECT 23.550 56.360 23.810 56.680 ;
        RECT 24.010 56.360 24.270 56.680 ;
        RECT 24.930 56.360 25.190 56.680 ;
        RECT 22.630 55.340 22.890 55.660 ;
        RECT 20.390 51.540 21.910 51.680 ;
        RECT 20.390 48.860 20.530 51.540 ;
        RECT 20.330 48.540 20.590 48.860 ;
        RECT 21.250 47.860 21.510 48.180 ;
        RECT 20.330 47.180 20.590 47.500 ;
        RECT 20.390 44.635 20.530 47.180 ;
        RECT 21.310 46.140 21.450 47.860 ;
        RECT 22.170 46.160 22.430 46.480 ;
        RECT 21.250 45.820 21.510 46.140 ;
        RECT 20.320 44.265 20.600 44.635 ;
        RECT 21.710 44.460 21.970 44.780 ;
        RECT 21.250 41.740 21.510 42.060 ;
        RECT 21.310 41.235 21.450 41.740 ;
        RECT 21.240 40.865 21.520 41.235 ;
        RECT 20.790 40.380 21.050 40.700 ;
        RECT 19.870 39.020 20.130 39.340 ;
        RECT 20.330 38.000 20.590 38.320 ;
        RECT 19.870 36.640 20.130 36.960 ;
        RECT 19.930 35.600 20.070 36.640 ;
        RECT 19.870 35.280 20.130 35.600 ;
        RECT 19.410 32.220 19.670 32.540 ;
        RECT 20.390 31.600 20.530 38.000 ;
        RECT 20.850 36.620 20.990 40.380 ;
        RECT 21.250 40.270 21.510 40.360 ;
        RECT 21.770 40.270 21.910 44.460 ;
        RECT 22.230 42.740 22.370 46.160 ;
        RECT 22.170 42.420 22.430 42.740 ;
        RECT 21.250 40.130 21.910 40.270 ;
        RECT 21.250 40.040 21.510 40.130 ;
        RECT 21.250 39.020 21.510 39.340 ;
        RECT 20.790 36.300 21.050 36.620 ;
        RECT 20.850 32.200 20.990 36.300 ;
        RECT 21.310 34.920 21.450 39.020 ;
        RECT 21.770 38.320 21.910 40.130 ;
        RECT 21.710 38.000 21.970 38.320 ;
        RECT 21.250 34.600 21.510 34.920 ;
        RECT 21.710 34.600 21.970 34.920 ;
        RECT 21.770 32.540 21.910 34.600 ;
        RECT 21.710 32.220 21.970 32.540 ;
        RECT 20.790 31.880 21.050 32.200 ;
        RECT 20.390 31.460 20.990 31.600 ;
        RECT 20.330 30.860 20.590 31.180 ;
        RECT 20.390 29.820 20.530 30.860 ;
        RECT 20.330 29.500 20.590 29.820 ;
        RECT 20.850 25.740 20.990 31.460 ;
        RECT 21.250 28.140 21.510 28.460 ;
        RECT 21.310 26.420 21.450 28.140 ;
        RECT 21.250 26.100 21.510 26.420 ;
        RECT 20.790 25.420 21.050 25.740 ;
        RECT 20.850 24.380 20.990 25.420 ;
        RECT 20.790 24.060 21.050 24.380 ;
        RECT 20.330 23.720 20.590 24.040 ;
        RECT 18.490 21.000 18.750 21.320 ;
        RECT 18.950 19.980 19.210 20.300 ;
        RECT 19.410 19.980 19.670 20.300 ;
        RECT 19.010 11.880 19.150 19.980 ;
        RECT 19.470 18.600 19.610 19.980 ;
        RECT 20.390 19.280 20.530 23.720 ;
        RECT 21.310 20.980 21.450 26.100 ;
        RECT 21.770 21.660 21.910 32.220 ;
        RECT 22.630 31.540 22.890 31.860 ;
        RECT 22.690 30.160 22.830 31.540 ;
        RECT 22.630 29.840 22.890 30.160 ;
        RECT 23.150 24.120 23.290 56.360 ;
        RECT 23.550 55.680 23.810 56.000 ;
        RECT 23.610 43.160 23.750 55.680 ;
        RECT 24.070 53.620 24.210 56.360 ;
        RECT 24.010 53.300 24.270 53.620 ;
        RECT 24.070 51.680 24.210 53.300 ;
        RECT 24.070 51.540 24.670 51.680 ;
        RECT 24.010 48.540 24.270 48.860 ;
        RECT 24.070 45.460 24.210 48.540 ;
        RECT 24.010 45.140 24.270 45.460 ;
        RECT 24.530 43.420 24.670 51.540 ;
        RECT 24.990 48.180 25.130 56.360 ;
        RECT 25.450 51.580 25.590 58.740 ;
        RECT 25.910 57.020 26.050 63.840 ;
        RECT 26.770 63.500 27.030 63.820 ;
        RECT 28.150 63.500 28.410 63.820 ;
        RECT 26.310 60.780 26.570 61.100 ;
        RECT 26.370 59.060 26.510 60.780 ;
        RECT 26.830 60.080 26.970 63.500 ;
        RECT 28.210 62.800 28.350 63.500 ;
        RECT 28.150 62.480 28.410 62.800 ;
        RECT 28.670 61.010 28.810 64.180 ;
        RECT 29.590 61.350 29.730 67.500 ;
        RECT 29.990 66.900 30.250 67.220 ;
        RECT 30.050 64.500 30.190 66.900 ;
        RECT 30.510 65.480 30.650 86.540 ;
        RECT 30.800 84.725 32.340 85.095 ;
        RECT 32.810 81.920 32.950 91.040 ;
        RECT 35.510 88.660 35.770 88.980 ;
        RECT 33.210 85.260 33.470 85.580 ;
        RECT 33.270 83.880 33.410 85.260 ;
        RECT 33.210 83.560 33.470 83.880 ;
        RECT 33.270 82.860 33.410 83.560 ;
        RECT 33.210 82.540 33.470 82.860 ;
        RECT 32.810 81.780 33.410 81.920 ;
        RECT 30.800 79.285 32.340 79.655 ;
        RECT 30.800 73.845 32.340 74.215 ;
        RECT 32.750 68.940 33.010 69.260 ;
        RECT 30.800 68.405 32.340 68.775 ;
        RECT 32.810 65.520 32.950 68.940 ;
        RECT 30.510 65.340 32.490 65.480 ;
        RECT 29.990 64.180 30.250 64.500 ;
        RECT 30.050 62.800 30.190 64.180 ;
        RECT 32.350 64.070 32.490 65.340 ;
        RECT 32.750 65.200 33.010 65.520 ;
        RECT 33.270 65.480 33.410 81.780 ;
        RECT 34.130 81.180 34.390 81.500 ;
        RECT 34.190 80.140 34.330 81.180 ;
        RECT 34.130 79.820 34.390 80.140 ;
        RECT 34.190 79.120 34.330 79.820 ;
        RECT 34.130 78.800 34.390 79.120 ;
        RECT 33.270 65.340 33.870 65.480 ;
        RECT 33.210 64.860 33.470 65.180 ;
        RECT 32.350 63.930 32.950 64.070 ;
        RECT 30.450 63.500 30.710 63.820 ;
        RECT 29.990 62.480 30.250 62.800 ;
        RECT 29.590 61.210 30.190 61.350 ;
        RECT 28.670 60.870 29.730 61.010 ;
        RECT 27.500 60.245 29.040 60.615 ;
        RECT 26.770 59.760 27.030 60.080 ;
        RECT 29.590 59.740 29.730 60.870 ;
        RECT 29.530 59.420 29.790 59.740 ;
        RECT 26.310 58.740 26.570 59.060 ;
        RECT 27.690 58.400 27.950 58.720 ;
        RECT 27.230 58.060 27.490 58.380 ;
        RECT 25.850 56.700 26.110 57.020 ;
        RECT 27.290 56.680 27.430 58.060 ;
        RECT 27.750 57.020 27.890 58.400 ;
        RECT 30.050 58.380 30.190 61.210 ;
        RECT 30.510 59.400 30.650 63.500 ;
        RECT 30.800 62.965 32.340 63.335 ;
        RECT 30.910 62.140 31.170 62.460 ;
        RECT 30.450 59.080 30.710 59.400 ;
        RECT 30.970 59.060 31.110 62.140 ;
        RECT 31.830 61.800 32.090 62.120 ;
        RECT 31.890 60.080 32.030 61.800 ;
        RECT 31.830 59.760 32.090 60.080 ;
        RECT 30.910 58.740 31.170 59.060 ;
        RECT 29.990 58.060 30.250 58.380 ;
        RECT 30.800 57.525 32.340 57.895 ;
        RECT 27.690 56.700 27.950 57.020 ;
        RECT 27.230 56.590 27.490 56.680 ;
        RECT 26.830 56.450 27.490 56.590 ;
        RECT 26.830 51.920 26.970 56.450 ;
        RECT 27.230 56.360 27.490 56.450 ;
        RECT 29.530 56.360 29.790 56.680 ;
        RECT 27.500 54.805 29.040 55.175 ;
        RECT 27.230 52.960 27.490 53.280 ;
        RECT 26.770 51.600 27.030 51.920 ;
        RECT 25.390 51.260 25.650 51.580 ;
        RECT 25.450 48.600 25.590 51.260 ;
        RECT 27.290 50.900 27.430 52.960 ;
        RECT 29.590 50.900 29.730 56.360 ;
        RECT 29.990 55.340 30.250 55.660 ;
        RECT 30.050 50.900 30.190 55.340 ;
        RECT 30.910 53.360 31.170 53.620 ;
        RECT 30.510 53.300 31.170 53.360 ;
        RECT 30.510 53.220 31.110 53.300 ;
        RECT 27.230 50.580 27.490 50.900 ;
        RECT 29.530 50.580 29.790 50.900 ;
        RECT 29.990 50.580 30.250 50.900 ;
        RECT 26.770 49.900 27.030 50.220 ;
        RECT 25.450 48.460 26.050 48.600 ;
        RECT 24.930 47.860 25.190 48.180 ;
        RECT 23.610 43.020 24.210 43.160 ;
        RECT 24.470 43.100 24.730 43.420 ;
        RECT 23.550 42.420 23.810 42.740 ;
        RECT 23.610 27.440 23.750 42.420 ;
        RECT 24.070 32.280 24.210 43.020 ;
        RECT 24.990 40.020 25.130 47.860 ;
        RECT 25.910 45.800 26.050 48.460 ;
        RECT 26.830 48.180 26.970 49.900 ;
        RECT 27.500 49.365 29.040 49.735 ;
        RECT 28.610 48.880 28.870 49.200 ;
        RECT 28.150 48.200 28.410 48.520 ;
        RECT 26.770 47.860 27.030 48.180 ;
        RECT 28.210 45.800 28.350 48.200 ;
        RECT 28.670 45.800 28.810 48.880 ;
        RECT 29.590 48.520 29.730 50.580 ;
        RECT 29.530 48.200 29.790 48.520 ;
        RECT 29.990 47.860 30.250 48.180 ;
        RECT 25.850 45.480 26.110 45.800 ;
        RECT 28.150 45.480 28.410 45.800 ;
        RECT 28.610 45.480 28.870 45.800 ;
        RECT 25.390 45.140 25.650 45.460 ;
        RECT 24.930 39.700 25.190 40.020 ;
        RECT 25.450 37.300 25.590 45.140 ;
        RECT 25.910 43.670 26.050 45.480 ;
        RECT 29.530 45.140 29.790 45.460 ;
        RECT 27.500 43.925 29.040 44.295 ;
        RECT 29.590 43.760 29.730 45.140 ;
        RECT 25.910 43.530 27.430 43.670 ;
        RECT 26.310 42.420 26.570 42.740 ;
        RECT 25.390 36.980 25.650 37.300 ;
        RECT 25.390 36.300 25.650 36.620 ;
        RECT 25.450 35.260 25.590 36.300 ;
        RECT 25.390 34.940 25.650 35.260 ;
        RECT 25.850 33.580 26.110 33.900 ;
        RECT 24.070 32.140 24.670 32.280 ;
        RECT 24.010 31.540 24.270 31.860 ;
        RECT 24.070 29.480 24.210 31.540 ;
        RECT 24.010 29.160 24.270 29.480 ;
        RECT 23.550 27.120 23.810 27.440 ;
        RECT 24.010 26.100 24.270 26.420 ;
        RECT 24.070 24.235 24.210 26.100 ;
        RECT 23.150 23.980 23.750 24.120 ;
        RECT 22.170 23.040 22.430 23.360 ;
        RECT 23.090 23.040 23.350 23.360 ;
        RECT 21.710 21.340 21.970 21.660 ;
        RECT 21.250 20.660 21.510 20.980 ;
        RECT 20.330 18.960 20.590 19.280 ;
        RECT 19.410 18.280 19.670 18.600 ;
        RECT 20.390 16.560 20.530 18.960 ;
        RECT 22.230 18.600 22.370 23.040 ;
        RECT 22.630 20.660 22.890 20.980 ;
        RECT 22.170 18.280 22.430 18.600 ;
        RECT 22.690 16.560 22.830 20.660 ;
        RECT 20.330 16.240 20.590 16.560 ;
        RECT 22.630 16.240 22.890 16.560 ;
        RECT 23.150 13.240 23.290 23.040 ;
        RECT 23.610 23.020 23.750 23.980 ;
        RECT 24.000 23.865 24.280 24.235 ;
        RECT 24.010 23.720 24.270 23.865 ;
        RECT 23.550 22.700 23.810 23.020 ;
        RECT 24.530 22.000 24.670 32.140 ;
        RECT 25.910 31.860 26.050 33.580 ;
        RECT 25.850 31.540 26.110 31.860 ;
        RECT 25.910 30.160 26.050 31.540 ;
        RECT 25.850 29.840 26.110 30.160 ;
        RECT 24.930 23.720 25.190 24.040 ;
        RECT 24.470 21.680 24.730 22.000 ;
        RECT 24.990 17.580 25.130 23.720 ;
        RECT 25.910 20.980 26.050 29.840 ;
        RECT 26.370 27.440 26.510 42.420 ;
        RECT 27.290 40.700 27.430 43.530 ;
        RECT 29.530 43.440 29.790 43.760 ;
        RECT 29.070 42.760 29.330 43.080 ;
        RECT 27.690 42.420 27.950 42.740 ;
        RECT 27.230 40.380 27.490 40.700 ;
        RECT 27.750 40.360 27.890 42.420 ;
        RECT 29.130 40.700 29.270 42.760 ;
        RECT 29.530 42.080 29.790 42.400 ;
        RECT 29.070 40.380 29.330 40.700 ;
        RECT 29.590 40.360 29.730 42.080 ;
        RECT 27.690 40.040 27.950 40.360 ;
        RECT 29.530 40.040 29.790 40.360 ;
        RECT 29.530 39.020 29.790 39.340 ;
        RECT 27.500 38.485 29.040 38.855 ;
        RECT 28.610 36.980 28.870 37.300 ;
        RECT 29.070 36.980 29.330 37.300 ;
        RECT 27.230 36.640 27.490 36.960 ;
        RECT 27.290 34.920 27.430 36.640 ;
        RECT 28.670 35.260 28.810 36.980 ;
        RECT 29.130 35.600 29.270 36.980 ;
        RECT 29.590 36.620 29.730 39.020 ;
        RECT 30.050 37.210 30.190 47.860 ;
        RECT 30.510 41.040 30.650 53.220 ;
        RECT 30.800 52.085 32.340 52.455 ;
        RECT 31.830 51.600 32.090 51.920 ;
        RECT 32.290 51.600 32.550 51.920 ;
        RECT 31.890 47.840 32.030 51.600 ;
        RECT 32.350 48.035 32.490 51.600 ;
        RECT 31.830 47.520 32.090 47.840 ;
        RECT 32.280 47.665 32.560 48.035 ;
        RECT 30.800 46.645 32.340 47.015 ;
        RECT 32.810 42.740 32.950 63.930 ;
        RECT 33.270 55.570 33.410 64.860 ;
        RECT 33.730 56.080 33.870 65.340 ;
        RECT 34.190 62.460 34.330 78.800 ;
        RECT 35.050 68.940 35.310 69.260 ;
        RECT 35.110 64.160 35.250 68.940 ;
        RECT 35.050 63.840 35.310 64.160 ;
        RECT 34.130 62.370 34.390 62.460 ;
        RECT 34.130 62.230 34.790 62.370 ;
        RECT 34.130 62.140 34.390 62.230 ;
        RECT 34.130 60.780 34.390 61.100 ;
        RECT 34.190 57.020 34.330 60.780 ;
        RECT 34.130 56.700 34.390 57.020 ;
        RECT 33.730 55.940 34.330 56.080 ;
        RECT 33.670 55.570 33.930 55.660 ;
        RECT 33.270 55.430 33.930 55.570 ;
        RECT 33.270 53.280 33.410 55.430 ;
        RECT 33.670 55.340 33.930 55.430 ;
        RECT 34.190 54.720 34.330 55.940 ;
        RECT 33.730 54.580 34.330 54.720 ;
        RECT 33.210 52.960 33.470 53.280 ;
        RECT 33.270 51.240 33.410 52.960 ;
        RECT 33.210 50.920 33.470 51.240 ;
        RECT 33.730 48.180 33.870 54.580 ;
        RECT 34.650 51.920 34.790 62.230 ;
        RECT 35.570 57.360 35.710 88.660 ;
        RECT 36.950 81.160 37.090 94.100 ;
        RECT 40.630 92.040 40.770 94.440 ;
        RECT 37.350 91.720 37.610 92.040 ;
        RECT 40.570 91.720 40.830 92.040 ;
        RECT 37.410 90.000 37.550 91.720 ;
        RECT 40.110 90.700 40.370 91.020 ;
        RECT 40.170 90.000 40.310 90.700 ;
        RECT 41.550 90.000 41.690 102.260 ;
        RECT 42.010 99.980 42.150 102.860 ;
        RECT 42.470 100.540 42.610 104.980 ;
        RECT 42.410 100.220 42.670 100.540 ;
        RECT 42.930 99.980 43.070 107.700 ;
        RECT 43.390 102.920 43.530 109.740 ;
        RECT 43.790 107.700 44.050 108.020 ;
        RECT 44.250 107.700 44.510 108.020 ;
        RECT 43.850 106.320 43.990 107.700 ;
        RECT 43.790 106.000 44.050 106.320 ;
        RECT 43.330 102.600 43.590 102.920 ;
        RECT 43.850 102.580 43.990 106.000 ;
        RECT 44.310 102.580 44.450 107.700 ;
        RECT 45.630 107.360 45.890 107.680 ;
        RECT 48.390 107.360 48.650 107.680 ;
        RECT 45.170 105.320 45.430 105.640 ;
        RECT 45.230 103.600 45.370 105.320 ;
        RECT 45.170 103.280 45.430 103.600 ;
        RECT 43.790 102.260 44.050 102.580 ;
        RECT 44.250 102.260 44.510 102.580 ;
        RECT 43.850 99.980 43.990 102.260 ;
        RECT 42.010 99.840 43.070 99.980 ;
        RECT 42.930 95.100 43.070 99.840 ;
        RECT 43.390 99.840 43.990 99.980 ;
        RECT 44.710 99.880 44.970 100.200 ;
        RECT 42.870 94.780 43.130 95.100 ;
        RECT 37.350 89.680 37.610 90.000 ;
        RECT 40.110 89.680 40.370 90.000 ;
        RECT 41.490 89.680 41.750 90.000 ;
        RECT 42.930 89.320 43.070 94.780 ;
        RECT 43.390 93.650 43.530 99.840 ;
        RECT 43.790 97.160 44.050 97.480 ;
        RECT 43.850 95.440 43.990 97.160 ;
        RECT 43.790 95.120 44.050 95.440 ;
        RECT 43.790 93.650 44.050 93.740 ;
        RECT 43.390 93.510 44.050 93.650 ;
        RECT 43.790 93.420 44.050 93.510 ;
        RECT 42.870 89.000 43.130 89.320 ;
        RECT 42.930 86.940 43.070 89.000 ;
        RECT 43.850 87.280 43.990 93.420 ;
        RECT 43.790 86.960 44.050 87.280 ;
        RECT 42.870 86.620 43.130 86.940 ;
        RECT 44.250 85.600 44.510 85.920 ;
        RECT 38.730 85.260 38.990 85.580 ;
        RECT 38.790 81.160 38.930 85.260 ;
        RECT 44.310 84.560 44.450 85.600 ;
        RECT 44.250 84.240 44.510 84.560 ;
        RECT 41.030 83.900 41.290 84.220 ;
        RECT 39.650 83.560 39.910 83.880 ;
        RECT 39.710 81.840 39.850 83.560 ;
        RECT 39.650 81.520 39.910 81.840 ;
        RECT 36.890 80.840 37.150 81.160 ;
        RECT 38.730 80.840 38.990 81.160 ;
        RECT 40.570 80.500 40.830 80.820 ;
        RECT 39.650 78.120 39.910 78.440 ;
        RECT 39.710 76.400 39.850 78.120 ;
        RECT 39.650 76.080 39.910 76.400 ;
        RECT 40.630 76.060 40.770 80.500 ;
        RECT 41.090 78.780 41.230 83.900 ;
        RECT 44.770 81.160 44.910 99.880 ;
        RECT 45.690 99.520 45.830 107.360 ;
        RECT 48.450 104.620 48.590 107.360 ;
        RECT 49.310 107.020 49.570 107.340 ;
        RECT 48.390 104.300 48.650 104.620 ;
        RECT 49.370 103.600 49.510 107.020 ;
        RECT 49.310 103.280 49.570 103.600 ;
        RECT 47.470 100.220 47.730 100.540 ;
        RECT 47.010 99.880 47.270 100.200 ;
        RECT 45.630 99.200 45.890 99.520 ;
        RECT 45.690 91.360 45.830 99.200 ;
        RECT 47.070 98.160 47.210 99.880 ;
        RECT 47.010 97.840 47.270 98.160 ;
        RECT 47.010 93.420 47.270 93.740 ;
        RECT 47.070 91.700 47.210 93.420 ;
        RECT 47.010 91.380 47.270 91.700 ;
        RECT 45.630 91.040 45.890 91.360 ;
        RECT 45.170 85.260 45.430 85.580 ;
        RECT 45.230 83.540 45.370 85.260 ;
        RECT 45.690 83.880 45.830 91.040 ;
        RECT 46.550 89.000 46.810 89.320 ;
        RECT 46.610 84.560 46.750 89.000 ;
        RECT 47.010 86.620 47.270 86.940 ;
        RECT 46.550 84.240 46.810 84.560 ;
        RECT 45.630 83.560 45.890 83.880 ;
        RECT 45.170 83.220 45.430 83.540 ;
        RECT 47.070 81.160 47.210 86.620 ;
        RECT 47.530 84.220 47.670 100.220 ;
        RECT 49.310 97.500 49.570 97.820 ;
        RECT 47.930 92.400 48.190 92.720 ;
        RECT 47.990 90.000 48.130 92.400 ;
        RECT 48.390 90.700 48.650 91.020 ;
        RECT 47.930 89.680 48.190 90.000 ;
        RECT 48.450 89.320 48.590 90.700 ;
        RECT 48.390 89.000 48.650 89.320 ;
        RECT 47.930 88.320 48.190 88.640 ;
        RECT 47.990 86.940 48.130 88.320 ;
        RECT 48.850 87.980 49.110 88.300 ;
        RECT 48.910 87.280 49.050 87.980 ;
        RECT 48.850 86.960 49.110 87.280 ;
        RECT 47.930 86.620 48.190 86.940 ;
        RECT 48.910 85.920 49.050 86.960 ;
        RECT 48.850 85.600 49.110 85.920 ;
        RECT 47.930 85.260 48.190 85.580 ;
        RECT 47.990 84.220 48.130 85.260 ;
        RECT 47.470 83.900 47.730 84.220 ;
        RECT 47.930 83.900 48.190 84.220 ;
        RECT 47.530 83.540 47.670 83.900 ;
        RECT 47.470 83.220 47.730 83.540 ;
        RECT 47.930 82.540 48.190 82.860 ;
        RECT 47.990 81.840 48.130 82.540 ;
        RECT 47.930 81.520 48.190 81.840 ;
        RECT 44.710 80.840 44.970 81.160 ;
        RECT 47.010 80.840 47.270 81.160 ;
        RECT 41.490 79.820 41.750 80.140 ;
        RECT 43.330 79.820 43.590 80.140 ;
        RECT 41.030 78.460 41.290 78.780 ;
        RECT 40.570 75.740 40.830 76.060 ;
        RECT 41.090 75.380 41.230 78.460 ;
        RECT 41.030 75.060 41.290 75.380 ;
        RECT 36.430 74.720 36.690 75.040 ;
        RECT 36.490 72.660 36.630 74.720 ;
        RECT 41.090 73.340 41.230 75.060 ;
        RECT 38.270 73.020 38.530 73.340 ;
        RECT 39.650 73.020 39.910 73.340 ;
        RECT 41.030 73.020 41.290 73.340 ;
        RECT 36.430 72.340 36.690 72.660 ;
        RECT 35.510 57.040 35.770 57.360 ;
        RECT 34.590 51.600 34.850 51.920 ;
        RECT 35.970 49.110 36.230 49.200 ;
        RECT 36.490 49.110 36.630 72.340 ;
        RECT 36.890 68.940 37.150 69.260 ;
        RECT 37.350 68.940 37.610 69.260 ;
        RECT 36.950 68.240 37.090 68.940 ;
        RECT 36.890 67.920 37.150 68.240 ;
        RECT 37.410 65.480 37.550 68.940 ;
        RECT 35.970 48.970 36.630 49.110 ;
        RECT 35.970 48.880 36.230 48.970 ;
        RECT 33.670 47.860 33.930 48.180 ;
        RECT 33.210 47.520 33.470 47.840 ;
        RECT 33.270 43.670 33.410 47.520 ;
        RECT 33.270 43.530 33.870 43.670 ;
        RECT 33.210 42.760 33.470 43.080 ;
        RECT 32.750 42.420 33.010 42.740 ;
        RECT 30.800 41.205 32.340 41.575 ;
        RECT 30.450 40.720 30.710 41.040 ;
        RECT 33.270 40.360 33.410 42.760 ;
        RECT 33.730 40.440 33.870 43.530 ;
        RECT 36.490 42.740 36.630 48.970 ;
        RECT 36.950 65.340 37.550 65.480 ;
        RECT 36.950 43.420 37.090 65.340 ;
        RECT 37.810 58.400 38.070 58.720 ;
        RECT 37.870 57.360 38.010 58.400 ;
        RECT 37.810 57.040 38.070 57.360 ;
        RECT 38.330 51.580 38.470 73.020 ;
        RECT 39.710 69.940 39.850 73.020 ;
        RECT 39.650 69.620 39.910 69.940 ;
        RECT 39.190 65.200 39.450 65.520 ;
        RECT 39.250 59.740 39.390 65.200 ;
        RECT 39.710 64.500 39.850 69.620 ;
        RECT 39.650 64.180 39.910 64.500 ;
        RECT 39.710 62.120 39.850 64.180 ;
        RECT 39.650 61.800 39.910 62.120 ;
        RECT 39.190 59.420 39.450 59.740 ;
        RECT 39.710 59.060 39.850 61.800 ;
        RECT 41.550 60.080 41.690 79.820 ;
        RECT 43.390 75.720 43.530 79.820 ;
        RECT 44.770 79.120 44.910 80.840 ;
        RECT 47.070 79.120 47.210 80.840 ;
        RECT 44.710 78.800 44.970 79.120 ;
        RECT 47.010 78.800 47.270 79.120 ;
        RECT 43.330 75.400 43.590 75.720 ;
        RECT 46.090 75.060 46.350 75.380 ;
        RECT 41.950 67.920 42.210 68.240 ;
        RECT 42.010 67.560 42.150 67.920 ;
        RECT 41.950 67.240 42.210 67.560 ;
        RECT 42.410 67.240 42.670 67.560 ;
        RECT 43.330 67.240 43.590 67.560 ;
        RECT 42.010 65.520 42.150 67.240 ;
        RECT 42.470 66.395 42.610 67.240 ;
        RECT 42.400 66.025 42.680 66.395 ;
        RECT 41.950 65.200 42.210 65.520 ;
        RECT 43.390 65.480 43.530 67.240 ;
        RECT 46.150 66.540 46.290 75.060 ;
        RECT 47.010 74.380 47.270 74.700 ;
        RECT 47.070 68.240 47.210 74.380 ;
        RECT 47.470 69.620 47.730 69.940 ;
        RECT 47.010 67.920 47.270 68.240 ;
        RECT 47.010 66.900 47.270 67.220 ;
        RECT 46.090 66.220 46.350 66.540 ;
        RECT 43.390 65.340 45.370 65.480 ;
        RECT 43.330 63.500 43.590 63.820 ;
        RECT 43.390 62.460 43.530 63.500 ;
        RECT 43.330 62.140 43.590 62.460 ;
        RECT 41.490 59.760 41.750 60.080 ;
        RECT 39.650 58.740 39.910 59.060 ;
        RECT 42.870 58.060 43.130 58.380 ;
        RECT 42.930 56.680 43.070 58.060 ;
        RECT 42.870 56.360 43.130 56.680 ;
        RECT 40.570 56.020 40.830 56.340 ;
        RECT 40.630 54.640 40.770 56.020 ;
        RECT 40.570 54.320 40.830 54.640 ;
        RECT 38.270 51.260 38.530 51.580 ;
        RECT 37.350 46.160 37.610 46.480 ;
        RECT 37.410 45.120 37.550 46.160 ;
        RECT 38.330 46.140 38.470 51.260 ;
        RECT 39.650 50.920 39.910 51.240 ;
        RECT 40.110 50.920 40.370 51.240 ;
        RECT 41.030 51.150 41.290 51.240 ;
        RECT 41.030 51.010 41.690 51.150 ;
        RECT 41.030 50.920 41.290 51.010 ;
        RECT 38.730 47.520 38.990 47.840 ;
        RECT 38.270 45.820 38.530 46.140 ;
        RECT 37.350 44.800 37.610 45.120 ;
        RECT 36.890 43.100 37.150 43.420 ;
        RECT 36.430 42.650 36.690 42.740 ;
        RECT 36.030 42.510 36.690 42.650 ;
        RECT 33.210 40.040 33.470 40.360 ;
        RECT 33.730 40.300 34.330 40.440 ;
        RECT 33.270 37.720 33.410 40.040 ;
        RECT 33.670 39.700 33.930 40.020 ;
        RECT 32.810 37.580 33.410 37.720 ;
        RECT 32.810 37.300 32.950 37.580 ;
        RECT 33.730 37.300 33.870 39.700 ;
        RECT 30.450 37.210 30.710 37.300 ;
        RECT 30.050 37.070 30.710 37.210 ;
        RECT 30.450 36.980 30.710 37.070 ;
        RECT 32.750 36.980 33.010 37.300 ;
        RECT 33.210 36.980 33.470 37.300 ;
        RECT 33.670 36.980 33.930 37.300 ;
        RECT 29.530 36.300 29.790 36.620 ;
        RECT 29.990 36.300 30.250 36.620 ;
        RECT 29.070 35.280 29.330 35.600 ;
        RECT 29.530 35.280 29.790 35.600 ;
        RECT 28.610 35.000 28.870 35.260 ;
        RECT 29.590 35.000 29.730 35.280 ;
        RECT 28.610 34.940 29.730 35.000 ;
        RECT 27.230 34.600 27.490 34.920 ;
        RECT 28.670 34.860 29.730 34.940 ;
        RECT 30.050 34.920 30.190 36.300 ;
        RECT 30.800 35.765 32.340 36.135 ;
        RECT 32.750 35.280 33.010 35.600 ;
        RECT 29.990 34.600 30.250 34.920 ;
        RECT 27.290 34.320 27.430 34.600 ;
        RECT 26.830 34.180 27.430 34.320 ;
        RECT 26.830 29.480 26.970 34.180 ;
        RECT 30.450 33.580 30.710 33.900 ;
        RECT 27.500 33.045 29.040 33.415 ;
        RECT 26.770 29.160 27.030 29.480 ;
        RECT 29.990 29.160 30.250 29.480 ;
        RECT 26.310 27.120 26.570 27.440 ;
        RECT 26.830 26.840 26.970 29.160 ;
        RECT 29.530 28.140 29.790 28.460 ;
        RECT 27.500 27.605 29.040 27.975 ;
        RECT 26.370 26.700 26.970 26.840 ;
        RECT 26.370 24.380 26.510 26.700 ;
        RECT 29.590 26.420 29.730 28.140 ;
        RECT 26.770 26.100 27.030 26.420 ;
        RECT 29.530 26.100 29.790 26.420 ;
        RECT 26.310 24.060 26.570 24.380 ;
        RECT 25.850 20.660 26.110 20.980 ;
        RECT 25.850 18.280 26.110 18.600 ;
        RECT 25.910 18.000 26.050 18.280 ;
        RECT 26.370 18.000 26.510 24.060 ;
        RECT 26.830 18.600 26.970 26.100 ;
        RECT 29.530 25.420 29.790 25.740 ;
        RECT 29.590 24.380 29.730 25.420 ;
        RECT 30.050 24.720 30.190 29.160 ;
        RECT 29.990 24.400 30.250 24.720 ;
        RECT 29.530 24.060 29.790 24.380 ;
        RECT 30.510 24.120 30.650 33.580 ;
        RECT 30.800 30.325 32.340 30.695 ;
        RECT 32.290 29.390 32.550 29.480 ;
        RECT 32.810 29.390 32.950 35.280 ;
        RECT 33.270 32.200 33.410 36.980 ;
        RECT 33.670 34.940 33.930 35.260 ;
        RECT 33.210 31.880 33.470 32.200 ;
        RECT 33.270 29.480 33.410 31.880 ;
        RECT 32.290 29.250 32.950 29.390 ;
        RECT 32.290 29.160 32.550 29.250 ;
        RECT 30.800 24.885 32.340 25.255 ;
        RECT 27.500 22.165 29.040 22.535 ;
        RECT 27.680 21.145 27.960 21.515 ;
        RECT 27.750 20.980 27.890 21.145 ;
        RECT 27.690 20.660 27.950 20.980 ;
        RECT 27.230 19.980 27.490 20.300 ;
        RECT 29.070 19.980 29.330 20.300 ;
        RECT 27.290 19.280 27.430 19.980 ;
        RECT 27.230 18.960 27.490 19.280 ;
        RECT 29.130 18.940 29.270 19.980 ;
        RECT 29.070 18.620 29.330 18.940 ;
        RECT 26.770 18.280 27.030 18.600 ;
        RECT 25.910 17.920 26.970 18.000 ;
        RECT 25.910 17.860 27.030 17.920 ;
        RECT 24.930 17.260 25.190 17.580 ;
        RECT 24.990 15.540 25.130 17.260 ;
        RECT 25.910 17.180 26.050 17.860 ;
        RECT 26.770 17.600 27.030 17.860 ;
        RECT 25.450 17.040 26.050 17.180 ;
        RECT 24.930 15.220 25.190 15.540 ;
        RECT 25.450 15.200 25.590 17.040 ;
        RECT 27.500 16.725 29.040 17.095 ;
        RECT 29.590 15.540 29.730 24.060 ;
        RECT 30.050 23.980 30.650 24.120 ;
        RECT 30.050 15.540 30.190 23.980 ;
        RECT 30.450 20.660 30.710 20.980 ;
        RECT 31.370 20.660 31.630 20.980 ;
        RECT 30.510 19.280 30.650 20.660 ;
        RECT 31.430 20.300 31.570 20.660 ;
        RECT 32.290 20.550 32.550 20.640 ;
        RECT 32.810 20.550 32.950 29.250 ;
        RECT 33.210 29.160 33.470 29.480 ;
        RECT 33.730 28.200 33.870 34.940 ;
        RECT 34.190 29.480 34.330 40.300 ;
        RECT 34.130 29.390 34.390 29.480 ;
        RECT 34.130 29.250 34.790 29.390 ;
        RECT 34.130 29.160 34.390 29.250 ;
        RECT 34.130 28.480 34.390 28.800 ;
        RECT 34.190 28.200 34.330 28.480 ;
        RECT 33.730 28.060 34.330 28.200 ;
        RECT 33.730 26.160 33.870 28.060 ;
        RECT 34.130 26.160 34.390 26.420 ;
        RECT 33.730 26.100 34.390 26.160 ;
        RECT 33.730 26.020 34.330 26.100 ;
        RECT 33.730 20.980 33.870 26.020 ;
        RECT 34.650 25.740 34.790 29.250 ;
        RECT 35.510 29.160 35.770 29.480 ;
        RECT 35.050 28.140 35.310 28.460 ;
        RECT 35.110 26.080 35.250 28.140 ;
        RECT 35.050 25.760 35.310 26.080 ;
        RECT 34.590 25.420 34.850 25.740 ;
        RECT 33.670 20.660 33.930 20.980 ;
        RECT 32.290 20.410 32.950 20.550 ;
        RECT 32.290 20.320 32.550 20.410 ;
        RECT 31.370 19.980 31.630 20.300 ;
        RECT 30.800 19.445 32.340 19.815 ;
        RECT 30.450 18.960 30.710 19.280 ;
        RECT 33.670 18.620 33.930 18.940 ;
        RECT 33.730 15.540 33.870 18.620 ;
        RECT 35.570 18.260 35.710 29.160 ;
        RECT 36.030 28.800 36.170 42.510 ;
        RECT 36.430 42.420 36.690 42.510 ;
        RECT 37.410 40.700 37.550 44.800 ;
        RECT 38.790 43.760 38.930 47.520 ;
        RECT 39.710 47.500 39.850 50.920 ;
        RECT 40.170 50.560 40.310 50.920 ;
        RECT 40.110 50.240 40.370 50.560 ;
        RECT 41.030 50.240 41.290 50.560 ;
        RECT 40.170 49.200 40.310 50.240 ;
        RECT 40.110 48.880 40.370 49.200 ;
        RECT 41.090 48.180 41.230 50.240 ;
        RECT 41.030 47.860 41.290 48.180 ;
        RECT 39.650 47.180 39.910 47.500 ;
        RECT 40.110 45.820 40.370 46.140 ;
        RECT 38.730 43.440 38.990 43.760 ;
        RECT 40.170 42.740 40.310 45.820 ;
        RECT 41.090 45.800 41.230 47.860 ;
        RECT 41.030 45.480 41.290 45.800 ;
        RECT 40.110 42.420 40.370 42.740 ;
        RECT 37.350 40.380 37.610 40.700 ;
        RECT 39.190 36.980 39.450 37.300 ;
        RECT 36.430 36.300 36.690 36.620 ;
        RECT 36.490 35.260 36.630 36.300 ;
        RECT 36.430 34.940 36.690 35.260 ;
        RECT 35.970 28.480 36.230 28.800 ;
        RECT 36.030 26.080 36.170 28.480 ;
        RECT 35.970 25.760 36.230 26.080 ;
        RECT 35.510 17.940 35.770 18.260 ;
        RECT 35.510 15.900 35.770 16.220 ;
        RECT 29.530 15.220 29.790 15.540 ;
        RECT 29.990 15.220 30.250 15.540 ;
        RECT 33.670 15.220 33.930 15.540 ;
        RECT 25.390 14.880 25.650 15.200 ;
        RECT 25.850 14.540 26.110 14.860 ;
        RECT 29.070 14.540 29.330 14.860 ;
        RECT 32.290 14.770 32.550 14.860 ;
        RECT 32.290 14.630 32.950 14.770 ;
        RECT 32.290 14.540 32.550 14.630 ;
        RECT 22.690 13.100 23.290 13.240 ;
        RECT 19.010 11.740 19.610 11.880 ;
        RECT 18.030 9.440 18.290 9.760 ;
        RECT 19.470 7.310 19.610 11.740 ;
        RECT 22.690 7.310 22.830 13.100 ;
        RECT 25.910 7.310 26.050 14.540 ;
        RECT 29.130 7.310 29.270 14.540 ;
        RECT 30.800 14.005 32.340 14.375 ;
        RECT 32.810 9.160 32.950 14.630 ;
        RECT 32.350 9.020 32.950 9.160 ;
        RECT 32.350 7.310 32.490 9.020 ;
        RECT 35.570 7.310 35.710 15.900 ;
        RECT 36.490 15.540 36.630 34.940 ;
        RECT 39.250 34.920 39.390 36.980 ;
        RECT 41.030 36.640 41.290 36.960 ;
        RECT 39.190 34.600 39.450 34.920 ;
        RECT 39.250 24.380 39.390 34.600 ;
        RECT 40.570 29.500 40.830 29.820 ;
        RECT 40.630 26.080 40.770 29.500 ;
        RECT 41.090 29.140 41.230 36.640 ;
        RECT 41.550 35.600 41.690 51.010 ;
        RECT 42.870 50.920 43.130 51.240 ;
        RECT 43.790 50.920 44.050 51.240 ;
        RECT 42.930 48.860 43.070 50.920 ;
        RECT 43.850 49.200 43.990 50.920 ;
        RECT 43.790 48.880 44.050 49.200 ;
        RECT 42.870 48.540 43.130 48.860 ;
        RECT 43.790 47.180 44.050 47.500 ;
        RECT 43.850 45.800 43.990 47.180 ;
        RECT 43.790 45.480 44.050 45.800 ;
        RECT 43.330 45.140 43.590 45.460 ;
        RECT 43.390 42.740 43.530 45.140 ;
        RECT 43.330 42.420 43.590 42.740 ;
        RECT 42.410 40.270 42.670 40.360 ;
        RECT 42.410 40.130 43.070 40.270 ;
        RECT 42.410 40.040 42.670 40.130 ;
        RECT 41.490 35.280 41.750 35.600 ;
        RECT 41.490 34.600 41.750 34.920 ;
        RECT 41.550 32.540 41.690 34.600 ;
        RECT 41.950 34.260 42.210 34.580 ;
        RECT 41.490 32.220 41.750 32.540 ;
        RECT 41.490 31.540 41.750 31.860 ;
        RECT 41.550 29.480 41.690 31.540 ;
        RECT 41.490 29.160 41.750 29.480 ;
        RECT 41.030 28.820 41.290 29.140 ;
        RECT 41.550 27.440 41.690 29.160 ;
        RECT 41.490 27.120 41.750 27.440 ;
        RECT 40.570 25.760 40.830 26.080 ;
        RECT 39.190 24.235 39.450 24.380 ;
        RECT 39.180 24.120 39.460 24.235 ;
        RECT 39.180 23.980 39.850 24.120 ;
        RECT 39.180 23.865 39.460 23.980 ;
        RECT 39.190 17.600 39.450 17.920 ;
        RECT 37.350 17.260 37.610 17.580 ;
        RECT 37.410 15.540 37.550 17.260 ;
        RECT 39.250 15.540 39.390 17.600 ;
        RECT 39.710 15.540 39.850 23.980 ;
        RECT 40.570 23.380 40.830 23.700 ;
        RECT 40.630 22.000 40.770 23.380 ;
        RECT 40.570 21.680 40.830 22.000 ;
        RECT 40.630 18.940 40.770 21.680 ;
        RECT 41.550 21.230 41.690 27.120 ;
        RECT 42.010 24.630 42.150 34.260 ;
        RECT 42.410 29.160 42.670 29.480 ;
        RECT 42.470 27.440 42.610 29.160 ;
        RECT 42.410 27.120 42.670 27.440 ;
        RECT 42.410 24.630 42.670 24.720 ;
        RECT 42.010 24.490 42.670 24.630 ;
        RECT 42.410 24.400 42.670 24.490 ;
        RECT 42.470 24.040 42.610 24.400 ;
        RECT 42.410 23.720 42.670 24.040 ;
        RECT 41.090 21.090 41.690 21.230 ;
        RECT 40.570 18.620 40.830 18.940 ;
        RECT 41.090 16.560 41.230 21.090 ;
        RECT 41.490 19.980 41.750 20.300 ;
        RECT 41.550 18.940 41.690 19.980 ;
        RECT 41.490 18.620 41.750 18.940 ;
        RECT 41.030 16.240 41.290 16.560 ;
        RECT 36.430 15.220 36.690 15.540 ;
        RECT 37.350 15.220 37.610 15.540 ;
        RECT 39.190 15.220 39.450 15.540 ;
        RECT 39.650 15.220 39.910 15.540 ;
        RECT 42.470 15.450 42.610 23.720 ;
        RECT 42.930 23.360 43.070 40.130 ;
        RECT 43.390 37.300 43.530 42.420 ;
        RECT 43.330 36.980 43.590 37.300 ;
        RECT 44.250 31.200 44.510 31.520 ;
        RECT 44.310 28.460 44.450 31.200 ;
        RECT 44.710 30.860 44.970 31.180 ;
        RECT 44.250 28.140 44.510 28.460 ;
        RECT 44.310 24.380 44.450 28.140 ;
        RECT 44.770 26.420 44.910 30.860 ;
        RECT 44.710 26.100 44.970 26.420 ;
        RECT 44.250 24.060 44.510 24.380 ;
        RECT 42.870 23.040 43.130 23.360 ;
        RECT 42.870 21.680 43.130 22.000 ;
        RECT 42.930 21.515 43.070 21.680 ;
        RECT 42.860 21.145 43.140 21.515 ;
        RECT 42.930 20.980 43.070 21.145 ;
        RECT 42.870 20.660 43.130 20.980 ;
        RECT 43.790 20.660 44.050 20.980 ;
        RECT 43.850 16.560 43.990 20.660 ;
        RECT 43.790 16.240 44.050 16.560 ;
        RECT 44.310 15.540 44.450 24.060 ;
        RECT 45.230 17.180 45.370 65.340 ;
        RECT 45.630 63.500 45.890 63.820 ;
        RECT 45.690 57.360 45.830 63.500 ;
        RECT 46.150 59.400 46.290 66.220 ;
        RECT 47.070 64.500 47.210 66.900 ;
        RECT 47.530 64.920 47.670 69.620 ;
        RECT 48.390 68.940 48.650 69.260 ;
        RECT 47.930 67.240 48.190 67.560 ;
        RECT 47.990 65.520 48.130 67.240 ;
        RECT 47.930 65.200 48.190 65.520 ;
        RECT 47.530 64.840 48.130 64.920 ;
        RECT 47.470 64.780 48.130 64.840 ;
        RECT 47.470 64.520 47.730 64.780 ;
        RECT 47.010 64.180 47.270 64.500 ;
        RECT 47.990 63.820 48.130 64.780 ;
        RECT 47.930 63.500 48.190 63.820 ;
        RECT 48.450 60.080 48.590 68.940 ;
        RECT 48.850 65.200 49.110 65.520 ;
        RECT 48.390 59.760 48.650 60.080 ;
        RECT 48.910 59.480 49.050 65.200 ;
        RECT 46.090 59.080 46.350 59.400 ;
        RECT 48.450 59.340 49.050 59.480 ;
        RECT 45.630 57.040 45.890 57.360 ;
        RECT 47.010 56.360 47.270 56.680 ;
        RECT 47.070 53.620 47.210 56.360 ;
        RECT 47.930 56.020 48.190 56.340 ;
        RECT 47.010 53.300 47.270 53.620 ;
        RECT 47.990 50.220 48.130 56.020 ;
        RECT 48.450 53.620 48.590 59.340 ;
        RECT 48.850 56.360 49.110 56.680 ;
        RECT 48.390 53.300 48.650 53.620 ;
        RECT 46.090 49.900 46.350 50.220 ;
        RECT 47.930 49.900 48.190 50.220 ;
        RECT 46.150 48.520 46.290 49.900 ;
        RECT 47.990 48.520 48.130 49.900 ;
        RECT 46.090 48.200 46.350 48.520 ;
        RECT 47.930 48.200 48.190 48.520 ;
        RECT 47.990 42.400 48.130 48.200 ;
        RECT 48.450 45.800 48.590 53.300 ;
        RECT 48.390 45.480 48.650 45.800 ;
        RECT 46.550 42.080 46.810 42.400 ;
        RECT 47.930 42.080 48.190 42.400 ;
        RECT 46.610 41.040 46.750 42.080 ;
        RECT 46.550 40.720 46.810 41.040 ;
        RECT 48.390 39.875 48.650 40.020 ;
        RECT 48.380 39.505 48.660 39.875 ;
        RECT 48.450 37.980 48.590 39.505 ;
        RECT 48.390 37.660 48.650 37.980 ;
        RECT 45.630 36.980 45.890 37.300 ;
        RECT 46.090 36.980 46.350 37.300 ;
        RECT 46.550 36.980 46.810 37.300 ;
        RECT 45.690 27.100 45.830 36.980 ;
        RECT 46.150 35.600 46.290 36.980 ;
        RECT 46.090 35.280 46.350 35.600 ;
        RECT 46.610 30.160 46.750 36.980 ;
        RECT 48.390 31.880 48.650 32.200 ;
        RECT 46.550 29.840 46.810 30.160 ;
        RECT 45.630 26.780 45.890 27.100 ;
        RECT 46.610 26.420 46.750 29.840 ;
        RECT 47.470 26.440 47.730 26.760 ;
        RECT 46.550 26.100 46.810 26.420 ;
        RECT 45.630 24.235 45.890 24.380 ;
        RECT 45.620 23.865 45.900 24.235 ;
        RECT 46.610 20.980 46.750 26.100 ;
        RECT 47.530 21.320 47.670 26.440 ;
        RECT 48.450 26.080 48.590 31.880 ;
        RECT 48.390 25.760 48.650 26.080 ;
        RECT 48.450 24.720 48.590 25.760 ;
        RECT 48.390 24.400 48.650 24.720 ;
        RECT 47.930 23.380 48.190 23.700 ;
        RECT 47.470 21.000 47.730 21.320 ;
        RECT 46.550 20.660 46.810 20.980 ;
        RECT 47.010 19.980 47.270 20.300 ;
        RECT 47.070 18.600 47.210 19.980 ;
        RECT 47.990 19.280 48.130 23.380 ;
        RECT 47.930 18.960 48.190 19.280 ;
        RECT 47.010 18.280 47.270 18.600 ;
        RECT 45.230 17.040 46.750 17.180 ;
        RECT 46.610 16.220 46.750 17.040 ;
        RECT 46.550 15.900 46.810 16.220 ;
        RECT 47.990 15.540 48.130 18.960 ;
        RECT 42.870 15.450 43.130 15.540 ;
        RECT 42.470 15.310 43.130 15.450 ;
        RECT 42.870 15.220 43.130 15.310 ;
        RECT 44.250 15.220 44.510 15.540 ;
        RECT 47.930 15.220 48.190 15.540 ;
        RECT 48.450 15.200 48.590 24.400 ;
        RECT 48.910 23.360 49.050 56.360 ;
        RECT 49.370 50.560 49.510 97.500 ;
        RECT 49.830 97.480 49.970 123.340 ;
        RECT 52.590 118.560 52.730 161.940 ;
        RECT 53.050 160.720 53.190 162.100 ;
        RECT 53.510 162.080 53.650 168.220 ;
        RECT 53.510 161.940 54.570 162.080 ;
        RECT 53.450 161.420 53.710 161.740 ;
        RECT 53.910 161.420 54.170 161.740 ;
        RECT 52.990 160.400 53.250 160.720 ;
        RECT 53.050 156.980 53.190 160.400 ;
        RECT 53.510 159.700 53.650 161.420 ;
        RECT 53.450 159.380 53.710 159.700 ;
        RECT 53.510 158.000 53.650 159.380 ;
        RECT 53.450 157.680 53.710 158.000 ;
        RECT 52.990 156.660 53.250 156.980 ;
        RECT 53.970 156.300 54.110 161.420 ;
        RECT 52.990 155.980 53.250 156.300 ;
        RECT 53.910 155.980 54.170 156.300 ;
        RECT 53.050 153.920 53.190 155.980 ;
        RECT 53.450 154.280 53.710 154.600 ;
        RECT 52.990 153.600 53.250 153.920 ;
        RECT 53.510 152.220 53.650 154.280 ;
        RECT 54.430 153.920 54.570 161.940 ;
        RECT 55.810 154.600 55.950 168.560 ;
        RECT 56.270 168.200 56.410 170.600 ;
        RECT 56.210 167.880 56.470 168.200 ;
        RECT 56.270 160.040 56.410 167.880 ;
        RECT 56.730 167.860 56.870 173.320 ;
        RECT 57.650 173.210 57.790 178.080 ;
        RECT 58.570 174.320 58.710 178.080 ;
        RECT 58.510 174.000 58.770 174.320 ;
        RECT 58.510 173.210 58.770 173.300 ;
        RECT 57.650 173.070 58.770 173.210 ;
        RECT 58.510 172.980 58.770 173.070 ;
        RECT 57.130 170.940 57.390 171.260 ;
        RECT 57.190 168.200 57.330 170.940 ;
        RECT 58.570 170.240 58.710 172.980 ;
        RECT 58.510 169.920 58.770 170.240 ;
        RECT 59.030 169.900 59.170 178.420 ;
        RECT 60.410 178.340 61.010 178.480 ;
        RECT 59.890 176.380 60.150 176.700 ;
        RECT 58.970 169.580 59.230 169.900 ;
        RECT 59.430 169.580 59.690 169.900 ;
        RECT 57.130 167.880 57.390 168.200 ;
        RECT 56.670 167.540 56.930 167.860 ;
        RECT 56.730 165.820 56.870 167.540 ;
        RECT 56.670 165.500 56.930 165.820 ;
        RECT 57.190 165.480 57.330 167.880 ;
        RECT 59.490 167.860 59.630 169.580 ;
        RECT 59.430 167.540 59.690 167.860 ;
        RECT 57.590 167.200 57.850 167.520 ;
        RECT 57.650 165.480 57.790 167.200 ;
        RECT 59.950 166.920 60.090 176.380 ;
        RECT 60.410 171.600 60.550 178.340 ;
        RECT 62.250 177.040 62.390 181.230 ;
        RECT 63.170 181.120 63.310 183.520 ;
        RECT 64.090 182.480 64.230 183.860 ;
        RECT 64.030 182.160 64.290 182.480 ;
        RECT 63.570 181.820 63.830 182.140 ;
        RECT 63.110 180.800 63.370 181.120 ;
        RECT 63.630 180.520 63.770 181.820 ;
        RECT 63.170 180.380 63.770 180.520 ;
        RECT 63.170 178.740 63.310 180.380 ;
        RECT 64.090 178.740 64.230 182.160 ;
        RECT 66.850 181.800 66.990 184.540 ;
        RECT 67.310 182.140 67.450 184.880 ;
        RECT 67.770 183.500 67.910 193.040 ;
        RECT 68.230 192.680 68.370 194.060 ;
        RECT 69.610 193.020 69.750 199.500 ;
        RECT 101.480 198.895 105.480 198.965 ;
        RECT 112.175 198.905 112.545 200.445 ;
        RECT 117.615 198.905 117.985 200.445 ;
        RECT 123.055 198.905 123.425 200.445 ;
        RECT 128.495 198.905 128.865 200.445 ;
        RECT 130.390 200.275 130.710 200.335 ;
        RECT 133.030 200.275 133.170 200.595 ;
        RECT 137.190 200.535 137.510 200.595 ;
        RECT 141.610 200.735 141.930 200.795 ;
        RECT 146.710 200.735 147.030 200.795 ;
        RECT 141.610 200.595 147.030 200.735 ;
        RECT 141.610 200.535 141.930 200.595 ;
        RECT 146.710 200.535 147.030 200.595 ;
        RECT 130.390 200.135 133.170 200.275 ;
        RECT 130.390 200.075 130.710 200.135 ;
        RECT 133.935 198.905 134.305 200.445 ;
        RECT 139.375 198.905 139.745 200.445 ;
        RECT 140.590 200.275 140.910 200.335 ;
        RECT 143.310 200.275 143.630 200.335 ;
        RECT 140.590 200.135 143.630 200.275 ;
        RECT 140.590 200.075 140.910 200.135 ;
        RECT 143.310 200.075 143.630 200.135 ;
        RECT 144.815 198.905 145.185 200.445 ;
        RECT 147.050 198.895 147.370 198.955 ;
        RECT 148.660 198.895 148.920 198.985 ;
        RECT 155.245 198.895 159.245 198.965 ;
        RECT 101.480 198.755 107.330 198.895 ;
        RECT 101.480 198.685 105.480 198.755 ;
        RECT 107.190 198.435 107.330 198.755 ;
        RECT 147.050 198.755 159.245 198.895 ;
        RECT 147.050 198.695 147.370 198.755 ;
        RECT 148.660 198.665 148.920 198.755 ;
        RECT 155.245 198.685 159.245 198.755 ;
        RECT 111.410 198.435 111.740 198.530 ;
        RECT 112.710 198.435 113.030 198.495 ;
        RECT 107.190 198.295 113.030 198.435 ;
        RECT 111.410 198.200 111.740 198.295 ;
        RECT 112.710 198.235 113.030 198.295 ;
        RECT 126.990 198.435 127.310 198.495 ;
        RECT 134.470 198.435 134.790 198.495 ;
        RECT 136.170 198.435 136.490 198.495 ;
        RECT 140.590 198.435 140.910 198.495 ;
        RECT 126.990 198.295 135.890 198.435 ;
        RECT 126.990 198.235 127.310 198.295 ;
        RECT 134.470 198.235 134.790 198.295 ;
        RECT 70.010 197.800 70.270 198.120 ;
        RECT 114.410 197.975 114.730 198.035 ;
        RECT 123.590 197.975 123.910 198.035 ;
        RECT 126.990 197.975 127.310 198.035 ;
        RECT 114.410 197.835 127.310 197.975 ;
        RECT 70.070 196.080 70.210 197.800 ;
        RECT 75.990 197.460 76.250 197.780 ;
        RECT 114.410 197.775 114.730 197.835 ;
        RECT 123.590 197.775 123.910 197.835 ;
        RECT 126.990 197.775 127.310 197.835 ;
        RECT 133.450 197.975 133.770 198.035 ;
        RECT 134.810 197.975 135.130 198.035 ;
        RECT 133.450 197.835 135.130 197.975 ;
        RECT 135.750 197.975 135.890 198.295 ;
        RECT 136.170 198.295 140.910 198.435 ;
        RECT 136.170 198.235 136.490 198.295 ;
        RECT 140.590 198.235 140.910 198.295 ;
        RECT 144.330 198.435 144.650 198.495 ;
        RECT 146.030 198.435 146.350 198.495 ;
        RECT 144.330 198.295 146.350 198.435 ;
        RECT 144.330 198.235 144.650 198.295 ;
        RECT 146.030 198.235 146.350 198.295 ;
        RECT 140.590 197.975 140.910 198.035 ;
        RECT 135.750 197.835 140.910 197.975 ;
        RECT 133.450 197.775 133.770 197.835 ;
        RECT 134.810 197.775 135.130 197.835 ;
        RECT 140.590 197.775 140.910 197.835 ;
        RECT 143.990 197.975 144.310 198.035 ;
        RECT 145.350 197.975 145.670 198.035 ;
        RECT 143.990 197.835 145.670 197.975 ;
        RECT 143.990 197.775 144.310 197.835 ;
        RECT 145.350 197.775 145.670 197.835 ;
        RECT 124.610 197.515 124.930 197.575 ;
        RECT 70.010 195.760 70.270 196.080 ;
        RECT 76.050 195.400 76.190 197.460 ;
        RECT 124.610 197.315 125.010 197.515 ;
        RECT 128.010 197.315 128.330 197.575 ;
        RECT 135.150 197.515 135.470 197.575 ;
        RECT 137.870 197.515 138.190 197.575 ;
        RECT 135.150 197.375 138.190 197.515 ;
        RECT 135.150 197.315 135.470 197.375 ;
        RECT 137.870 197.315 138.190 197.375 ;
        RECT 140.930 197.515 141.250 197.575 ;
        RECT 142.630 197.515 142.950 197.575 ;
        RECT 140.930 197.375 142.950 197.515 ;
        RECT 140.930 197.315 141.250 197.375 ;
        RECT 142.630 197.315 142.950 197.375 ;
        RECT 124.870 197.055 125.010 197.315 ;
        RECT 128.100 197.055 128.240 197.315 ;
        RECT 130.050 197.055 130.370 197.115 ;
        RECT 135.830 197.055 136.150 197.115 ;
        RECT 124.870 196.915 136.150 197.055 ;
        RECT 130.050 196.855 130.370 196.915 ;
        RECT 135.830 196.855 136.150 196.915 ;
        RECT 140.590 197.055 140.910 197.115 ;
        RECT 143.650 197.055 143.970 197.115 ;
        RECT 140.590 196.915 143.970 197.055 ;
        RECT 140.590 196.855 140.910 196.915 ;
        RECT 143.650 196.855 143.970 196.915 ;
        RECT 124.950 196.595 125.270 196.655 ;
        RECT 134.810 196.595 135.130 196.655 ;
        RECT 124.950 196.455 135.130 196.595 ;
        RECT 124.950 196.395 125.270 196.455 ;
        RECT 134.810 196.395 135.130 196.455 ;
        RECT 117.130 196.135 117.450 196.195 ;
        RECT 122.230 196.135 122.550 196.195 ;
        RECT 126.650 196.135 126.970 196.195 ;
        RECT 117.130 195.995 126.970 196.135 ;
        RECT 117.130 195.935 117.450 195.995 ;
        RECT 122.230 195.935 122.550 195.995 ;
        RECT 126.650 195.935 126.970 195.995 ;
        RECT 130.390 196.135 130.710 196.195 ;
        RECT 131.750 196.135 132.070 196.195 ;
        RECT 138.550 196.135 138.870 196.195 ;
        RECT 143.310 196.135 143.630 196.195 ;
        RECT 130.390 195.995 143.630 196.135 ;
        RECT 130.390 195.935 130.710 195.995 ;
        RECT 131.750 195.935 132.070 195.995 ;
        RECT 138.550 195.935 138.870 195.995 ;
        RECT 143.310 195.935 143.630 195.995 ;
        RECT 133.450 195.675 133.770 195.735 ;
        RECT 137.530 195.675 137.850 195.735 ;
        RECT 140.250 195.675 140.570 195.735 ;
        RECT 141.610 195.675 141.930 195.735 ;
        RECT 143.650 195.675 143.970 195.735 ;
        RECT 133.450 195.535 140.570 195.675 ;
        RECT 133.450 195.475 133.770 195.535 ;
        RECT 137.530 195.475 137.850 195.535 ;
        RECT 140.250 195.475 140.570 195.535 ;
        RECT 141.190 195.535 143.970 195.675 ;
        RECT 75.990 195.080 76.250 195.400 ;
        RECT 116.110 195.215 116.430 195.275 ;
        RECT 121.890 195.215 122.210 195.275 ;
        RECT 125.290 195.215 125.610 195.275 ;
        RECT 141.190 195.215 141.330 195.535 ;
        RECT 141.610 195.475 141.930 195.535 ;
        RECT 143.650 195.475 143.970 195.535 ;
        RECT 146.030 195.675 146.350 195.735 ;
        RECT 148.050 195.675 148.470 195.800 ;
        RECT 155.245 195.675 159.245 195.745 ;
        RECT 146.030 195.535 159.245 195.675 ;
        RECT 146.030 195.475 146.350 195.535 ;
        RECT 148.050 195.410 148.470 195.535 ;
        RECT 155.245 195.465 159.245 195.535 ;
        RECT 71.850 194.400 72.110 194.720 ;
        RECT 71.910 193.360 72.050 194.400 ;
        RECT 71.850 193.040 72.110 193.360 ;
        RECT 69.550 192.700 69.810 193.020 ;
        RECT 68.170 192.360 68.430 192.680 ;
        RECT 70.470 192.360 70.730 192.680 ;
        RECT 73.230 192.360 73.490 192.680 ;
        RECT 68.230 189.960 68.370 192.360 ;
        RECT 69.550 192.020 69.810 192.340 ;
        RECT 68.170 189.640 68.430 189.960 ;
        RECT 69.610 189.620 69.750 192.020 ;
        RECT 70.530 190.640 70.670 192.360 ;
        RECT 70.470 190.320 70.730 190.640 ;
        RECT 73.290 189.620 73.430 192.360 ;
        RECT 69.550 189.300 69.810 189.620 ;
        RECT 73.230 189.300 73.490 189.620 ;
        RECT 71.390 188.960 71.650 189.280 ;
        RECT 70.470 183.520 70.730 183.840 ;
        RECT 67.710 183.180 67.970 183.500 ;
        RECT 68.630 183.180 68.890 183.500 ;
        RECT 67.250 181.820 67.510 182.140 ;
        RECT 66.790 181.480 67.050 181.800 ;
        RECT 63.110 178.420 63.370 178.740 ;
        RECT 64.030 178.420 64.290 178.740 ;
        RECT 64.490 178.420 64.750 178.740 ;
        RECT 62.190 176.720 62.450 177.040 ;
        RECT 62.250 173.300 62.390 176.720 ;
        RECT 63.170 176.700 63.310 178.420 ;
        RECT 63.110 176.380 63.370 176.700 ;
        RECT 62.190 172.980 62.450 173.300 ;
        RECT 62.650 172.980 62.910 173.300 ;
        RECT 60.350 171.280 60.610 171.600 ;
        RECT 60.410 170.920 60.550 171.280 ;
        RECT 60.350 170.600 60.610 170.920 ;
        RECT 60.410 169.900 60.550 170.600 ;
        RECT 60.350 169.580 60.610 169.900 ;
        RECT 62.250 168.790 62.390 172.980 ;
        RECT 62.710 170.580 62.850 172.980 ;
        RECT 64.550 171.600 64.690 178.420 ;
        RECT 66.850 178.400 66.990 181.480 ;
        RECT 67.770 180.780 67.910 183.180 ;
        RECT 68.170 181.820 68.430 182.140 ;
        RECT 68.690 182.050 68.830 183.180 ;
        RECT 69.090 182.050 69.350 182.140 ;
        RECT 68.690 181.910 69.350 182.050 ;
        RECT 69.090 181.820 69.350 181.910 ;
        RECT 67.710 180.460 67.970 180.780 ;
        RECT 67.770 179.080 67.910 180.460 ;
        RECT 68.230 179.760 68.370 181.820 ;
        RECT 68.630 181.140 68.890 181.460 ;
        RECT 69.550 181.140 69.810 181.460 ;
        RECT 68.170 179.440 68.430 179.760 ;
        RECT 67.710 178.760 67.970 179.080 ;
        RECT 66.790 178.080 67.050 178.400 ;
        RECT 66.850 172.620 66.990 178.080 ;
        RECT 68.690 178.060 68.830 181.140 ;
        RECT 68.630 177.740 68.890 178.060 ;
        RECT 67.710 176.040 67.970 176.360 ;
        RECT 67.770 173.300 67.910 176.040 ;
        RECT 68.690 176.020 68.830 177.740 ;
        RECT 69.090 176.040 69.350 176.360 ;
        RECT 68.630 175.700 68.890 176.020 ;
        RECT 68.170 175.020 68.430 175.340 ;
        RECT 67.710 172.980 67.970 173.300 ;
        RECT 66.790 172.300 67.050 172.620 ;
        RECT 64.490 171.280 64.750 171.600 ;
        RECT 64.950 171.280 65.210 171.600 ;
        RECT 62.650 170.260 62.910 170.580 ;
        RECT 62.250 168.650 62.850 168.790 ;
        RECT 60.810 167.880 61.070 168.200 ;
        RECT 62.190 167.880 62.450 168.200 ;
        RECT 59.030 166.780 60.090 166.920 ;
        RECT 59.030 166.160 59.170 166.780 ;
        RECT 58.970 165.840 59.230 166.160 ;
        RECT 57.130 165.160 57.390 165.480 ;
        RECT 57.590 165.160 57.850 165.480 ;
        RECT 57.650 162.420 57.790 165.160 ;
        RECT 57.590 162.100 57.850 162.420 ;
        RECT 56.210 159.720 56.470 160.040 ;
        RECT 57.650 157.400 57.790 162.100 ;
        RECT 57.650 157.260 58.250 157.400 ;
        RECT 56.210 156.660 56.470 156.980 ;
        RECT 57.590 156.660 57.850 156.980 ;
        RECT 56.270 155.280 56.410 156.660 ;
        RECT 56.210 154.960 56.470 155.280 ;
        RECT 55.750 154.280 56.010 154.600 ;
        RECT 54.370 153.600 54.630 153.920 ;
        RECT 53.910 153.260 54.170 153.580 ;
        RECT 53.450 151.900 53.710 152.220 ;
        RECT 53.510 149.840 53.650 151.900 ;
        RECT 53.970 151.540 54.110 153.260 ;
        RECT 53.910 151.220 54.170 151.540 ;
        RECT 57.650 151.200 57.790 156.660 ;
        RECT 57.590 150.880 57.850 151.200 ;
        RECT 53.450 149.520 53.710 149.840 ;
        RECT 57.590 148.840 57.850 149.160 ;
        RECT 57.650 147.120 57.790 148.840 ;
        RECT 57.590 146.800 57.850 147.120 ;
        RECT 58.110 144.060 58.250 157.260 ;
        RECT 58.510 152.240 58.770 152.560 ;
        RECT 58.570 151.880 58.710 152.240 ;
        RECT 58.510 151.560 58.770 151.880 ;
        RECT 58.050 143.740 58.310 144.060 ;
        RECT 58.570 143.720 58.710 151.560 ;
        RECT 59.030 146.100 59.170 165.840 ;
        RECT 60.870 160.380 61.010 167.880 ;
        RECT 62.250 165.480 62.390 167.880 ;
        RECT 62.710 165.480 62.850 168.650 ;
        RECT 65.010 166.160 65.150 171.280 ;
        RECT 66.330 170.830 66.590 170.920 ;
        RECT 66.850 170.830 66.990 172.300 ;
        RECT 67.770 170.920 67.910 172.980 ;
        RECT 68.230 172.960 68.370 175.020 ;
        RECT 69.150 174.320 69.290 176.040 ;
        RECT 69.090 174.000 69.350 174.320 ;
        RECT 68.620 173.465 68.900 173.835 ;
        RECT 68.630 173.320 68.890 173.465 ;
        RECT 68.170 172.640 68.430 172.960 ;
        RECT 69.610 171.260 69.750 181.140 ;
        RECT 70.530 180.780 70.670 183.520 ;
        RECT 70.470 180.460 70.730 180.780 ;
        RECT 71.450 178.740 71.590 188.960 ;
        RECT 76.050 184.520 76.190 195.080 ;
        RECT 116.110 195.075 141.330 195.215 ;
        RECT 116.110 195.015 116.430 195.075 ;
        RECT 121.890 195.015 122.210 195.075 ;
        RECT 125.290 195.015 125.610 195.075 ;
        RECT 113.390 194.755 113.710 194.815 ;
        RECT 114.070 194.755 114.390 194.815 ;
        RECT 116.110 194.755 116.430 194.815 ;
        RECT 113.390 194.615 116.430 194.755 ;
        RECT 113.390 194.555 113.710 194.615 ;
        RECT 114.070 194.555 114.390 194.615 ;
        RECT 116.110 194.555 116.430 194.615 ;
        RECT 140.590 194.755 140.910 194.815 ;
        RECT 142.630 194.755 142.950 194.815 ;
        RECT 140.590 194.615 142.950 194.755 ;
        RECT 140.590 194.555 140.910 194.615 ;
        RECT 142.630 194.555 142.950 194.615 ;
        RECT 120.870 194.295 121.190 194.355 ;
        RECT 121.550 194.295 121.870 194.355 ;
        RECT 129.030 194.295 129.350 194.355 ;
        RECT 120.870 194.155 129.350 194.295 ;
        RECT 120.870 194.095 121.190 194.155 ;
        RECT 121.550 194.095 121.870 194.155 ;
        RECT 129.030 194.095 129.350 194.155 ;
        RECT 115.235 193.835 115.605 193.905 ;
        RECT 118.830 193.835 119.150 193.895 ;
        RECT 115.235 193.695 119.150 193.835 ;
        RECT 115.235 193.625 115.605 193.695 ;
        RECT 118.830 193.635 119.150 193.695 ;
        RECT 127.330 193.835 127.650 193.895 ;
        RECT 130.730 193.835 131.050 193.895 ;
        RECT 137.190 193.835 137.510 193.895 ;
        RECT 127.330 193.695 137.510 193.835 ;
        RECT 127.330 193.635 127.650 193.695 ;
        RECT 130.730 193.635 131.050 193.695 ;
        RECT 137.190 193.635 137.510 193.695 ;
        RECT 143.650 193.835 143.970 193.895 ;
        RECT 146.710 193.835 147.030 193.895 ;
        RECT 143.650 193.695 147.030 193.835 ;
        RECT 143.650 193.635 143.970 193.695 ;
        RECT 146.710 193.635 147.030 193.695 ;
        RECT 132.770 192.915 133.090 192.975 ;
        RECT 134.470 192.915 134.790 192.975 ;
        RECT 132.770 192.775 134.790 192.915 ;
        RECT 132.770 192.715 133.090 192.775 ;
        RECT 134.470 192.715 134.790 192.775 ;
        RECT 101.480 192.455 105.480 192.525 ;
        RECT 109.920 192.455 110.240 192.515 ;
        RECT 112.710 192.455 113.030 192.515 ;
        RECT 101.480 192.315 113.030 192.455 ;
        RECT 101.480 192.245 105.480 192.315 ;
        RECT 109.920 192.255 110.240 192.315 ;
        RECT 112.710 192.255 113.030 192.315 ;
        RECT 118.830 192.455 119.150 192.515 ;
        RECT 125.435 192.455 125.805 192.525 ;
        RECT 118.830 192.315 125.805 192.455 ;
        RECT 118.830 192.255 119.150 192.315 ;
        RECT 125.435 192.245 125.805 192.315 ;
        RECT 147.050 192.455 147.370 192.515 ;
        RECT 148.570 192.455 148.900 192.550 ;
        RECT 155.245 192.455 159.245 192.525 ;
        RECT 147.050 192.315 159.245 192.455 ;
        RECT 147.050 192.255 147.370 192.315 ;
        RECT 148.570 192.220 148.900 192.315 ;
        RECT 155.245 192.245 159.245 192.315 ;
        RECT 113.390 191.995 113.710 192.055 ;
        RECT 120.870 191.995 121.190 192.055 ;
        RECT 124.270 191.995 124.590 192.055 ;
        RECT 113.390 191.855 124.590 191.995 ;
        RECT 113.390 191.795 113.710 191.855 ;
        RECT 120.870 191.795 121.190 191.855 ;
        RECT 124.270 191.795 124.590 191.855 ;
        RECT 132.770 191.995 133.090 192.055 ;
        RECT 138.210 191.995 138.530 192.055 ;
        RECT 145.350 191.995 145.670 192.055 ;
        RECT 132.770 191.855 145.670 191.995 ;
        RECT 132.770 191.795 133.090 191.855 ;
        RECT 138.210 191.795 138.530 191.855 ;
        RECT 145.350 191.795 145.670 191.855 ;
        RECT 127.330 191.535 127.650 191.595 ;
        RECT 129.030 191.535 129.350 191.595 ;
        RECT 127.330 191.395 129.350 191.535 ;
        RECT 127.330 191.335 127.650 191.395 ;
        RECT 129.030 191.335 129.350 191.395 ;
        RECT 138.550 191.535 138.870 191.595 ;
        RECT 138.550 191.395 143.880 191.535 ;
        RECT 138.550 191.335 138.870 191.395 ;
        RECT 143.740 191.145 143.880 191.395 ;
        RECT 118.635 191.135 119.005 191.145 ;
        RECT 143.740 191.135 144.165 191.145 ;
        RECT 118.635 190.875 119.150 191.135 ;
        RECT 122.570 191.075 122.890 191.135 ;
        RECT 123.590 191.075 123.910 191.135 ;
        RECT 122.570 190.935 123.910 191.075 ;
        RECT 122.570 190.875 122.890 190.935 ;
        RECT 123.590 190.875 123.910 190.935 ;
        RECT 129.710 191.075 130.030 191.135 ;
        RECT 135.150 191.075 135.470 191.135 ;
        RECT 137.530 191.075 137.850 191.135 ;
        RECT 138.550 191.075 138.870 191.135 ;
        RECT 129.710 190.935 130.450 191.075 ;
        RECT 129.710 190.875 130.030 190.935 ;
        RECT 118.635 190.865 119.005 190.875 ;
        RECT 128.835 190.155 129.205 190.225 ;
        RECT 129.710 190.155 130.030 190.215 ;
        RECT 128.835 190.015 130.030 190.155 ;
        RECT 130.310 190.155 130.450 190.935 ;
        RECT 135.150 190.935 138.870 191.075 ;
        RECT 135.150 190.875 135.470 190.935 ;
        RECT 137.530 190.875 137.850 190.935 ;
        RECT 138.550 190.875 138.870 190.935 ;
        RECT 143.650 190.875 144.165 191.135 ;
        RECT 143.795 190.865 144.165 190.875 ;
        RECT 141.610 190.615 141.930 190.675 ;
        RECT 142.970 190.615 143.290 190.675 ;
        RECT 146.030 190.615 146.350 190.675 ;
        RECT 141.610 190.475 146.350 190.615 ;
        RECT 141.610 190.415 141.930 190.475 ;
        RECT 142.970 190.415 143.290 190.475 ;
        RECT 146.030 190.415 146.350 190.475 ;
        RECT 135.830 190.155 136.150 190.215 ;
        RECT 130.310 190.015 136.150 190.155 ;
        RECT 128.835 189.945 129.205 190.015 ;
        RECT 129.710 189.955 130.030 190.015 ;
        RECT 135.830 189.955 136.150 190.015 ;
        RECT 113.730 189.695 114.050 189.755 ;
        RECT 116.110 189.695 116.430 189.755 ;
        RECT 118.150 189.695 118.470 189.755 ;
        RECT 113.730 189.555 118.470 189.695 ;
        RECT 113.730 189.495 114.050 189.555 ;
        RECT 116.110 189.495 116.430 189.555 ;
        RECT 118.150 189.495 118.470 189.555 ;
        RECT 124.610 189.695 124.930 189.755 ;
        RECT 127.670 189.695 127.990 189.755 ;
        RECT 129.370 189.695 129.690 189.755 ;
        RECT 131.750 189.695 132.070 189.755 ;
        RECT 124.610 189.555 132.070 189.695 ;
        RECT 124.610 189.495 124.930 189.555 ;
        RECT 127.670 189.495 127.990 189.555 ;
        RECT 129.370 189.495 129.690 189.555 ;
        RECT 131.750 189.495 132.070 189.555 ;
        RECT 111.835 189.235 112.205 189.305 ;
        RECT 113.390 189.235 113.710 189.295 ;
        RECT 111.835 189.095 113.710 189.235 ;
        RECT 111.835 189.025 112.205 189.095 ;
        RECT 113.390 189.035 113.710 189.095 ;
        RECT 116.450 189.235 116.770 189.295 ;
        RECT 118.150 189.235 118.470 189.295 ;
        RECT 116.450 189.095 118.470 189.235 ;
        RECT 116.450 189.035 116.770 189.095 ;
        RECT 118.150 189.035 118.470 189.095 ;
        RECT 119.850 189.235 120.170 189.295 ;
        RECT 121.550 189.235 121.870 189.295 ;
        RECT 124.270 189.235 124.590 189.295 ;
        RECT 119.850 189.095 124.590 189.235 ;
        RECT 119.850 189.035 120.170 189.095 ;
        RECT 121.550 189.035 121.870 189.095 ;
        RECT 124.270 189.035 124.590 189.095 ;
        RECT 125.290 189.235 125.610 189.295 ;
        RECT 135.490 189.235 135.810 189.295 ;
        RECT 125.290 189.095 135.810 189.235 ;
        RECT 125.290 189.035 125.610 189.095 ;
        RECT 135.490 189.035 135.810 189.095 ;
        RECT 122.035 188.835 122.405 188.845 ;
        RECT 114.070 188.775 114.390 188.835 ;
        RECT 119.510 188.775 119.830 188.835 ;
        RECT 114.070 188.635 119.830 188.775 ;
        RECT 114.070 188.575 114.390 188.635 ;
        RECT 119.510 188.575 119.830 188.635 ;
        RECT 121.890 188.575 122.405 188.835 ;
        RECT 140.590 188.775 140.910 188.835 ;
        RECT 142.630 188.775 142.950 188.835 ;
        RECT 140.590 188.635 142.950 188.775 ;
        RECT 140.590 188.575 140.910 188.635 ;
        RECT 142.630 188.575 142.950 188.635 ;
        RECT 122.035 188.565 122.405 188.575 ;
        RECT 114.410 188.315 114.730 188.375 ;
        RECT 118.830 188.315 119.150 188.375 ;
        RECT 120.870 188.315 121.190 188.375 ;
        RECT 127.330 188.315 127.650 188.375 ;
        RECT 114.410 188.175 127.650 188.315 ;
        RECT 114.410 188.115 114.730 188.175 ;
        RECT 118.830 188.115 119.150 188.175 ;
        RECT 120.870 188.115 121.190 188.175 ;
        RECT 127.330 188.115 127.650 188.175 ;
        RECT 135.150 188.315 135.470 188.375 ;
        RECT 138.210 188.315 138.530 188.375 ;
        RECT 138.890 188.315 139.210 188.375 ;
        RECT 145.350 188.315 145.670 188.375 ;
        RECT 135.150 188.175 145.670 188.315 ;
        RECT 135.150 188.115 135.470 188.175 ;
        RECT 138.210 188.115 138.530 188.175 ;
        RECT 138.890 188.115 139.210 188.175 ;
        RECT 145.350 188.115 145.670 188.175 ;
        RECT 119.850 187.855 120.170 187.915 ;
        RECT 127.330 187.855 127.650 187.915 ;
        RECT 119.850 187.715 127.650 187.855 ;
        RECT 119.850 187.655 120.170 187.715 ;
        RECT 127.330 187.655 127.650 187.715 ;
        RECT 128.010 187.855 128.330 187.915 ;
        RECT 129.710 187.855 130.030 187.915 ;
        RECT 128.010 187.715 130.030 187.855 ;
        RECT 128.010 187.655 128.330 187.715 ;
        RECT 129.710 187.655 130.030 187.715 ;
        RECT 130.390 187.855 130.710 187.915 ;
        RECT 135.150 187.855 135.470 187.915 ;
        RECT 141.610 187.855 141.930 187.915 ;
        RECT 143.650 187.855 143.970 187.915 ;
        RECT 130.390 187.715 141.330 187.855 ;
        RECT 130.390 187.655 130.710 187.715 ;
        RECT 135.150 187.655 135.470 187.715 ;
        RECT 118.830 187.395 119.150 187.455 ;
        RECT 121.890 187.395 122.210 187.455 ;
        RECT 118.830 187.255 122.210 187.395 ;
        RECT 118.830 187.195 119.150 187.255 ;
        RECT 121.890 187.195 122.210 187.255 ;
        RECT 122.570 187.395 122.890 187.455 ;
        RECT 126.990 187.395 127.310 187.455 ;
        RECT 122.570 187.255 127.310 187.395 ;
        RECT 122.570 187.195 122.890 187.255 ;
        RECT 126.990 187.195 127.310 187.255 ;
        RECT 129.710 187.395 130.030 187.455 ;
        RECT 132.770 187.395 133.090 187.455 ;
        RECT 129.710 187.255 133.090 187.395 ;
        RECT 129.710 187.195 130.030 187.255 ;
        RECT 132.770 187.195 133.090 187.255 ;
        RECT 135.635 187.395 136.005 187.465 ;
        RECT 140.590 187.395 140.910 187.455 ;
        RECT 135.635 187.255 140.910 187.395 ;
        RECT 141.190 187.395 141.330 187.715 ;
        RECT 141.610 187.715 143.970 187.855 ;
        RECT 141.610 187.655 141.930 187.715 ;
        RECT 143.650 187.655 143.970 187.715 ;
        RECT 146.030 187.855 146.350 187.915 ;
        RECT 149.235 187.855 149.605 187.925 ;
        RECT 146.030 187.715 149.605 187.855 ;
        RECT 146.030 187.655 146.350 187.715 ;
        RECT 149.235 187.645 149.605 187.715 ;
        RECT 142.970 187.395 143.290 187.455 ;
        RECT 141.190 187.255 143.290 187.395 ;
        RECT 135.635 187.185 136.005 187.255 ;
        RECT 140.590 187.195 140.910 187.255 ;
        RECT 142.970 187.195 143.290 187.255 ;
        RECT 122.230 186.935 122.550 186.995 ;
        RECT 124.270 186.935 124.590 186.995 ;
        RECT 129.370 186.935 129.690 186.995 ;
        RECT 122.230 186.795 129.690 186.935 ;
        RECT 122.230 186.735 122.550 186.795 ;
        RECT 124.270 186.735 124.590 186.795 ;
        RECT 129.370 186.735 129.690 186.795 ;
        RECT 136.170 186.935 136.490 186.995 ;
        RECT 138.210 186.935 138.530 186.995 ;
        RECT 136.170 186.795 138.530 186.935 ;
        RECT 136.170 186.735 136.490 186.795 ;
        RECT 138.210 186.735 138.530 186.795 ;
        RECT 145.835 186.535 146.205 186.545 ;
        RECT 117.130 186.475 117.450 186.535 ;
        RECT 124.270 186.475 124.590 186.535 ;
        RECT 117.130 186.335 124.590 186.475 ;
        RECT 117.130 186.275 117.450 186.335 ;
        RECT 124.270 186.275 124.590 186.335 ;
        RECT 130.730 186.475 131.050 186.535 ;
        RECT 135.150 186.475 135.470 186.535 ;
        RECT 139.910 186.475 140.230 186.535 ;
        RECT 130.730 186.335 135.470 186.475 ;
        RECT 130.730 186.275 131.050 186.335 ;
        RECT 135.150 186.275 135.470 186.335 ;
        RECT 135.750 186.335 140.230 186.475 ;
        RECT 114.410 186.015 114.730 186.075 ;
        RECT 118.830 186.015 119.150 186.075 ;
        RECT 114.410 185.875 119.150 186.015 ;
        RECT 114.410 185.815 114.730 185.875 ;
        RECT 118.830 185.815 119.150 185.875 ;
        RECT 121.550 186.015 121.870 186.075 ;
        RECT 127.330 186.015 127.650 186.075 ;
        RECT 121.550 185.875 127.650 186.015 ;
        RECT 121.550 185.815 121.870 185.875 ;
        RECT 127.330 185.815 127.650 185.875 ;
        RECT 132.770 186.015 133.090 186.075 ;
        RECT 135.150 186.015 135.470 186.075 ;
        RECT 135.750 186.015 135.890 186.335 ;
        RECT 139.910 186.275 140.230 186.335 ;
        RECT 145.835 186.275 146.350 186.535 ;
        RECT 145.835 186.265 146.205 186.275 ;
        RECT 132.770 185.875 135.890 186.015 ;
        RECT 138.890 186.015 139.210 186.075 ;
        RECT 139.910 186.015 140.230 186.075 ;
        RECT 138.890 185.875 140.230 186.015 ;
        RECT 132.770 185.815 133.090 185.875 ;
        RECT 135.150 185.815 135.470 185.875 ;
        RECT 138.890 185.815 139.210 185.875 ;
        RECT 139.910 185.815 140.230 185.875 ;
        RECT 108.435 185.555 108.805 185.625 ;
        RECT 119.170 185.555 119.490 185.615 ;
        RECT 108.435 185.415 119.490 185.555 ;
        RECT 108.435 185.345 108.805 185.415 ;
        RECT 119.170 185.355 119.490 185.415 ;
        RECT 135.830 185.555 136.150 185.615 ;
        RECT 138.210 185.555 138.530 185.615 ;
        RECT 145.350 185.555 145.670 185.615 ;
        RECT 135.830 185.415 145.670 185.555 ;
        RECT 135.830 185.355 136.150 185.415 ;
        RECT 138.210 185.355 138.530 185.415 ;
        RECT 145.350 185.355 145.670 185.415 ;
        RECT 116.110 185.095 116.430 185.155 ;
        RECT 118.830 185.095 119.150 185.155 ;
        RECT 121.210 185.095 121.530 185.155 ;
        RECT 116.110 184.955 121.530 185.095 ;
        RECT 116.110 184.895 116.430 184.955 ;
        RECT 118.830 184.895 119.150 184.955 ;
        RECT 121.210 184.895 121.530 184.955 ;
        RECT 132.235 185.095 132.605 185.165 ;
        RECT 132.770 185.095 133.090 185.155 ;
        RECT 132.235 184.955 133.090 185.095 ;
        RECT 132.235 184.885 132.605 184.955 ;
        RECT 132.770 184.895 133.090 184.955 ;
        RECT 139.035 185.095 139.405 185.165 ;
        RECT 140.590 185.095 140.910 185.155 ;
        RECT 139.035 184.955 140.910 185.095 ;
        RECT 139.035 184.885 139.405 184.955 ;
        RECT 140.590 184.895 140.910 184.955 ;
        RECT 142.435 185.095 142.805 185.165 ;
        RECT 143.650 185.095 143.970 185.155 ;
        RECT 142.435 184.955 143.970 185.095 ;
        RECT 142.435 184.885 142.805 184.955 ;
        RECT 143.650 184.895 143.970 184.955 ;
        RECT 146.030 185.095 146.350 185.155 ;
        RECT 152.635 185.095 153.005 185.165 ;
        RECT 146.030 184.955 153.005 185.095 ;
        RECT 146.030 184.895 146.350 184.955 ;
        RECT 152.635 184.885 153.005 184.955 ;
        RECT 75.990 184.200 76.250 184.520 ;
        RECT 71.850 183.860 72.110 184.180 ;
        RECT 71.910 182.480 72.050 183.860 ;
        RECT 71.850 182.160 72.110 182.480 ;
        RECT 71.390 178.420 71.650 178.740 ;
        RECT 70.010 177.740 70.270 178.060 ;
        RECT 70.070 176.360 70.210 177.740 ;
        RECT 70.010 176.040 70.270 176.360 ;
        RECT 70.470 176.040 70.730 176.360 ;
        RECT 70.530 175.680 70.670 176.040 ;
        RECT 70.930 175.700 71.190 176.020 ;
        RECT 70.470 175.360 70.730 175.680 ;
        RECT 70.010 175.020 70.270 175.340 ;
        RECT 70.070 173.980 70.210 175.020 ;
        RECT 70.010 173.660 70.270 173.980 ;
        RECT 70.530 173.300 70.670 175.360 ;
        RECT 70.470 172.980 70.730 173.300 ;
        RECT 69.550 170.940 69.810 171.260 ;
        RECT 66.330 170.690 66.990 170.830 ;
        RECT 66.330 170.600 66.590 170.690 ;
        RECT 67.710 170.600 67.970 170.920 ;
        RECT 70.470 170.600 70.730 170.920 ;
        RECT 67.250 170.260 67.510 170.580 ;
        RECT 67.310 168.200 67.450 170.260 ;
        RECT 70.010 169.580 70.270 169.900 ;
        RECT 67.250 167.880 67.510 168.200 ;
        RECT 64.950 165.840 65.210 166.160 ;
        RECT 62.190 165.160 62.450 165.480 ;
        RECT 62.650 165.160 62.910 165.480 ;
        RECT 63.570 164.140 63.830 164.460 ;
        RECT 63.630 162.420 63.770 164.140 ;
        RECT 63.570 162.100 63.830 162.420 ;
        RECT 64.030 162.100 64.290 162.420 ;
        RECT 61.730 161.420 61.990 161.740 ;
        RECT 60.810 160.060 61.070 160.380 ;
        RECT 59.890 158.700 60.150 159.020 ;
        RECT 60.350 158.700 60.610 159.020 ;
        RECT 59.950 156.980 60.090 158.700 ;
        RECT 60.410 157.660 60.550 158.700 ;
        RECT 61.790 158.000 61.930 161.420 ;
        RECT 64.090 160.040 64.230 162.100 ;
        RECT 64.030 159.720 64.290 160.040 ;
        RECT 61.730 157.680 61.990 158.000 ;
        RECT 60.350 157.340 60.610 157.660 ;
        RECT 59.890 156.660 60.150 156.980 ;
        RECT 61.270 156.890 61.530 156.980 ;
        RECT 61.790 156.890 61.930 157.680 ;
        RECT 65.010 157.320 65.150 165.840 ;
        RECT 65.870 165.500 66.130 165.820 ;
        RECT 62.190 157.000 62.450 157.320 ;
        RECT 64.950 157.000 65.210 157.320 ;
        RECT 61.270 156.750 61.930 156.890 ;
        RECT 61.270 156.660 61.530 156.750 ;
        RECT 60.350 155.980 60.610 156.300 ;
        RECT 60.410 151.540 60.550 155.980 ;
        RECT 61.730 154.280 61.990 154.600 ;
        RECT 59.890 151.220 60.150 151.540 ;
        RECT 60.350 151.220 60.610 151.540 ;
        RECT 59.430 150.540 59.690 150.860 ;
        RECT 59.490 149.840 59.630 150.540 ;
        RECT 59.950 149.840 60.090 151.220 ;
        RECT 60.810 151.110 61.070 151.200 ;
        RECT 61.790 151.110 61.930 154.280 ;
        RECT 62.250 152.640 62.390 157.000 ;
        RECT 63.110 156.660 63.370 156.980 ;
        RECT 62.650 155.980 62.910 156.300 ;
        RECT 62.710 153.580 62.850 155.980 ;
        RECT 63.170 154.600 63.310 156.660 ;
        RECT 63.110 154.280 63.370 154.600 ;
        RECT 62.650 153.260 62.910 153.580 ;
        RECT 63.570 153.260 63.830 153.580 ;
        RECT 62.250 152.560 62.850 152.640 ;
        RECT 62.250 152.500 62.910 152.560 ;
        RECT 62.650 152.240 62.910 152.500 ;
        RECT 60.810 150.970 61.930 151.110 ;
        RECT 60.810 150.880 61.070 150.970 ;
        RECT 59.430 149.520 59.690 149.840 ;
        RECT 59.890 149.520 60.150 149.840 ;
        RECT 59.430 148.840 59.690 149.160 ;
        RECT 59.490 146.100 59.630 148.840 ;
        RECT 61.790 147.120 61.930 150.970 ;
        RECT 63.630 149.500 63.770 153.260 ;
        RECT 64.490 150.880 64.750 151.200 ;
        RECT 63.570 149.180 63.830 149.500 ;
        RECT 61.730 146.800 61.990 147.120 ;
        RECT 58.970 145.780 59.230 146.100 ;
        RECT 59.430 145.780 59.690 146.100 ;
        RECT 64.030 145.780 64.290 146.100 ;
        RECT 59.030 143.720 59.170 145.780 ;
        RECT 59.490 144.400 59.630 145.780 ;
        RECT 59.890 145.440 60.150 145.760 ;
        RECT 63.570 145.440 63.830 145.760 ;
        RECT 59.430 144.080 59.690 144.400 ;
        RECT 59.950 143.720 60.090 145.440 ;
        RECT 55.750 143.400 56.010 143.720 ;
        RECT 58.510 143.400 58.770 143.720 ;
        RECT 58.970 143.400 59.230 143.720 ;
        RECT 59.890 143.400 60.150 143.720 ;
        RECT 53.970 141.680 55.490 141.760 ;
        RECT 55.810 141.680 55.950 143.400 ;
        RECT 57.130 143.060 57.390 143.380 ;
        RECT 53.910 141.620 55.490 141.680 ;
        RECT 53.910 141.360 54.170 141.620 ;
        RECT 54.830 141.020 55.090 141.340 ;
        RECT 52.990 140.515 53.250 140.660 ;
        RECT 52.980 140.145 53.260 140.515 ;
        RECT 54.370 140.000 54.630 140.320 ;
        RECT 52.990 139.660 53.250 139.980 ;
        RECT 53.050 136.240 53.190 139.660 ;
        RECT 54.430 137.940 54.570 140.000 ;
        RECT 54.890 138.280 55.030 141.020 ;
        RECT 55.350 139.980 55.490 141.620 ;
        RECT 55.750 141.360 56.010 141.680 ;
        RECT 57.190 141.000 57.330 143.060 ;
        RECT 58.570 142.440 58.710 143.400 ;
        RECT 58.110 142.300 58.710 142.440 ;
        RECT 57.130 140.680 57.390 141.000 ;
        RECT 55.290 139.660 55.550 139.980 ;
        RECT 54.830 137.960 55.090 138.280 ;
        RECT 54.370 137.620 54.630 137.940 ;
        RECT 55.350 137.260 55.490 139.660 ;
        RECT 57.190 138.280 57.330 140.680 ;
        RECT 57.590 140.000 57.850 140.320 ;
        RECT 57.650 138.620 57.790 140.000 ;
        RECT 57.590 138.300 57.850 138.620 ;
        RECT 57.130 137.960 57.390 138.280 ;
        RECT 55.290 136.940 55.550 137.260 ;
        RECT 52.990 135.920 53.250 136.240 ;
        RECT 53.050 133.520 53.190 135.920 ;
        RECT 52.990 133.200 53.250 133.520 ;
        RECT 53.050 129.100 53.190 133.200 ;
        RECT 57.190 132.920 57.330 137.960 ;
        RECT 56.730 132.840 57.330 132.920 ;
        RECT 56.670 132.780 57.330 132.840 ;
        RECT 56.670 132.520 56.930 132.780 ;
        RECT 53.910 131.500 54.170 131.820 ;
        RECT 53.970 129.440 54.110 131.500 ;
        RECT 56.730 129.780 56.870 132.520 ;
        RECT 56.670 129.460 56.930 129.780 ;
        RECT 53.910 129.120 54.170 129.440 ;
        RECT 52.990 128.780 53.250 129.100 ;
        RECT 55.290 123.340 55.550 123.660 ;
        RECT 55.350 121.960 55.490 123.340 ;
        RECT 56.730 122.300 56.870 129.460 ;
        RECT 56.670 121.980 56.930 122.300 ;
        RECT 55.290 121.640 55.550 121.960 ;
        RECT 56.730 118.900 56.870 121.980 ;
        RECT 56.670 118.580 56.930 118.900 ;
        RECT 52.530 118.240 52.790 118.560 ;
        RECT 55.750 117.900 56.010 118.220 ;
        RECT 50.230 116.200 50.490 116.520 ;
        RECT 50.290 107.340 50.430 116.200 ;
        RECT 55.810 113.120 55.950 117.900 ;
        RECT 56.210 114.160 56.470 114.480 ;
        RECT 55.750 112.800 56.010 113.120 ;
        RECT 54.830 112.460 55.090 112.780 ;
        RECT 54.890 111.080 55.030 112.460 ;
        RECT 55.810 111.080 55.950 112.800 ;
        RECT 56.270 111.080 56.410 114.160 ;
        RECT 56.730 113.800 56.870 118.580 ;
        RECT 56.670 113.480 56.930 113.800 ;
        RECT 54.830 110.760 55.090 111.080 ;
        RECT 55.750 110.760 56.010 111.080 ;
        RECT 56.210 110.760 56.470 111.080 ;
        RECT 50.230 107.020 50.490 107.340 ;
        RECT 49.770 97.160 50.030 97.480 ;
        RECT 50.290 93.650 50.430 107.020 ;
        RECT 54.890 105.980 55.030 110.760 ;
        RECT 55.290 110.420 55.550 110.740 ;
        RECT 55.350 107.680 55.490 110.420 ;
        RECT 57.650 109.040 57.790 138.300 ;
        RECT 58.110 135.560 58.250 142.300 ;
        RECT 59.430 139.720 59.690 139.980 ;
        RECT 59.950 139.720 60.090 143.400 ;
        RECT 60.350 140.680 60.610 141.000 ;
        RECT 59.430 139.660 60.090 139.720 ;
        RECT 59.490 139.580 60.090 139.660 ;
        RECT 58.510 138.640 58.770 138.960 ;
        RECT 58.570 135.560 58.710 138.640 ;
        RECT 58.050 135.240 58.310 135.560 ;
        RECT 58.510 135.240 58.770 135.560 ;
        RECT 59.490 130.800 59.630 139.580 ;
        RECT 59.890 138.300 60.150 138.620 ;
        RECT 59.950 135.220 60.090 138.300 ;
        RECT 60.410 135.220 60.550 140.680 ;
        RECT 62.190 140.340 62.450 140.660 ;
        RECT 62.250 135.220 62.390 140.340 ;
        RECT 63.630 140.320 63.770 145.440 ;
        RECT 64.090 144.400 64.230 145.780 ;
        RECT 64.030 144.080 64.290 144.400 ;
        RECT 63.570 140.000 63.830 140.320 ;
        RECT 64.550 139.980 64.690 150.880 ;
        RECT 65.010 149.500 65.150 157.000 ;
        RECT 65.410 156.660 65.670 156.980 ;
        RECT 65.470 154.600 65.610 156.660 ;
        RECT 65.410 154.280 65.670 154.600 ;
        RECT 64.950 149.180 65.210 149.500 ;
        RECT 65.470 149.160 65.610 154.280 ;
        RECT 65.410 148.840 65.670 149.160 ;
        RECT 65.930 145.760 66.070 165.500 ;
        RECT 67.310 157.320 67.450 167.880 ;
        RECT 68.630 162.100 68.890 162.420 ;
        RECT 69.550 162.100 69.810 162.420 ;
        RECT 68.690 157.400 68.830 162.100 ;
        RECT 69.610 159.360 69.750 162.100 ;
        RECT 69.550 159.040 69.810 159.360 ;
        RECT 67.250 157.000 67.510 157.320 ;
        RECT 68.690 157.260 69.750 157.400 ;
        RECT 67.310 154.600 67.450 157.000 ;
        RECT 68.630 156.660 68.890 156.980 ;
        RECT 68.690 154.600 68.830 156.660 ;
        RECT 69.610 154.940 69.750 157.260 ;
        RECT 69.550 154.620 69.810 154.940 ;
        RECT 67.250 154.280 67.510 154.600 ;
        RECT 68.630 154.280 68.890 154.600 ;
        RECT 68.690 153.920 68.830 154.280 ;
        RECT 68.630 153.600 68.890 153.920 ;
        RECT 69.610 153.580 69.750 154.620 ;
        RECT 68.170 153.260 68.430 153.580 ;
        RECT 69.550 153.260 69.810 153.580 ;
        RECT 68.230 151.540 68.370 153.260 ;
        RECT 66.330 151.220 66.590 151.540 ;
        RECT 68.170 151.220 68.430 151.540 ;
        RECT 66.390 149.160 66.530 151.220 ;
        RECT 67.250 150.880 67.510 151.200 ;
        RECT 67.310 149.160 67.450 150.880 ;
        RECT 66.330 148.840 66.590 149.160 ;
        RECT 67.250 148.840 67.510 149.160 ;
        RECT 66.790 148.500 67.050 148.820 ;
        RECT 65.870 145.440 66.130 145.760 ;
        RECT 66.850 143.720 66.990 148.500 ;
        RECT 68.230 146.520 68.370 151.220 ;
        RECT 70.070 149.500 70.210 169.580 ;
        RECT 70.530 168.880 70.670 170.600 ;
        RECT 70.470 168.560 70.730 168.880 ;
        RECT 70.990 167.520 71.130 175.700 ;
        RECT 71.450 175.340 71.590 178.420 ;
        RECT 71.910 176.360 72.050 182.160 ;
        RECT 72.310 176.380 72.570 176.700 ;
        RECT 71.850 176.040 72.110 176.360 ;
        RECT 71.390 175.020 71.650 175.340 ;
        RECT 71.910 174.320 72.050 176.040 ;
        RECT 71.850 174.000 72.110 174.320 ;
        RECT 71.390 173.660 71.650 173.980 ;
        RECT 71.910 173.835 72.050 174.000 ;
        RECT 71.450 172.620 71.590 173.660 ;
        RECT 71.840 173.465 72.120 173.835 ;
        RECT 72.370 173.300 72.510 176.380 ;
        RECT 73.230 176.040 73.490 176.360 ;
        RECT 73.290 173.980 73.430 176.040 ;
        RECT 75.070 174.000 75.330 174.320 ;
        RECT 73.230 173.660 73.490 173.980 ;
        RECT 72.310 172.980 72.570 173.300 ;
        RECT 73.290 172.620 73.430 173.660 ;
        RECT 75.130 172.960 75.270 174.000 ;
        RECT 76.050 173.640 76.190 184.200 ;
        RECT 100.970 182.410 102.630 184.070 ;
        RECT 123.240 180.480 125.770 180.490 ;
        RECT 100.360 180.380 108.770 180.390 ;
        RECT 100.360 180.100 108.805 180.380 ;
        RECT 123.240 180.200 125.805 180.480 ;
        RECT 123.240 180.190 125.770 180.200 ;
        RECT 100.360 180.090 108.770 180.100 ;
        RECT 75.990 173.320 76.250 173.640 ;
        RECT 75.070 172.640 75.330 172.960 ;
        RECT 71.390 172.300 71.650 172.620 ;
        RECT 71.850 172.300 72.110 172.620 ;
        RECT 72.310 172.300 72.570 172.620 ;
        RECT 73.230 172.300 73.490 172.620 ;
        RECT 71.910 168.880 72.050 172.300 ;
        RECT 71.850 168.560 72.110 168.880 ;
        RECT 72.370 167.520 72.510 172.300 ;
        RECT 76.050 170.920 76.190 173.320 ;
        RECT 75.990 170.600 76.250 170.920 ;
        RECT 76.050 167.860 76.190 170.600 ;
        RECT 75.990 167.540 76.250 167.860 ;
        RECT 70.930 167.200 71.190 167.520 ;
        RECT 72.310 167.200 72.570 167.520 ;
        RECT 76.050 165.820 76.190 167.540 ;
        RECT 75.990 165.500 76.250 165.820 ;
        RECT 70.930 162.100 71.190 162.420 ;
        RECT 71.390 162.100 71.650 162.420 ;
        RECT 70.470 159.040 70.730 159.360 ;
        RECT 70.530 158.000 70.670 159.040 ;
        RECT 70.470 157.680 70.730 158.000 ;
        RECT 70.470 156.660 70.730 156.980 ;
        RECT 70.530 155.280 70.670 156.660 ;
        RECT 70.470 154.960 70.730 155.280 ;
        RECT 70.990 152.220 71.130 162.100 ;
        RECT 71.450 159.700 71.590 162.100 ;
        RECT 76.050 162.080 76.190 165.500 ;
        RECT 76.050 161.940 77.110 162.080 ;
        RECT 73.230 161.420 73.490 161.740 ;
        RECT 73.290 160.380 73.430 161.420 ;
        RECT 72.310 160.060 72.570 160.380 ;
        RECT 73.230 160.060 73.490 160.380 ;
        RECT 74.150 160.060 74.410 160.380 ;
        RECT 71.390 159.380 71.650 159.700 ;
        RECT 71.390 158.700 71.650 159.020 ;
        RECT 71.450 157.660 71.590 158.700 ;
        RECT 71.390 157.340 71.650 157.660 ;
        RECT 70.930 151.900 71.190 152.220 ;
        RECT 70.930 150.540 71.190 150.860 ;
        RECT 70.010 149.180 70.270 149.500 ;
        RECT 70.470 148.840 70.730 149.160 ;
        RECT 70.010 148.500 70.270 148.820 ;
        RECT 67.770 146.380 68.370 146.520 ;
        RECT 64.950 143.400 65.210 143.720 ;
        RECT 66.790 143.400 67.050 143.720 ;
        RECT 65.010 140.660 65.150 143.400 ;
        RECT 64.950 140.340 65.210 140.660 ;
        RECT 65.410 140.000 65.670 140.320 ;
        RECT 64.490 139.660 64.750 139.980 ;
        RECT 64.550 138.870 64.690 139.660 ;
        RECT 64.550 138.730 65.150 138.870 ;
        RECT 64.490 137.960 64.750 138.280 ;
        RECT 64.550 136.240 64.690 137.960 ;
        RECT 65.010 137.600 65.150 138.730 ;
        RECT 64.950 137.280 65.210 137.600 ;
        RECT 65.010 136.240 65.150 137.280 ;
        RECT 64.490 135.920 64.750 136.240 ;
        RECT 64.950 135.920 65.210 136.240 ;
        RECT 63.570 135.580 63.830 135.900 ;
        RECT 59.890 134.900 60.150 135.220 ;
        RECT 60.350 134.900 60.610 135.220 ;
        RECT 62.190 134.900 62.450 135.220 ;
        RECT 59.890 134.220 60.150 134.540 ;
        RECT 59.950 133.180 60.090 134.220 ;
        RECT 62.250 133.520 62.390 134.900 ;
        RECT 62.190 133.200 62.450 133.520 ;
        RECT 59.890 132.860 60.150 133.180 ;
        RECT 59.430 130.480 59.690 130.800 ;
        RECT 63.630 129.780 63.770 135.580 ;
        RECT 65.470 134.880 65.610 140.000 ;
        RECT 66.850 139.980 66.990 143.400 ;
        RECT 67.770 140.320 67.910 146.380 ;
        RECT 68.170 145.440 68.430 145.760 ;
        RECT 69.550 145.440 69.810 145.760 ;
        RECT 68.230 143.380 68.370 145.440 ;
        RECT 68.170 143.060 68.430 143.380 ;
        RECT 67.710 140.000 67.970 140.320 ;
        RECT 66.790 139.890 67.050 139.980 ;
        RECT 66.390 139.750 67.050 139.890 ;
        RECT 66.390 134.880 66.530 139.750 ;
        RECT 66.790 139.660 67.050 139.750 ;
        RECT 66.790 137.960 67.050 138.280 ;
        RECT 66.850 136.240 66.990 137.960 ;
        RECT 67.250 136.940 67.510 137.260 ;
        RECT 66.790 135.920 67.050 136.240 ;
        RECT 65.410 134.560 65.670 134.880 ;
        RECT 66.330 134.560 66.590 134.880 ;
        RECT 66.390 133.520 66.530 134.560 ;
        RECT 66.330 133.200 66.590 133.520 ;
        RECT 66.330 132.520 66.590 132.840 ;
        RECT 66.390 130.800 66.530 132.520 ;
        RECT 66.330 130.480 66.590 130.800 ;
        RECT 67.310 130.120 67.450 136.940 ;
        RECT 67.770 136.240 67.910 140.000 ;
        RECT 67.710 135.920 67.970 136.240 ;
        RECT 68.230 133.180 68.370 143.060 ;
        RECT 69.610 138.960 69.750 145.440 ;
        RECT 69.550 138.640 69.810 138.960 ;
        RECT 70.070 138.620 70.210 148.500 ;
        RECT 70.530 140.515 70.670 148.840 ;
        RECT 70.990 148.820 71.130 150.540 ;
        RECT 71.450 149.840 71.590 157.340 ;
        RECT 71.850 155.980 72.110 156.300 ;
        RECT 71.390 149.520 71.650 149.840 ;
        RECT 71.910 149.160 72.050 155.980 ;
        RECT 72.370 154.940 72.510 160.060 ;
        RECT 72.770 157.680 73.030 158.000 ;
        RECT 72.830 156.980 72.970 157.680 ;
        RECT 73.690 157.340 73.950 157.660 ;
        RECT 73.750 156.980 73.890 157.340 ;
        RECT 72.770 156.660 73.030 156.980 ;
        RECT 73.690 156.660 73.950 156.980 ;
        RECT 72.310 154.620 72.570 154.940 ;
        RECT 72.370 154.260 72.510 154.620 ;
        RECT 72.310 153.940 72.570 154.260 ;
        RECT 72.310 151.900 72.570 152.220 ;
        RECT 71.850 148.840 72.110 149.160 ;
        RECT 70.930 148.500 71.190 148.820 ;
        RECT 72.370 146.100 72.510 151.900 ;
        RECT 72.830 151.280 72.970 156.660 ;
        RECT 73.230 154.960 73.490 155.280 ;
        RECT 73.290 154.000 73.430 154.960 ;
        RECT 73.290 153.860 73.890 154.000 ;
        RECT 73.750 151.540 73.890 153.860 ;
        RECT 72.830 151.140 73.430 151.280 ;
        RECT 73.690 151.220 73.950 151.540 ;
        RECT 73.290 146.780 73.430 151.140 ;
        RECT 73.690 148.500 73.950 148.820 ;
        RECT 73.230 146.460 73.490 146.780 ;
        RECT 73.750 146.440 73.890 148.500 ;
        RECT 73.690 146.120 73.950 146.440 ;
        RECT 72.310 145.780 72.570 146.100 ;
        RECT 74.210 145.760 74.350 160.060 ;
        RECT 76.970 159.020 77.110 161.940 ;
        RECT 76.910 158.700 77.170 159.020 ;
        RECT 78.750 158.700 79.010 159.020 ;
        RECT 76.970 157.320 77.110 158.700 ;
        RECT 76.450 157.000 76.710 157.320 ;
        RECT 76.910 157.000 77.170 157.320 ;
        RECT 75.070 153.940 75.330 154.260 ;
        RECT 74.610 153.600 74.870 153.920 ;
        RECT 74.670 151.540 74.810 153.600 ;
        RECT 74.610 151.220 74.870 151.540 ;
        RECT 75.130 145.760 75.270 153.940 ;
        RECT 76.510 153.920 76.650 157.000 ;
        RECT 76.910 155.980 77.170 156.300 ;
        RECT 76.970 154.940 77.110 155.980 ;
        RECT 76.910 154.620 77.170 154.940 ;
        RECT 78.810 154.600 78.950 158.700 ;
        RECT 78.750 154.280 79.010 154.600 ;
        RECT 76.450 153.600 76.710 153.920 ;
        RECT 80.590 151.220 80.850 151.540 ;
        RECT 80.650 149.840 80.790 151.220 ;
        RECT 80.590 149.520 80.850 149.840 ;
        RECT 75.530 145.780 75.790 146.100 ;
        RECT 74.150 145.440 74.410 145.760 ;
        RECT 75.070 145.440 75.330 145.760 ;
        RECT 70.930 145.100 71.190 145.420 ;
        RECT 70.990 144.060 71.130 145.100 ;
        RECT 75.130 144.400 75.270 145.440 ;
        RECT 75.070 144.080 75.330 144.400 ;
        RECT 70.930 143.740 71.190 144.060 ;
        RECT 70.460 140.145 70.740 140.515 ;
        RECT 68.630 138.300 68.890 138.620 ;
        RECT 70.010 138.300 70.270 138.620 ;
        RECT 68.690 137.940 68.830 138.300 ;
        RECT 68.630 137.620 68.890 137.940 ;
        RECT 70.010 137.680 70.270 137.940 ;
        RECT 70.530 137.680 70.670 140.145 ;
        RECT 75.590 138.280 75.730 145.780 ;
        RECT 75.530 137.960 75.790 138.280 ;
        RECT 75.990 137.960 76.250 138.280 ;
        RECT 70.010 137.620 70.670 137.680 ;
        RECT 71.850 137.620 72.110 137.940 ;
        RECT 68.170 132.860 68.430 133.180 ;
        RECT 68.690 130.460 68.830 137.620 ;
        RECT 70.070 137.540 70.670 137.620 ;
        RECT 71.910 136.240 72.050 137.620 ;
        RECT 71.850 135.920 72.110 136.240 ;
        RECT 76.050 134.790 76.190 137.960 ;
        RECT 75.130 134.650 76.190 134.790 ;
        RECT 75.130 133.180 75.270 134.650 ;
        RECT 72.770 132.860 73.030 133.180 ;
        RECT 75.070 132.860 75.330 133.180 ;
        RECT 68.630 130.140 68.890 130.460 ;
        RECT 67.250 129.800 67.510 130.120 ;
        RECT 63.570 129.460 63.830 129.780 ;
        RECT 58.510 124.020 58.770 124.340 ;
        RECT 66.330 124.020 66.590 124.340 ;
        RECT 66.790 124.020 67.050 124.340 ;
        RECT 67.710 124.250 67.970 124.340 ;
        RECT 67.310 124.110 67.970 124.250 ;
        RECT 58.570 117.200 58.710 124.020 ;
        RECT 64.490 123.680 64.750 124.000 ;
        RECT 60.350 123.340 60.610 123.660 ;
        RECT 60.410 118.900 60.550 123.340 ;
        RECT 60.350 118.580 60.610 118.900 ;
        RECT 58.510 116.880 58.770 117.200 ;
        RECT 64.550 116.520 64.690 123.680 ;
        RECT 65.870 121.640 66.130 121.960 ;
        RECT 65.930 119.920 66.070 121.640 ;
        RECT 66.390 119.920 66.530 124.020 ;
        RECT 65.870 119.600 66.130 119.920 ;
        RECT 66.330 119.600 66.590 119.920 ;
        RECT 64.950 118.240 65.210 118.560 ;
        RECT 65.010 117.200 65.150 118.240 ;
        RECT 66.850 117.200 66.990 124.020 ;
        RECT 67.310 120.940 67.450 124.110 ;
        RECT 67.710 124.020 67.970 124.110 ;
        RECT 72.830 121.960 72.970 132.860 ;
        RECT 72.310 121.640 72.570 121.960 ;
        RECT 72.770 121.640 73.030 121.960 ;
        RECT 75.530 121.640 75.790 121.960 ;
        RECT 67.250 120.620 67.510 120.940 ;
        RECT 67.310 118.900 67.450 120.620 ;
        RECT 72.370 119.920 72.510 121.640 ;
        RECT 72.310 119.600 72.570 119.920 ;
        RECT 67.250 118.580 67.510 118.900 ;
        RECT 70.470 118.580 70.730 118.900 ;
        RECT 71.850 118.580 72.110 118.900 ;
        RECT 64.950 116.880 65.210 117.200 ;
        RECT 66.790 116.880 67.050 117.200 ;
        RECT 64.490 116.200 64.750 116.520 ;
        RECT 67.250 116.200 67.510 116.520 ;
        RECT 68.630 116.200 68.890 116.520 ;
        RECT 64.550 113.780 64.690 116.200 ;
        RECT 63.630 113.640 64.690 113.780 ;
        RECT 63.110 113.140 63.370 113.460 ;
        RECT 63.170 111.760 63.310 113.140 ;
        RECT 63.630 112.780 63.770 113.640 ;
        RECT 67.310 112.780 67.450 116.200 ;
        RECT 68.690 114.140 68.830 116.200 ;
        RECT 70.530 116.180 70.670 118.580 ;
        RECT 71.390 118.240 71.650 118.560 ;
        RECT 70.470 115.860 70.730 116.180 ;
        RECT 68.630 113.820 68.890 114.140 ;
        RECT 63.570 112.460 63.830 112.780 ;
        RECT 65.410 112.460 65.670 112.780 ;
        RECT 67.250 112.460 67.510 112.780 ;
        RECT 67.710 112.460 67.970 112.780 ;
        RECT 63.630 111.760 63.770 112.460 ;
        RECT 63.110 111.440 63.370 111.760 ;
        RECT 63.570 111.440 63.830 111.760 ;
        RECT 62.190 110.760 62.450 111.080 ;
        RECT 62.250 109.040 62.390 110.760 ;
        RECT 65.470 110.740 65.610 112.460 ;
        RECT 65.410 110.420 65.670 110.740 ;
        RECT 66.330 110.420 66.590 110.740 ;
        RECT 62.650 110.080 62.910 110.400 ;
        RECT 57.590 108.720 57.850 109.040 ;
        RECT 62.190 108.720 62.450 109.040 ;
        RECT 55.750 108.380 56.010 108.700 ;
        RECT 55.290 107.360 55.550 107.680 ;
        RECT 54.830 105.660 55.090 105.980 ;
        RECT 52.530 104.980 52.790 105.300 ;
        RECT 53.910 104.980 54.170 105.300 ;
        RECT 50.690 104.300 50.950 104.620 ;
        RECT 50.750 97.140 50.890 104.300 ;
        RECT 52.590 100.880 52.730 104.980 ;
        RECT 53.970 103.600 54.110 104.980 ;
        RECT 53.910 103.280 54.170 103.600 ;
        RECT 52.530 100.560 52.790 100.880 ;
        RECT 50.690 96.820 50.950 97.140 ;
        RECT 53.970 96.800 54.110 103.280 ;
        RECT 54.370 101.920 54.630 102.240 ;
        RECT 54.430 99.180 54.570 101.920 ;
        RECT 54.890 100.200 55.030 105.660 ;
        RECT 55.350 104.620 55.490 107.360 ;
        RECT 55.810 106.320 55.950 108.380 ;
        RECT 55.750 106.000 56.010 106.320 ;
        RECT 55.290 104.300 55.550 104.620 ;
        RECT 55.350 100.540 55.490 104.300 ;
        RECT 55.750 102.260 56.010 102.580 ;
        RECT 55.290 100.220 55.550 100.540 ;
        RECT 54.830 99.880 55.090 100.200 ;
        RECT 55.810 99.520 55.950 102.260 ;
        RECT 55.750 99.200 56.010 99.520 ;
        RECT 54.370 98.860 54.630 99.180 ;
        RECT 54.430 97.480 54.570 98.860 ;
        RECT 54.370 97.160 54.630 97.480 ;
        RECT 53.910 96.480 54.170 96.800 ;
        RECT 54.430 94.420 54.570 97.160 ;
        RECT 54.370 94.100 54.630 94.420 ;
        RECT 55.810 93.740 55.950 99.200 ;
        RECT 57.130 97.160 57.390 97.480 ;
        RECT 49.830 93.510 50.430 93.650 ;
        RECT 49.830 86.940 49.970 93.510 ;
        RECT 55.750 93.420 56.010 93.740 ;
        RECT 51.150 91.040 51.410 91.360 ;
        RECT 51.210 90.000 51.350 91.040 ;
        RECT 50.690 89.680 50.950 90.000 ;
        RECT 51.150 89.680 51.410 90.000 ;
        RECT 50.750 89.320 50.890 89.680 ;
        RECT 55.290 89.340 55.550 89.660 ;
        RECT 50.690 89.000 50.950 89.320 ;
        RECT 49.770 86.620 50.030 86.940 ;
        RECT 49.830 75.120 49.970 86.620 ;
        RECT 50.750 80.480 50.890 89.000 ;
        RECT 52.070 88.320 52.330 88.640 ;
        RECT 51.610 85.600 51.870 85.920 ;
        RECT 51.150 85.260 51.410 85.580 ;
        RECT 51.210 84.220 51.350 85.260 ;
        RECT 51.150 83.900 51.410 84.220 ;
        RECT 51.670 81.840 51.810 85.600 ;
        RECT 51.610 81.520 51.870 81.840 ;
        RECT 50.690 80.160 50.950 80.480 ;
        RECT 50.230 79.820 50.490 80.140 ;
        RECT 50.290 75.720 50.430 79.820 ;
        RECT 50.690 78.460 50.950 78.780 ;
        RECT 50.750 76.400 50.890 78.460 ;
        RECT 51.610 78.120 51.870 78.440 ;
        RECT 51.150 77.100 51.410 77.420 ;
        RECT 50.690 76.080 50.950 76.400 ;
        RECT 50.230 75.400 50.490 75.720 ;
        RECT 49.830 74.980 50.430 75.120 ;
        RECT 49.770 66.900 50.030 67.220 ;
        RECT 49.830 62.800 49.970 66.900 ;
        RECT 50.290 64.500 50.430 74.980 ;
        RECT 50.750 70.280 50.890 76.080 ;
        RECT 51.210 75.380 51.350 77.100 ;
        RECT 51.670 76.400 51.810 78.120 ;
        RECT 51.610 76.080 51.870 76.400 ;
        RECT 51.150 75.060 51.410 75.380 ;
        RECT 50.690 69.960 50.950 70.280 ;
        RECT 51.210 64.840 51.350 75.060 ;
        RECT 52.130 73.340 52.270 88.320 ;
        RECT 54.370 86.280 54.630 86.600 ;
        RECT 52.990 85.260 53.250 85.580 ;
        RECT 53.050 81.840 53.190 85.260 ;
        RECT 52.990 81.520 53.250 81.840 ;
        RECT 53.910 79.820 54.170 80.140 ;
        RECT 52.990 74.380 53.250 74.700 ;
        RECT 52.070 73.020 52.330 73.340 ;
        RECT 52.130 72.660 52.270 73.020 ;
        RECT 52.070 72.340 52.330 72.660 ;
        RECT 53.050 68.240 53.190 74.380 ;
        RECT 53.970 70.280 54.110 79.820 ;
        RECT 54.430 78.780 54.570 86.280 ;
        RECT 55.350 84.560 55.490 89.340 ;
        RECT 55.810 88.980 55.950 93.420 ;
        RECT 55.750 88.660 56.010 88.980 ;
        RECT 55.810 86.600 55.950 88.660 ;
        RECT 55.750 86.280 56.010 86.600 ;
        RECT 55.290 84.240 55.550 84.560 ;
        RECT 54.370 78.460 54.630 78.780 ;
        RECT 54.430 75.720 54.570 78.460 ;
        RECT 54.370 75.400 54.630 75.720 ;
        RECT 54.430 72.230 54.570 75.400 ;
        RECT 55.810 75.380 55.950 86.280 ;
        RECT 56.210 85.260 56.470 85.580 ;
        RECT 56.270 84.560 56.410 85.260 ;
        RECT 56.210 84.240 56.470 84.560 ;
        RECT 57.190 81.160 57.330 97.160 ;
        RECT 57.130 80.840 57.390 81.160 ;
        RECT 56.670 80.500 56.930 80.820 ;
        RECT 56.730 79.120 56.870 80.500 ;
        RECT 56.670 78.800 56.930 79.120 ;
        RECT 55.750 75.060 56.010 75.380 ;
        RECT 56.210 72.680 56.470 73.000 ;
        RECT 54.830 72.230 55.090 72.320 ;
        RECT 54.430 72.090 55.090 72.230 ;
        RECT 54.830 72.000 55.090 72.090 ;
        RECT 53.910 69.960 54.170 70.280 ;
        RECT 55.750 69.280 56.010 69.600 ;
        RECT 55.810 68.240 55.950 69.280 ;
        RECT 52.990 67.920 53.250 68.240 ;
        RECT 55.750 67.920 56.010 68.240 ;
        RECT 51.610 66.560 51.870 66.880 ;
        RECT 51.150 64.520 51.410 64.840 ;
        RECT 50.230 64.180 50.490 64.500 ;
        RECT 51.150 63.500 51.410 63.820 ;
        RECT 49.770 62.480 50.030 62.800 ;
        RECT 49.830 59.060 49.970 62.480 ;
        RECT 51.210 61.780 51.350 63.500 ;
        RECT 51.670 62.800 51.810 66.560 ;
        RECT 53.910 63.840 54.170 64.160 ;
        RECT 53.970 62.800 54.110 63.840 ;
        RECT 51.610 62.480 51.870 62.800 ;
        RECT 53.910 62.480 54.170 62.800 ;
        RECT 51.150 61.460 51.410 61.780 ;
        RECT 54.370 61.460 54.630 61.780 ;
        RECT 49.770 58.740 50.030 59.060 ;
        RECT 53.910 58.400 54.170 58.720 ;
        RECT 53.970 57.020 54.110 58.400 ;
        RECT 53.910 56.700 54.170 57.020 ;
        RECT 52.070 56.020 52.330 56.340 ;
        RECT 53.450 56.020 53.710 56.340 ;
        RECT 51.150 55.340 51.410 55.660 ;
        RECT 50.230 53.300 50.490 53.620 ;
        RECT 49.310 50.240 49.570 50.560 ;
        RECT 49.370 48.520 49.510 50.240 ;
        RECT 49.310 48.200 49.570 48.520 ;
        RECT 49.770 42.080 50.030 42.400 ;
        RECT 49.830 40.020 49.970 42.080 ;
        RECT 49.770 39.700 50.030 40.020 ;
        RECT 49.310 39.020 49.570 39.340 ;
        RECT 49.370 31.600 49.510 39.020 ;
        RECT 49.830 37.640 49.970 39.700 ;
        RECT 49.770 37.320 50.030 37.640 ;
        RECT 49.770 35.280 50.030 35.600 ;
        RECT 49.830 32.280 49.970 35.280 ;
        RECT 50.290 32.880 50.430 53.300 ;
        RECT 51.210 51.580 51.350 55.340 ;
        RECT 51.150 51.260 51.410 51.580 ;
        RECT 51.610 48.880 51.870 49.200 ;
        RECT 51.670 45.800 51.810 48.880 ;
        RECT 50.690 45.480 50.950 45.800 ;
        RECT 51.610 45.480 51.870 45.800 ;
        RECT 50.750 42.740 50.890 45.480 ;
        RECT 51.670 43.760 51.810 45.480 ;
        RECT 51.610 43.440 51.870 43.760 ;
        RECT 50.690 42.420 50.950 42.740 ;
        RECT 50.750 34.920 50.890 42.420 ;
        RECT 51.670 41.040 51.810 43.440 ;
        RECT 51.610 40.720 51.870 41.040 ;
        RECT 51.670 39.340 51.810 40.720 ;
        RECT 51.150 39.020 51.410 39.340 ;
        RECT 51.610 39.020 51.870 39.340 ;
        RECT 50.690 34.600 50.950 34.920 ;
        RECT 51.210 34.240 51.350 39.020 ;
        RECT 51.670 34.920 51.810 39.020 ;
        RECT 51.610 34.600 51.870 34.920 ;
        RECT 51.150 33.920 51.410 34.240 ;
        RECT 50.230 32.560 50.490 32.880 ;
        RECT 49.830 32.140 50.430 32.280 ;
        RECT 50.290 31.860 50.430 32.140 ;
        RECT 50.690 31.880 50.950 32.200 ;
        RECT 49.370 31.520 49.970 31.600 ;
        RECT 50.230 31.540 50.490 31.860 ;
        RECT 49.370 31.460 50.030 31.520 ;
        RECT 49.770 31.200 50.030 31.460 ;
        RECT 50.290 24.380 50.430 31.540 ;
        RECT 50.750 25.740 50.890 31.880 ;
        RECT 51.210 31.180 51.350 33.920 ;
        RECT 51.150 30.860 51.410 31.180 ;
        RECT 51.150 29.160 51.410 29.480 ;
        RECT 51.210 27.100 51.350 29.160 ;
        RECT 51.150 26.780 51.410 27.100 ;
        RECT 50.690 25.420 50.950 25.740 ;
        RECT 50.230 24.060 50.490 24.380 ;
        RECT 48.850 23.040 49.110 23.360 ;
        RECT 49.310 20.660 49.570 20.980 ;
        RECT 49.370 16.560 49.510 20.660 ;
        RECT 52.130 17.580 52.270 56.020 ;
        RECT 53.510 54.640 53.650 56.020 ;
        RECT 53.970 54.640 54.110 56.700 ;
        RECT 54.430 56.340 54.570 61.460 ;
        RECT 56.270 60.080 56.410 72.680 ;
        RECT 57.190 66.540 57.330 80.840 ;
        RECT 57.650 73.680 57.790 108.720 ;
        RECT 62.710 106.320 62.850 110.080 ;
        RECT 64.490 109.740 64.750 110.060 ;
        RECT 64.030 108.720 64.290 109.040 ;
        RECT 62.650 106.000 62.910 106.320 ;
        RECT 64.090 105.640 64.230 108.720 ;
        RECT 64.030 105.320 64.290 105.640 ;
        RECT 64.550 105.040 64.690 109.740 ;
        RECT 65.470 108.020 65.610 110.420 ;
        RECT 65.410 107.700 65.670 108.020 ;
        RECT 65.870 106.000 66.130 106.320 ;
        RECT 65.410 105.660 65.670 105.980 ;
        RECT 64.090 104.900 64.690 105.040 ;
        RECT 64.090 104.620 64.230 104.900 ;
        RECT 60.350 104.300 60.610 104.620 ;
        RECT 64.030 104.300 64.290 104.620 ;
        RECT 60.410 102.920 60.550 104.300 ;
        RECT 60.350 102.600 60.610 102.920 ;
        RECT 63.570 102.260 63.830 102.580 ;
        RECT 63.630 100.880 63.770 102.260 ;
        RECT 63.570 100.560 63.830 100.880 ;
        RECT 60.350 96.820 60.610 97.140 ;
        RECT 60.410 95.440 60.550 96.820 ;
        RECT 60.350 95.120 60.610 95.440 ;
        RECT 63.630 88.300 63.770 100.560 ;
        RECT 64.090 97.480 64.230 104.300 ;
        RECT 65.470 102.580 65.610 105.660 ;
        RECT 65.930 102.580 66.070 106.000 ;
        RECT 66.390 105.980 66.530 110.420 ;
        RECT 67.250 110.080 67.510 110.400 ;
        RECT 67.310 108.700 67.450 110.080 ;
        RECT 67.770 109.040 67.910 112.460 ;
        RECT 68.170 110.760 68.430 111.080 ;
        RECT 67.710 108.720 67.970 109.040 ;
        RECT 67.250 108.380 67.510 108.700 ;
        RECT 67.250 107.700 67.510 108.020 ;
        RECT 68.230 107.760 68.370 110.760 ;
        RECT 68.690 110.480 68.830 113.820 ;
        RECT 69.090 113.140 69.350 113.460 ;
        RECT 69.150 111.760 69.290 113.140 ;
        RECT 69.550 112.800 69.810 113.120 ;
        RECT 69.090 111.440 69.350 111.760 ;
        RECT 69.610 111.420 69.750 112.800 ;
        RECT 69.550 111.100 69.810 111.420 ;
        RECT 68.690 110.400 69.290 110.480 ;
        RECT 68.690 110.340 69.350 110.400 ;
        RECT 69.090 110.080 69.350 110.340 ;
        RECT 70.530 108.700 70.670 115.860 ;
        RECT 71.450 113.460 71.590 118.240 ;
        RECT 71.390 113.140 71.650 113.460 ;
        RECT 71.910 111.420 72.050 118.580 ;
        RECT 75.590 113.460 75.730 121.640 ;
        RECT 87.030 116.200 87.290 116.520 ;
        RECT 77.830 115.180 78.090 115.500 ;
        RECT 75.530 113.140 75.790 113.460 ;
        RECT 73.230 112.800 73.490 113.120 ;
        RECT 72.770 112.460 73.030 112.780 ;
        RECT 71.850 111.100 72.110 111.420 ;
        RECT 72.830 110.740 72.970 112.460 ;
        RECT 72.770 110.420 73.030 110.740 ;
        RECT 70.930 110.080 71.190 110.400 ;
        RECT 70.990 109.040 71.130 110.080 ;
        RECT 73.290 110.060 73.430 112.800 ;
        RECT 73.690 110.760 73.950 111.080 ;
        RECT 73.230 109.740 73.490 110.060 ;
        RECT 73.750 109.040 73.890 110.760 ;
        RECT 77.370 110.080 77.630 110.400 ;
        RECT 70.930 108.720 71.190 109.040 ;
        RECT 71.850 108.720 72.110 109.040 ;
        RECT 73.690 108.720 73.950 109.040 ;
        RECT 70.470 108.380 70.730 108.700 ;
        RECT 66.330 105.660 66.590 105.980 ;
        RECT 66.330 104.300 66.590 104.620 ;
        RECT 65.410 102.260 65.670 102.580 ;
        RECT 65.870 102.260 66.130 102.580 ;
        RECT 64.950 101.580 65.210 101.900 ;
        RECT 64.490 100.560 64.750 100.880 ;
        RECT 64.030 97.160 64.290 97.480 ;
        RECT 64.550 88.980 64.690 100.560 ;
        RECT 65.010 100.200 65.150 101.580 ;
        RECT 66.390 100.880 66.530 104.300 ;
        RECT 66.790 102.940 67.050 103.260 ;
        RECT 66.330 100.560 66.590 100.880 ;
        RECT 64.950 99.880 65.210 100.200 ;
        RECT 65.010 89.320 65.150 99.880 ;
        RECT 66.850 99.860 66.990 102.940 ;
        RECT 66.790 99.540 67.050 99.860 ;
        RECT 66.790 96.820 67.050 97.140 ;
        RECT 65.870 96.370 66.130 96.460 ;
        RECT 65.870 96.230 66.530 96.370 ;
        RECT 65.870 96.140 66.130 96.230 ;
        RECT 65.400 95.265 65.680 95.635 ;
        RECT 65.470 95.100 65.610 95.265 ;
        RECT 65.410 94.780 65.670 95.100 ;
        RECT 65.870 93.420 66.130 93.740 ;
        RECT 65.930 91.360 66.070 93.420 ;
        RECT 65.870 91.040 66.130 91.360 ;
        RECT 64.950 89.000 65.210 89.320 ;
        RECT 65.410 89.000 65.670 89.320 ;
        RECT 64.490 88.660 64.750 88.980 ;
        RECT 63.570 87.980 63.830 88.300 ;
        RECT 64.550 86.680 64.690 88.660 ;
        RECT 64.090 86.540 64.690 86.680 ;
        RECT 64.090 86.260 64.230 86.540 ;
        RECT 64.030 85.940 64.290 86.260 ;
        RECT 64.950 85.940 65.210 86.260 ;
        RECT 64.490 85.260 64.750 85.580 ;
        RECT 58.050 79.820 58.310 80.140 ;
        RECT 57.590 73.360 57.850 73.680 ;
        RECT 57.650 69.940 57.790 73.360 ;
        RECT 57.590 69.620 57.850 69.940 ;
        RECT 57.590 67.240 57.850 67.560 ;
        RECT 57.130 66.220 57.390 66.540 ;
        RECT 56.670 64.180 56.930 64.500 ;
        RECT 56.730 62.800 56.870 64.180 ;
        RECT 56.670 62.480 56.930 62.800 ;
        RECT 56.210 59.760 56.470 60.080 ;
        RECT 56.730 59.400 56.870 62.480 ;
        RECT 56.670 59.080 56.930 59.400 ;
        RECT 57.650 56.340 57.790 67.240 ;
        RECT 58.110 65.520 58.250 79.820 ;
        RECT 62.650 78.120 62.910 78.440 ;
        RECT 62.710 75.380 62.850 78.120 ;
        RECT 64.550 75.380 64.690 85.260 ;
        RECT 65.010 83.880 65.150 85.940 ;
        RECT 65.470 84.560 65.610 89.000 ;
        RECT 65.410 84.240 65.670 84.560 ;
        RECT 64.950 83.560 65.210 83.880 ;
        RECT 65.010 80.480 65.150 83.560 ;
        RECT 64.950 80.160 65.210 80.480 ;
        RECT 65.930 78.440 66.070 91.040 ;
        RECT 66.390 86.260 66.530 96.230 ;
        RECT 66.850 94.760 66.990 96.820 ;
        RECT 67.310 96.800 67.450 107.700 ;
        RECT 68.230 107.620 68.830 107.760 ;
        RECT 68.690 107.340 68.830 107.620 ;
        RECT 67.710 107.020 67.970 107.340 ;
        RECT 68.630 107.020 68.890 107.340 ;
        RECT 67.770 105.640 67.910 107.020 ;
        RECT 67.710 105.320 67.970 105.640 ;
        RECT 67.770 100.200 67.910 105.320 ;
        RECT 67.710 99.880 67.970 100.200 ;
        RECT 67.770 98.160 67.910 99.880 ;
        RECT 69.090 99.540 69.350 99.860 ;
        RECT 71.910 99.715 72.050 108.720 ;
        RECT 74.150 108.380 74.410 108.700 ;
        RECT 73.690 105.320 73.950 105.640 ;
        RECT 72.310 104.980 72.570 105.300 ;
        RECT 72.370 104.620 72.510 104.980 ;
        RECT 73.750 104.620 73.890 105.320 ;
        RECT 72.310 104.300 72.570 104.620 ;
        RECT 73.690 104.300 73.950 104.620 ;
        RECT 67.710 97.840 67.970 98.160 ;
        RECT 67.770 97.420 68.830 97.560 ;
        RECT 67.250 96.480 67.510 96.800 ;
        RECT 66.790 94.440 67.050 94.760 ;
        RECT 67.770 94.420 67.910 97.420 ;
        RECT 68.170 96.820 68.430 97.140 ;
        RECT 67.710 94.100 67.970 94.420 ;
        RECT 68.230 93.740 68.370 96.820 ;
        RECT 68.690 96.460 68.830 97.420 ;
        RECT 69.150 97.140 69.290 99.540 ;
        RECT 71.390 99.200 71.650 99.520 ;
        RECT 71.840 99.345 72.120 99.715 ;
        RECT 71.450 97.140 71.590 99.200 ;
        RECT 69.090 96.820 69.350 97.140 ;
        RECT 71.390 96.820 71.650 97.140 ;
        RECT 68.630 96.140 68.890 96.460 ;
        RECT 69.150 94.760 69.290 96.820 ;
        RECT 70.930 96.480 71.190 96.800 ;
        RECT 68.630 94.440 68.890 94.760 ;
        RECT 69.090 94.440 69.350 94.760 ;
        RECT 70.470 94.440 70.730 94.760 ;
        RECT 68.170 93.420 68.430 93.740 ;
        RECT 67.250 91.720 67.510 92.040 ;
        RECT 67.310 90.000 67.450 91.720 ;
        RECT 68.690 91.020 68.830 94.440 ;
        RECT 69.150 91.360 69.290 94.440 ;
        RECT 70.530 93.740 70.670 94.440 ;
        RECT 70.470 93.420 70.730 93.740 ;
        RECT 69.090 91.270 69.350 91.360 ;
        RECT 69.090 91.130 69.750 91.270 ;
        RECT 69.090 91.040 69.350 91.130 ;
        RECT 68.630 90.700 68.890 91.020 ;
        RECT 67.250 89.680 67.510 90.000 ;
        RECT 67.310 89.320 67.450 89.680 ;
        RECT 68.170 89.340 68.430 89.660 ;
        RECT 67.250 89.000 67.510 89.320 ;
        RECT 67.250 87.980 67.510 88.300 ;
        RECT 66.790 86.960 67.050 87.280 ;
        RECT 66.330 85.940 66.590 86.260 ;
        RECT 65.870 78.120 66.130 78.440 ;
        RECT 65.870 77.440 66.130 77.760 ;
        RECT 65.930 76.060 66.070 77.440 ;
        RECT 65.870 75.740 66.130 76.060 ;
        RECT 62.650 75.060 62.910 75.380 ;
        RECT 64.490 75.060 64.750 75.380 ;
        RECT 62.710 73.000 62.850 75.060 ;
        RECT 65.930 73.680 66.070 75.740 ;
        RECT 65.870 73.360 66.130 73.680 ;
        RECT 64.950 73.020 65.210 73.340 ;
        RECT 62.650 72.680 62.910 73.000 ;
        RECT 62.710 70.280 62.850 72.680 ;
        RECT 62.650 69.960 62.910 70.280 ;
        RECT 64.030 69.620 64.290 69.940 ;
        RECT 63.110 66.900 63.370 67.220 ;
        RECT 58.970 66.220 59.230 66.540 ;
        RECT 58.050 65.200 58.310 65.520 ;
        RECT 58.510 63.500 58.770 63.820 ;
        RECT 58.570 62.460 58.710 63.500 ;
        RECT 58.510 62.140 58.770 62.460 ;
        RECT 59.030 59.400 59.170 66.220 ;
        RECT 63.170 62.120 63.310 66.900 ;
        RECT 64.090 64.160 64.230 69.620 ;
        RECT 64.490 64.180 64.750 64.500 ;
        RECT 64.030 63.840 64.290 64.160 ;
        RECT 64.550 62.120 64.690 64.180 ;
        RECT 63.110 61.800 63.370 62.120 ;
        RECT 64.490 61.800 64.750 62.120 ;
        RECT 65.010 62.030 65.150 73.020 ;
        RECT 65.410 71.660 65.670 71.980 ;
        RECT 65.470 69.600 65.610 71.660 ;
        RECT 65.410 69.280 65.670 69.600 ;
        RECT 65.870 68.940 66.130 69.260 ;
        RECT 65.930 68.240 66.070 68.940 ;
        RECT 65.870 67.920 66.130 68.240 ;
        RECT 66.390 64.840 66.530 85.940 ;
        RECT 66.850 82.860 66.990 86.960 ;
        RECT 67.310 86.260 67.450 87.980 ;
        RECT 68.230 87.280 68.370 89.340 ;
        RECT 69.090 89.000 69.350 89.320 ;
        RECT 68.170 86.960 68.430 87.280 ;
        RECT 69.150 86.260 69.290 89.000 ;
        RECT 67.250 85.940 67.510 86.260 ;
        RECT 69.090 86.170 69.350 86.260 ;
        RECT 68.690 86.030 69.350 86.170 ;
        RECT 67.710 84.240 67.970 84.560 ;
        RECT 66.790 82.540 67.050 82.860 ;
        RECT 66.850 81.840 66.990 82.540 ;
        RECT 66.790 81.520 67.050 81.840 ;
        RECT 67.770 80.480 67.910 84.240 ;
        RECT 68.690 83.200 68.830 86.030 ;
        RECT 69.090 85.940 69.350 86.030 ;
        RECT 69.090 85.260 69.350 85.580 ;
        RECT 69.150 84.560 69.290 85.260 ;
        RECT 69.090 84.240 69.350 84.560 ;
        RECT 68.630 82.880 68.890 83.200 ;
        RECT 68.620 82.600 68.900 82.715 ;
        RECT 68.230 82.460 68.900 82.600 ;
        RECT 67.710 80.160 67.970 80.480 ;
        RECT 67.710 75.060 67.970 75.380 ;
        RECT 67.240 72.825 67.520 73.195 ;
        RECT 67.250 72.680 67.510 72.825 ;
        RECT 67.770 72.515 67.910 75.060 ;
        RECT 67.700 72.145 67.980 72.515 ;
        RECT 66.790 69.960 67.050 70.280 ;
        RECT 66.330 64.520 66.590 64.840 ;
        RECT 66.850 64.500 66.990 69.960 ;
        RECT 67.250 67.240 67.510 67.560 ;
        RECT 66.790 64.180 67.050 64.500 ;
        RECT 66.330 63.840 66.590 64.160 ;
        RECT 65.410 63.500 65.670 63.820 ;
        RECT 65.870 63.500 66.130 63.820 ;
        RECT 65.470 62.800 65.610 63.500 ;
        RECT 65.410 62.480 65.670 62.800 ;
        RECT 65.930 62.460 66.070 63.500 ;
        RECT 65.870 62.140 66.130 62.460 ;
        RECT 65.410 62.030 65.670 62.120 ;
        RECT 65.010 61.890 65.670 62.030 ;
        RECT 65.410 61.800 65.670 61.890 ;
        RECT 64.030 59.420 64.290 59.740 ;
        RECT 58.970 59.080 59.230 59.400 ;
        RECT 63.110 58.740 63.370 59.060 ;
        RECT 58.970 58.060 59.230 58.380 ;
        RECT 59.030 56.340 59.170 58.060 ;
        RECT 54.370 56.020 54.630 56.340 ;
        RECT 57.590 56.020 57.850 56.340 ;
        RECT 58.970 56.020 59.230 56.340 ;
        RECT 53.450 54.320 53.710 54.640 ;
        RECT 53.910 54.320 54.170 54.640 ;
        RECT 52.530 52.960 52.790 53.280 ;
        RECT 52.590 51.240 52.730 52.960 ;
        RECT 52.530 50.920 52.790 51.240 ;
        RECT 52.590 45.800 52.730 50.920 ;
        RECT 54.430 50.220 54.570 56.020 ;
        RECT 57.130 52.960 57.390 53.280 ;
        RECT 57.190 51.920 57.330 52.960 ;
        RECT 57.130 51.600 57.390 51.920 ;
        RECT 57.650 50.560 57.790 56.020 ;
        RECT 59.030 54.640 59.170 56.020 ;
        RECT 59.430 55.340 59.690 55.660 ;
        RECT 58.970 54.320 59.230 54.640 ;
        RECT 59.490 51.920 59.630 55.340 ;
        RECT 63.170 54.640 63.310 58.740 ;
        RECT 63.110 54.320 63.370 54.640 ;
        RECT 59.890 53.300 60.150 53.620 ;
        RECT 59.950 51.920 60.090 53.300 ;
        RECT 60.810 52.620 61.070 52.940 ;
        RECT 59.430 51.600 59.690 51.920 ;
        RECT 59.890 51.600 60.150 51.920 ;
        RECT 59.430 50.580 59.690 50.900 ;
        RECT 57.590 50.240 57.850 50.560 ;
        RECT 54.370 49.900 54.630 50.220 ;
        RECT 54.370 48.200 54.630 48.520 ;
        RECT 54.430 46.140 54.570 48.200 ;
        RECT 54.830 47.520 55.090 47.840 ;
        RECT 54.370 45.820 54.630 46.140 ;
        RECT 52.530 45.480 52.790 45.800 ;
        RECT 53.910 42.080 54.170 42.400 ;
        RECT 52.990 41.740 53.250 42.060 ;
        RECT 53.050 40.700 53.190 41.740 ;
        RECT 53.450 40.720 53.710 41.040 ;
        RECT 52.990 40.380 53.250 40.700 ;
        RECT 53.510 34.920 53.650 40.720 ;
        RECT 53.970 38.320 54.110 42.080 ;
        RECT 54.890 42.060 55.030 47.520 ;
        RECT 55.750 47.180 56.010 47.500 ;
        RECT 55.290 45.480 55.550 45.800 ;
        RECT 55.350 42.740 55.490 45.480 ;
        RECT 55.810 45.120 55.950 47.180 ;
        RECT 58.970 45.140 59.230 45.460 ;
        RECT 55.750 44.800 56.010 45.120 ;
        RECT 55.290 42.420 55.550 42.740 ;
        RECT 54.830 41.740 55.090 42.060 ;
        RECT 55.810 40.360 55.950 44.800 ;
        RECT 57.130 42.080 57.390 42.400 ;
        RECT 55.750 40.040 56.010 40.360 ;
        RECT 57.190 40.020 57.330 42.080 ;
        RECT 57.130 39.700 57.390 40.020 ;
        RECT 53.910 38.000 54.170 38.320 ;
        RECT 56.670 36.300 56.930 36.620 ;
        RECT 54.370 34.940 54.630 35.260 ;
        RECT 53.450 34.600 53.710 34.920 ;
        RECT 54.430 31.860 54.570 34.940 ;
        RECT 55.750 34.600 56.010 34.920 ;
        RECT 55.810 32.880 55.950 34.600 ;
        RECT 55.750 32.560 56.010 32.880 ;
        RECT 52.530 31.540 52.790 31.860 ;
        RECT 54.370 31.540 54.630 31.860 ;
        RECT 52.590 29.480 52.730 31.540 ;
        RECT 52.530 29.160 52.790 29.480 ;
        RECT 54.430 28.880 54.570 31.540 ;
        RECT 56.210 31.200 56.470 31.520 ;
        RECT 52.590 28.740 54.570 28.880 ;
        RECT 54.830 28.820 55.090 29.140 ;
        RECT 52.590 26.420 52.730 28.740 ;
        RECT 54.370 28.200 54.630 28.460 ;
        RECT 53.970 28.140 54.630 28.200 ;
        RECT 53.970 28.060 54.570 28.140 ;
        RECT 52.530 26.100 52.790 26.420 ;
        RECT 53.970 25.740 54.110 28.060 ;
        RECT 54.890 27.520 55.030 28.820 ;
        RECT 54.430 27.380 55.030 27.520 ;
        RECT 54.430 25.740 54.570 27.380 ;
        RECT 54.830 25.760 55.090 26.080 ;
        RECT 53.910 25.420 54.170 25.740 ;
        RECT 54.370 25.420 54.630 25.740 ;
        RECT 52.070 17.260 52.330 17.580 ;
        RECT 49.310 16.240 49.570 16.560 ;
        RECT 53.970 15.880 54.110 25.420 ;
        RECT 54.430 24.380 54.570 25.420 ;
        RECT 54.890 24.720 55.030 25.760 ;
        RECT 54.830 24.400 55.090 24.720 ;
        RECT 54.370 24.060 54.630 24.380 ;
        RECT 54.430 20.980 54.570 24.060 ;
        RECT 55.290 23.380 55.550 23.700 ;
        RECT 54.830 23.040 55.090 23.360 ;
        RECT 54.890 20.980 55.030 23.040 ;
        RECT 55.350 20.980 55.490 23.380 ;
        RECT 54.370 20.660 54.630 20.980 ;
        RECT 54.830 20.660 55.090 20.980 ;
        RECT 55.290 20.660 55.550 20.980 ;
        RECT 55.750 20.660 56.010 20.980 ;
        RECT 54.370 19.980 54.630 20.300 ;
        RECT 54.430 18.600 54.570 19.980 ;
        RECT 55.810 19.280 55.950 20.660 ;
        RECT 55.750 18.960 56.010 19.280 ;
        RECT 54.370 18.280 54.630 18.600 ;
        RECT 53.910 15.560 54.170 15.880 ;
        RECT 56.270 15.540 56.410 31.200 ;
        RECT 56.730 24.040 56.870 36.300 ;
        RECT 57.190 33.900 57.330 39.700 ;
        RECT 59.030 39.340 59.170 45.140 ;
        RECT 59.490 39.680 59.630 50.580 ;
        RECT 60.870 49.200 61.010 52.620 ;
        RECT 60.810 48.880 61.070 49.200 ;
        RECT 61.730 48.880 61.990 49.200 ;
        RECT 61.790 48.180 61.930 48.880 ;
        RECT 61.730 47.860 61.990 48.180 ;
        RECT 63.570 47.860 63.830 48.180 ;
        RECT 61.270 47.520 61.530 47.840 ;
        RECT 61.330 45.800 61.470 47.520 ;
        RECT 59.890 45.480 60.150 45.800 ;
        RECT 61.270 45.480 61.530 45.800 ;
        RECT 59.950 43.760 60.090 45.480 ;
        RECT 59.890 43.440 60.150 43.760 ;
        RECT 59.950 40.020 60.090 43.440 ;
        RECT 60.810 41.740 61.070 42.060 ;
        RECT 60.870 40.360 61.010 41.740 ;
        RECT 61.330 40.360 61.470 45.480 ;
        RECT 63.110 40.720 63.370 41.040 ;
        RECT 60.810 40.040 61.070 40.360 ;
        RECT 61.270 40.040 61.530 40.360 ;
        RECT 59.890 39.700 60.150 40.020 ;
        RECT 59.430 39.360 59.690 39.680 ;
        RECT 58.970 39.020 59.230 39.340 ;
        RECT 57.130 33.580 57.390 33.900 ;
        RECT 57.590 33.580 57.850 33.900 ;
        RECT 57.190 32.200 57.330 33.580 ;
        RECT 57.130 31.880 57.390 32.200 ;
        RECT 57.190 29.820 57.330 31.880 ;
        RECT 57.650 31.520 57.790 33.580 ;
        RECT 57.590 31.200 57.850 31.520 ;
        RECT 58.510 31.200 58.770 31.520 ;
        RECT 57.130 29.500 57.390 29.820 ;
        RECT 56.670 23.720 56.930 24.040 ;
        RECT 56.730 22.000 56.870 23.720 ;
        RECT 56.670 21.680 56.930 22.000 ;
        RECT 56.730 20.300 56.870 21.680 ;
        RECT 57.190 20.980 57.330 29.500 ;
        RECT 58.570 28.800 58.710 31.200 ;
        RECT 59.030 31.180 59.170 39.020 ;
        RECT 60.870 37.640 61.010 40.040 ;
        RECT 60.810 37.320 61.070 37.640 ;
        RECT 58.970 30.860 59.230 31.180 ;
        RECT 59.030 29.390 59.170 30.860 ;
        RECT 59.430 29.390 59.690 29.480 ;
        RECT 59.030 29.250 59.690 29.390 ;
        RECT 59.430 29.160 59.690 29.250 ;
        RECT 58.510 28.480 58.770 28.800 ;
        RECT 59.490 24.040 59.630 29.160 ;
        RECT 61.330 28.800 61.470 40.040 ;
        RECT 61.730 39.020 61.990 39.340 ;
        RECT 61.790 31.860 61.930 39.020 ;
        RECT 62.190 36.640 62.450 36.960 ;
        RECT 62.250 35.600 62.390 36.640 ;
        RECT 62.650 36.300 62.910 36.620 ;
        RECT 62.190 35.280 62.450 35.600 ;
        RECT 62.710 34.920 62.850 36.300 ;
        RECT 62.650 34.600 62.910 34.920 ;
        RECT 61.730 31.540 61.990 31.860 ;
        RECT 62.650 31.540 62.910 31.860 ;
        RECT 61.730 30.860 61.990 31.180 ;
        RECT 61.790 29.480 61.930 30.860 ;
        RECT 62.710 29.480 62.850 31.540 ;
        RECT 63.170 30.160 63.310 40.720 ;
        RECT 63.630 33.900 63.770 47.860 ;
        RECT 64.090 43.160 64.230 59.420 ;
        RECT 64.550 56.340 64.690 61.800 ;
        RECT 65.470 60.080 65.610 61.800 ;
        RECT 66.390 61.520 66.530 63.840 ;
        RECT 67.310 62.120 67.450 67.240 ;
        RECT 68.230 67.220 68.370 82.460 ;
        RECT 68.620 82.345 68.900 82.460 ;
        RECT 69.610 81.240 69.750 91.130 ;
        RECT 70.990 90.000 71.130 96.480 ;
        RECT 71.450 94.760 71.590 96.820 ;
        RECT 71.390 94.440 71.650 94.760 ;
        RECT 71.450 92.720 71.590 94.440 ;
        RECT 71.910 94.420 72.050 99.345 ;
        RECT 71.850 94.100 72.110 94.420 ;
        RECT 71.390 92.400 71.650 92.720 ;
        RECT 71.390 91.380 71.650 91.700 ;
        RECT 70.930 89.910 71.190 90.000 ;
        RECT 70.530 89.770 71.190 89.910 ;
        RECT 70.010 84.240 70.270 84.560 ;
        RECT 69.150 81.100 69.750 81.240 ;
        RECT 68.630 79.820 68.890 80.140 ;
        RECT 68.690 78.780 68.830 79.820 ;
        RECT 69.150 79.120 69.290 81.100 ;
        RECT 69.550 80.500 69.810 80.820 ;
        RECT 69.090 78.800 69.350 79.120 ;
        RECT 68.630 78.460 68.890 78.780 ;
        RECT 69.610 78.440 69.750 80.500 ;
        RECT 69.550 78.120 69.810 78.440 ;
        RECT 70.070 78.100 70.210 84.240 ;
        RECT 70.530 78.440 70.670 89.770 ;
        RECT 70.930 89.680 71.190 89.770 ;
        RECT 71.450 89.320 71.590 91.380 ;
        RECT 71.390 89.000 71.650 89.320 ;
        RECT 71.450 86.260 71.590 89.000 ;
        RECT 71.910 86.600 72.050 94.100 ;
        RECT 71.850 86.280 72.110 86.600 ;
        RECT 71.390 85.940 71.650 86.260 ;
        RECT 71.450 84.220 71.590 85.940 ;
        RECT 71.390 83.900 71.650 84.220 ;
        RECT 70.930 83.220 71.190 83.540 ;
        RECT 70.470 78.120 70.730 78.440 ;
        RECT 69.090 78.010 69.350 78.100 ;
        RECT 68.690 77.870 69.350 78.010 ;
        RECT 68.690 73.680 68.830 77.870 ;
        RECT 69.090 77.780 69.350 77.870 ;
        RECT 70.010 77.780 70.270 78.100 ;
        RECT 70.530 77.330 70.670 78.120 ;
        RECT 69.610 77.190 70.670 77.330 ;
        RECT 69.090 75.400 69.350 75.720 ;
        RECT 69.150 75.040 69.290 75.400 ;
        RECT 69.090 74.720 69.350 75.040 ;
        RECT 69.150 73.680 69.290 74.720 ;
        RECT 69.610 73.680 69.750 77.190 ;
        RECT 70.010 75.400 70.270 75.720 ;
        RECT 68.630 73.360 68.890 73.680 ;
        RECT 69.090 73.360 69.350 73.680 ;
        RECT 69.550 73.360 69.810 73.680 ;
        RECT 68.630 72.910 68.890 73.000 ;
        RECT 68.630 72.770 69.750 72.910 ;
        RECT 68.630 72.680 68.890 72.770 ;
        RECT 69.090 72.000 69.350 72.320 ;
        RECT 69.150 69.940 69.290 72.000 ;
        RECT 69.610 69.940 69.750 72.770 ;
        RECT 69.090 69.620 69.350 69.940 ;
        RECT 69.550 69.620 69.810 69.940 ;
        RECT 69.610 67.560 69.750 69.620 ;
        RECT 70.070 69.600 70.210 75.400 ;
        RECT 70.990 75.380 71.130 83.220 ;
        RECT 71.390 82.715 71.650 82.860 ;
        RECT 71.380 82.345 71.660 82.715 ;
        RECT 72.370 81.500 72.510 104.300 ;
        RECT 73.690 102.600 73.950 102.920 ;
        RECT 73.230 101.920 73.490 102.240 ;
        RECT 73.290 100.880 73.430 101.920 ;
        RECT 73.750 101.900 73.890 102.600 ;
        RECT 73.690 101.580 73.950 101.900 ;
        RECT 73.230 100.560 73.490 100.880 ;
        RECT 72.770 99.880 73.030 100.200 ;
        RECT 72.830 97.820 72.970 99.880 ;
        RECT 73.230 99.540 73.490 99.860 ;
        RECT 73.290 98.160 73.430 99.540 ;
        RECT 73.750 98.160 73.890 101.580 ;
        RECT 74.210 100.200 74.350 108.380 ;
        RECT 77.430 108.020 77.570 110.080 ;
        RECT 77.370 107.700 77.630 108.020 ;
        RECT 75.530 107.020 75.790 107.340 ;
        RECT 74.610 106.000 74.870 106.320 ;
        RECT 74.670 100.200 74.810 106.000 ;
        RECT 75.590 105.640 75.730 107.020 ;
        RECT 75.070 105.320 75.330 105.640 ;
        RECT 75.530 105.320 75.790 105.640 ;
        RECT 75.130 100.880 75.270 105.320 ;
        RECT 75.530 104.300 75.790 104.620 ;
        RECT 75.590 102.920 75.730 104.300 ;
        RECT 75.990 102.940 76.250 103.260 ;
        RECT 75.530 102.600 75.790 102.920 ;
        RECT 75.070 100.560 75.330 100.880 ;
        RECT 74.150 99.880 74.410 100.200 ;
        RECT 74.610 99.880 74.870 100.200 ;
        RECT 74.150 99.200 74.410 99.520 ;
        RECT 75.070 99.200 75.330 99.520 ;
        RECT 73.230 97.840 73.490 98.160 ;
        RECT 73.690 97.840 73.950 98.160 ;
        RECT 72.770 97.500 73.030 97.820 ;
        RECT 72.830 88.980 72.970 97.500 ;
        RECT 73.230 96.820 73.490 97.140 ;
        RECT 73.290 90.000 73.430 96.820 ;
        RECT 74.210 95.635 74.350 99.200 ;
        RECT 75.130 96.460 75.270 99.200 ;
        RECT 75.070 96.140 75.330 96.460 ;
        RECT 74.140 95.265 74.420 95.635 ;
        RECT 73.230 89.680 73.490 90.000 ;
        RECT 72.770 88.660 73.030 88.980 ;
        RECT 72.770 87.980 73.030 88.300 ;
        RECT 72.830 84.560 72.970 87.980 ;
        RECT 73.290 86.260 73.430 89.680 ;
        RECT 73.690 88.660 73.950 88.980 ;
        RECT 73.230 85.940 73.490 86.260 ;
        RECT 72.770 84.240 73.030 84.560 ;
        RECT 73.230 82.880 73.490 83.200 ;
        RECT 72.310 81.180 72.570 81.500 ;
        RECT 72.370 80.820 72.510 81.180 ;
        RECT 72.310 80.500 72.570 80.820 ;
        RECT 71.850 78.800 72.110 79.120 ;
        RECT 72.300 78.945 72.580 79.315 ;
        RECT 71.390 76.080 71.650 76.400 ;
        RECT 70.930 75.290 71.190 75.380 ;
        RECT 70.530 75.150 71.190 75.290 ;
        RECT 70.010 69.280 70.270 69.600 ;
        RECT 69.550 67.240 69.810 67.560 ;
        RECT 68.170 66.900 68.430 67.220 ;
        RECT 70.530 66.880 70.670 75.150 ;
        RECT 70.930 75.060 71.190 75.150 ;
        RECT 70.920 72.145 71.200 72.515 ;
        RECT 70.990 71.980 71.130 72.145 ;
        RECT 70.930 71.660 71.190 71.980 ;
        RECT 70.930 70.300 71.190 70.620 ;
        RECT 70.990 67.560 71.130 70.300 ;
        RECT 70.930 67.240 71.190 67.560 ;
        RECT 70.470 66.560 70.730 66.880 ;
        RECT 69.090 64.520 69.350 64.840 ;
        RECT 67.250 61.800 67.510 62.120 ;
        RECT 65.930 61.380 66.530 61.520 ;
        RECT 65.410 59.760 65.670 60.080 ;
        RECT 65.470 59.060 65.610 59.760 ;
        RECT 65.410 58.740 65.670 59.060 ;
        RECT 64.950 58.060 65.210 58.380 ;
        RECT 64.490 56.020 64.750 56.340 ;
        RECT 65.010 53.620 65.150 58.060 ;
        RECT 64.950 53.300 65.210 53.620 ;
        RECT 64.950 47.520 65.210 47.840 ;
        RECT 65.010 45.800 65.150 47.520 ;
        RECT 65.930 46.140 66.070 61.380 ;
        RECT 66.320 60.585 66.600 60.955 ;
        RECT 68.630 60.780 68.890 61.100 ;
        RECT 66.390 59.400 66.530 60.585 ;
        RECT 66.330 59.080 66.590 59.400 ;
        RECT 67.250 58.740 67.510 59.060 ;
        RECT 67.710 58.800 67.970 59.060 ;
        RECT 68.690 58.800 68.830 60.780 ;
        RECT 69.150 59.060 69.290 64.520 ;
        RECT 69.550 62.480 69.810 62.800 ;
        RECT 69.610 59.060 69.750 62.480 ;
        RECT 67.710 58.740 68.830 58.800 ;
        RECT 69.090 58.740 69.350 59.060 ;
        RECT 69.550 58.740 69.810 59.060 ;
        RECT 70.010 58.740 70.270 59.060 ;
        RECT 66.330 58.400 66.590 58.720 ;
        RECT 66.390 56.000 66.530 58.400 ;
        RECT 67.310 57.360 67.450 58.740 ;
        RECT 67.770 58.660 68.830 58.740 ;
        RECT 67.710 58.060 67.970 58.380 ;
        RECT 67.250 57.040 67.510 57.360 ;
        RECT 67.770 56.680 67.910 58.060 ;
        RECT 67.710 56.360 67.970 56.680 ;
        RECT 66.330 55.680 66.590 56.000 ;
        RECT 68.690 55.660 68.830 58.660 ;
        RECT 70.070 58.380 70.210 58.740 ;
        RECT 69.550 58.060 69.810 58.380 ;
        RECT 70.010 58.060 70.270 58.380 ;
        RECT 69.610 56.340 69.750 58.060 ;
        RECT 70.010 56.700 70.270 57.020 ;
        RECT 69.550 56.020 69.810 56.340 ;
        RECT 68.630 55.340 68.890 55.660 ;
        RECT 70.070 53.280 70.210 56.700 ;
        RECT 70.530 56.680 70.670 66.560 ;
        RECT 71.450 66.540 71.590 76.080 ;
        RECT 71.910 75.720 72.050 78.800 ;
        RECT 72.370 78.780 72.510 78.945 ;
        RECT 72.310 78.460 72.570 78.780 ;
        RECT 72.770 78.120 73.030 78.440 ;
        RECT 72.830 77.760 72.970 78.120 ;
        RECT 72.770 77.440 73.030 77.760 ;
        RECT 71.850 75.400 72.110 75.720 ;
        RECT 73.290 75.380 73.430 82.880 ;
        RECT 73.750 75.380 73.890 88.660 ;
        RECT 74.210 88.300 74.350 95.265 ;
        RECT 75.130 94.760 75.270 96.140 ;
        RECT 75.070 94.440 75.330 94.760 ;
        RECT 75.590 94.420 75.730 102.600 ;
        RECT 76.050 99.520 76.190 102.940 ;
        RECT 77.890 100.110 78.030 115.180 ;
        RECT 87.090 114.480 87.230 116.200 ;
        RECT 88.400 115.665 88.680 116.035 ;
        RECT 88.410 115.520 88.670 115.665 ;
        RECT 87.030 114.160 87.290 114.480 ;
        RECT 78.290 113.140 78.550 113.460 ;
        RECT 86.110 113.140 86.370 113.460 ;
        RECT 87.030 113.140 87.290 113.460 ;
        RECT 78.350 111.080 78.490 113.140 ;
        RECT 78.290 110.760 78.550 111.080 ;
        RECT 79.670 110.760 79.930 111.080 ;
        RECT 79.730 109.040 79.870 110.760 ;
        RECT 86.170 110.740 86.310 113.140 ;
        RECT 86.110 110.420 86.370 110.740 ;
        RECT 85.650 109.740 85.910 110.060 ;
        RECT 79.670 108.720 79.930 109.040 ;
        RECT 83.350 108.040 83.610 108.360 ;
        RECT 81.510 107.020 81.770 107.340 ;
        RECT 78.750 104.640 79.010 104.960 ;
        RECT 78.290 100.110 78.550 100.200 ;
        RECT 77.430 99.970 78.550 100.110 ;
        RECT 76.910 99.540 77.170 99.860 ;
        RECT 75.990 99.200 76.250 99.520 ;
        RECT 76.450 98.860 76.710 99.180 ;
        RECT 76.510 97.820 76.650 98.860 ;
        RECT 76.970 98.160 77.110 99.540 ;
        RECT 76.910 97.840 77.170 98.160 ;
        RECT 76.450 97.500 76.710 97.820 ;
        RECT 76.450 94.440 76.710 94.760 ;
        RECT 75.530 94.100 75.790 94.420 ;
        RECT 76.510 94.080 76.650 94.440 ;
        RECT 76.450 93.760 76.710 94.080 ;
        RECT 76.510 91.020 76.650 93.760 ;
        RECT 77.430 93.740 77.570 99.970 ;
        RECT 78.290 99.880 78.550 99.970 ;
        RECT 77.820 99.345 78.100 99.715 ;
        RECT 77.890 99.180 78.030 99.345 ;
        RECT 77.830 98.860 78.090 99.180 ;
        RECT 78.810 97.480 78.950 104.640 ;
        RECT 79.210 102.260 79.470 102.580 ;
        RECT 78.750 97.160 79.010 97.480 ;
        RECT 78.750 94.440 79.010 94.760 ;
        RECT 77.830 94.100 78.090 94.420 ;
        RECT 77.370 93.420 77.630 93.740 ;
        RECT 77.430 91.700 77.570 93.420 ;
        RECT 77.890 91.700 78.030 94.100 ;
        RECT 78.810 92.040 78.950 94.440 ;
        RECT 78.750 91.720 79.010 92.040 ;
        RECT 77.370 91.380 77.630 91.700 ;
        RECT 77.830 91.380 78.090 91.700 ;
        RECT 76.450 90.700 76.710 91.020 ;
        RECT 74.150 87.980 74.410 88.300 ;
        RECT 74.150 86.960 74.410 87.280 ;
        RECT 74.210 81.240 74.350 86.960 ;
        RECT 76.510 86.940 76.650 90.700 ;
        RECT 77.890 89.910 78.030 91.380 ;
        RECT 77.890 89.770 78.490 89.910 ;
        RECT 77.370 89.340 77.630 89.660 ;
        RECT 76.450 86.620 76.710 86.940 ;
        RECT 75.530 86.280 75.790 86.600 ;
        RECT 75.070 85.600 75.330 85.920 ;
        RECT 74.610 85.260 74.870 85.580 ;
        RECT 74.670 82.860 74.810 85.260 ;
        RECT 74.610 82.540 74.870 82.860 ;
        RECT 74.210 81.100 74.810 81.240 ;
        RECT 74.670 80.820 74.810 81.100 ;
        RECT 74.150 80.500 74.410 80.820 ;
        RECT 74.610 80.500 74.870 80.820 ;
        RECT 74.210 79.315 74.350 80.500 ;
        RECT 74.140 78.945 74.420 79.315 ;
        RECT 74.150 77.440 74.410 77.760 ;
        RECT 73.230 75.060 73.490 75.380 ;
        RECT 73.690 75.060 73.950 75.380 ;
        RECT 71.850 74.720 72.110 75.040 ;
        RECT 71.910 69.940 72.050 74.720 ;
        RECT 72.310 74.380 72.570 74.700 ;
        RECT 72.770 74.380 73.030 74.700 ;
        RECT 72.370 73.680 72.510 74.380 ;
        RECT 72.310 73.360 72.570 73.680 ;
        RECT 72.310 72.680 72.570 73.000 ;
        RECT 72.370 70.960 72.510 72.680 ;
        RECT 72.830 72.660 72.970 74.380 ;
        RECT 72.770 72.340 73.030 72.660 ;
        RECT 72.310 70.640 72.570 70.960 ;
        RECT 72.770 70.300 73.030 70.620 ;
        RECT 71.850 69.620 72.110 69.940 ;
        RECT 72.310 69.280 72.570 69.600 ;
        RECT 72.370 67.560 72.510 69.280 ;
        RECT 72.310 67.240 72.570 67.560 ;
        RECT 71.390 66.220 71.650 66.540 ;
        RECT 71.450 64.500 71.590 66.220 ;
        RECT 72.370 64.840 72.510 67.240 ;
        RECT 72.310 64.520 72.570 64.840 ;
        RECT 71.390 64.180 71.650 64.500 ;
        RECT 71.450 60.955 71.590 64.180 ;
        RECT 72.370 61.780 72.510 64.520 ;
        RECT 72.310 61.460 72.570 61.780 ;
        RECT 71.380 60.585 71.660 60.955 ;
        RECT 72.310 60.780 72.570 61.100 ;
        RECT 70.930 59.760 71.190 60.080 ;
        RECT 71.390 59.760 71.650 60.080 ;
        RECT 70.990 59.060 71.130 59.760 ;
        RECT 71.450 59.060 71.590 59.760 ;
        RECT 71.850 59.420 72.110 59.740 ;
        RECT 70.930 58.740 71.190 59.060 ;
        RECT 71.390 58.740 71.650 59.060 ;
        RECT 70.990 57.360 71.130 58.740 ;
        RECT 71.910 58.720 72.050 59.420 ;
        RECT 72.370 59.060 72.510 60.780 ;
        RECT 72.830 59.400 72.970 70.300 ;
        RECT 73.290 62.460 73.430 75.060 ;
        RECT 74.210 74.700 74.350 77.440 ;
        RECT 74.150 74.610 74.410 74.700 ;
        RECT 73.750 74.470 74.410 74.610 ;
        RECT 73.750 73.195 73.890 74.470 ;
        RECT 74.150 74.380 74.410 74.470 ;
        RECT 74.670 73.760 74.810 80.500 ;
        RECT 75.130 76.400 75.270 85.600 ;
        RECT 75.590 84.220 75.730 86.280 ;
        RECT 75.990 85.600 76.250 85.920 ;
        RECT 75.530 83.900 75.790 84.220 ;
        RECT 75.530 81.240 75.790 81.500 ;
        RECT 76.050 81.240 76.190 85.600 ;
        RECT 75.530 81.180 76.190 81.240 ;
        RECT 75.590 81.100 76.190 81.180 ;
        RECT 75.070 76.080 75.330 76.400 ;
        RECT 75.530 75.400 75.790 75.720 ;
        RECT 75.590 74.440 75.730 75.400 ;
        RECT 74.210 73.620 74.810 73.760 ;
        RECT 75.130 74.300 75.730 74.440 ;
        RECT 73.680 72.825 73.960 73.195 ;
        RECT 73.750 70.280 73.890 72.825 ;
        RECT 74.210 71.980 74.350 73.620 ;
        RECT 74.610 73.080 74.870 73.340 ;
        RECT 75.130 73.080 75.270 74.300 ;
        RECT 75.530 73.360 75.790 73.680 ;
        RECT 74.610 73.020 75.270 73.080 ;
        RECT 74.670 72.940 75.270 73.020 ;
        RECT 74.610 72.570 74.870 72.660 ;
        RECT 75.590 72.570 75.730 73.360 ;
        RECT 76.050 73.000 76.190 81.100 ;
        RECT 76.510 78.520 76.650 86.620 ;
        RECT 77.430 80.820 77.570 89.340 ;
        RECT 78.350 89.320 78.490 89.770 ;
        RECT 78.810 89.660 78.950 91.720 ;
        RECT 78.750 89.340 79.010 89.660 ;
        RECT 79.270 89.320 79.410 102.260 ;
        RECT 81.050 101.920 81.310 102.240 ;
        RECT 81.110 100.880 81.250 101.920 ;
        RECT 81.050 100.560 81.310 100.880 ;
        RECT 80.130 99.200 80.390 99.520 ;
        RECT 79.670 96.140 79.930 96.460 ;
        RECT 79.730 95.440 79.870 96.140 ;
        RECT 79.670 95.120 79.930 95.440 ;
        RECT 77.830 89.000 78.090 89.320 ;
        RECT 78.290 89.000 78.550 89.320 ;
        RECT 79.210 89.000 79.470 89.320 ;
        RECT 77.890 83.880 78.030 89.000 ;
        RECT 78.350 85.830 78.490 89.000 ;
        RECT 78.350 85.690 78.950 85.830 ;
        RECT 77.830 83.560 78.090 83.880 ;
        RECT 78.810 80.820 78.950 85.690 ;
        RECT 79.270 81.160 79.410 89.000 ;
        RECT 80.190 86.260 80.330 99.200 ;
        RECT 81.570 95.440 81.710 107.020 ;
        RECT 83.410 106.320 83.550 108.040 ;
        RECT 85.710 108.020 85.850 109.740 ;
        RECT 87.090 109.040 87.230 113.140 ;
        RECT 88.410 112.635 88.670 112.780 ;
        RECT 88.400 112.265 88.680 112.635 ;
        RECT 87.030 108.720 87.290 109.040 ;
        RECT 85.650 107.700 85.910 108.020 ;
        RECT 86.110 107.700 86.370 108.020 ;
        RECT 83.350 106.000 83.610 106.320 ;
        RECT 86.170 105.300 86.310 107.700 ;
        RECT 100.360 105.820 100.660 180.090 ;
        RECT 100.860 179.630 118.970 179.640 ;
        RECT 100.860 179.350 119.005 179.630 ;
        RECT 100.860 179.340 118.970 179.350 ;
        RECT 100.860 120.760 101.160 179.340 ;
        RECT 101.580 178.940 122.370 178.950 ;
        RECT 101.580 178.660 122.405 178.940 ;
        RECT 101.580 178.650 122.370 178.660 ;
        RECT 101.580 135.760 101.880 178.650 ;
        RECT 102.210 178.350 115.570 178.360 ;
        RECT 102.210 178.070 115.605 178.350 ;
        RECT 102.210 178.060 115.570 178.070 ;
        RECT 102.210 150.840 102.510 178.060 ;
        RECT 102.770 177.660 112.170 177.670 ;
        RECT 102.770 177.380 112.205 177.660 ;
        RECT 102.770 177.370 112.170 177.380 ;
        RECT 102.790 165.570 103.090 177.370 ;
        RECT 106.840 176.770 107.540 176.780 ;
        RECT 106.500 176.030 107.850 176.770 ;
        RECT 106.840 166.600 107.540 176.030 ;
        RECT 117.980 174.620 118.880 176.640 ;
        RECT 116.255 172.705 116.575 172.760 ;
        RECT 116.255 172.550 118.860 172.705 ;
        RECT 116.255 172.500 116.575 172.550 ;
        RECT 108.890 171.080 116.880 171.470 ;
        RECT 108.820 168.770 109.400 169.400 ;
        RECT 111.430 168.020 114.090 171.080 ;
        RECT 108.930 167.570 116.870 168.020 ;
        RECT 106.750 165.810 107.610 166.600 ;
        RECT 106.840 161.770 107.540 161.780 ;
        RECT 106.500 161.030 107.850 161.770 ;
        RECT 106.840 151.600 107.540 161.030 ;
        RECT 116.160 157.690 116.480 157.750 ;
        RECT 116.160 157.550 118.510 157.690 ;
        RECT 116.160 157.490 116.480 157.550 ;
        RECT 108.890 156.080 116.880 156.470 ;
        RECT 108.790 153.690 109.370 154.320 ;
        RECT 111.430 153.020 114.090 156.080 ;
        RECT 108.930 152.570 116.870 153.020 ;
        RECT 102.210 150.540 103.050 150.840 ;
        RECT 106.750 150.810 107.610 151.600 ;
        RECT 106.840 146.720 107.540 146.730 ;
        RECT 106.500 145.980 107.850 146.720 ;
        RECT 106.840 136.550 107.540 145.980 ;
        RECT 116.400 142.635 116.720 142.690 ;
        RECT 116.400 142.485 118.115 142.635 ;
        RECT 116.400 142.430 116.720 142.485 ;
        RECT 108.890 141.030 116.880 141.420 ;
        RECT 108.790 138.740 109.370 139.370 ;
        RECT 111.430 137.970 114.090 141.030 ;
        RECT 108.930 137.520 116.870 137.970 ;
        RECT 106.750 135.760 107.610 136.550 ;
        RECT 101.580 135.460 103.130 135.760 ;
        RECT 106.840 131.720 107.540 131.730 ;
        RECT 106.500 130.980 107.850 131.720 ;
        RECT 106.840 121.550 107.540 130.980 ;
        RECT 116.290 127.640 116.610 127.680 ;
        RECT 116.290 127.460 117.690 127.640 ;
        RECT 116.290 127.420 116.610 127.460 ;
        RECT 108.890 126.030 116.880 126.420 ;
        RECT 108.790 123.740 109.370 124.370 ;
        RECT 111.430 122.970 114.090 126.030 ;
        RECT 108.930 122.520 116.870 122.970 ;
        RECT 106.750 120.760 107.610 121.550 ;
        RECT 100.860 120.460 103.170 120.760 ;
        RECT 106.790 116.780 107.490 116.790 ;
        RECT 106.450 116.040 107.800 116.780 ;
        RECT 106.790 106.610 107.490 116.040 ;
        RECT 116.510 112.675 116.830 112.720 ;
        RECT 116.510 112.505 117.195 112.675 ;
        RECT 116.510 112.460 116.830 112.505 ;
        RECT 108.840 111.090 116.830 111.480 ;
        RECT 108.750 108.700 109.330 109.330 ;
        RECT 111.380 108.030 114.040 111.090 ;
        RECT 108.880 107.580 116.820 108.030 ;
        RECT 106.700 105.820 107.560 106.610 ;
        RECT 100.360 105.520 103.080 105.820 ;
        RECT 86.110 104.980 86.370 105.300 ;
        RECT 82.890 104.300 83.150 104.620 ;
        RECT 82.950 100.880 83.090 104.300 ;
        RECT 86.170 103.600 86.310 104.980 ;
        RECT 100.180 103.665 112.290 103.900 ;
        RECT 86.110 103.280 86.370 103.600 ;
        RECT 100.180 103.175 110.620 103.390 ;
        RECT 100.180 102.760 109.045 102.970 ;
        RECT 100.180 102.210 107.455 102.480 ;
        RECT 83.810 101.580 84.070 101.900 ;
        RECT 100.180 101.665 105.905 101.930 ;
        RECT 82.890 100.560 83.150 100.880 ;
        RECT 83.870 99.860 84.010 101.580 ;
        RECT 100.180 101.075 104.305 101.360 ;
        RECT 100.180 100.400 102.800 100.700 ;
        RECT 83.350 99.540 83.610 99.860 ;
        RECT 83.810 99.540 84.070 99.860 ;
        RECT 100.180 99.790 101.275 100.035 ;
        RECT 83.410 98.160 83.550 99.540 ;
        RECT 83.350 97.840 83.610 98.160 ;
        RECT 81.510 95.120 81.770 95.440 ;
        RECT 101.030 92.875 101.275 99.790 ;
        RECT 102.500 92.925 102.800 100.400 ;
        RECT 104.020 92.925 104.305 101.075 ;
        RECT 105.640 92.955 105.905 101.665 ;
        RECT 100.620 92.615 101.680 92.875 ;
        RECT 102.120 92.625 103.180 92.925 ;
        RECT 103.630 92.640 104.690 92.925 ;
        RECT 105.240 92.690 106.300 92.955 ;
        RECT 107.185 92.925 107.455 102.210 ;
        RECT 108.835 92.955 109.045 102.760 ;
        RECT 106.790 92.655 107.850 92.925 ;
        RECT 108.410 92.695 109.470 92.955 ;
        RECT 110.405 92.925 110.620 103.175 ;
        RECT 112.055 92.945 112.290 103.665 ;
        RECT 117.025 101.605 117.195 112.505 ;
        RECT 117.510 102.010 117.690 127.460 ;
        RECT 117.965 102.335 118.115 142.485 ;
        RECT 118.370 102.640 118.510 157.550 ;
        RECT 118.705 102.965 118.860 172.550 ;
        RECT 123.240 169.890 123.540 180.190 ;
        RECT 120.480 169.590 123.540 169.890 ;
        RECT 123.830 179.710 129.170 179.720 ;
        RECT 123.830 179.430 129.205 179.710 ;
        RECT 152.680 179.480 152.960 179.515 ;
        RECT 123.830 179.420 129.170 179.430 ;
        RECT 120.480 105.740 120.780 169.590 ;
        RECT 123.830 168.770 124.130 179.420 ;
        RECT 143.320 179.180 152.970 179.480 ;
        RECT 121.150 168.470 124.130 168.770 ;
        RECT 124.430 179.000 132.570 179.010 ;
        RECT 124.430 178.720 132.605 179.000 ;
        RECT 124.430 178.710 132.570 178.720 ;
        RECT 121.150 120.900 121.450 168.470 ;
        RECT 124.430 167.820 124.730 178.710 ;
        RECT 121.750 167.520 124.730 167.820 ;
        RECT 124.920 178.280 135.970 178.290 ;
        RECT 124.920 178.000 136.005 178.280 ;
        RECT 124.920 177.990 135.970 178.000 ;
        RECT 121.750 135.710 122.050 167.520 ;
        RECT 124.920 166.810 125.220 177.990 ;
        RECT 122.310 166.510 125.220 166.810 ;
        RECT 125.540 177.560 142.770 177.570 ;
        RECT 125.540 177.280 142.805 177.560 ;
        RECT 125.540 177.270 142.770 177.280 ;
        RECT 122.310 150.820 122.610 166.510 ;
        RECT 125.540 166.000 125.840 177.270 ;
        RECT 126.720 176.720 127.420 176.730 ;
        RECT 126.380 175.980 127.730 176.720 ;
        RECT 126.720 166.550 127.420 175.980 ;
        RECT 137.800 174.600 138.700 176.620 ;
        RECT 136.460 172.635 136.780 172.690 ;
        RECT 136.460 172.485 138.465 172.635 ;
        RECT 136.460 172.430 136.780 172.485 ;
        RECT 128.770 171.030 136.760 171.420 ;
        RECT 128.680 168.760 129.260 169.390 ;
        RECT 131.310 167.970 133.970 171.030 ;
        RECT 128.810 167.520 136.750 167.970 ;
        RECT 122.900 165.700 125.840 166.000 ;
        RECT 126.630 165.760 127.490 166.550 ;
        RECT 126.720 161.770 127.420 161.780 ;
        RECT 126.380 161.030 127.730 161.770 ;
        RECT 126.720 151.600 127.420 161.030 ;
        RECT 136.270 157.695 136.590 157.720 ;
        RECT 136.270 157.485 138.095 157.695 ;
        RECT 136.270 157.460 136.590 157.485 ;
        RECT 128.770 156.080 136.760 156.470 ;
        RECT 128.680 153.800 129.260 154.430 ;
        RECT 131.310 153.020 133.970 156.080 ;
        RECT 128.810 152.570 136.750 153.020 ;
        RECT 122.310 150.520 122.980 150.820 ;
        RECT 126.630 150.810 127.490 151.600 ;
        RECT 126.720 146.720 127.420 146.730 ;
        RECT 126.380 145.980 127.730 146.720 ;
        RECT 126.720 136.550 127.420 145.980 ;
        RECT 136.150 142.705 136.470 142.750 ;
        RECT 136.150 142.535 137.715 142.705 ;
        RECT 136.150 142.490 136.470 142.535 ;
        RECT 128.770 141.030 136.760 141.420 ;
        RECT 128.680 138.730 129.260 139.360 ;
        RECT 131.310 137.970 133.970 141.030 ;
        RECT 128.810 137.520 136.750 137.970 ;
        RECT 126.630 135.760 127.490 136.550 ;
        RECT 121.750 135.410 122.980 135.710 ;
        RECT 126.720 131.780 127.420 131.790 ;
        RECT 126.380 131.040 127.730 131.780 ;
        RECT 126.720 121.610 127.420 131.040 ;
        RECT 136.335 127.700 136.655 127.760 ;
        RECT 136.335 127.555 137.375 127.700 ;
        RECT 136.335 127.500 136.655 127.555 ;
        RECT 128.770 126.090 136.760 126.480 ;
        RECT 128.610 123.790 129.190 124.420 ;
        RECT 131.310 123.030 133.970 126.090 ;
        RECT 128.810 122.580 136.750 123.030 ;
        RECT 121.150 120.600 123.010 120.900 ;
        RECT 126.630 120.820 127.490 121.610 ;
        RECT 126.720 116.780 127.420 116.790 ;
        RECT 126.380 116.040 127.730 116.780 ;
        RECT 126.720 106.610 127.420 116.040 ;
        RECT 136.160 112.690 136.480 112.750 ;
        RECT 136.160 112.550 137.090 112.690 ;
        RECT 136.160 112.490 136.480 112.550 ;
        RECT 128.770 111.090 136.760 111.480 ;
        RECT 128.730 108.760 129.310 109.390 ;
        RECT 131.310 108.030 133.970 111.090 ;
        RECT 128.810 107.580 136.750 108.030 ;
        RECT 126.630 105.820 127.490 106.610 ;
        RECT 120.480 105.440 123.040 105.740 ;
        RECT 136.950 103.450 137.090 112.550 ;
        RECT 137.230 103.740 137.375 127.555 ;
        RECT 137.545 104.065 137.715 142.535 ;
        RECT 137.885 104.455 138.095 157.485 ;
        RECT 138.315 104.825 138.465 172.485 ;
        RECT 143.320 169.390 143.620 179.180 ;
        RECT 152.680 179.145 152.960 179.180 ;
        RECT 140.280 169.090 143.620 169.390 ;
        RECT 144.050 178.740 146.170 178.750 ;
        RECT 144.050 178.460 146.205 178.740 ;
        RECT 144.050 178.450 146.170 178.460 ;
        RECT 140.280 105.820 140.580 169.090 ;
        RECT 144.050 168.490 144.350 178.450 ;
        RECT 145.290 178.030 149.570 178.040 ;
        RECT 145.290 177.750 149.605 178.030 ;
        RECT 145.290 177.740 149.570 177.750 ;
        RECT 144.680 176.850 144.960 176.885 ;
        RECT 140.940 168.190 144.350 168.490 ;
        RECT 140.940 120.830 141.240 168.190 ;
        RECT 144.670 167.700 144.970 176.850 ;
        RECT 141.710 167.400 144.970 167.700 ;
        RECT 141.710 135.850 142.010 167.400 ;
        RECT 145.290 166.930 145.590 177.740 ;
        RECT 142.350 166.630 145.590 166.930 ;
        RECT 145.960 177.370 148.420 177.380 ;
        RECT 145.960 177.090 148.455 177.370 ;
        RECT 145.960 177.080 148.420 177.090 ;
        RECT 142.350 150.730 142.650 166.630 ;
        RECT 145.960 166.020 146.260 177.080 ;
        RECT 146.750 176.770 147.450 176.780 ;
        RECT 146.410 176.030 147.760 176.770 ;
        RECT 146.750 166.600 147.450 176.030 ;
        RECT 157.570 174.580 158.470 176.600 ;
        RECT 156.415 172.650 156.735 172.710 ;
        RECT 156.415 172.505 158.350 172.650 ;
        RECT 156.415 172.450 156.735 172.505 ;
        RECT 148.800 171.080 156.790 171.470 ;
        RECT 148.880 168.740 149.460 169.370 ;
        RECT 151.340 168.020 154.000 171.080 ;
        RECT 148.840 167.570 156.780 168.020 ;
        RECT 142.960 165.720 146.260 166.020 ;
        RECT 146.660 165.810 147.520 166.600 ;
        RECT 146.800 161.720 147.500 161.730 ;
        RECT 146.460 160.980 147.810 161.720 ;
        RECT 146.800 151.550 147.500 160.980 ;
        RECT 156.500 157.640 156.820 157.700 ;
        RECT 156.500 157.500 158.030 157.640 ;
        RECT 156.500 157.440 156.820 157.500 ;
        RECT 148.850 156.030 156.840 156.420 ;
        RECT 148.920 153.710 149.500 154.340 ;
        RECT 151.390 152.970 154.050 156.030 ;
        RECT 148.890 152.520 156.830 152.970 ;
        RECT 146.710 150.760 147.570 151.550 ;
        RECT 142.350 150.430 142.970 150.730 ;
        RECT 146.750 146.720 147.450 146.730 ;
        RECT 146.410 145.980 147.760 146.720 ;
        RECT 146.750 136.550 147.450 145.980 ;
        RECT 156.330 142.625 156.590 142.710 ;
        RECT 156.330 142.475 157.705 142.625 ;
        RECT 156.330 142.390 156.590 142.475 ;
        RECT 148.800 141.030 156.790 141.420 ;
        RECT 148.830 138.670 149.410 139.300 ;
        RECT 151.340 137.970 154.000 141.030 ;
        RECT 148.840 137.520 156.780 137.970 ;
        RECT 141.710 135.550 143.010 135.850 ;
        RECT 146.660 135.760 147.520 136.550 ;
        RECT 146.750 131.780 147.450 131.790 ;
        RECT 146.410 131.040 147.760 131.780 ;
        RECT 146.750 121.610 147.450 131.040 ;
        RECT 156.410 127.660 156.730 127.720 ;
        RECT 156.410 127.520 157.410 127.660 ;
        RECT 156.410 127.460 156.730 127.520 ;
        RECT 148.800 126.090 156.790 126.480 ;
        RECT 148.950 123.750 149.530 124.380 ;
        RECT 151.340 123.030 154.000 126.090 ;
        RECT 148.840 122.580 156.780 123.030 ;
        RECT 140.940 120.530 142.990 120.830 ;
        RECT 146.660 120.820 147.520 121.610 ;
        RECT 146.750 116.780 147.450 116.790 ;
        RECT 146.410 116.040 147.760 116.780 ;
        RECT 146.750 106.610 147.450 116.040 ;
        RECT 156.000 112.715 156.320 112.770 ;
        RECT 156.000 112.565 157.115 112.715 ;
        RECT 156.000 112.510 156.320 112.565 ;
        RECT 148.800 111.090 156.790 111.480 ;
        RECT 148.910 108.790 149.490 109.420 ;
        RECT 151.340 108.030 154.000 111.090 ;
        RECT 148.840 107.580 156.780 108.030 ;
        RECT 146.660 105.820 147.520 106.610 ;
        RECT 140.280 105.520 143.020 105.820 ;
        RECT 138.315 104.675 149.650 104.825 ;
        RECT 137.885 104.245 147.750 104.455 ;
        RECT 137.545 103.895 146.220 104.065 ;
        RECT 137.230 103.595 144.785 103.740 ;
        RECT 136.950 103.310 143.320 103.450 ;
        RECT 118.705 102.810 141.785 102.965 ;
        RECT 118.370 102.500 140.290 102.640 ;
        RECT 117.965 102.185 138.860 102.335 ;
        RECT 117.510 101.970 137.340 102.010 ;
        RECT 117.510 101.830 137.730 101.970 ;
        RECT 137.160 101.620 137.730 101.830 ;
        RECT 117.025 101.435 135.840 101.605 ;
        RECT 137.210 101.500 137.730 101.620 ;
        RECT 135.670 99.200 135.840 101.435 ;
        RECT 138.710 99.390 138.860 102.185 ;
        RECT 140.150 101.990 140.290 102.500 ;
        RECT 140.150 101.620 140.700 101.990 ;
        RECT 140.180 101.520 140.700 101.620 ;
        RECT 135.670 98.995 136.300 99.200 ;
        RECT 138.710 99.015 139.270 99.390 ;
        RECT 135.690 98.720 136.300 98.995 ;
        RECT 138.750 98.920 139.270 99.015 ;
        RECT 141.630 99.310 141.785 102.810 ;
        RECT 143.180 102.050 143.320 103.310 ;
        RECT 143.180 101.580 143.700 102.050 ;
        RECT 144.640 99.340 144.785 103.595 ;
        RECT 146.050 102.080 146.220 103.895 ;
        RECT 146.050 101.950 146.610 102.080 ;
        RECT 146.090 101.610 146.610 101.950 ;
        RECT 147.540 99.390 147.750 104.245 ;
        RECT 149.500 101.940 149.650 104.675 ;
        RECT 156.965 103.015 157.115 112.565 ;
        RECT 149.120 101.705 149.650 101.940 ;
        RECT 150.960 102.865 157.115 103.015 ;
        RECT 149.120 101.470 149.640 101.705 ;
        RECT 141.630 98.955 142.180 99.310 ;
        RECT 141.660 98.840 142.180 98.955 ;
        RECT 144.640 98.870 145.160 99.340 ;
        RECT 147.540 99.075 148.230 99.390 ;
        RECT 150.960 99.310 151.110 102.865 ;
        RECT 157.270 102.720 157.410 127.520 ;
        RECT 152.470 102.580 157.410 102.720 ;
        RECT 152.470 102.060 152.610 102.580 ;
        RECT 157.555 102.375 157.705 142.475 ;
        RECT 152.090 101.590 152.610 102.060 ;
        RECT 153.960 102.225 157.705 102.375 ;
        RECT 147.560 98.860 148.230 99.075 ;
        RECT 150.570 99.055 151.110 99.310 ;
        RECT 153.960 99.280 154.110 102.225 ;
        RECT 155.040 101.990 155.560 102.050 ;
        RECT 157.890 101.990 158.030 157.500 ;
        RECT 155.040 101.850 158.030 101.990 ;
        RECT 155.040 101.580 155.560 101.850 ;
        RECT 158.205 99.285 158.350 172.505 ;
        RECT 153.580 99.115 154.110 99.280 ;
        RECT 156.480 99.140 158.350 99.285 ;
        RECT 150.570 98.840 151.090 99.055 ;
        RECT 153.580 98.810 154.100 99.115 ;
        RECT 156.510 98.780 157.030 99.140 ;
        RECT 109.980 92.665 111.040 92.925 ;
        RECT 111.640 92.685 112.700 92.945 ;
        RECT 80.590 91.380 80.850 91.700 ;
        RECT 88.410 91.380 88.670 91.700 ;
        RECT 80.130 85.940 80.390 86.260 ;
        RECT 79.210 80.840 79.470 81.160 ;
        RECT 76.910 80.500 77.170 80.820 ;
        RECT 77.370 80.500 77.630 80.820 ;
        RECT 78.750 80.500 79.010 80.820 ;
        RECT 76.970 79.120 77.110 80.500 ;
        RECT 76.910 78.800 77.170 79.120 ;
        RECT 76.510 78.440 77.110 78.520 ;
        RECT 76.510 78.380 77.170 78.440 ;
        RECT 76.910 78.120 77.170 78.380 ;
        RECT 75.990 72.680 76.250 73.000 ;
        RECT 76.450 72.680 76.710 73.000 ;
        RECT 74.610 72.430 75.730 72.570 ;
        RECT 74.610 72.340 74.870 72.430 ;
        RECT 74.150 71.660 74.410 71.980 ;
        RECT 74.210 70.960 74.350 71.660 ;
        RECT 74.150 70.640 74.410 70.960 ;
        RECT 75.530 70.300 75.790 70.620 ;
        RECT 73.690 69.960 73.950 70.280 ;
        RECT 75.590 67.560 75.730 70.300 ;
        RECT 76.050 67.900 76.190 72.680 ;
        RECT 76.510 70.960 76.650 72.680 ;
        RECT 76.450 70.640 76.710 70.960 ;
        RECT 76.970 70.360 77.110 78.120 ;
        RECT 77.430 75.720 77.570 80.500 ;
        RECT 77.830 79.820 78.090 80.140 ;
        RECT 77.370 75.400 77.630 75.720 ;
        RECT 76.510 70.220 77.110 70.360 ;
        RECT 75.990 67.580 76.250 67.900 ;
        RECT 75.070 67.240 75.330 67.560 ;
        RECT 75.530 67.240 75.790 67.560 ;
        RECT 75.130 66.880 75.270 67.240 ;
        RECT 75.070 66.560 75.330 66.880 ;
        RECT 75.590 65.480 75.730 67.240 ;
        RECT 76.050 66.880 76.190 67.580 ;
        RECT 75.990 66.560 76.250 66.880 ;
        RECT 75.130 65.340 75.730 65.480 ;
        RECT 73.230 62.140 73.490 62.460 ;
        RECT 72.770 59.080 73.030 59.400 ;
        RECT 73.290 59.310 73.430 62.140 ;
        RECT 74.150 59.310 74.410 59.400 ;
        RECT 73.290 59.170 74.410 59.310 ;
        RECT 74.150 59.080 74.410 59.170 ;
        RECT 72.310 58.740 72.570 59.060 ;
        RECT 71.850 58.400 72.110 58.720 ;
        RECT 70.930 57.040 71.190 57.360 ;
        RECT 70.470 56.360 70.730 56.680 ;
        RECT 70.990 56.590 71.130 57.040 ;
        RECT 72.830 57.020 72.970 59.080 ;
        RECT 75.130 59.060 75.270 65.340 ;
        RECT 75.530 64.520 75.790 64.840 ;
        RECT 75.590 62.120 75.730 64.520 ;
        RECT 76.510 64.500 76.650 70.220 ;
        RECT 77.430 69.600 77.570 75.400 ;
        RECT 77.890 73.000 78.030 79.820 ;
        RECT 78.290 77.780 78.550 78.100 ;
        RECT 77.830 72.680 78.090 73.000 ;
        RECT 77.890 70.620 78.030 72.680 ;
        RECT 78.350 72.660 78.490 77.780 ;
        RECT 78.810 73.680 78.950 80.500 ;
        RECT 79.270 75.720 79.410 80.840 ;
        RECT 80.190 80.480 80.330 85.940 ;
        RECT 80.130 80.160 80.390 80.480 ;
        RECT 79.210 75.400 79.470 75.720 ;
        RECT 80.130 75.400 80.390 75.720 ;
        RECT 79.670 74.720 79.930 75.040 ;
        RECT 78.750 73.360 79.010 73.680 ;
        RECT 78.290 72.340 78.550 72.660 ;
        RECT 77.830 70.300 78.090 70.620 ;
        RECT 78.810 70.280 78.950 73.360 ;
        RECT 78.750 69.960 79.010 70.280 ;
        RECT 77.830 69.620 78.090 69.940 ;
        RECT 77.370 69.280 77.630 69.600 ;
        RECT 77.430 69.000 77.570 69.280 ;
        RECT 76.970 68.860 77.570 69.000 ;
        RECT 76.450 64.180 76.710 64.500 ;
        RECT 75.530 61.800 75.790 62.120 ;
        RECT 76.450 61.800 76.710 62.120 ;
        RECT 75.990 61.120 76.250 61.440 ;
        RECT 76.050 60.080 76.190 61.120 ;
        RECT 75.530 59.760 75.790 60.080 ;
        RECT 75.990 59.760 76.250 60.080 ;
        RECT 74.610 58.740 74.870 59.060 ;
        RECT 75.070 58.740 75.330 59.060 ;
        RECT 74.670 58.380 74.810 58.740 ;
        RECT 74.610 58.060 74.870 58.380 ;
        RECT 72.770 56.700 73.030 57.020 ;
        RECT 71.390 56.590 71.650 56.680 ;
        RECT 70.990 56.450 71.650 56.590 ;
        RECT 71.390 56.360 71.650 56.450 ;
        RECT 74.150 55.340 74.410 55.660 ;
        RECT 74.210 53.620 74.350 55.340 ;
        RECT 74.670 54.300 74.810 58.060 ;
        RECT 75.130 56.680 75.270 58.740 ;
        RECT 75.590 57.440 75.730 59.760 ;
        RECT 75.590 57.300 76.190 57.440 ;
        RECT 76.510 57.360 76.650 61.800 ;
        RECT 76.970 58.970 77.110 68.860 ;
        RECT 77.370 67.240 77.630 67.560 ;
        RECT 77.430 65.520 77.570 67.240 ;
        RECT 77.370 65.200 77.630 65.520 ;
        RECT 77.890 62.800 78.030 69.620 ;
        RECT 78.290 69.280 78.550 69.600 ;
        RECT 78.350 67.900 78.490 69.280 ;
        RECT 78.290 67.580 78.550 67.900 ;
        RECT 78.810 67.470 78.950 69.960 ;
        RECT 79.210 67.470 79.470 67.560 ;
        RECT 78.810 67.330 79.470 67.470 ;
        RECT 78.290 64.180 78.550 64.500 ;
        RECT 77.830 62.480 78.090 62.800 ;
        RECT 77.370 58.970 77.630 59.060 ;
        RECT 76.970 58.830 77.630 58.970 ;
        RECT 77.370 58.740 77.630 58.830 ;
        RECT 75.530 56.700 75.790 57.020 ;
        RECT 75.070 56.360 75.330 56.680 ;
        RECT 74.610 53.980 74.870 54.300 ;
        RECT 75.590 53.620 75.730 56.700 ;
        RECT 74.150 53.300 74.410 53.620 ;
        RECT 75.530 53.300 75.790 53.620 ;
        RECT 70.010 52.960 70.270 53.280 ;
        RECT 76.050 51.580 76.190 57.300 ;
        RECT 76.450 57.040 76.710 57.360 ;
        RECT 78.350 57.020 78.490 64.180 ;
        RECT 78.810 59.060 78.950 67.330 ;
        RECT 79.210 67.240 79.470 67.330 ;
        RECT 79.210 66.560 79.470 66.880 ;
        RECT 79.270 61.100 79.410 66.560 ;
        RECT 79.730 62.120 79.870 74.720 ;
        RECT 80.190 67.560 80.330 75.400 ;
        RECT 80.650 74.700 80.790 91.380 ;
        RECT 85.650 90.700 85.910 91.020 ;
        RECT 81.510 89.000 81.770 89.320 ;
        RECT 81.570 87.280 81.710 89.000 ;
        RECT 83.350 87.980 83.610 88.300 ;
        RECT 81.510 86.960 81.770 87.280 ;
        RECT 83.410 85.920 83.550 87.980 ;
        RECT 85.710 86.260 85.850 90.700 ;
        RECT 88.470 90.000 88.610 91.380 ;
        RECT 100.150 90.045 100.470 90.915 ;
        RECT 86.110 89.680 86.370 90.000 ;
        RECT 88.410 89.680 88.670 90.000 ;
        RECT 86.170 86.260 86.310 89.680 ;
        RECT 87.490 89.000 87.750 89.320 ;
        RECT 100.140 89.015 100.470 90.045 ;
        RECT 101.820 90.025 102.140 90.905 ;
        RECT 87.550 87.280 87.690 89.000 ;
        RECT 88.400 88.465 88.680 88.835 ;
        RECT 88.410 88.320 88.670 88.465 ;
        RECT 87.490 86.960 87.750 87.280 ;
        RECT 100.140 87.255 100.450 89.015 ;
        RECT 101.800 89.005 102.140 90.025 ;
        RECT 103.380 89.005 103.700 90.905 ;
        RECT 104.920 90.015 105.240 90.915 ;
        RECT 104.900 89.015 105.240 90.015 ;
        RECT 106.510 89.825 106.830 90.935 ;
        RECT 101.800 87.365 102.110 89.005 ;
        RECT 100.140 87.095 100.360 87.255 ;
        RECT 100.610 87.095 101.150 87.235 ;
        RECT 85.650 85.940 85.910 86.260 ;
        RECT 86.110 85.940 86.370 86.260 ;
        RECT 83.350 85.600 83.610 85.920 ;
        RECT 100.140 85.005 101.150 87.095 ;
        RECT 100.180 84.985 101.150 85.005 ;
        RECT 101.800 87.045 102.610 87.365 ;
        RECT 103.380 87.235 103.690 89.005 ;
        RECT 101.800 84.985 102.530 87.045 ;
        RECT 100.540 84.895 101.150 84.985 ;
        RECT 102.080 84.955 102.530 84.985 ;
        RECT 102.110 84.925 102.480 84.955 ;
        RECT 103.380 84.945 104.050 87.235 ;
        RECT 104.900 87.215 105.210 89.015 ;
        RECT 106.470 87.245 106.840 89.825 ;
        RECT 108.070 89.815 108.390 90.905 ;
        RECT 109.660 89.855 109.980 90.925 ;
        RECT 111.260 90.165 111.540 90.915 ;
        RECT 108.050 87.275 108.420 89.815 ;
        RECT 104.900 84.975 105.560 87.215 ;
        RECT 103.500 84.885 104.050 84.945 ;
        RECT 105.010 84.865 105.560 84.975 ;
        RECT 106.470 84.895 107.020 87.245 ;
        RECT 107.950 84.925 108.500 87.275 ;
        RECT 109.660 87.265 110.010 89.855 ;
        RECT 111.240 87.275 111.540 90.165 ;
        RECT 109.400 85.015 110.010 87.265 ;
        RECT 109.400 84.915 109.950 85.015 ;
        RECT 110.900 84.985 111.540 87.275 ;
        RECT 122.930 88.730 123.320 91.520 ;
        RECT 126.380 88.730 126.830 91.510 ;
        RECT 122.930 86.070 126.830 88.730 ;
        RECT 110.900 84.925 111.450 84.985 ;
        RECT 87.030 83.560 87.290 83.880 ;
        RECT 85.190 82.540 85.450 82.860 ;
        RECT 85.650 82.540 85.910 82.860 ;
        RECT 84.730 81.520 84.990 81.840 ;
        RECT 81.970 80.160 82.230 80.480 ;
        RECT 82.030 79.120 82.170 80.160 ;
        RECT 84.270 79.820 84.530 80.140 ;
        RECT 81.970 78.800 82.230 79.120 ;
        RECT 84.330 78.780 84.470 79.820 ;
        RECT 84.270 78.460 84.530 78.780 ;
        RECT 84.790 78.100 84.930 81.520 ;
        RECT 85.250 80.820 85.390 82.540 ;
        RECT 85.190 80.500 85.450 80.820 ;
        RECT 85.710 79.120 85.850 82.540 ;
        RECT 87.090 81.840 87.230 83.560 ;
        RECT 122.930 83.530 123.320 86.070 ;
        RECT 126.380 83.570 126.830 86.070 ;
        RECT 135.870 84.040 138.500 84.390 ;
        RECT 135.870 83.840 136.140 84.040 ;
        RECT 117.630 82.180 118.370 82.490 ;
        RECT 127.800 82.180 128.590 82.250 ;
        RECT 87.030 81.520 87.290 81.840 ;
        RECT 88.400 81.665 88.680 82.035 ;
        RECT 88.410 81.520 88.670 81.665 ;
        RECT 117.620 81.480 128.590 82.180 ;
        RECT 117.630 81.140 118.370 81.480 ;
        RECT 127.800 81.390 128.590 81.480 ;
        RECT 135.460 79.960 136.140 83.840 ;
        RECT 135.850 79.740 136.130 79.960 ;
        RECT 135.850 79.420 138.990 79.740 ;
        RECT 136.730 79.410 137.060 79.420 ;
        RECT 137.690 79.410 138.020 79.420 ;
        RECT 138.650 79.410 138.980 79.420 ;
        RECT 85.650 78.800 85.910 79.120 ;
        RECT 87.030 78.120 87.290 78.440 ;
        RECT 134.410 78.430 135.590 79.090 ;
        RECT 84.730 77.780 84.990 78.100 ;
        RECT 87.090 76.400 87.230 78.120 ;
        RECT 134.410 78.090 136.250 78.430 ;
        RECT 134.410 78.080 135.590 78.090 ;
        RECT 135.980 77.880 136.210 78.090 ;
        RECT 135.980 77.560 138.490 77.880 ;
        RECT 87.490 77.100 87.750 77.420 ;
        RECT 87.030 76.080 87.290 76.400 ;
        RECT 86.570 75.060 86.830 75.380 ;
        RECT 81.510 74.720 81.770 75.040 ;
        RECT 80.590 74.380 80.850 74.700 ;
        RECT 81.570 73.680 81.710 74.720 ;
        RECT 81.510 73.360 81.770 73.680 ;
        RECT 86.110 69.620 86.370 69.940 ;
        RECT 81.510 69.280 81.770 69.600 ;
        RECT 80.130 67.240 80.390 67.560 ;
        RECT 81.050 67.240 81.310 67.560 ;
        RECT 80.190 64.840 80.330 67.240 ;
        RECT 80.130 64.520 80.390 64.840 ;
        RECT 79.670 61.800 79.930 62.120 ;
        RECT 79.210 60.780 79.470 61.100 ;
        RECT 78.750 58.740 79.010 59.060 ;
        RECT 78.290 56.700 78.550 57.020 ;
        RECT 78.750 56.250 79.010 56.340 ;
        RECT 79.270 56.250 79.410 60.780 ;
        RECT 80.190 59.400 80.330 64.520 ;
        RECT 80.130 59.310 80.390 59.400 ;
        RECT 79.730 59.170 80.390 59.310 ;
        RECT 79.730 56.680 79.870 59.170 ;
        RECT 80.130 59.080 80.390 59.170 ;
        RECT 79.670 56.360 79.930 56.680 ;
        RECT 80.590 56.360 80.850 56.680 ;
        RECT 78.750 56.110 79.410 56.250 ;
        RECT 78.750 56.020 79.010 56.110 ;
        RECT 79.730 54.300 79.870 56.360 ;
        RECT 80.650 54.640 80.790 56.360 ;
        RECT 80.590 54.320 80.850 54.640 ;
        RECT 79.670 53.980 79.930 54.300 ;
        RECT 76.910 52.620 77.170 52.940 ;
        RECT 76.450 51.600 76.710 51.920 ;
        RECT 75.990 51.260 76.250 51.580 ;
        RECT 70.470 48.880 70.730 49.200 ;
        RECT 70.530 48.180 70.670 48.880 ;
        RECT 72.770 48.200 73.030 48.520 ;
        RECT 67.250 47.860 67.510 48.180 ;
        RECT 69.090 48.090 69.350 48.180 ;
        RECT 70.470 48.090 70.730 48.180 ;
        RECT 69.090 47.950 69.750 48.090 ;
        RECT 69.090 47.860 69.350 47.950 ;
        RECT 67.310 47.500 67.450 47.860 ;
        RECT 67.250 47.180 67.510 47.500 ;
        RECT 65.870 45.820 66.130 46.140 ;
        RECT 64.950 45.480 65.210 45.800 ;
        RECT 65.870 45.140 66.130 45.460 ;
        RECT 64.090 43.020 64.690 43.160 ;
        RECT 64.030 42.080 64.290 42.400 ;
        RECT 64.090 41.040 64.230 42.080 ;
        RECT 64.030 40.720 64.290 41.040 ;
        RECT 63.570 33.580 63.830 33.900 ;
        RECT 63.110 29.840 63.370 30.160 ;
        RECT 61.730 29.160 61.990 29.480 ;
        RECT 62.650 29.160 62.910 29.480 ;
        RECT 61.270 28.480 61.530 28.800 ;
        RECT 59.430 23.720 59.690 24.040 ;
        RECT 57.590 22.700 57.850 23.020 ;
        RECT 57.650 20.980 57.790 22.700 ;
        RECT 57.130 20.660 57.390 20.980 ;
        RECT 57.590 20.660 57.850 20.980 ;
        RECT 56.670 19.980 56.930 20.300 ;
        RECT 57.190 18.940 57.330 20.660 ;
        RECT 61.270 19.980 61.530 20.300 ;
        RECT 57.130 18.620 57.390 18.940 ;
        RECT 61.330 17.920 61.470 19.980 ;
        RECT 61.270 17.600 61.530 17.920 ;
        RECT 56.210 15.220 56.470 15.540 ;
        RECT 61.790 15.200 61.930 29.160 ;
        RECT 62.710 24.040 62.850 29.160 ;
        RECT 64.550 24.720 64.690 43.020 ;
        RECT 65.930 42.740 66.070 45.140 ;
        RECT 67.310 42.740 67.450 47.180 ;
        RECT 67.710 45.480 67.970 45.800 ;
        RECT 65.870 42.420 66.130 42.740 ;
        RECT 67.250 42.420 67.510 42.740 ;
        RECT 67.310 40.360 67.450 42.420 ;
        RECT 67.770 40.700 67.910 45.480 ;
        RECT 68.630 42.080 68.890 42.400 ;
        RECT 67.710 40.380 67.970 40.700 ;
        RECT 65.410 40.040 65.670 40.360 ;
        RECT 67.250 40.040 67.510 40.360 ;
        RECT 68.170 40.040 68.430 40.360 ;
        RECT 65.470 39.340 65.610 40.040 ;
        RECT 65.410 39.020 65.670 39.340 ;
        RECT 65.470 37.300 65.610 39.020 ;
        RECT 65.410 36.980 65.670 37.300 ;
        RECT 65.870 35.280 66.130 35.600 ;
        RECT 65.930 29.480 66.070 35.280 ;
        RECT 66.330 31.540 66.590 31.860 ;
        RECT 66.390 29.820 66.530 31.540 ;
        RECT 66.330 29.500 66.590 29.820 ;
        RECT 65.870 29.390 66.130 29.480 ;
        RECT 65.010 29.250 66.130 29.390 ;
        RECT 64.490 24.400 64.750 24.720 ;
        RECT 62.650 23.720 62.910 24.040 ;
        RECT 62.710 18.940 62.850 23.720 ;
        RECT 64.550 23.700 64.690 24.400 ;
        RECT 65.010 24.040 65.150 29.250 ;
        RECT 65.870 29.160 66.130 29.250 ;
        RECT 66.790 29.160 67.050 29.480 ;
        RECT 66.850 28.880 66.990 29.160 ;
        RECT 65.930 28.800 66.990 28.880 ;
        RECT 65.870 28.740 66.990 28.800 ;
        RECT 65.870 28.480 66.130 28.740 ;
        RECT 65.930 24.040 66.070 28.480 ;
        RECT 67.310 26.420 67.450 40.040 ;
        RECT 68.230 39.680 68.370 40.040 ;
        RECT 68.170 39.360 68.430 39.680 ;
        RECT 68.170 34.940 68.430 35.260 ;
        RECT 68.230 32.960 68.370 34.940 ;
        RECT 68.690 32.960 68.830 42.080 ;
        RECT 69.610 42.060 69.750 47.950 ;
        RECT 70.070 47.950 70.730 48.090 ;
        RECT 69.550 41.740 69.810 42.060 ;
        RECT 69.610 40.360 69.750 41.740 ;
        RECT 70.070 40.700 70.210 47.950 ;
        RECT 70.470 47.860 70.730 47.950 ;
        RECT 72.830 47.840 72.970 48.200 ;
        RECT 70.930 47.520 71.190 47.840 ;
        RECT 72.770 47.520 73.030 47.840 ;
        RECT 73.690 47.520 73.950 47.840 ;
        RECT 70.990 44.520 71.130 47.520 ;
        RECT 71.850 47.180 72.110 47.500 ;
        RECT 70.990 44.380 71.590 44.520 ;
        RECT 70.930 43.440 71.190 43.760 ;
        RECT 70.470 42.420 70.730 42.740 ;
        RECT 70.530 42.060 70.670 42.420 ;
        RECT 70.470 41.740 70.730 42.060 ;
        RECT 70.010 40.380 70.270 40.700 ;
        RECT 70.990 40.360 71.130 43.440 ;
        RECT 71.450 42.740 71.590 44.380 ;
        RECT 71.910 43.080 72.050 47.180 ;
        RECT 72.830 46.480 72.970 47.520 ;
        RECT 72.770 46.160 73.030 46.480 ;
        RECT 72.310 45.480 72.570 45.800 ;
        RECT 72.370 43.760 72.510 45.480 ;
        RECT 72.310 43.440 72.570 43.760 ;
        RECT 71.850 42.760 72.110 43.080 ;
        RECT 71.390 42.420 71.650 42.740 ;
        RECT 71.850 41.740 72.110 42.060 ;
        RECT 73.230 41.970 73.490 42.060 ;
        RECT 73.750 41.970 73.890 47.520 ;
        RECT 73.230 41.830 73.890 41.970 ;
        RECT 73.230 41.740 73.490 41.830 ;
        RECT 69.550 40.040 69.810 40.360 ;
        RECT 70.930 40.270 71.190 40.360 ;
        RECT 70.530 40.130 71.190 40.270 ;
        RECT 68.230 32.820 68.830 32.960 ;
        RECT 68.630 30.860 68.890 31.180 ;
        RECT 68.170 29.840 68.430 30.160 ;
        RECT 68.230 28.800 68.370 29.840 ;
        RECT 68.690 29.480 68.830 30.860 ;
        RECT 68.630 29.160 68.890 29.480 ;
        RECT 68.170 28.480 68.430 28.800 ;
        RECT 67.250 26.100 67.510 26.420 ;
        RECT 64.950 23.720 65.210 24.040 ;
        RECT 65.870 23.950 66.130 24.040 ;
        RECT 65.470 23.810 66.130 23.950 ;
        RECT 64.020 23.185 64.300 23.555 ;
        RECT 64.490 23.380 64.750 23.700 ;
        RECT 64.030 23.040 64.290 23.185 ;
        RECT 62.650 18.620 62.910 18.940 ;
        RECT 65.010 18.600 65.150 23.720 ;
        RECT 65.470 18.850 65.610 23.810 ;
        RECT 65.870 23.720 66.130 23.810 ;
        RECT 66.330 23.720 66.590 24.040 ;
        RECT 65.870 22.700 66.130 23.020 ;
        RECT 65.930 20.640 66.070 22.700 ;
        RECT 65.870 20.320 66.130 20.640 ;
        RECT 66.390 20.300 66.530 23.720 ;
        RECT 67.710 23.380 67.970 23.700 ;
        RECT 66.330 19.980 66.590 20.300 ;
        RECT 65.870 18.850 66.130 18.940 ;
        RECT 65.470 18.710 66.130 18.850 ;
        RECT 65.870 18.620 66.130 18.710 ;
        RECT 64.950 18.280 65.210 18.600 ;
        RECT 63.570 17.940 63.830 18.260 ;
        RECT 63.630 15.540 63.770 17.940 ;
        RECT 66.390 15.540 66.530 19.980 ;
        RECT 67.770 15.880 67.910 23.380 ;
        RECT 69.090 23.270 69.350 23.360 ;
        RECT 68.230 23.130 69.350 23.270 ;
        RECT 68.230 22.000 68.370 23.130 ;
        RECT 69.090 23.040 69.350 23.130 ;
        RECT 68.170 21.680 68.430 22.000 ;
        RECT 68.630 20.660 68.890 20.980 ;
        RECT 68.690 18.260 68.830 20.660 ;
        RECT 68.630 17.940 68.890 18.260 ;
        RECT 67.710 15.560 67.970 15.880 ;
        RECT 69.610 15.540 69.750 40.040 ;
        RECT 70.530 34.580 70.670 40.130 ;
        RECT 70.930 40.040 71.190 40.130 ;
        RECT 71.910 40.020 72.050 41.740 ;
        RECT 71.850 39.700 72.110 40.020 ;
        RECT 70.930 39.250 71.190 39.340 ;
        RECT 71.910 39.250 72.050 39.700 ;
        RECT 73.750 39.340 73.890 41.830 ;
        RECT 74.150 40.040 74.410 40.360 ;
        RECT 70.930 39.110 72.050 39.250 ;
        RECT 70.930 39.020 71.190 39.110 ;
        RECT 73.690 39.020 73.950 39.340 ;
        RECT 70.470 34.260 70.730 34.580 ;
        RECT 70.470 29.730 70.730 29.820 ;
        RECT 70.990 29.730 71.130 39.020 ;
        RECT 73.230 37.660 73.490 37.980 ;
        RECT 72.770 36.300 73.030 36.620 ;
        RECT 72.830 34.580 72.970 36.300 ;
        RECT 72.770 34.260 73.030 34.580 ;
        RECT 71.850 31.540 72.110 31.860 ;
        RECT 71.390 31.200 71.650 31.520 ;
        RECT 71.450 30.160 71.590 31.200 ;
        RECT 71.390 29.840 71.650 30.160 ;
        RECT 71.910 29.820 72.050 31.540 ;
        RECT 70.470 29.590 71.130 29.730 ;
        RECT 70.470 29.500 70.730 29.590 ;
        RECT 71.850 29.500 72.110 29.820 ;
        RECT 70.530 24.720 70.670 29.500 ;
        RECT 72.830 26.760 72.970 34.260 ;
        RECT 72.770 26.440 73.030 26.760 ;
        RECT 70.470 24.400 70.730 24.720 ;
        RECT 71.850 23.720 72.110 24.040 ;
        RECT 71.910 22.000 72.050 23.720 ;
        RECT 71.850 21.910 72.110 22.000 ;
        RECT 71.450 21.770 72.110 21.910 ;
        RECT 71.450 19.280 71.590 21.770 ;
        RECT 71.850 21.680 72.110 21.770 ;
        RECT 72.830 21.320 72.970 26.440 ;
        RECT 73.290 22.000 73.430 37.660 ;
        RECT 73.750 36.960 73.890 39.020 ;
        RECT 73.690 36.640 73.950 36.960 ;
        RECT 73.750 31.520 73.890 36.640 ;
        RECT 74.210 35.260 74.350 40.040 ;
        RECT 74.150 34.940 74.410 35.260 ;
        RECT 73.690 31.200 73.950 31.520 ;
        RECT 73.750 24.380 73.890 31.200 ;
        RECT 74.210 24.380 74.350 34.940 ;
        RECT 75.980 34.745 76.260 35.115 ;
        RECT 75.990 34.600 76.250 34.745 ;
        RECT 76.510 34.240 76.650 51.600 ;
        RECT 76.970 51.240 77.110 52.620 ;
        RECT 76.910 50.920 77.170 51.240 ;
        RECT 77.830 47.860 78.090 48.180 ;
        RECT 78.290 47.860 78.550 48.180 ;
        RECT 78.750 47.860 79.010 48.180 ;
        RECT 76.910 45.820 77.170 46.140 ;
        RECT 76.970 42.740 77.110 45.820 ;
        RECT 77.890 43.760 78.030 47.860 ;
        RECT 77.830 43.440 78.090 43.760 ;
        RECT 76.910 42.420 77.170 42.740 ;
        RECT 77.830 40.040 78.090 40.360 ;
        RECT 77.890 37.300 78.030 40.040 ;
        RECT 78.350 40.020 78.490 47.860 ;
        RECT 78.290 39.700 78.550 40.020 ;
        RECT 78.810 39.680 78.950 47.860 ;
        RECT 80.130 47.180 80.390 47.500 ;
        RECT 80.190 42.400 80.330 47.180 ;
        RECT 80.130 42.080 80.390 42.400 ;
        RECT 81.110 40.360 81.250 67.240 ;
        RECT 79.670 40.040 79.930 40.360 ;
        RECT 81.050 40.040 81.310 40.360 ;
        RECT 78.750 39.360 79.010 39.680 ;
        RECT 79.730 38.320 79.870 40.040 ;
        RECT 79.670 38.000 79.930 38.320 ;
        RECT 81.110 37.640 81.250 40.040 ;
        RECT 81.050 37.320 81.310 37.640 ;
        RECT 77.830 36.980 78.090 37.300 ;
        RECT 78.750 36.980 79.010 37.300 ;
        RECT 75.530 33.920 75.790 34.240 ;
        RECT 76.450 33.920 76.710 34.240 ;
        RECT 75.590 26.330 75.730 33.920 ;
        RECT 77.890 29.560 78.030 36.980 ;
        RECT 78.290 36.640 78.550 36.960 ;
        RECT 78.350 35.260 78.490 36.640 ;
        RECT 78.810 35.600 78.950 36.980 ;
        RECT 78.750 35.280 79.010 35.600 ;
        RECT 78.290 34.940 78.550 35.260 ;
        RECT 78.750 34.600 79.010 34.920 ;
        RECT 79.670 34.600 79.930 34.920 ;
        RECT 80.580 34.745 80.860 35.115 ;
        RECT 80.590 34.600 80.850 34.745 ;
        RECT 78.810 34.240 78.950 34.600 ;
        RECT 78.750 33.920 79.010 34.240 ;
        RECT 79.730 33.900 79.870 34.600 ;
        RECT 81.050 33.920 81.310 34.240 ;
        RECT 79.670 33.580 79.930 33.900 ;
        RECT 78.290 31.200 78.550 31.520 ;
        RECT 78.350 30.160 78.490 31.200 ;
        RECT 79.210 30.860 79.470 31.180 ;
        RECT 78.290 29.840 78.550 30.160 ;
        RECT 76.910 29.160 77.170 29.480 ;
        RECT 77.370 29.160 77.630 29.480 ;
        RECT 77.890 29.420 78.950 29.560 ;
        RECT 76.970 27.440 77.110 29.160 ;
        RECT 76.910 27.120 77.170 27.440 ;
        RECT 76.910 26.440 77.170 26.760 ;
        RECT 75.990 26.330 76.250 26.420 ;
        RECT 75.590 26.190 76.250 26.330 ;
        RECT 75.990 26.100 76.250 26.190 ;
        RECT 73.690 24.060 73.950 24.380 ;
        RECT 74.150 24.060 74.410 24.380 ;
        RECT 73.230 21.680 73.490 22.000 ;
        RECT 72.770 21.000 73.030 21.320 ;
        RECT 73.290 20.980 73.430 21.680 ;
        RECT 73.230 20.660 73.490 20.980 ;
        RECT 71.850 19.980 72.110 20.300 ;
        RECT 71.390 18.960 71.650 19.280 ;
        RECT 71.450 15.540 71.590 18.960 ;
        RECT 71.910 18.600 72.050 19.980 ;
        RECT 71.850 18.280 72.110 18.600 ;
        RECT 73.750 17.180 73.890 24.060 ;
        RECT 75.530 23.720 75.790 24.040 ;
        RECT 75.590 21.320 75.730 23.720 ;
        RECT 75.530 21.000 75.790 21.320 ;
        RECT 74.150 20.660 74.410 20.980 ;
        RECT 74.210 19.280 74.350 20.660 ;
        RECT 74.150 18.960 74.410 19.280 ;
        RECT 76.050 18.600 76.190 26.100 ;
        RECT 76.970 24.720 77.110 26.440 ;
        RECT 76.910 24.400 77.170 24.720 ;
        RECT 76.970 23.020 77.110 24.400 ;
        RECT 77.430 24.040 77.570 29.160 ;
        RECT 77.830 26.100 78.090 26.420 ;
        RECT 78.290 26.100 78.550 26.420 ;
        RECT 77.890 24.720 78.030 26.100 ;
        RECT 78.350 24.720 78.490 26.100 ;
        RECT 77.830 24.400 78.090 24.720 ;
        RECT 78.290 24.400 78.550 24.720 ;
        RECT 78.810 24.040 78.950 29.420 ;
        RECT 79.270 26.420 79.410 30.860 ;
        RECT 79.730 29.140 79.870 33.580 ;
        RECT 81.110 29.480 81.250 33.920 ;
        RECT 81.050 29.160 81.310 29.480 ;
        RECT 79.670 28.820 79.930 29.140 ;
        RECT 81.570 28.880 81.710 69.280 ;
        RECT 83.350 68.940 83.610 69.260 ;
        RECT 84.270 68.940 84.530 69.260 ;
        RECT 85.650 68.940 85.910 69.260 ;
        RECT 82.430 67.580 82.690 67.900 ;
        RECT 82.490 65.520 82.630 67.580 ;
        RECT 82.430 65.200 82.690 65.520 ;
        RECT 81.970 60.780 82.230 61.100 ;
        RECT 82.030 59.060 82.170 60.780 ;
        RECT 81.970 58.740 82.230 59.060 ;
        RECT 82.430 56.360 82.690 56.680 ;
        RECT 82.490 46.480 82.630 56.360 ;
        RECT 83.410 53.960 83.550 68.940 ;
        RECT 84.330 68.435 84.470 68.940 ;
        RECT 84.260 68.065 84.540 68.435 ;
        RECT 85.190 67.920 85.450 68.240 ;
        RECT 84.270 66.220 84.530 66.540 ;
        RECT 84.330 64.840 84.470 66.220 ;
        RECT 85.250 64.840 85.390 67.920 ;
        RECT 84.270 64.520 84.530 64.840 ;
        RECT 85.190 64.520 85.450 64.840 ;
        RECT 85.710 64.160 85.850 68.940 ;
        RECT 85.650 63.840 85.910 64.160 ;
        RECT 83.810 63.500 84.070 63.820 ;
        RECT 83.870 62.800 84.010 63.500 ;
        RECT 86.170 62.800 86.310 69.620 ;
        RECT 86.630 66.880 86.770 75.060 ;
        RECT 87.090 73.000 87.230 76.080 ;
        RECT 87.550 75.380 87.690 77.100 ;
        RECT 135.980 76.240 136.210 77.560 ;
        RECT 137.200 77.550 137.530 77.560 ;
        RECT 138.160 77.550 138.490 77.560 ;
        RECT 135.980 75.900 138.980 76.240 ;
        RECT 87.490 75.060 87.750 75.380 ;
        RECT 88.400 74.865 88.680 75.235 ;
        RECT 88.470 74.700 88.610 74.865 ;
        RECT 88.410 74.380 88.670 74.700 ;
        RECT 87.030 72.680 87.290 73.000 ;
        RECT 88.860 71.465 89.140 71.835 ;
        RECT 88.410 69.620 88.670 69.940 ;
        RECT 88.470 68.240 88.610 69.620 ;
        RECT 87.030 67.920 87.290 68.240 ;
        RECT 88.410 67.920 88.670 68.240 ;
        RECT 86.570 66.560 86.830 66.880 ;
        RECT 86.570 64.180 86.830 64.500 ;
        RECT 83.810 62.480 84.070 62.800 ;
        RECT 86.110 62.480 86.370 62.800 ;
        RECT 84.270 61.460 84.530 61.780 ;
        RECT 84.330 60.080 84.470 61.460 ;
        RECT 86.630 60.080 86.770 64.180 ;
        RECT 87.090 62.120 87.230 67.920 ;
        RECT 88.930 67.560 89.070 71.465 ;
        RECT 88.870 67.240 89.130 67.560 ;
        RECT 88.410 65.035 88.670 65.180 ;
        RECT 88.400 64.665 88.680 65.035 ;
        RECT 87.950 64.180 88.210 64.500 ;
        RECT 87.030 61.800 87.290 62.120 ;
        RECT 87.490 61.800 87.750 62.120 ;
        RECT 84.270 59.760 84.530 60.080 ;
        RECT 86.570 59.760 86.830 60.080 ;
        RECT 83.810 55.340 84.070 55.660 ;
        RECT 86.110 55.340 86.370 55.660 ;
        RECT 83.870 53.960 84.010 55.340 ;
        RECT 86.170 53.960 86.310 55.340 ;
        RECT 83.350 53.640 83.610 53.960 ;
        RECT 83.810 53.640 84.070 53.960 ;
        RECT 86.110 53.640 86.370 53.960 ;
        RECT 87.550 50.560 87.690 61.800 ;
        RECT 88.010 60.080 88.150 64.180 ;
        RECT 88.400 61.265 88.680 61.635 ;
        RECT 88.410 61.120 88.670 61.265 ;
        RECT 87.950 59.760 88.210 60.080 ;
        RECT 88.410 55.340 88.670 55.660 ;
        RECT 88.470 54.835 88.610 55.340 ;
        RECT 88.400 54.465 88.680 54.835 ;
        RECT 88.870 53.640 89.130 53.960 ;
        RECT 88.930 51.240 89.070 53.640 ;
        RECT 88.870 50.920 89.130 51.240 ;
        RECT 87.490 50.240 87.750 50.560 ;
        RECT 83.350 47.520 83.610 47.840 ;
        RECT 82.430 46.160 82.690 46.480 ;
        RECT 81.970 42.420 82.230 42.740 ;
        RECT 82.030 37.300 82.170 42.420 ;
        RECT 83.410 40.360 83.550 47.520 ;
        RECT 87.490 45.480 87.750 45.800 ;
        RECT 87.550 42.060 87.690 45.480 ;
        RECT 89.330 44.800 89.590 45.120 ;
        RECT 89.390 44.635 89.530 44.800 ;
        RECT 89.320 44.265 89.600 44.635 ;
        RECT 87.490 41.740 87.750 42.060 ;
        RECT 83.350 40.040 83.610 40.360 ;
        RECT 83.350 39.360 83.610 39.680 ;
        RECT 81.970 36.980 82.230 37.300 ;
        RECT 82.030 34.580 82.170 36.980 ;
        RECT 83.410 35.260 83.550 39.360 ;
        RECT 85.650 36.300 85.910 36.620 ;
        RECT 83.350 34.940 83.610 35.260 ;
        RECT 85.710 34.920 85.850 36.300 ;
        RECT 87.490 35.280 87.750 35.600 ;
        RECT 85.650 34.600 85.910 34.920 ;
        RECT 81.970 34.260 82.230 34.580 ;
        RECT 82.030 29.820 82.170 34.260 ;
        RECT 82.430 32.220 82.690 32.540 ;
        RECT 81.970 29.500 82.230 29.820 ;
        RECT 81.110 28.740 81.710 28.880 ;
        RECT 80.130 28.140 80.390 28.460 ;
        RECT 79.670 26.440 79.930 26.760 ;
        RECT 79.210 26.100 79.470 26.420 ;
        RECT 79.210 25.420 79.470 25.740 ;
        RECT 79.270 24.040 79.410 25.420 ;
        RECT 77.370 23.720 77.630 24.040 ;
        RECT 77.830 23.720 78.090 24.040 ;
        RECT 78.750 23.950 79.010 24.040 ;
        RECT 78.350 23.810 79.010 23.950 ;
        RECT 76.910 22.700 77.170 23.020 ;
        RECT 77.370 20.660 77.630 20.980 ;
        RECT 77.430 20.300 77.570 20.660 ;
        RECT 77.370 19.980 77.630 20.300 ;
        RECT 77.890 18.600 78.030 23.720 ;
        RECT 78.350 21.660 78.490 23.810 ;
        RECT 78.750 23.720 79.010 23.810 ;
        RECT 79.210 23.720 79.470 24.040 ;
        RECT 78.750 22.700 79.010 23.020 ;
        RECT 78.290 21.340 78.550 21.660 ;
        RECT 78.810 20.980 78.950 22.700 ;
        RECT 78.290 20.660 78.550 20.980 ;
        RECT 78.750 20.660 79.010 20.980 ;
        RECT 79.210 20.660 79.470 20.980 ;
        RECT 75.990 18.280 76.250 18.600 ;
        RECT 77.830 18.280 78.090 18.600 ;
        RECT 75.990 17.600 76.250 17.920 ;
        RECT 72.830 17.040 73.890 17.180 ;
        RECT 63.570 15.220 63.830 15.540 ;
        RECT 66.330 15.220 66.590 15.540 ;
        RECT 69.550 15.220 69.810 15.540 ;
        RECT 71.390 15.220 71.650 15.540 ;
        RECT 72.830 15.200 72.970 17.040 ;
        RECT 76.050 15.540 76.190 17.600 ;
        RECT 78.350 16.560 78.490 20.660 ;
        RECT 78.750 18.960 79.010 19.280 ;
        RECT 78.290 16.240 78.550 16.560 ;
        RECT 78.810 15.880 78.950 18.960 ;
        RECT 79.270 17.580 79.410 20.660 ;
        RECT 79.730 18.940 79.870 26.440 ;
        RECT 80.190 26.420 80.330 28.140 ;
        RECT 80.130 26.100 80.390 26.420 ;
        RECT 80.190 20.980 80.330 26.100 ;
        RECT 81.110 24.380 81.250 28.740 ;
        RECT 81.510 28.140 81.770 28.460 ;
        RECT 81.570 27.100 81.710 28.140 ;
        RECT 81.510 26.780 81.770 27.100 ;
        RECT 82.030 26.760 82.170 29.500 ;
        RECT 81.970 26.440 82.230 26.760 ;
        RECT 81.970 25.760 82.230 26.080 ;
        RECT 81.050 24.060 81.310 24.380 ;
        RECT 82.030 23.700 82.170 25.760 ;
        RECT 81.970 23.380 82.230 23.700 ;
        RECT 80.130 20.660 80.390 20.980 ;
        RECT 80.190 20.300 80.330 20.660 ;
        RECT 80.130 19.980 80.390 20.300 ;
        RECT 81.050 19.980 81.310 20.300 ;
        RECT 81.970 19.980 82.230 20.300 ;
        RECT 79.670 18.620 79.930 18.940 ;
        RECT 79.730 18.260 79.870 18.620 ;
        RECT 81.110 18.600 81.250 19.980 ;
        RECT 81.050 18.280 81.310 18.600 ;
        RECT 79.670 17.940 79.930 18.260 ;
        RECT 79.210 17.260 79.470 17.580 ;
        RECT 79.730 15.880 79.870 17.940 ;
        RECT 82.030 16.560 82.170 19.980 ;
        RECT 82.490 18.600 82.630 32.220 ;
        RECT 84.730 29.500 84.990 29.820 ;
        RECT 84.270 29.160 84.530 29.480 ;
        RECT 84.330 25.740 84.470 29.160 ;
        RECT 84.270 25.420 84.530 25.740 ;
        RECT 84.270 23.720 84.530 24.040 ;
        RECT 83.810 21.340 84.070 21.660 ;
        RECT 83.350 19.980 83.610 20.300 ;
        RECT 82.430 18.280 82.690 18.600 ;
        RECT 81.970 16.240 82.230 16.560 ;
        RECT 78.750 15.560 79.010 15.880 ;
        RECT 79.670 15.560 79.930 15.880 ;
        RECT 83.410 15.540 83.550 19.980 ;
        RECT 75.990 15.220 76.250 15.540 ;
        RECT 83.350 15.220 83.610 15.540 ;
        RECT 38.730 14.880 38.990 15.200 ;
        RECT 48.390 14.880 48.650 15.200 ;
        RECT 61.730 14.880 61.990 15.200 ;
        RECT 72.770 14.880 73.030 15.200 ;
        RECT 38.790 7.310 38.930 14.880 ;
        RECT 41.490 14.540 41.750 14.860 ;
        RECT 45.170 14.540 45.430 14.860 ;
        RECT 47.930 14.540 48.190 14.860 ;
        RECT 51.610 14.540 51.870 14.860 ;
        RECT 54.830 14.540 55.090 14.860 ;
        RECT 58.050 14.540 58.310 14.860 ;
        RECT 61.270 14.540 61.530 14.860 ;
        RECT 64.490 14.540 64.750 14.860 ;
        RECT 67.710 14.540 67.970 14.860 ;
        RECT 70.930 14.540 71.190 14.860 ;
        RECT 74.150 14.540 74.410 14.860 ;
        RECT 41.550 8.480 41.690 14.540 ;
        RECT 41.550 8.340 42.150 8.480 ;
        RECT 42.010 7.310 42.150 8.340 ;
        RECT 45.230 7.310 45.370 14.540 ;
        RECT 47.990 9.160 48.130 14.540 ;
        RECT 47.990 9.020 48.590 9.160 ;
        RECT 48.450 7.310 48.590 9.020 ;
        RECT 51.670 7.310 51.810 14.540 ;
        RECT 54.890 7.310 55.030 14.540 ;
        RECT 58.110 7.310 58.250 14.540 ;
        RECT 61.330 7.310 61.470 14.540 ;
        RECT 64.550 7.310 64.690 14.540 ;
        RECT 67.770 7.310 67.910 14.540 ;
        RECT 70.990 7.310 71.130 14.540 ;
        RECT 74.210 7.310 74.350 14.540 ;
        RECT 77.370 9.780 77.630 10.100 ;
        RECT 77.430 7.310 77.570 9.780 ;
        RECT 80.590 8.760 80.850 9.080 ;
        RECT 80.650 7.310 80.790 8.760 ;
        RECT 83.870 7.310 84.010 21.340 ;
        RECT 84.330 15.200 84.470 23.720 ;
        RECT 84.790 20.980 84.930 29.500 ;
        RECT 85.710 24.040 85.850 34.600 ;
        RECT 87.550 31.860 87.690 35.280 ;
        RECT 87.490 31.540 87.750 31.860 ;
        RECT 89.330 31.035 89.590 31.180 ;
        RECT 89.320 30.665 89.600 31.035 ;
        RECT 88.870 25.420 89.130 25.740 ;
        RECT 88.930 24.040 89.070 25.420 ;
        RECT 85.650 23.720 85.910 24.040 ;
        RECT 88.870 23.720 89.130 24.040 ;
        RECT 93.470 23.380 93.730 23.700 ;
        RECT 90.250 23.040 90.510 23.360 ;
        RECT 87.030 22.700 87.290 23.020 ;
        RECT 84.730 20.660 84.990 20.980 ;
        RECT 86.570 20.660 86.830 20.980 ;
        RECT 85.650 19.980 85.910 20.300 ;
        RECT 84.270 14.880 84.530 15.200 ;
        RECT 85.710 9.080 85.850 19.980 ;
        RECT 86.630 19.280 86.770 20.660 ;
        RECT 86.570 18.960 86.830 19.280 ;
        RECT 85.650 8.760 85.910 9.080 ;
        RECT 87.090 7.310 87.230 22.700 ;
        RECT 87.950 17.260 88.210 17.580 ;
        RECT 88.010 10.100 88.150 17.260 ;
        RECT 87.950 9.780 88.210 10.100 ;
        RECT 90.310 7.310 90.450 23.040 ;
        RECT 93.530 7.310 93.670 23.380 ;
        RECT 6.520 3.310 6.800 7.310 ;
        RECT 9.740 3.310 10.020 7.310 ;
        RECT 12.960 3.310 13.240 7.310 ;
        RECT 16.180 3.310 16.460 7.310 ;
        RECT 19.400 3.310 19.680 7.310 ;
        RECT 22.620 3.310 22.900 7.310 ;
        RECT 25.840 3.310 26.120 7.310 ;
        RECT 29.060 3.310 29.340 7.310 ;
        RECT 32.280 3.310 32.560 7.310 ;
        RECT 35.500 3.310 35.780 7.310 ;
        RECT 38.720 3.310 39.000 7.310 ;
        RECT 41.940 3.310 42.220 7.310 ;
        RECT 45.160 3.310 45.440 7.310 ;
        RECT 48.380 3.310 48.660 7.310 ;
        RECT 51.600 3.310 51.880 7.310 ;
        RECT 54.820 3.310 55.100 7.310 ;
        RECT 58.040 3.310 58.320 7.310 ;
        RECT 61.260 3.310 61.540 7.310 ;
        RECT 64.480 3.310 64.760 7.310 ;
        RECT 67.700 3.310 67.980 7.310 ;
        RECT 70.920 3.310 71.200 7.310 ;
        RECT 74.140 3.310 74.420 7.310 ;
        RECT 77.360 3.310 77.640 7.310 ;
        RECT 80.580 3.310 80.860 7.310 ;
        RECT 83.800 3.310 84.080 7.310 ;
        RECT 87.020 3.310 87.300 7.310 ;
        RECT 90.240 3.310 90.520 7.310 ;
        RECT 93.460 3.310 93.740 7.310 ;
      LAYER met3 ;
        RECT 63.690 224.960 64.010 225.340 ;
        RECT 63.700 218.305 64.000 224.960 ;
        RECT 66.520 224.940 66.840 225.320 ;
        RECT 69.240 224.980 69.560 225.360 ;
        RECT 72.110 225.020 72.430 225.400 ;
        RECT 66.530 218.835 66.830 224.940 ;
        RECT 69.250 222.665 69.550 224.980 ;
        RECT 69.225 222.315 69.575 222.665 ;
        RECT 72.120 222.195 72.420 225.020 ;
        RECT 74.805 224.950 75.125 225.330 ;
        RECT 77.570 224.970 77.890 225.350 ;
        RECT 72.095 221.845 72.445 222.195 ;
        RECT 74.815 221.810 75.115 224.950 ;
        RECT 74.790 221.460 75.140 221.810 ;
        RECT 77.580 219.195 77.880 224.970 ;
        RECT 80.310 224.890 80.630 225.270 ;
        RECT 83.120 224.920 83.440 225.300 ;
        RECT 85.820 225.000 86.140 225.380 ;
        RECT 80.320 221.330 80.620 224.890 ;
        RECT 80.295 220.980 80.645 221.330 ;
        RECT 83.130 221.005 83.430 224.920 ;
        RECT 83.105 220.655 83.455 221.005 ;
        RECT 85.830 220.620 86.130 225.000 ;
        RECT 88.590 224.930 88.910 225.310 ;
        RECT 91.315 224.960 91.635 225.340 ;
        RECT 93.990 224.990 94.310 225.370 ;
        RECT 142.460 225.130 142.780 225.440 ;
        RECT 85.805 220.270 86.155 220.620 ;
        RECT 88.600 219.595 88.900 224.930 ;
        RECT 91.325 220.245 91.625 224.960 ;
        RECT 91.300 219.895 91.650 220.245 ;
        RECT 94.000 219.905 94.300 224.990 ;
        RECT 142.400 224.815 142.840 225.130 ;
        RECT 115.120 220.825 115.720 224.815 ;
        RECT 115.120 220.815 116.250 220.825 ;
        RECT 125.320 220.815 125.920 224.815 ;
        RECT 132.120 220.815 132.720 224.815 ;
        RECT 138.920 220.815 139.520 224.815 ;
        RECT 142.320 220.815 142.920 224.815 ;
        RECT 115.270 220.610 116.250 220.815 ;
        RECT 115.270 220.525 116.265 220.610 ;
        RECT 115.935 220.280 116.265 220.525 ;
        RECT 88.575 219.245 88.925 219.595 ;
        RECT 93.975 219.555 94.325 219.905 ;
        RECT 77.555 218.845 77.905 219.195 ;
        RECT 66.505 218.485 66.855 218.835 ;
        RECT 125.470 218.310 125.770 220.815 ;
        RECT 132.270 220.455 132.570 220.815 ;
        RECT 132.255 220.125 132.585 220.455 ;
        RECT 132.270 218.310 132.570 220.125 ;
        RECT 139.070 218.310 139.370 220.815 ;
        RECT 63.675 217.955 64.025 218.305 ;
        RECT 125.455 217.980 125.785 218.310 ;
        RECT 132.255 217.980 132.585 218.310 ;
        RECT 139.055 217.980 139.385 218.310 ;
        RECT 142.470 207.270 142.770 220.815 ;
        RECT 143.815 208.320 144.145 208.650 ;
        RECT 142.455 206.940 142.785 207.270 ;
        RECT 143.830 204.510 144.130 208.320 ;
        RECT 143.815 204.180 144.145 204.510 ;
        RECT 8.180 203.770 9.760 203.795 ;
        RECT 1.125 202.180 9.765 203.770 ;
        RECT 103.875 203.765 105.465 203.770 ;
        RECT 103.850 202.185 105.490 203.765 ;
        RECT 114.915 202.185 115.245 203.765 ;
        RECT 120.355 202.185 120.685 203.765 ;
        RECT 125.795 202.185 126.125 203.765 ;
        RECT 131.235 202.185 131.565 203.765 ;
        RECT 136.675 202.185 137.005 203.765 ;
        RECT 142.115 202.185 142.445 203.765 ;
        RECT 8.180 202.155 9.760 202.180 ;
        RECT 27.480 201.705 29.060 202.035 ;
        RECT 100.980 199.740 102.620 200.510 ;
        RECT 30.780 198.985 32.360 199.315 ;
        RECT 6.955 198.960 7.285 198.975 ;
        RECT 6.955 198.660 11.640 198.960 ;
        RECT 6.955 198.645 7.285 198.660 ;
        RECT 6.430 197.600 10.430 197.750 ;
        RECT 11.340 197.600 11.640 198.660 ;
        RECT 6.430 197.300 11.640 197.600 ;
        RECT 6.430 197.150 10.430 197.300 ;
        RECT 27.480 196.265 29.060 196.595 ;
        RECT 30.780 193.545 32.360 193.875 ;
        RECT 44.675 192.840 45.005 192.855 ;
        RECT 50.195 192.840 50.525 192.855 ;
        RECT 44.675 192.540 50.525 192.840 ;
        RECT 44.675 192.525 45.005 192.540 ;
        RECT 50.195 192.525 50.525 192.540 ;
        RECT 27.480 190.825 29.060 191.155 ;
        RECT 30.780 188.105 32.360 188.435 ;
        RECT 27.480 185.385 29.060 185.715 ;
        RECT 101.005 184.070 102.595 199.740 ;
        RECT 59.395 184.000 59.725 184.015 ;
        RECT 62.155 184.000 62.485 184.015 ;
        RECT 59.395 183.700 62.485 184.000 ;
        RECT 59.395 183.685 59.725 183.700 ;
        RECT 62.155 183.685 62.485 183.700 ;
        RECT 30.780 182.665 32.360 182.995 ;
        RECT 100.970 182.410 102.630 184.070 ;
        RECT 27.480 179.945 29.060 180.275 ;
        RECT 30.780 177.225 32.360 177.555 ;
        RECT 103.875 176.485 105.465 202.185 ;
        RECT 109.840 198.890 113.500 200.480 ;
        RECT 112.195 198.885 112.525 198.890 ;
        RECT 117.635 198.885 117.965 200.465 ;
        RECT 123.075 198.885 123.405 200.465 ;
        RECT 128.515 198.885 128.845 200.465 ;
        RECT 133.955 198.885 134.285 200.465 ;
        RECT 139.395 198.885 139.725 200.465 ;
        RECT 115.255 193.600 115.585 193.930 ;
        RECT 111.855 189.000 112.185 189.330 ;
        RECT 108.455 185.320 108.785 185.650 ;
        RECT 108.470 181.770 108.770 185.320 ;
        RECT 111.870 181.770 112.170 189.000 ;
        RECT 115.270 181.770 115.570 193.600 ;
        RECT 125.455 192.220 125.785 192.550 ;
        RECT 118.655 190.840 118.985 191.170 ;
        RECT 118.670 181.770 118.970 190.840 ;
        RECT 122.055 188.540 122.385 188.870 ;
        RECT 122.070 181.770 122.370 188.540 ;
        RECT 125.470 181.770 125.770 192.220 ;
        RECT 143.830 191.170 144.130 204.180 ;
        RECT 147.555 202.185 147.885 203.765 ;
        RECT 144.835 198.885 145.165 200.465 ;
        RECT 148.095 195.430 148.445 195.780 ;
        RECT 143.815 190.840 144.145 191.170 ;
        RECT 128.855 189.920 129.185 190.250 ;
        RECT 128.870 181.770 129.170 189.920 ;
        RECT 135.655 187.160 135.985 187.490 ;
        RECT 132.255 184.860 132.585 185.190 ;
        RECT 132.270 181.770 132.570 184.860 ;
        RECT 135.670 181.770 135.970 187.160 ;
        RECT 145.855 186.240 146.185 186.570 ;
        RECT 139.055 184.860 139.385 185.190 ;
        RECT 142.455 184.860 142.785 185.190 ;
        RECT 139.070 181.770 139.370 184.860 ;
        RECT 142.470 181.770 142.770 184.860 ;
        RECT 145.870 181.770 146.170 186.240 ;
        RECT 108.320 177.770 108.920 181.770 ;
        RECT 111.720 177.770 112.320 181.770 ;
        RECT 115.120 177.770 115.720 181.770 ;
        RECT 118.520 177.770 119.120 181.770 ;
        RECT 121.920 177.770 122.520 181.770 ;
        RECT 125.320 177.770 125.920 181.770 ;
        RECT 128.720 177.770 129.320 181.770 ;
        RECT 132.120 177.770 132.720 181.770 ;
        RECT 135.520 177.770 136.120 181.770 ;
        RECT 138.920 177.770 139.520 181.770 ;
        RECT 142.320 177.770 142.920 181.770 ;
        RECT 145.720 177.770 146.320 181.770 ;
        RECT 111.850 177.430 112.190 177.770 ;
        RECT 111.855 177.355 112.185 177.430 ;
        RECT 139.070 176.850 139.370 177.770 ;
        RECT 142.450 177.440 142.790 177.770 ;
        RECT 142.455 177.255 142.785 177.440 ;
        RECT 148.120 177.395 148.420 195.430 ;
        RECT 149.255 187.620 149.585 187.950 ;
        RECT 149.270 181.770 149.570 187.620 ;
        RECT 152.655 184.860 152.985 185.190 ;
        RECT 152.670 181.770 152.970 184.860 ;
        RECT 149.120 177.770 149.720 181.770 ;
        RECT 152.520 177.770 153.120 181.770 ;
        RECT 149.255 177.725 149.585 177.770 ;
        RECT 148.105 177.065 148.435 177.395 ;
        RECT 144.655 176.850 144.985 176.865 ;
        RECT 117.980 176.485 118.880 176.640 ;
        RECT 137.800 176.485 138.700 176.620 ;
        RECT 139.070 176.550 144.985 176.850 ;
        RECT 144.655 176.535 144.985 176.550 ;
        RECT 103.865 176.250 138.700 176.485 ;
        RECT 157.570 176.250 158.470 176.600 ;
        RECT 103.865 176.230 144.350 176.250 ;
        RECT 145.300 176.230 158.470 176.250 ;
        RECT 103.865 175.110 158.470 176.230 ;
        RECT 103.865 174.875 138.700 175.110 ;
        RECT 27.480 174.505 29.060 174.835 ;
        RECT 117.980 174.620 118.880 174.875 ;
        RECT 137.800 174.600 138.700 174.875 ;
        RECT 157.570 174.580 158.470 175.110 ;
        RECT 68.595 173.800 68.925 173.815 ;
        RECT 71.815 173.800 72.145 173.815 ;
        RECT 68.595 173.500 72.145 173.800 ;
        RECT 68.595 173.485 68.925 173.500 ;
        RECT 71.815 173.485 72.145 173.500 ;
        RECT 30.780 171.785 32.360 172.115 ;
        RECT 27.480 169.065 29.060 169.395 ;
        RECT 108.820 169.350 109.400 169.400 ;
        RECT 128.680 169.350 129.260 169.390 ;
        RECT 148.880 169.350 149.460 169.370 ;
        RECT 108.800 168.720 149.480 169.350 ;
        RECT 30.780 166.345 32.360 166.675 ;
        RECT 27.480 163.625 29.060 163.955 ;
        RECT 30.780 160.905 32.360 161.235 ;
        RECT 27.480 158.185 29.060 158.515 ;
        RECT 30.780 155.465 32.360 155.795 ;
        RECT 128.680 154.340 129.260 154.430 ;
        RECT 139.065 154.340 139.695 168.720 ;
        RECT 108.740 153.710 149.500 154.340 ;
        RECT 108.790 153.690 109.370 153.710 ;
        RECT 27.480 152.745 29.060 153.075 ;
        RECT 30.780 150.025 32.360 150.355 ;
        RECT 27.480 147.305 29.060 147.635 ;
        RECT 30.780 144.585 32.360 144.915 ;
        RECT 27.480 141.865 29.060 142.195 ;
        RECT 52.955 140.480 53.285 140.495 ;
        RECT 70.435 140.480 70.765 140.495 ;
        RECT 52.955 140.180 70.765 140.480 ;
        RECT 52.955 140.165 53.285 140.180 ;
        RECT 70.435 140.165 70.765 140.180 ;
        RECT 30.780 139.145 32.360 139.475 ;
        RECT 108.790 139.340 109.370 139.370 ;
        RECT 128.680 139.340 129.260 139.360 ;
        RECT 139.065 139.340 139.695 153.710 ;
        RECT 108.790 138.740 149.490 139.340 ;
        RECT 108.810 138.710 149.490 138.740 ;
        RECT 10.635 137.080 10.965 137.095 ;
        RECT 10.420 136.765 10.965 137.080 ;
        RECT 10.420 136.550 10.720 136.765 ;
        RECT 6.430 136.100 10.720 136.550 ;
        RECT 27.480 136.425 29.060 136.755 ;
        RECT 6.430 135.950 10.430 136.100 ;
        RECT 30.780 133.705 32.360 134.035 ;
        RECT 27.480 130.985 29.060 131.315 ;
        RECT 30.780 128.265 32.360 128.595 ;
        RECT 27.480 125.545 29.060 125.875 ;
        RECT 128.610 124.380 129.190 124.420 ;
        RECT 139.065 124.380 139.695 138.710 ;
        RECT 148.830 138.670 149.410 138.710 ;
        RECT 108.800 124.370 149.530 124.380 ;
        RECT 108.790 123.750 149.530 124.370 ;
        RECT 108.790 123.740 109.370 123.750 ;
        RECT 30.780 122.825 32.360 123.155 ;
        RECT 27.480 120.105 29.060 120.435 ;
        RECT 30.780 117.385 32.360 117.715 ;
        RECT 10.635 116.680 10.965 116.695 ;
        RECT 10.420 116.365 10.965 116.680 ;
        RECT 10.420 116.150 10.720 116.365 ;
        RECT 6.430 115.700 10.720 116.150 ;
        RECT 88.375 116.000 88.705 116.015 ;
        RECT 92.430 116.000 96.430 116.150 ;
        RECT 88.375 115.700 96.430 116.000 ;
        RECT 6.430 115.550 10.430 115.700 ;
        RECT 88.375 115.685 88.705 115.700 ;
        RECT 92.430 115.550 96.430 115.700 ;
        RECT 27.480 114.665 29.060 114.995 ;
        RECT 10.635 113.280 10.965 113.295 ;
        RECT 10.420 112.965 10.965 113.280 ;
        RECT 10.420 112.750 10.720 112.965 ;
        RECT 6.430 112.300 10.720 112.750 ;
        RECT 88.375 112.600 88.705 112.615 ;
        RECT 92.430 112.600 96.430 112.750 ;
        RECT 88.375 112.300 96.430 112.600 ;
        RECT 6.430 112.150 10.430 112.300 ;
        RECT 88.375 112.285 88.705 112.300 ;
        RECT 30.780 111.945 32.360 112.275 ;
        RECT 92.430 112.150 96.430 112.300 ;
        RECT 6.430 109.200 10.430 109.350 ;
        RECT 27.480 109.225 29.060 109.555 ;
        RECT 128.730 109.330 129.310 109.390 ;
        RECT 139.065 109.330 139.695 123.750 ;
        RECT 148.910 109.330 149.490 109.420 ;
        RECT 12.935 109.200 13.265 109.215 ;
        RECT 6.430 108.900 13.265 109.200 ;
        RECT 6.430 108.750 10.430 108.900 ;
        RECT 12.935 108.885 13.265 108.900 ;
        RECT 108.740 108.790 149.490 109.330 ;
        RECT 108.740 108.700 149.420 108.790 ;
        RECT 30.780 106.505 32.360 106.835 ;
        RECT 6.430 105.800 10.430 105.950 ;
        RECT 21.675 105.800 22.005 105.815 ;
        RECT 6.430 105.500 22.005 105.800 ;
        RECT 6.430 105.350 10.430 105.500 ;
        RECT 21.675 105.485 22.005 105.500 ;
        RECT 27.480 103.785 29.060 104.115 ;
        RECT 10.635 103.080 10.965 103.095 ;
        RECT 10.420 102.765 10.965 103.080 ;
        RECT 10.420 102.550 10.720 102.765 ;
        RECT 6.430 102.100 10.720 102.550 ;
        RECT 139.065 102.305 139.695 108.700 ;
        RECT 6.430 101.950 10.430 102.100 ;
        RECT 139.065 101.675 158.365 102.305 ;
        RECT 30.780 101.065 32.360 101.395 ;
        RECT 71.815 99.680 72.145 99.695 ;
        RECT 77.795 99.680 78.125 99.695 ;
        RECT 71.815 99.380 78.125 99.680 ;
        RECT 71.815 99.365 72.145 99.380 ;
        RECT 77.795 99.365 78.125 99.380 ;
        RECT 27.480 98.345 29.060 98.675 ;
        RECT 157.735 96.565 158.365 101.675 ;
        RECT 30.780 95.625 32.360 95.955 ;
        RECT 65.375 95.600 65.705 95.615 ;
        RECT 74.115 95.600 74.445 95.615 ;
        RECT 65.375 95.300 74.445 95.600 ;
        RECT 65.375 95.285 65.705 95.300 ;
        RECT 74.115 95.285 74.445 95.300 ;
        RECT 27.480 92.905 29.060 93.235 ;
        RECT 30.780 90.185 32.360 90.515 ;
        RECT 88.375 88.800 88.705 88.815 ;
        RECT 92.430 88.800 96.430 88.950 ;
        RECT 88.375 88.500 96.430 88.800 ;
        RECT 88.375 88.485 88.705 88.500 ;
        RECT 92.430 88.350 96.430 88.500 ;
        RECT 27.480 87.465 29.060 87.795 ;
        RECT 30.780 84.745 32.360 85.075 ;
        RECT 68.595 82.680 68.925 82.695 ;
        RECT 71.355 82.680 71.685 82.695 ;
        RECT 68.595 82.380 71.685 82.680 ;
        RECT 68.595 82.365 68.925 82.380 ;
        RECT 71.355 82.365 71.685 82.380 ;
        RECT 27.480 82.025 29.060 82.355 ;
        RECT 88.375 82.000 88.705 82.015 ;
        RECT 92.430 82.000 96.430 82.150 ;
        RECT 88.375 81.700 96.430 82.000 ;
        RECT 88.375 81.685 88.705 81.700 ;
        RECT 92.430 81.550 96.430 81.700 ;
        RECT 30.780 79.305 32.360 79.635 ;
        RECT 72.275 79.280 72.605 79.295 ;
        RECT 74.115 79.280 74.445 79.295 ;
        RECT 72.275 78.980 74.445 79.280 ;
        RECT 72.275 78.965 72.605 78.980 ;
        RECT 74.115 78.965 74.445 78.980 ;
        RECT 27.480 76.585 29.060 76.915 ;
        RECT 88.375 75.200 88.705 75.215 ;
        RECT 92.430 75.200 96.430 75.350 ;
        RECT 88.375 74.900 96.430 75.200 ;
        RECT 88.375 74.885 88.705 74.900 ;
        RECT 92.430 74.750 96.430 74.900 ;
        RECT 30.780 73.865 32.360 74.195 ;
        RECT 67.215 73.160 67.545 73.175 ;
        RECT 73.655 73.160 73.985 73.175 ;
        RECT 67.215 72.860 73.985 73.160 ;
        RECT 67.215 72.845 67.545 72.860 ;
        RECT 73.655 72.845 73.985 72.860 ;
        RECT 67.675 72.480 68.005 72.495 ;
        RECT 70.895 72.480 71.225 72.495 ;
        RECT 67.675 72.180 71.225 72.480 ;
        RECT 67.675 72.165 68.005 72.180 ;
        RECT 70.895 72.165 71.225 72.180 ;
        RECT 88.835 71.800 89.165 71.815 ;
        RECT 92.430 71.800 96.430 71.950 ;
        RECT 88.835 71.500 96.430 71.800 ;
        RECT 88.835 71.485 89.165 71.500 ;
        RECT 27.480 71.145 29.060 71.475 ;
        RECT 92.430 71.350 96.430 71.500 ;
        RECT 6.430 68.400 10.430 68.550 ;
        RECT 30.780 68.425 32.360 68.755 ;
        RECT 12.935 68.400 13.265 68.415 ;
        RECT 6.430 68.100 13.265 68.400 ;
        RECT 6.430 67.950 10.430 68.100 ;
        RECT 12.935 68.085 13.265 68.100 ;
        RECT 84.235 68.400 84.565 68.415 ;
        RECT 92.430 68.400 96.430 68.550 ;
        RECT 84.235 68.100 96.430 68.400 ;
        RECT 84.235 68.085 84.565 68.100 ;
        RECT 92.430 67.950 96.430 68.100 ;
        RECT 42.375 66.370 42.705 66.375 ;
        RECT 42.375 66.360 42.960 66.370 ;
        RECT 42.375 66.060 43.160 66.360 ;
        RECT 42.375 66.050 42.960 66.060 ;
        RECT 42.375 66.045 42.705 66.050 ;
        RECT 27.480 65.705 29.060 66.035 ;
        RECT 6.430 65.000 10.430 65.150 ;
        RECT 88.375 65.000 88.705 65.015 ;
        RECT 92.430 65.000 96.430 65.150 ;
        RECT 6.430 64.550 10.720 65.000 ;
        RECT 88.375 64.700 96.430 65.000 ;
        RECT 88.375 64.685 88.705 64.700 ;
        RECT 92.430 64.550 96.430 64.700 ;
        RECT 10.420 64.335 10.720 64.550 ;
        RECT 10.420 64.020 10.965 64.335 ;
        RECT 10.635 64.005 10.965 64.020 ;
        RECT 30.780 62.985 32.360 63.315 ;
        RECT 6.430 61.600 10.430 61.750 ;
        RECT 12.015 61.600 12.345 61.615 ;
        RECT 6.430 61.300 12.345 61.600 ;
        RECT 6.430 61.150 10.430 61.300 ;
        RECT 12.015 61.285 12.345 61.300 ;
        RECT 88.375 61.600 88.705 61.615 ;
        RECT 92.430 61.600 96.430 61.750 ;
        RECT 88.375 61.300 96.430 61.600 ;
        RECT 88.375 61.285 88.705 61.300 ;
        RECT 92.430 61.150 96.430 61.300 ;
        RECT 66.295 60.920 66.625 60.935 ;
        RECT 71.355 60.920 71.685 60.935 ;
        RECT 66.295 60.620 71.685 60.920 ;
        RECT 66.295 60.605 66.625 60.620 ;
        RECT 71.355 60.605 71.685 60.620 ;
        RECT 27.480 60.265 29.060 60.595 ;
        RECT 6.430 58.200 10.430 58.350 ;
        RECT 15.695 58.200 16.025 58.215 ;
        RECT 6.430 57.900 16.025 58.200 ;
        RECT 6.430 57.750 10.430 57.900 ;
        RECT 15.695 57.885 16.025 57.900 ;
        RECT 30.780 57.545 32.360 57.875 ;
        RECT 19.375 56.840 19.705 56.855 ;
        RECT 20.295 56.840 20.625 56.855 ;
        RECT 19.375 56.540 20.625 56.840 ;
        RECT 19.375 56.525 19.705 56.540 ;
        RECT 20.295 56.525 20.625 56.540 ;
        RECT 6.430 54.800 10.430 54.950 ;
        RECT 27.480 54.825 29.060 55.155 ;
        RECT 12.935 54.800 13.265 54.815 ;
        RECT 6.430 54.500 13.265 54.800 ;
        RECT 6.430 54.350 10.430 54.500 ;
        RECT 12.935 54.485 13.265 54.500 ;
        RECT 88.375 54.800 88.705 54.815 ;
        RECT 92.430 54.800 96.430 54.950 ;
        RECT 88.375 54.500 96.430 54.800 ;
        RECT 88.375 54.485 88.705 54.500 ;
        RECT 92.430 54.350 96.430 54.500 ;
        RECT 30.780 52.105 32.360 52.435 ;
        RECT 6.430 51.400 10.430 51.550 ;
        RECT 11.555 51.400 11.885 51.415 ;
        RECT 6.430 51.100 11.885 51.400 ;
        RECT 6.430 50.950 10.430 51.100 ;
        RECT 11.555 51.085 11.885 51.100 ;
        RECT 27.480 49.385 29.060 49.715 ;
        RECT 10.635 48.680 10.965 48.695 ;
        RECT 10.420 48.365 10.965 48.680 ;
        RECT 10.420 48.150 10.720 48.365 ;
        RECT 6.430 47.700 10.720 48.150 ;
        RECT 29.700 48.000 30.080 48.010 ;
        RECT 32.255 48.000 32.585 48.015 ;
        RECT 29.700 47.700 32.585 48.000 ;
        RECT 6.430 47.550 10.430 47.700 ;
        RECT 29.700 47.690 30.080 47.700 ;
        RECT 32.255 47.685 32.585 47.700 ;
        RECT 30.780 46.665 32.360 46.995 ;
        RECT 6.430 44.600 10.430 44.750 ;
        RECT 20.295 44.600 20.625 44.615 ;
        RECT 6.430 44.300 20.625 44.600 ;
        RECT 6.430 44.150 10.430 44.300 ;
        RECT 20.295 44.285 20.625 44.300 ;
        RECT 89.295 44.600 89.625 44.615 ;
        RECT 92.430 44.600 96.430 44.750 ;
        RECT 89.295 44.300 96.430 44.600 ;
        RECT 89.295 44.285 89.625 44.300 ;
        RECT 27.480 43.945 29.060 44.275 ;
        RECT 92.430 44.150 96.430 44.300 ;
        RECT 6.430 41.200 10.430 41.350 ;
        RECT 30.780 41.225 32.360 41.555 ;
        RECT 21.215 41.200 21.545 41.215 ;
        RECT 6.430 40.900 21.545 41.200 ;
        RECT 6.430 40.750 10.430 40.900 ;
        RECT 21.215 40.885 21.545 40.900 ;
        RECT 18.455 39.840 18.785 39.855 ;
        RECT 48.355 39.840 48.685 39.855 ;
        RECT 18.455 39.540 48.685 39.840 ;
        RECT 18.455 39.525 18.785 39.540 ;
        RECT 48.355 39.525 48.685 39.540 ;
        RECT 27.480 38.505 29.060 38.835 ;
        RECT 30.780 35.785 32.360 36.115 ;
        RECT 75.955 35.080 76.285 35.095 ;
        RECT 80.555 35.080 80.885 35.095 ;
        RECT 75.955 34.780 80.885 35.080 ;
        RECT 75.955 34.765 76.285 34.780 ;
        RECT 80.555 34.765 80.885 34.780 ;
        RECT 27.480 33.065 29.060 33.395 ;
        RECT 89.295 31.000 89.625 31.015 ;
        RECT 92.430 31.000 96.430 31.150 ;
        RECT 89.295 30.700 96.430 31.000 ;
        RECT 89.295 30.685 89.625 30.700 ;
        RECT 30.780 30.345 32.360 30.675 ;
        RECT 92.430 30.550 96.430 30.700 ;
        RECT 27.480 27.625 29.060 27.955 ;
        RECT 30.780 24.905 32.360 25.235 ;
        RECT 23.975 24.200 24.305 24.215 ;
        RECT 39.155 24.200 39.485 24.215 ;
        RECT 45.595 24.200 45.925 24.215 ;
        RECT 23.975 23.900 45.925 24.200 ;
        RECT 23.975 23.885 24.305 23.900 ;
        RECT 39.155 23.885 39.485 23.900 ;
        RECT 45.595 23.885 45.925 23.900 ;
        RECT 42.580 23.520 42.960 23.530 ;
        RECT 63.995 23.520 64.325 23.535 ;
        RECT 42.580 23.220 64.325 23.520 ;
        RECT 42.580 23.210 42.960 23.220 ;
        RECT 63.995 23.205 64.325 23.220 ;
        RECT 27.480 22.185 29.060 22.515 ;
        RECT 27.655 21.480 27.985 21.495 ;
        RECT 29.700 21.480 30.080 21.490 ;
        RECT 42.835 21.480 43.165 21.495 ;
        RECT 27.655 21.180 43.165 21.480 ;
        RECT 27.655 21.165 27.985 21.180 ;
        RECT 29.700 21.170 30.080 21.180 ;
        RECT 42.835 21.165 43.165 21.180 ;
        RECT 30.780 19.465 32.360 19.795 ;
        RECT 27.480 16.745 29.060 17.075 ;
        RECT 30.780 14.025 32.360 14.355 ;
      LAYER met4 ;
        RECT 63.685 224.985 63.790 225.315 ;
        RECT 66.515 224.965 66.550 225.295 ;
        RECT 69.235 225.005 69.310 225.335 ;
        RECT 72.370 225.045 72.435 225.375 ;
        RECT 74.800 224.975 74.830 225.305 ;
        RECT 77.565 224.995 77.590 225.325 ;
        RECT 77.890 224.995 77.895 225.325 ;
        RECT 80.305 224.915 80.350 225.245 ;
        RECT 83.410 224.945 83.445 225.275 ;
        RECT 85.815 225.025 85.870 225.355 ;
        RECT 88.585 224.955 88.630 225.285 ;
        RECT 91.310 224.985 91.390 225.315 ;
        RECT 93.985 225.015 94.150 225.345 ;
        RECT 118.795 224.760 118.990 225.215 ;
        RECT 119.290 224.760 119.455 225.215 ;
        RECT 121.530 224.805 121.750 225.455 ;
        RECT 122.050 224.805 122.190 225.455 ;
        RECT 124.275 224.945 124.510 225.595 ;
        RECT 124.810 224.945 124.935 225.595 ;
        RECT 127.145 224.965 127.270 225.615 ;
        RECT 127.570 224.965 127.805 225.615 ;
        RECT 129.605 224.960 130.030 225.610 ;
        RECT 133.090 224.945 133.645 225.595 ;
        RECT 134.915 225.075 135.550 225.725 ;
        RECT 137.630 224.895 138.310 225.575 ;
        RECT 142.455 225.400 142.785 225.415 ;
        RECT 142.455 225.100 143.830 225.400 ;
        RECT 142.455 225.085 142.785 225.100 ;
        RECT 118.795 224.565 119.455 224.760 ;
        RECT 112.120 203.770 147.960 203.775 ;
        RECT 98.780 202.180 147.960 203.770 ;
        RECT 112.120 202.175 147.960 202.180 ;
        RECT 6.000 198.890 6.020 200.480 ;
        RECT 27.470 13.950 29.070 202.110 ;
        RECT 29.725 47.685 30.055 48.015 ;
        RECT 29.740 21.495 30.040 47.685 ;
        RECT 29.725 21.165 30.055 21.495 ;
        RECT 30.770 13.950 32.370 202.110 ;
        RECT 98.780 200.475 113.500 200.480 ;
        RECT 98.780 198.890 147.960 200.475 ;
        RECT 112.120 198.875 147.960 198.890 ;
        RECT 157.730 96.590 158.370 97.230 ;
        RECT 42.605 66.045 42.935 66.375 ;
        RECT 42.620 23.535 42.920 66.045 ;
        RECT 42.605 23.205 42.935 23.535 ;
        RECT 157.735 1.065 158.365 96.590 ;
        RECT 16.570 1.000 17.470 1.040 ;
        RECT 35.890 1.000 36.790 1.040 ;
        RECT 55.210 1.000 56.110 1.030 ;
        RECT 132.490 1.000 133.390 1.010 ;
        RECT 152.045 1.000 158.365 1.065 ;
        RECT 152.710 0.435 158.365 1.000 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

