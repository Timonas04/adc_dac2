magic
tech sky130A
magscale 1 2
timestamp 1730635755
<< pwell >>
rect 1336 -2940 1368 -2886
rect 1002 -3120 3340 -2940
rect 1336 -4190 1368 -3120
rect 1336 -4220 1400 -4190
<< psubdiff >>
rect 1336 -4190 1368 -2886
rect 1336 -4220 1400 -4190
<< locali >>
rect 1046 -370 3588 -358
rect 1054 -2698 3592 -2688
rect 1054 -2886 3592 -2878
rect 1336 -4190 1368 -2886
rect 1336 -4220 1400 -4190
<< viali >>
rect 1046 -358 3588 -208
rect 1054 -2878 3592 -2698
<< metal1 >>
rect 1038 -196 3600 -192
rect 1034 -208 3602 -196
rect 1034 -358 1046 -208
rect 3588 -358 3602 -208
rect 1038 -370 3600 -358
rect 1066 -452 1112 -446
rect 1066 -1630 1184 -452
rect 1238 -1630 1326 -370
rect 1554 -392 1786 -370
rect 1400 -1626 1502 -456
rect 1554 -1626 1642 -392
rect 1702 -1374 1824 -456
rect 1400 -1630 1432 -1626
rect 1474 -1630 1502 -1626
rect 1066 -1686 1114 -1630
rect 1182 -1640 1184 -1630
rect 1402 -1678 1432 -1630
rect 1698 -1632 1824 -1374
rect 1872 -1624 1960 -370
rect 2014 -1632 2128 -452
rect 2190 -1626 2278 -370
rect 1066 -2172 1142 -1686
rect 1180 -1834 1244 -1688
rect 1170 -2034 1370 -1834
rect 1180 -2172 1244 -2034
rect 1066 -2234 1114 -2172
rect 1190 -2180 1244 -2172
rect 1402 -2184 1442 -1678
rect 1496 -1824 1564 -1684
rect 1470 -2024 1670 -1824
rect 1496 -2178 1564 -2024
rect 1066 -2236 1186 -2234
rect 1060 -2596 1070 -2236
rect 1134 -2596 1186 -2236
rect 1242 -2590 1346 -2228
rect 1402 -2236 1432 -2184
rect 1482 -2236 1502 -2226
rect 1402 -2238 1502 -2236
rect 1066 -2600 1112 -2596
rect 1242 -2600 1256 -2590
rect 1312 -2654 1346 -2590
rect 1394 -2598 1404 -2238
rect 1468 -2248 1502 -2238
rect 1558 -2230 1652 -2224
rect 1468 -2598 1504 -2248
rect 1404 -2600 1504 -2598
rect 1558 -2592 1658 -2230
rect 1698 -2234 1736 -1632
rect 1808 -1824 1880 -1682
rect 1772 -2024 1972 -1824
rect 1808 -2182 1880 -2024
rect 1698 -2238 1818 -2234
rect 1698 -2368 1716 -2238
rect 1558 -2600 1584 -2592
rect 1624 -2638 1658 -2592
rect 1702 -2598 1716 -2368
rect 1780 -2598 1818 -2238
rect 1702 -2608 1818 -2598
rect 1872 -2600 1974 -2224
rect 2018 -2228 2052 -1632
rect 2326 -1634 2448 -458
rect 2128 -1818 2196 -1684
rect 2094 -2018 2294 -1818
rect 2128 -2180 2196 -2018
rect 2018 -2236 2136 -2228
rect 2014 -2596 2024 -2236
rect 2088 -2596 2136 -2236
rect 2020 -2600 2136 -2596
rect 1872 -2602 1906 -2600
rect 1040 -2682 1240 -2680
rect 1296 -2682 1346 -2654
rect 1622 -2682 1658 -2638
rect 1940 -2648 1974 -2600
rect 2188 -2604 2290 -2228
rect 2328 -2230 2366 -1634
rect 2494 -1636 2582 -370
rect 2634 -1632 2768 -446
rect 2818 -1630 2906 -370
rect 2950 -1632 3078 -450
rect 2442 -1824 2514 -1684
rect 2404 -2024 2604 -1824
rect 2442 -2182 2514 -2024
rect 2636 -2222 2688 -1632
rect 2756 -1818 2824 -1684
rect 2728 -2018 2928 -1818
rect 2756 -2182 2824 -2018
rect 2328 -2232 2448 -2230
rect 2328 -2592 2342 -2232
rect 2406 -2592 2448 -2232
rect 2328 -2600 2448 -2592
rect 2504 -2600 2606 -2224
rect 1938 -2682 1974 -2648
rect 2256 -2682 2290 -2604
rect 2572 -2682 2606 -2600
rect 2636 -2238 2768 -2222
rect 2636 -2598 2654 -2238
rect 2718 -2598 2768 -2238
rect 2636 -2606 2768 -2598
rect 2822 -2602 2924 -2226
rect 2960 -2230 3012 -1632
rect 3136 -1634 3224 -370
rect 3270 -1628 3398 -450
rect 3452 -1624 3540 -370
rect 3270 -1632 3322 -1628
rect 3370 -1632 3398 -1628
rect 3272 -1674 3322 -1632
rect 3076 -1824 3142 -1684
rect 3042 -2024 3242 -1824
rect 3076 -2182 3142 -2024
rect 3272 -2094 3332 -1674
rect 3390 -1820 3462 -1684
rect 3374 -2020 3574 -1820
rect 3288 -2184 3332 -2094
rect 3390 -2182 3462 -2020
rect 2956 -2234 3082 -2230
rect 2956 -2594 2972 -2234
rect 3036 -2594 3082 -2234
rect 2956 -2600 3082 -2594
rect 2892 -2682 2924 -2602
rect 3134 -2604 3240 -2226
rect 3288 -2232 3324 -2184
rect 3366 -2232 3400 -2228
rect 3288 -2236 3400 -2232
rect 3288 -2262 3292 -2236
rect 3282 -2596 3292 -2262
rect 3348 -2596 3400 -2236
rect 3284 -2602 3400 -2596
rect 3452 -2596 3584 -2226
rect 3452 -2602 3476 -2596
rect 3206 -2682 3240 -2604
rect 3522 -2646 3584 -2596
rect 3518 -2654 3584 -2646
rect 3518 -2682 3616 -2654
rect 1040 -2688 3616 -2682
rect 1036 -2698 3616 -2688
rect 1036 -2878 1054 -2698
rect 3592 -2878 3616 -2698
rect 1036 -2886 3616 -2878
rect 1040 -2894 3616 -2886
rect 1148 -2978 1270 -2962
rect 1148 -3418 1164 -2978
rect 1240 -3418 1270 -2978
rect 1436 -3000 1568 -2936
rect 1148 -3430 1270 -3418
rect 1446 -3120 1464 -3000
rect 1446 -3414 1462 -3120
rect 1536 -3414 1568 -3000
rect 1446 -3424 1568 -3414
rect 1536 -3430 1568 -3424
rect 1740 -2984 1850 -2962
rect 1740 -3120 1760 -2984
rect 1824 -3120 1850 -2984
rect 1740 -3416 1756 -3120
rect 1830 -3416 1850 -3120
rect 1740 -3432 1850 -3416
rect 2042 -2980 2152 -2966
rect 2042 -3120 2058 -2980
rect 2122 -3120 2152 -2980
rect 2042 -3414 2054 -3120
rect 2128 -3414 2152 -3120
rect 2042 -3436 2152 -3414
rect 2334 -2984 2444 -2960
rect 2334 -3120 2356 -2984
rect 2420 -3120 2444 -2984
rect 2334 -3414 2350 -3120
rect 2424 -3414 2444 -3120
rect 2334 -3430 2444 -3414
rect 2630 -2984 2740 -2954
rect 2630 -3120 2654 -2984
rect 2718 -3120 2740 -2984
rect 2630 -3414 2646 -3120
rect 2720 -3414 2740 -3120
rect 2630 -3424 2740 -3414
rect 2920 -2984 3030 -2956
rect 2920 -3120 2950 -2984
rect 3014 -3120 3030 -2984
rect 2920 -3414 2944 -3120
rect 3018 -3414 3030 -3120
rect 2920 -3426 3030 -3414
rect 3220 -2984 3330 -2954
rect 3220 -3120 3242 -2984
rect 3306 -3120 3330 -2984
rect 3220 -3414 3240 -3120
rect 3314 -3414 3330 -3120
rect 3220 -3424 3330 -3414
rect 3504 -2982 3616 -2894
rect 3504 -3414 3618 -2982
rect 3504 -3416 3616 -3414
rect 1036 -3666 1114 -3664
rect 1036 -4098 1240 -3666
rect 1036 -4862 1114 -4098
rect 1332 -4146 1532 -3666
rect 1630 -4092 1830 -3662
rect 1282 -4192 1532 -4146
rect 1170 -4224 1532 -4192
rect 1584 -4220 1830 -4092
rect 1926 -4094 2126 -3664
rect 2218 -4094 2418 -3666
rect 1170 -4284 1426 -4224
rect 1170 -4660 1370 -4284
rect 1584 -4314 1720 -4220
rect 1882 -4222 2126 -4094
rect 1882 -4314 2018 -4222
rect 2180 -4224 2418 -4094
rect 2518 -4100 2718 -3662
rect 3106 -3666 3568 -3664
rect 2470 -4220 2718 -4100
rect 2820 -4102 3020 -3666
rect 3106 -4100 3602 -3666
rect 2180 -4314 2316 -4224
rect 2470 -4314 2606 -4220
rect 1460 -4408 1720 -4314
rect 1460 -4642 1668 -4408
rect 1762 -4410 2018 -4314
rect 2056 -4410 2316 -4314
rect 1762 -4642 1970 -4410
rect 2056 -4642 2264 -4410
rect 2354 -4416 2606 -4314
rect 2770 -4224 3020 -4102
rect 3072 -4222 3602 -4100
rect 2770 -4316 2906 -4224
rect 3072 -4314 3208 -4222
rect 3402 -4224 3602 -4222
rect 1170 -4750 1416 -4660
rect 1460 -4750 1726 -4642
rect 1762 -4750 2024 -4642
rect 2056 -4750 2322 -4642
rect 2354 -4644 2562 -4416
rect 2650 -4418 2906 -4316
rect 2946 -4416 3208 -4314
rect 2650 -4644 2858 -4418
rect 2354 -4750 2608 -4644
rect 1280 -4862 1416 -4750
rect 1590 -4860 1726 -4750
rect 1888 -4858 2024 -4750
rect 2186 -4858 2322 -4750
rect 2472 -4858 2608 -4750
rect 2650 -4752 2910 -4644
rect 2946 -4750 3154 -4416
rect 2774 -4858 2910 -4752
rect 1036 -5292 1240 -4862
rect 1280 -4976 1542 -4862
rect 1590 -4958 1832 -4860
rect 1888 -4958 2134 -4858
rect 2186 -4958 2428 -4858
rect 1334 -5294 1542 -4976
rect 1624 -5296 1832 -4958
rect 1926 -5294 2134 -4958
rect 2220 -5294 2428 -4958
rect 2472 -4960 2726 -4858
rect 2774 -4960 3020 -4858
rect 2518 -5294 2726 -4960
rect 2812 -5294 3020 -4960
<< via1 >>
rect 1070 -2596 1134 -2236
rect 1404 -2598 1468 -2238
rect 1716 -2598 1780 -2238
rect 2024 -2596 2088 -2236
rect 2342 -2592 2406 -2232
rect 2654 -2598 2718 -2238
rect 2972 -2594 3036 -2234
rect 3292 -2596 3348 -2236
rect 1164 -3418 1240 -2978
rect 1464 -3120 1536 -3000
rect 1462 -3414 1536 -3120
rect 1760 -3120 1824 -2984
rect 1756 -3416 1830 -3120
rect 2058 -3120 2122 -2980
rect 2054 -3414 2128 -3120
rect 2356 -3120 2420 -2984
rect 2350 -3414 2424 -3120
rect 2654 -3120 2718 -2984
rect 2646 -3414 2720 -3120
rect 2950 -3120 3014 -2984
rect 2944 -3414 3018 -3120
rect 3242 -3120 3306 -2984
rect 3240 -3414 3314 -3120
<< metal2 >>
rect 1070 -2236 1134 -2226
rect 1068 -2596 1070 -2400
rect 1404 -2238 1468 -2228
rect 1068 -2606 1134 -2596
rect 1400 -2598 1404 -2404
rect 1068 -2958 1130 -2606
rect 1400 -2608 1468 -2598
rect 1716 -2238 1780 -2228
rect 2024 -2236 2088 -2226
rect 1716 -2608 1780 -2598
rect 2020 -2596 2024 -2406
rect 2342 -2232 2406 -2222
rect 2020 -2606 2088 -2596
rect 2334 -2592 2342 -2444
rect 2654 -2238 2718 -2228
rect 2406 -2592 2408 -2444
rect 1400 -2936 1462 -2608
rect 1068 -2990 1112 -2958
rect 1162 -2978 1270 -2962
rect 1162 -2990 1164 -2978
rect 1068 -3408 1164 -2990
rect 1076 -3412 1164 -3408
rect 1148 -3418 1164 -3412
rect 1240 -3418 1270 -2978
rect 1400 -3000 1562 -2936
rect 1716 -2962 1778 -2608
rect 1716 -2984 1850 -2962
rect 1400 -3120 1464 -3000
rect 1400 -3412 1462 -3120
rect 1456 -3414 1462 -3412
rect 1536 -3414 1546 -3000
rect 1456 -3418 1546 -3414
rect 1716 -3120 1760 -2984
rect 1824 -3120 1850 -2984
rect 1716 -3416 1756 -3120
rect 1830 -3416 1850 -3120
rect 2020 -2966 2082 -2606
rect 2334 -2960 2408 -2592
rect 2650 -2598 2654 -2446
rect 2972 -2234 3036 -2224
rect 2718 -2598 2724 -2446
rect 2650 -2954 2724 -2598
rect 3292 -2236 3348 -2226
rect 3036 -2594 3042 -2438
rect 2020 -2980 2152 -2966
rect 2020 -3120 2058 -2980
rect 2122 -3120 2152 -2980
rect 2020 -3414 2054 -3120
rect 2128 -3414 2152 -3120
rect 1148 -3430 1270 -3418
rect 1462 -3424 1536 -3418
rect 1716 -3420 1850 -3416
rect 1740 -3432 1850 -3420
rect 2042 -3436 2152 -3414
rect 2334 -2984 2444 -2960
rect 2334 -3120 2356 -2984
rect 2420 -3120 2444 -2984
rect 2334 -3414 2350 -3120
rect 2424 -3414 2444 -3120
rect 2334 -3430 2444 -3414
rect 2630 -2984 2740 -2954
rect 2972 -2956 3042 -2594
rect 3288 -2596 3292 -2376
rect 3288 -2954 3348 -2596
rect 2630 -3120 2654 -2984
rect 2718 -3120 2740 -2984
rect 2630 -3414 2646 -3120
rect 2720 -3414 2740 -3120
rect 2630 -3424 2740 -3414
rect 2920 -2984 3042 -2956
rect 2920 -3120 2950 -2984
rect 3014 -3120 3042 -2984
rect 2920 -3414 2944 -3120
rect 3018 -3406 3042 -3120
rect 3220 -2984 3348 -2954
rect 3220 -3120 3242 -2984
rect 3306 -3120 3348 -2984
rect 3018 -3414 3030 -3406
rect 2920 -3426 3030 -3414
rect 3220 -3414 3240 -3120
rect 3314 -3412 3348 -3120
rect 3314 -3414 3330 -3412
rect 3220 -3424 3330 -3414
<< rmetal2 >>
rect 1112 -2990 1162 -2958
use sky130_fd_pr__nfet_01v8_ATMSL9  sky130_fd_pr__nfet_01v8_ATMSL9_0
timestamp 1730493024
transform 1 0 3109 0 1 -2383
box -211 -379 211 379
use sky130_fd_pr__pfet_01v8_LGA5KQ  sky130_fd_pr__pfet_01v8_LGA5KQ_0
timestamp 1730493024
transform 1 0 1211 0 1 -1078
box -211 -784 211 784
use sky130_fd_pr__nfet_01v8_ATMSL9  XM1
timestamp 1730493024
transform 1 0 1213 0 1 -2383
box -211 -379 211 379
use sky130_fd_pr__nfet_01v8_ATMSL9  XM3
timestamp 1730493024
transform 1 0 1529 0 1 -2383
box -211 -379 211 379
use sky130_fd_pr__pfet_01v8_MGA5KJ  XM4
timestamp 1730493024
transform -1 0 1527 0 -1 -1078
box -211 -784 211 784
use sky130_fd_pr__nfet_01v8_ATMSL9  XM5
timestamp 1730493024
transform 1 0 1845 0 1 -2383
box -211 -379 211 379
use sky130_fd_pr__pfet_01v8_LGA5KQ  XM6
timestamp 1730493024
transform 1 0 1843 0 1 -1078
box -211 -784 211 784
use sky130_fd_pr__nfet_01v8_ATMSL9  XM7
timestamp 1730493024
transform 1 0 2161 0 1 -2383
box -211 -379 211 379
use sky130_fd_pr__pfet_01v8_LGA5KQ  XM8
timestamp 1730493024
transform 1 0 2159 0 1 -1078
box -211 -784 211 784
use sky130_fd_pr__nfet_01v8_ATMSL9  XM9
timestamp 1730493024
transform 1 0 2477 0 1 -2383
box -211 -379 211 379
use sky130_fd_pr__pfet_01v8_LGA5KQ  XM10
timestamp 1730493024
transform 1 0 2475 0 1 -1078
box -211 -784 211 784
use sky130_fd_pr__nfet_01v8_ATMSL9  XM11
timestamp 1730493024
transform 1 0 2793 0 1 -2383
box -211 -379 211 379
use sky130_fd_pr__pfet_01v8_LGA5KQ  XM12
timestamp 1730493024
transform 1 0 2791 0 1 -1078
box -211 -784 211 784
use sky130_fd_pr__pfet_01v8_LGA5KQ  XM14
timestamp 1730493024
transform 1 0 3107 0 1 -1078
box -211 -784 211 784
use sky130_fd_pr__nfet_01v8_ATMSL9  XM15
timestamp 1730493024
transform 1 0 3425 0 1 -2383
box -211 -379 211 379
use sky130_fd_pr__pfet_01v8_LGA5KQ  XM16
timestamp 1730493024
transform 1 0 3423 0 1 -1078
box -211 -784 211 784
use sky130_fd_pr__res_xhigh_po_0p35_ABVTW2  XR1
timestamp 1730493024
transform 1 0 1499 0 1 -3538
box -201 -722 201 722
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR2
timestamp 1730493024
transform 1 0 1203 0 1 -4806
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_ABVTW2  XR3
timestamp 1730493024
transform 1 0 1203 0 1 -3538
box -201 -722 201 722
use sky130_fd_pr__res_xhigh_po_0p35_ABVTW2  XR5
timestamp 1730493024
transform 1 0 3571 0 1 -3538
box -201 -722 201 722
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR6
timestamp 1730493024
transform 1 0 1499 0 1 -4806
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_ABVTW2  XR7
timestamp 1730493024
transform 1 0 1795 0 1 -3538
box -201 -722 201 722
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR8
timestamp 1730493024
transform 1 0 1795 0 1 -4806
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_ABVTW2  XR9
timestamp 1730493024
transform 1 0 2091 0 1 -3538
box -201 -722 201 722
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR10
timestamp 1730493024
transform 1 0 2091 0 1 -4806
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_ABVTW2  XR11
timestamp 1730493024
transform 1 0 2387 0 1 -3538
box -201 -722 201 722
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR12
timestamp 1730493024
transform 1 0 2387 0 1 -4806
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_ABVTW2  XR13
timestamp 1730493024
transform 1 0 2683 0 1 -3538
box -201 -722 201 722
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR14
timestamp 1730493024
transform 1 0 2683 0 1 -4806
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_ABVTW2  XR15
timestamp 1730493024
transform 1 0 2979 0 1 -3538
box -201 -722 201 722
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR16
timestamp 1730493024
transform 1 0 2979 0 1 -4806
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_ABVTW2  XR17
timestamp 1730493024
transform -1 0 3275 0 1 -3538
box -201 -722 201 722
<< labels >>
flabel metal1 3374 -2034 3574 -1834 0 FreeSans 256 0 0 0 b0
port 2 nsew
flabel metal1 3042 -2024 3242 -1824 0 FreeSans 256 0 0 0 b1
port 3 nsew
flabel metal1 2728 -2024 2928 -1824 0 FreeSans 256 0 0 0 b2
port 4 nsew
flabel metal1 2404 -2018 2604 -1818 0 FreeSans 256 0 0 0 b3
port 5 nsew
flabel metal1 2094 -2024 2294 -1824 0 FreeSans 256 0 0 0 b4
port 6 nsew
flabel metal1 1772 -2018 1972 -1818 0 FreeSans 256 0 0 0 b5
port 7 nsew
flabel metal1 1470 -2024 1670 -1824 0 FreeSans 256 0 0 0 b6
port 8 nsew
flabel metal1 1170 -2020 1370 -1820 0 FreeSans 256 0 0 0 b7
port 9 nsew
flabel metal1 1586 -392 1786 -192 0 FreeSans 256 0 0 0 vdd
port 1 nsew
flabel metal1 1040 -2880 1240 -2680 0 FreeSans 256 0 0 0 vss
port 10 nsew
flabel metal1 1040 -4080 1240 -3880 0 FreeSans 256 0 0 0 out
port 0 nsew
<< end >>
