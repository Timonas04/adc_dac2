magic
tech sky130A
magscale 1 2
timestamp 1730901241
<< pwell >>
rect 30680 18340 31040 18740
rect 28020 17760 28380 18160
<< locali >>
rect 25210 17291 25389 17652
<< metal1 >>
rect 25360 18420 25720 18720
rect 25360 18360 25480 18420
rect 25560 18360 25720 18420
rect 25360 18320 25720 18360
rect 25940 18420 26300 18720
rect 25940 18360 26080 18420
rect 26140 18360 26300 18420
rect 25940 18320 26300 18360
rect 26540 18420 26900 18720
rect 26540 18360 26680 18420
rect 26740 18360 26900 18420
rect 26540 18320 26900 18360
rect 27140 18400 27500 18720
rect 27140 18340 27260 18400
rect 27320 18340 27500 18400
rect 27140 18320 27500 18340
rect 27720 18400 28080 18720
rect 27720 18340 27860 18400
rect 27920 18340 28080 18400
rect 27720 18320 28080 18340
rect 28320 18400 28680 18720
rect 28320 18340 28460 18400
rect 28520 18340 28680 18400
rect 28320 18320 28680 18340
rect 28900 18400 29260 18720
rect 28900 18340 29060 18400
rect 29120 18340 29260 18400
rect 28900 18320 29260 18340
rect 29500 18400 29860 18720
rect 29500 18340 29640 18400
rect 29700 18340 29860 18400
rect 29500 18320 29860 18340
rect 30080 18320 30440 18720
rect 30680 18340 31040 18740
rect 31280 18320 31640 18720
rect 25207 17285 25402 18190
rect 25640 17880 26000 18160
rect 25640 17820 25780 17880
rect 25840 17820 26000 17880
rect 25640 17760 26000 17820
rect 26240 17840 26600 18160
rect 26240 17780 26380 17840
rect 26440 17780 26600 17840
rect 26840 17880 27200 18180
rect 26840 17820 26980 17880
rect 27040 17820 27200 17880
rect 26840 17780 27200 17820
rect 27420 17860 27780 18160
rect 27420 17800 27560 17860
rect 27620 17800 27780 17860
rect 26240 17760 26600 17780
rect 27420 17760 27780 17800
rect 28020 17840 28380 18160
rect 28020 17780 28160 17840
rect 28220 17780 28380 17840
rect 28600 17860 28960 18180
rect 28600 17800 28760 17860
rect 28820 17800 28960 17860
rect 28600 17780 28960 17800
rect 29200 17860 29560 18180
rect 29200 17800 29340 17860
rect 29400 17800 29560 17860
rect 29200 17780 29560 17800
rect 28020 17760 28380 17780
rect 29800 17760 30160 18160
rect 30380 17760 30740 18160
rect 30980 17760 31340 18160
rect 31580 17360 31720 18180
rect 9216 11996 9222 12048
rect 9274 12047 9280 12048
rect 15958 12047 16008 12125
rect 9274 11997 16008 12047
rect 9274 11996 9280 11997
rect 12019 11888 12071 11894
rect 12143 11879 12149 11931
rect 12201 11925 12207 11931
rect 19363 11925 19404 12121
rect 12201 11884 19404 11925
rect 12201 11879 12207 11884
rect 22769 11847 22798 12115
rect 12071 11836 22798 11847
rect 12019 11830 22798 11836
rect 12030 11818 22798 11830
rect 11866 11734 11872 11786
rect 11924 11780 11930 11786
rect 26163 11780 26203 12120
rect 11924 11740 26203 11780
rect 11924 11734 11930 11740
rect 11733 11661 11739 11713
rect 11791 11706 11797 11713
rect 29564 11706 29603 12120
rect 11791 11667 29603 11706
rect 11791 11661 11797 11667
rect 12521 6238 12573 6244
rect 12658 6224 12664 6276
rect 12716 6268 12722 6276
rect 15965 6268 16001 6318
rect 12716 6232 16001 6268
rect 12716 6224 12722 6232
rect 12573 6186 12576 6208
rect 12521 6180 12576 6186
rect 12530 6171 12576 6180
rect 19367 6171 19400 6317
rect 12530 6138 19400 6171
rect 12390 6064 12396 6116
rect 12448 6113 12454 6116
rect 22760 6113 22806 6323
rect 12448 6110 12498 6113
rect 19618 6110 22806 6113
rect 12448 6067 22806 6110
rect 12448 6064 12454 6067
rect 12211 5967 12217 6019
rect 12269 6017 12275 6019
rect 26159 6017 26208 6325
rect 12269 5968 26208 6017
rect 12269 5967 12275 5968
rect 12054 5878 12060 5930
rect 12112 5927 12118 5930
rect 29560 5927 29606 6323
rect 12112 5881 29606 5927
rect 12112 5878 12118 5881
rect 12170 390 12176 442
rect 12228 438 12234 442
rect 15961 438 16005 522
rect 12228 394 16005 438
rect 12228 390 12234 394
rect 11791 379 11843 385
rect 11217 360 11269 366
rect 12049 354 12125 387
rect 11791 321 11843 327
rect 12045 348 12125 354
rect 11217 302 11269 308
rect 11224 102 11262 302
rect 11800 175 11834 321
rect 12097 327 12125 348
rect 19363 327 19404 521
rect 12097 296 19404 327
rect 11915 289 11967 295
rect 12045 290 19404 296
rect 12049 286 19404 290
rect 22765 243 22802 519
rect 11967 237 22802 243
rect 11915 231 22802 237
rect 11922 206 22802 231
rect 26166 175 26200 517
rect 11800 141 26200 175
rect 29564 102 29602 519
rect 11224 64 29602 102
<< via1 >>
rect 25480 18360 25560 18420
rect 26080 18360 26140 18420
rect 26680 18360 26740 18420
rect 27260 18340 27320 18400
rect 27860 18340 27920 18400
rect 28460 18340 28520 18400
rect 29060 18340 29120 18400
rect 29640 18340 29700 18400
rect 25780 17820 25840 17880
rect 26380 17780 26440 17840
rect 26980 17820 27040 17880
rect 27560 17800 27620 17860
rect 28160 17780 28220 17840
rect 28760 17800 28820 17860
rect 29340 17800 29400 17860
rect 9222 11996 9274 12048
rect 12019 11836 12071 11888
rect 12149 11879 12201 11931
rect 11872 11734 11924 11786
rect 11739 11661 11791 11713
rect 12521 6186 12573 6238
rect 12664 6224 12716 6276
rect 12396 6064 12448 6116
rect 12217 5967 12269 6019
rect 12060 5878 12112 5930
rect 12176 390 12228 442
rect 11217 308 11269 360
rect 11791 327 11843 379
rect 12045 296 12097 348
rect 11915 237 11967 289
<< metal2 >>
rect 25460 18420 25580 18440
rect 25460 18360 25480 18420
rect 25560 18360 25580 18420
rect 25460 18340 25580 18360
rect 26060 18420 26160 18440
rect 26060 18360 26080 18420
rect 26140 18360 26160 18420
rect 26060 18340 26160 18360
rect 26660 18420 26760 18440
rect 26660 18360 26680 18420
rect 26740 18360 26760 18420
rect 26660 18340 26760 18360
rect 27240 18400 27340 18420
rect 27240 18340 27260 18400
rect 27320 18340 27340 18400
rect 27240 18320 27340 18340
rect 27840 18400 27940 18420
rect 27840 18340 27860 18400
rect 27920 18340 27940 18400
rect 27840 18320 27940 18340
rect 28440 18400 28540 18420
rect 28440 18340 28460 18400
rect 28520 18340 28540 18400
rect 28440 18320 28540 18340
rect 29040 18400 29140 18420
rect 29040 18340 29060 18400
rect 29120 18340 29140 18400
rect 29040 18320 29140 18340
rect 29620 18400 29720 18420
rect 29620 18340 29640 18400
rect 29700 18340 29720 18400
rect 29620 18320 29720 18340
rect 25760 17880 25860 17900
rect 25760 17820 25780 17880
rect 25840 17820 25860 17880
rect 26960 17880 27060 17900
rect 25760 17800 25860 17820
rect 26360 17840 26460 17860
rect 26360 17780 26380 17840
rect 26440 17780 26460 17840
rect 26960 17820 26980 17880
rect 27040 17820 27060 17880
rect 26960 17800 27060 17820
rect 27540 17860 27640 17880
rect 28740 17860 28840 17880
rect 27540 17800 27560 17860
rect 27620 17800 27640 17860
rect 27540 17780 27640 17800
rect 28140 17840 28240 17860
rect 28140 17780 28160 17840
rect 28220 17780 28240 17840
rect 28740 17800 28760 17860
rect 28820 17800 28840 17860
rect 28740 17780 28840 17800
rect 29320 17860 29420 17880
rect 29320 17800 29340 17860
rect 29400 17800 29420 17860
rect 29320 17780 29420 17800
rect 26360 17760 26460 17780
rect 28140 17760 28240 17780
rect 12146 12220 12206 12229
rect 12146 12151 12206 12160
rect 9222 12048 9274 12054
rect 9222 11990 9274 11996
rect 11345 11918 11785 11957
rect 12155 11937 12196 12151
rect 11746 11719 11785 11918
rect 12149 11931 12201 11937
rect 12013 11836 12019 11888
rect 12071 11836 12077 11888
rect 12149 11873 12201 11879
rect 11872 11786 11924 11792
rect 11872 11728 11924 11734
rect 11739 11713 11791 11719
rect 11739 11655 11791 11661
rect 11878 11543 11918 11728
rect 11868 11534 11928 11543
rect 11868 11465 11928 11474
rect 12031 10182 12060 11836
rect 12660 10858 12720 10867
rect 12660 10789 12720 10798
rect 12016 10173 12076 10182
rect 12016 10104 12076 10113
rect 12518 9494 12578 9503
rect 12518 9425 12578 9434
rect 12392 8820 12452 8829
rect 12392 8751 12452 8760
rect 12214 8138 12274 8147
rect 12214 8069 12274 8078
rect 12056 7462 12116 7471
rect 12056 7393 12116 7402
rect 11912 6777 11972 6786
rect 11912 6708 11972 6717
rect 11787 6098 11847 6107
rect 11787 6029 11847 6038
rect 11224 360 11262 4201
rect 11800 379 11834 6029
rect 11211 308 11217 360
rect 11269 308 11275 360
rect 11785 327 11791 379
rect 11843 327 11849 379
rect 11923 289 11960 6708
rect 12063 5936 12109 7393
rect 12219 6025 12268 8069
rect 12399 6122 12445 8751
rect 12531 6238 12564 9425
rect 12672 6282 12708 10789
rect 12664 6276 12716 6282
rect 12515 6186 12521 6238
rect 12573 6186 12579 6238
rect 12664 6218 12716 6224
rect 12396 6116 12448 6122
rect 12396 6058 12448 6064
rect 12217 6019 12269 6025
rect 12217 5961 12269 5967
rect 12060 5930 12112 5936
rect 12060 5872 12112 5878
rect 12042 5419 12102 5428
rect 12042 5350 12102 5359
rect 12051 348 12092 5350
rect 12172 4737 12232 4746
rect 12172 4668 12232 4677
rect 12180 448 12224 4668
rect 12176 442 12228 448
rect 12176 384 12228 390
rect 12039 296 12045 348
rect 12097 296 12103 348
rect 11909 237 11915 289
rect 11967 237 11973 289
<< via2 >>
rect 12146 12160 12206 12220
rect 11868 11474 11928 11534
rect 12660 10798 12720 10858
rect 12016 10113 12076 10173
rect 12518 9434 12578 9494
rect 12392 8760 12452 8820
rect 12214 8078 12274 8138
rect 12056 7402 12116 7462
rect 11912 6717 11972 6777
rect 11787 6038 11847 6098
rect 12042 5359 12102 5419
rect 12172 4677 12232 4737
<< metal3 >>
rect 12141 12220 12211 12225
rect 12141 12160 12146 12220
rect 12206 12160 12211 12220
rect 12141 12155 12211 12160
rect 11863 11534 11933 11539
rect 11863 11474 11868 11534
rect 11928 11474 11933 11534
rect 11863 11469 11933 11474
rect 12655 10858 12725 10863
rect 12655 10798 12660 10858
rect 12720 10798 12725 10858
rect 12655 10793 12725 10798
rect 12011 10173 12081 10178
rect 12011 10113 12016 10173
rect 12076 10113 12081 10173
rect 12011 10108 12081 10113
rect 12513 9494 12583 9499
rect 12513 9434 12518 9494
rect 12578 9434 12583 9494
rect 12513 9429 12583 9434
rect 12387 8820 12457 8825
rect 12387 8760 12392 8820
rect 12452 8760 12457 8820
rect 12387 8755 12457 8760
rect 12209 8138 12279 8143
rect 12209 8078 12214 8138
rect 12274 8078 12279 8138
rect 12209 8073 12279 8078
rect 12051 7462 12121 7467
rect 12051 7402 12056 7462
rect 12116 7402 12121 7462
rect 12051 7397 12121 7402
rect 11879 6777 12054 6811
rect 11879 6717 11912 6777
rect 11972 6717 12054 6777
rect 11879 6683 12039 6717
rect 11782 6098 11852 6103
rect 11782 6038 11787 6098
rect 11847 6038 11852 6098
rect 11782 6033 11852 6038
rect 12037 5419 12107 5424
rect 12037 5359 12042 5419
rect 12102 5359 12107 5419
rect 12037 5354 12107 5359
rect 12167 4737 12237 4742
rect 12167 4677 12172 4737
rect 12232 4677 12237 4737
rect 12167 4672 12237 4677
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 45077 12818 45152
rect 12758 45011 12829 45077
rect 13310 45059 13370 45152
rect 13862 45093 13922 45152
rect 12758 44952 12818 45011
rect 13291 44993 13370 45059
rect 13861 45027 13927 45093
rect 14414 45045 14474 45152
rect 14966 45055 15026 45152
rect 13310 44952 13370 44993
rect 13862 44952 13922 45027
rect 14399 44979 14474 45045
rect 14957 44989 15026 45055
rect 15518 45017 15578 45152
rect 16070 45051 16130 45152
rect 14414 44952 14474 44979
rect 14966 44952 15026 44989
rect 15503 44952 15578 45017
rect 16059 44985 16130 45051
rect 16622 45017 16682 45152
rect 17174 45049 17234 45152
rect 17726 45049 17786 45152
rect 16070 44952 16130 44985
rect 16605 44952 16682 45017
rect 17159 44983 17234 45049
rect 17707 44983 17786 45049
rect 18278 45033 18338 45152
rect 17174 44952 17234 44983
rect 17726 44952 17786 44983
rect 18270 44967 18338 45033
rect 18830 45029 18890 45152
rect 18278 44952 18338 44967
rect 18825 44963 18891 45029
rect 18830 44952 18890 44963
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 15503 44951 15569 44952
rect 16605 44951 16671 44952
rect 200 1000 600 44152
rect 800 39832 1200 44152
rect 800 39512 1228 39832
rect 800 1000 1200 39512
rect 3314 0 3494 204
rect 7178 0 7358 204
rect 11042 0 11222 204
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use bit4_encoder  bit4_encoder_0 ~/Documents/github_project/adc_dac2/mag
timestamp 1730889744
transform 1 0 3400 0 1 2600
box 0 0 9409 11553
use compr2  compr2_0
timestamp 1730896912
transform 0 1 30003 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_1
timestamp 1730896912
transform 0 1 26603 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_2
timestamp 1730896912
transform 0 1 23203 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_3
timestamp 1730896912
transform 0 1 19803 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_4
timestamp 1730896912
transform 0 1 16403 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_5
timestamp 1730896912
transform 0 1 30003 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_6
timestamp 1730896912
transform 0 1 26603 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_7
timestamp 1730896912
transform 0 1 23203 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_8
timestamp 1730896912
transform 0 1 19803 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_9
timestamp 1730896912
transform 0 1 16403 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_10
timestamp 1730896912
transform 0 1 30003 -1 0 17975
box 510 -1403 5975 1713
use compr2  compr2_11
timestamp 1730896912
transform 0 1 26603 -1 0 17975
box 510 -1403 5975 1713
use compr2  compr2_12
timestamp 1730896912
transform 0 1 23203 -1 0 17975
box 510 -1403 5975 1713
use compr2  compr2_13
timestamp 1730896912
transform 0 1 19803 -1 0 17975
box 510 -1403 5975 1713
use compr2  compr2_14
timestamp 1730896912
transform 0 1 16403 -1 0 17975
box 510 -1403 5975 1713
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR1
timestamp 1730882523
transform 1 0 28049 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR2
timestamp 1730882523
transform 1 0 26273 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR3
timestamp 1730882523
transform 1 0 26865 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR4
timestamp 1730882523
transform 1 0 27753 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR5
timestamp 1730882523
transform 1 0 27457 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR6
timestamp 1730882523
transform 1 0 30417 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR7
timestamp 1730882523
transform 1 0 27161 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR8
timestamp 1730882523
transform 1 0 29529 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR9
timestamp 1730882523
transform 1 0 28345 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR10
timestamp 1730882523
transform 1 0 29233 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR11
timestamp 1730882523
transform 1 0 28641 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR12
timestamp 1730882523
transform 1 0 28937 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR13
timestamp 1730882523
transform 1 0 29825 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR14
timestamp 1730882523
transform 1 0 26569 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR15
timestamp 1730882523
transform 1 0 25977 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR16
timestamp 1730882523
transform 1 0 30121 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR17
timestamp 1730882523
transform 1 0 30713 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR18
timestamp 1730882523
transform 1 0 31305 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR19
timestamp 1730882523
transform 1 0 31009 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR20
timestamp 1730882523
transform 1 0 31601 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR21
timestamp 1730882523
transform 1 0 25681 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR22
timestamp 1730882523
transform 1 0 25385 0 1 18252
box -201 -652 201 652
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
