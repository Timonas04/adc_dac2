magic
tech sky130A
magscale 1 2
timestamp 1730847319
<< locali >>
rect 24000 20548 24192 21250
rect 24000 20494 26910 20548
rect 24000 20384 24044 20494
rect 26474 20384 26910 20494
rect 24000 20344 26910 20384
rect 27186 20344 27214 20548
rect 24000 20330 24192 20344
<< viali >>
rect 24044 20384 26474 20494
<< metal1 >>
rect 29942 44424 29994 44430
rect 29942 44366 29994 44372
rect 29830 44212 29882 44218
rect 29830 44154 29882 44160
rect 29726 44010 29732 44062
rect 29784 44010 29790 44062
rect 29628 43972 29680 43978
rect 29628 43914 29680 43920
rect 22190 41320 22242 41326
rect 22190 41262 22242 41268
rect 21990 41230 22042 41236
rect 21990 41172 22042 41178
rect 22002 38509 22030 41172
rect 22202 40306 22230 41262
rect 22272 41224 22324 41230
rect 22272 41166 22324 41172
rect 22284 40527 22312 41166
rect 22266 40475 22272 40527
rect 22324 40475 22330 40527
rect 22202 40278 22328 40306
rect 22300 39706 22328 40278
rect 29640 40258 29668 43914
rect 29622 40251 29688 40258
rect 29622 40199 29628 40251
rect 29680 40199 29688 40251
rect 29622 40192 29688 40199
rect 29744 39791 29772 44010
rect 29726 39739 29732 39791
rect 29784 39739 29790 39791
rect 22282 39699 22348 39706
rect 22282 39647 22288 39699
rect 22340 39647 22348 39699
rect 22282 39640 22348 39647
rect 29842 39612 29870 44154
rect 29954 41086 29982 44366
rect 29936 41079 30000 41086
rect 29936 41027 29942 41079
rect 29994 41027 30000 41079
rect 29936 41020 30000 41027
rect 29734 39584 29870 39612
rect 29734 38510 29762 39584
rect 21990 38503 22042 38509
rect 21990 38445 22042 38451
rect 29714 38503 29780 38510
rect 29714 38451 29722 38503
rect 29774 38451 29780 38503
rect 29714 38444 29780 38451
rect 20194 36807 20526 36814
rect 20194 36489 20201 36807
rect 20519 36489 20526 36807
rect 20194 36482 20526 36489
rect 20201 35624 20519 36482
rect 20020 35620 28074 35624
rect 20020 35616 28172 35620
rect 19998 35410 28172 35616
rect 19998 35052 20154 35410
rect 23596 35296 23776 35328
rect 23596 34946 23624 35296
rect 23754 34946 23776 35296
rect 24006 35052 24162 35410
rect 27560 35294 27740 35324
rect 23596 34924 23776 34946
rect 27560 34944 27592 35294
rect 27722 34944 27740 35294
rect 28016 35056 28172 35410
rect 31514 35294 31694 35320
rect 27560 34920 27740 34944
rect 31514 34944 31540 35294
rect 31670 34944 31694 35294
rect 31514 34916 31694 34944
rect 23257 34552 23309 34558
rect 23257 34494 23309 34500
rect 27298 34538 27350 34544
rect 27298 34480 27350 34486
rect 31289 34542 31341 34548
rect 31289 34484 31341 34490
rect 20002 21320 20156 33448
rect 20552 33120 20558 33180
rect 20618 33120 20624 33180
rect 23238 31550 23290 31556
rect 23238 31492 23290 31498
rect 20544 30168 20604 30174
rect 20544 30102 20604 30108
rect 23286 28538 23338 28544
rect 23248 28486 23286 28534
rect 23248 28480 23338 28486
rect 23248 28470 23300 28480
rect 20560 27152 20620 27158
rect 20560 27086 20620 27092
rect 23236 25542 23288 25544
rect 23236 25536 23316 25542
rect 23236 25484 23264 25536
rect 23236 25480 23316 25484
rect 23264 25478 23316 25480
rect 20568 24152 20628 24158
rect 20568 24086 20628 24092
rect 23264 22544 23360 22550
rect 23264 22492 23308 22544
rect 23264 22486 23360 22492
rect 20550 21164 20610 21170
rect 20550 21098 20610 21104
rect 21243 20694 21493 20955
rect 23540 20808 23712 33188
rect 24000 21326 24154 33454
rect 24586 33200 24646 33206
rect 24586 33134 24646 33140
rect 27260 31544 27312 31550
rect 27260 31486 27312 31492
rect 24530 30164 24590 30170
rect 24530 30098 24590 30104
rect 27236 28550 27288 28556
rect 27236 28492 27288 28498
rect 24530 27142 24590 27148
rect 24530 27076 24590 27082
rect 27273 25552 27325 25558
rect 27273 25494 27325 25500
rect 24536 24180 24596 24186
rect 24536 24114 24596 24120
rect 27238 22550 27290 22556
rect 27238 22492 27290 22498
rect 21239 20595 21493 20694
rect 21239 20088 21491 20595
rect 23980 20552 24198 21176
rect 24542 21148 24602 21154
rect 24542 21082 24602 21088
rect 27520 20808 27692 33188
rect 27986 21326 28140 33454
rect 28598 33204 28658 33210
rect 28598 33138 28658 33144
rect 31306 31540 31358 31546
rect 31306 31482 31358 31488
rect 28528 30146 28588 30152
rect 28528 30080 28588 30086
rect 31260 28484 31266 28536
rect 31318 28484 31324 28536
rect 28536 27170 28596 27176
rect 28536 27104 28596 27110
rect 31288 25544 31340 25550
rect 31288 25486 31340 25492
rect 28532 24166 28592 24172
rect 28532 24100 28592 24106
rect 31206 22554 31258 22560
rect 31206 22496 31258 22502
rect 28538 21164 28598 21170
rect 28538 21098 28598 21104
rect 31528 20970 31700 33192
rect 31454 20812 31700 20970
rect 22608 20539 23346 20542
rect 23980 20539 27090 20552
rect 22608 20494 27090 20539
rect 22608 20384 24044 20494
rect 26474 20384 27090 20494
rect 22608 20342 27090 20384
rect 27326 20384 27690 20412
rect 22608 20338 26474 20342
rect 22608 20335 24672 20338
rect 22608 20332 23346 20335
rect 21054 18591 21254 18597
rect 21688 18591 21888 18597
rect 20430 18585 20630 18591
rect 20130 18575 20330 18581
rect 20130 18517 20330 18523
rect 20430 18519 20630 18525
rect 20732 18585 20932 18591
rect 21054 18532 21254 18538
rect 21364 18585 21564 18591
rect 20732 18522 20932 18528
rect 21688 18533 21888 18539
rect 22002 18585 22202 18591
rect 21364 18525 21564 18531
rect 22002 18527 22202 18533
rect 22334 18589 22534 18595
rect 22334 18531 22534 18537
rect 22614 17710 22740 20332
rect 23980 20330 24198 20335
rect 26896 19990 27086 20342
rect 27326 20318 27458 20384
rect 27534 20318 27690 20384
rect 27326 19992 27690 20318
rect 27914 20384 28278 20412
rect 27914 20318 28052 20384
rect 28128 20318 28278 20384
rect 27914 19992 28278 20318
rect 28494 20392 28860 20418
rect 28494 20326 28648 20392
rect 28714 20326 28860 20392
rect 28494 19992 28860 20326
rect 29088 20398 29454 20418
rect 29088 20332 29232 20398
rect 29298 20332 29454 20398
rect 29088 19992 29454 20332
rect 29684 20372 30050 20420
rect 29684 20306 29836 20372
rect 29902 20306 30050 20372
rect 29684 19994 30050 20306
rect 30274 20396 30640 20418
rect 30274 20330 30428 20396
rect 30494 20330 30640 20396
rect 30274 19992 30640 20330
rect 30868 20398 31234 20416
rect 30868 20332 31026 20398
rect 31092 20332 31234 20398
rect 30868 19990 31234 20332
rect 31454 19996 31692 20812
rect 27020 19860 27382 19868
rect 27618 19866 27982 19874
rect 27020 19832 27388 19860
rect 27020 19758 27164 19832
rect 27240 19758 27388 19832
rect 27020 19454 27388 19758
rect 27618 19800 27764 19866
rect 27840 19800 27982 19866
rect 27618 19454 27982 19800
rect 28206 19850 28570 19876
rect 28206 19784 28350 19850
rect 28426 19784 28570 19850
rect 28206 19456 28570 19784
rect 28792 19852 29158 19872
rect 28792 19786 28942 19852
rect 29008 19786 29158 19852
rect 27020 19448 27382 19454
rect 28792 19446 29158 19786
rect 29388 19856 29754 19874
rect 29388 19790 29546 19856
rect 29612 19790 29754 19856
rect 29388 19448 29754 19790
rect 29986 19846 30352 19874
rect 29986 19780 30130 19846
rect 30196 19780 30352 19846
rect 29986 19448 30352 19780
rect 30570 19840 30936 19872
rect 30570 19774 30728 19840
rect 30794 19774 30936 19840
rect 30570 19446 30936 19774
rect 31164 19838 31530 19874
rect 31164 19772 31318 19838
rect 31384 19772 31530 19838
rect 31164 19448 31530 19772
rect 23588 18626 23724 18632
rect 23588 18484 23724 18490
rect 22479 17529 23434 17710
rect 20142 16352 20148 16556
rect 20200 16352 20206 16556
rect 23253 15125 23434 17529
rect 26022 16910 26918 17110
rect 25042 16820 25048 16872
rect 25100 16820 25106 16872
rect 27848 15751 27978 15772
rect 27848 15673 27869 15751
rect 27947 15673 27978 15751
rect 27848 15660 27978 15673
rect 23253 14944 23602 15125
rect 25727 14982 27032 15110
rect 25784 14961 25798 14982
<< via1 >>
rect 29942 44372 29994 44424
rect 29830 44160 29882 44212
rect 29732 44010 29784 44062
rect 29628 43920 29680 43972
rect 22190 41268 22242 41320
rect 21990 41178 22042 41230
rect 22272 41172 22324 41224
rect 22272 40475 22324 40527
rect 29628 40199 29680 40251
rect 29732 39739 29784 39791
rect 22288 39647 22340 39699
rect 29942 41027 29994 41079
rect 21990 38451 22042 38503
rect 29722 38451 29774 38503
rect 20201 36489 20519 36807
rect 23624 34946 23754 35296
rect 27592 34944 27722 35294
rect 31540 34944 31670 35294
rect 23257 34500 23309 34552
rect 27298 34486 27350 34538
rect 31289 34490 31341 34542
rect 21782 33766 21866 33854
rect 25754 33768 25838 33856
rect 29792 33764 29876 33852
rect 20558 33120 20618 33180
rect 23238 31498 23290 31550
rect 21776 30760 21860 30848
rect 20544 30108 20604 30168
rect 23286 28486 23338 28538
rect 21774 27762 21858 27850
rect 20560 27092 20620 27152
rect 23264 25484 23316 25536
rect 21776 24762 21860 24850
rect 20568 24092 20628 24152
rect 23308 22492 23360 22544
rect 21766 21760 21850 21848
rect 20550 21104 20610 21164
rect 22582 20838 22792 20914
rect 24586 33140 24646 33200
rect 27260 31492 27312 31544
rect 25748 30774 25832 30862
rect 24530 30104 24590 30164
rect 27236 28498 27288 28550
rect 25756 27760 25840 27848
rect 24530 27082 24590 27142
rect 27273 25500 27325 25552
rect 25736 24772 25820 24860
rect 24536 24120 24596 24180
rect 27238 22498 27290 22550
rect 25766 21768 25850 21856
rect 24542 21088 24602 21148
rect 28598 33144 28658 33204
rect 31306 31488 31358 31540
rect 29796 30756 29880 30844
rect 28528 30086 28588 30146
rect 31266 28484 31318 28536
rect 29784 27754 29868 27842
rect 28536 27110 28596 27170
rect 31288 25492 31340 25544
rect 29802 24762 29886 24850
rect 28532 24106 28592 24166
rect 31206 22502 31258 22554
rect 29798 21770 29882 21858
rect 28538 21104 28598 21164
rect 20130 18523 20330 18575
rect 20430 18525 20630 18585
rect 20732 18528 20932 18585
rect 21054 18538 21254 18591
rect 21364 18531 21564 18585
rect 21688 18539 21888 18591
rect 22002 18533 22202 18585
rect 22334 18537 22534 18589
rect 27458 20318 27534 20384
rect 28052 20318 28128 20384
rect 28648 20326 28714 20392
rect 29232 20332 29298 20398
rect 29836 20306 29902 20372
rect 30428 20330 30494 20396
rect 31026 20332 31092 20398
rect 27164 19758 27240 19832
rect 27764 19800 27840 19866
rect 28350 19784 28426 19850
rect 28942 19786 29008 19852
rect 29546 19790 29612 19856
rect 30130 19780 30196 19846
rect 30728 19774 30794 19840
rect 31318 19772 31384 19838
rect 23588 18490 23724 18626
rect 20148 16352 20200 16556
rect 24329 16771 24407 16849
rect 25048 16820 25100 16872
rect 27408 15702 27468 15762
rect 27869 15673 27947 15751
<< metal2 >>
rect 13841 44468 13850 44528
rect 13910 44512 13919 44528
rect 13910 44484 25532 44512
rect 13910 44468 13919 44484
rect 14424 44434 14484 44443
rect 14484 44390 25384 44418
rect 14424 44365 14484 44374
rect 14954 44297 14963 44357
rect 15023 44345 15032 44357
rect 25048 44354 25154 44356
rect 25048 44345 25096 44354
rect 15023 44308 25096 44345
rect 15023 44297 15032 44308
rect 25048 44298 25096 44308
rect 25152 44298 25161 44354
rect 25356 44324 25384 44390
rect 25504 44412 25532 44484
rect 29936 44412 29942 44424
rect 25504 44384 29942 44412
rect 29936 44372 29942 44384
rect 29994 44372 30000 44424
rect 25048 44296 25154 44298
rect 25356 44296 28040 44324
rect 27776 44262 27874 44264
rect 16055 44201 16064 44261
rect 16124 44248 16133 44261
rect 16554 44248 16768 44256
rect 16124 44232 23510 44248
rect 27776 44232 27816 44262
rect 16124 44224 27816 44232
rect 16124 44214 16588 44224
rect 16724 44214 27816 44224
rect 16124 44201 16133 44214
rect 23411 44206 27816 44214
rect 27872 44206 27881 44262
rect 23411 44204 27874 44206
rect 16617 44136 16626 44196
rect 16686 44180 16695 44196
rect 23411 44193 27826 44204
rect 28012 44200 28040 44296
rect 29824 44200 29830 44212
rect 16686 44160 23352 44180
rect 28012 44172 29830 44200
rect 29824 44160 29830 44172
rect 29882 44160 29888 44212
rect 16686 44152 26674 44160
rect 16686 44136 16695 44152
rect 23324 44132 26674 44152
rect 17157 44059 17166 44119
rect 17226 44105 17235 44119
rect 23114 44105 23192 44116
rect 17226 44073 23192 44105
rect 17226 44059 17235 44073
rect 23114 44062 23192 44073
rect 26444 44086 26522 44096
rect 18256 43984 18265 44044
rect 18325 44028 18334 44044
rect 26444 44042 26456 44086
rect 18734 44028 18930 44032
rect 23369 44030 26456 44042
rect 26512 44030 26522 44086
rect 23369 44028 26522 44030
rect 18325 44008 26522 44028
rect 26646 44050 26674 44132
rect 29732 44062 29784 44068
rect 26646 44022 29732 44050
rect 18325 44007 26502 44008
rect 18325 44004 23401 44007
rect 29732 44004 29784 44010
rect 18325 43999 18762 44004
rect 18898 44000 23401 44004
rect 18898 43999 23372 44000
rect 18325 43984 18334 43999
rect 17720 43914 17780 43923
rect 18791 43916 18800 43976
rect 18860 43960 18869 43976
rect 29622 43960 29628 43972
rect 18860 43932 29628 43960
rect 18860 43916 18869 43932
rect 29622 43920 29628 43932
rect 29680 43920 29686 43972
rect 17780 43888 18762 43898
rect 18898 43888 22390 43898
rect 17780 43870 22390 43888
rect 18712 43862 18946 43870
rect 18734 43858 18922 43862
rect 17720 43845 17780 43854
rect 15507 43774 15516 43834
rect 15576 43818 15585 43834
rect 19218 43818 22312 43836
rect 15576 43816 17688 43818
rect 17814 43816 22312 43818
rect 15576 43808 22312 43816
rect 15576 43790 19246 43808
rect 15576 43774 15585 43790
rect 17666 43788 17838 43790
rect 13297 43702 13306 43762
rect 13366 43746 13375 43762
rect 19350 43746 22230 43766
rect 13366 43738 22230 43746
rect 13366 43718 19378 43738
rect 13366 43702 13375 43718
rect 12731 43596 12740 43656
rect 12800 43640 12809 43656
rect 12800 43612 22030 43640
rect 12800 43596 12809 43612
rect 22002 41230 22030 43612
rect 22202 41320 22230 43738
rect 22184 41268 22190 41320
rect 22242 41268 22248 41320
rect 21984 41178 21990 41230
rect 22042 41178 22048 41230
rect 22284 41224 22312 43808
rect 22266 41172 22272 41224
rect 22324 41172 22330 41224
rect 22362 41039 22390 43870
rect 29936 41079 30000 41086
rect 29936 41027 29942 41079
rect 29994 41027 30000 41079
rect 29936 41020 30000 41027
rect 22272 40527 22324 40533
rect 22272 40469 22324 40475
rect 29622 40251 29688 40258
rect 29622 40199 29628 40251
rect 29680 40199 29688 40251
rect 29622 40192 29688 40199
rect 29732 39791 29784 39797
rect 29732 39733 29784 39739
rect 22282 39699 22348 39706
rect 22282 39647 22288 39699
rect 22340 39647 22348 39699
rect 22282 39640 22348 39647
rect 29610 39151 29694 39160
rect 29610 39091 29624 39151
rect 29684 39091 29694 39151
rect 29610 39082 29694 39091
rect 29714 38503 29780 38510
rect 21984 38451 21990 38503
rect 22042 38451 22048 38503
rect 29714 38451 29722 38503
rect 29774 38451 29780 38503
rect 29714 38444 29780 38451
rect 20194 36807 20526 36814
rect 20194 36489 20201 36807
rect 20519 36489 20526 36807
rect 20194 36482 20526 36489
rect 24648 36096 25154 36098
rect 20072 36076 21754 36078
rect 20072 36020 21696 36076
rect 21752 36020 21761 36076
rect 24648 36040 25096 36096
rect 25152 36040 25161 36096
rect 24648 36038 25154 36040
rect 20072 36018 21754 36020
rect 20072 21164 20132 36018
rect 20172 35926 23794 35928
rect 20172 35870 23736 35926
rect 23792 35870 23801 35926
rect 20172 35868 23794 35870
rect 20172 24152 20232 35868
rect 20316 35788 24474 35790
rect 20316 35732 24416 35788
rect 24472 35732 24481 35788
rect 20316 35730 24474 35732
rect 20316 27152 20376 35730
rect 20442 35670 23114 35672
rect 20442 35614 23056 35670
rect 23112 35614 23121 35670
rect 20442 35612 23114 35614
rect 20442 30168 20502 35612
rect 20554 35532 22434 35534
rect 20554 35476 22376 35532
rect 22432 35476 22441 35532
rect 20554 35474 22434 35476
rect 20558 33180 20618 35474
rect 23596 35296 23776 35328
rect 23596 34946 23624 35296
rect 23754 34946 23776 35296
rect 23596 34924 23776 34946
rect 23251 34500 23257 34552
rect 23309 34541 23315 34552
rect 23309 34510 23772 34541
rect 23309 34500 23315 34510
rect 21764 33854 21880 33880
rect 21764 33766 21782 33854
rect 21866 33766 21880 33854
rect 21764 33754 21880 33766
rect 20558 33114 20618 33120
rect 23232 31498 23238 31550
rect 23290 31538 23296 31550
rect 23290 31510 23702 31538
rect 23290 31498 23296 31510
rect 21758 30848 21874 30864
rect 21758 30760 21776 30848
rect 21860 30760 21874 30848
rect 21758 30738 21874 30760
rect 20442 30108 20544 30168
rect 20604 30108 20610 30168
rect 23280 28486 23286 28538
rect 23338 28527 23344 28538
rect 23338 28497 23623 28527
rect 23338 28486 23344 28497
rect 21758 27850 21874 27874
rect 21758 27762 21774 27850
rect 21858 27762 21874 27850
rect 21758 27748 21874 27762
rect 20316 27092 20560 27152
rect 20620 27092 20626 27152
rect 23258 25484 23264 25536
rect 23316 25528 23322 25536
rect 23316 25492 23538 25528
rect 23316 25484 23322 25492
rect 21758 24850 21874 24874
rect 21758 24762 21776 24850
rect 21860 24762 21874 24850
rect 21758 24748 21874 24762
rect 20172 24092 20568 24152
rect 20628 24092 20634 24152
rect 23302 22492 23308 22544
rect 23360 22535 23366 22544
rect 23360 22501 23439 22535
rect 23360 22492 23366 22501
rect 21750 21848 21866 21866
rect 21750 21760 21766 21848
rect 21850 21760 21866 21848
rect 21750 21740 21866 21760
rect 20072 21104 20550 21164
rect 20610 21104 20616 21164
rect 22562 20914 22812 20936
rect 22562 20838 22582 20914
rect 22792 20838 22812 20914
rect 22562 20812 22812 20838
rect 20036 20733 22458 20780
rect 20036 20635 22124 20678
rect 20036 20552 21809 20594
rect 20036 20442 21491 20496
rect 20036 20333 21181 20386
rect 20036 20215 20861 20272
rect 20036 20080 20560 20140
rect 20036 19958 20255 20007
rect 20206 18575 20255 19958
rect 20500 18585 20560 20080
rect 20804 18585 20861 20215
rect 21128 18591 21181 20333
rect 20124 18523 20130 18575
rect 20330 18523 20336 18575
rect 20424 18525 20430 18585
rect 20630 18525 20636 18585
rect 20726 18528 20732 18585
rect 20932 18528 20938 18585
rect 21048 18538 21054 18591
rect 21254 18538 21260 18591
rect 21437 18585 21491 20442
rect 21767 18591 21809 20552
rect 21358 18531 21364 18585
rect 21564 18531 21570 18585
rect 21682 18539 21688 18591
rect 21888 18539 21894 18591
rect 22081 18585 22124 20635
rect 22411 18589 22458 20733
rect 22616 18626 22752 20812
rect 23405 20321 23439 22501
rect 23502 20402 23538 25492
rect 23593 20467 23623 28497
rect 23674 20528 23702 31510
rect 23741 20593 23772 34510
rect 24648 33978 24708 36038
rect 24096 33918 24708 33978
rect 24766 35942 25834 35944
rect 24766 35886 25776 35942
rect 25832 35886 25841 35942
rect 30536 35896 30592 35903
rect 28664 35894 30594 35896
rect 24766 35884 25834 35886
rect 24096 21148 24156 33918
rect 24766 33754 24826 35884
rect 28664 35838 30536 35894
rect 30592 35838 30594 35894
rect 28664 35836 30594 35838
rect 24230 33694 24826 33754
rect 24886 35800 26514 35802
rect 24886 35744 26456 35800
rect 26512 35744 26521 35800
rect 24886 35742 26514 35744
rect 24230 24180 24290 33694
rect 24886 33564 24946 35742
rect 24350 33504 24946 33564
rect 24984 35656 27194 35658
rect 24984 35600 27136 35656
rect 27192 35600 27201 35656
rect 24984 35598 27194 35600
rect 24350 27142 24410 33504
rect 24984 33362 25044 35598
rect 24462 33302 25044 33362
rect 25108 35512 28554 35514
rect 25108 35456 28496 35512
rect 28552 35456 28561 35512
rect 25108 35454 28554 35456
rect 24462 30164 24522 33302
rect 25108 33200 25168 35454
rect 27560 35294 27740 35324
rect 27560 34944 27592 35294
rect 27722 34944 27740 35294
rect 27560 34920 27740 34944
rect 27292 34486 27298 34538
rect 27350 34527 27356 34538
rect 27350 34497 27693 34527
rect 27350 34486 27356 34497
rect 25736 33856 25852 33878
rect 25736 33768 25754 33856
rect 25838 33768 25852 33856
rect 25736 33752 25852 33768
rect 24580 33140 24586 33200
rect 24646 33140 25168 33200
rect 27254 31492 27260 31544
rect 27312 31539 27318 31544
rect 27312 31497 27619 31539
rect 27312 31492 27318 31497
rect 25736 30862 25852 30886
rect 25736 30774 25748 30862
rect 25832 30774 25852 30862
rect 25736 30760 25852 30774
rect 24462 30104 24530 30164
rect 24590 30104 24596 30164
rect 27230 28498 27236 28550
rect 27288 28541 27294 28550
rect 27288 28507 27543 28541
rect 27288 28498 27294 28507
rect 25736 27848 25852 27872
rect 25736 27760 25756 27848
rect 25840 27760 25852 27848
rect 25736 27746 25852 27760
rect 24350 27082 24530 27142
rect 24590 27082 24596 27142
rect 27267 25500 27273 25552
rect 27325 25540 27331 25552
rect 27325 25511 27475 25540
rect 27325 25500 27331 25511
rect 25722 24860 25838 24884
rect 25722 24772 25736 24860
rect 25820 24772 25838 24860
rect 25722 24758 25838 24772
rect 24230 24120 24536 24180
rect 24596 24120 24602 24180
rect 27232 22498 27238 22550
rect 27290 22538 27296 22550
rect 27290 22510 27418 22538
rect 27290 22498 27296 22510
rect 25746 21856 25862 21878
rect 25746 21768 25766 21856
rect 25850 21768 25862 21856
rect 25746 21752 25862 21768
rect 24096 21088 24542 21148
rect 24602 21088 24608 21148
rect 27390 20690 27418 22510
rect 27446 20748 27475 25511
rect 27509 20813 27543 28507
rect 27577 20891 27619 31497
rect 27663 20965 27693 34497
rect 28664 33878 28724 35836
rect 30536 35829 30592 35836
rect 28056 33818 28724 33878
rect 28810 35748 29234 35750
rect 28810 35692 29176 35748
rect 29232 35692 29241 35748
rect 28810 35690 29234 35692
rect 28056 21164 28116 33818
rect 28810 33698 28870 35690
rect 29058 35606 29914 35608
rect 29058 35550 29856 35606
rect 29912 35550 29921 35606
rect 29058 35548 29914 35550
rect 28936 35370 28992 35377
rect 28188 33638 28870 33698
rect 28934 35368 28994 35370
rect 28934 35312 28936 35368
rect 28992 35312 28994 35368
rect 28188 24166 28248 33638
rect 28934 33540 28994 35312
rect 28342 33480 28994 33540
rect 28342 27170 28402 33480
rect 29058 33386 29118 35548
rect 28470 33326 29118 33386
rect 29192 35474 29684 35476
rect 29192 35418 29626 35474
rect 29682 35418 29691 35474
rect 29192 35416 29684 35418
rect 28470 30146 28530 33326
rect 29192 33204 29252 35416
rect 31514 35294 31694 35320
rect 31514 34944 31540 35294
rect 31670 34944 31694 35294
rect 31514 34916 31694 34944
rect 31283 34490 31289 34542
rect 31341 34530 31347 34542
rect 31341 34501 31670 34530
rect 31341 34490 31347 34501
rect 29776 33852 29892 33874
rect 29776 33764 29792 33852
rect 29876 33764 29892 33852
rect 29776 33748 29892 33764
rect 28592 33144 28598 33204
rect 28658 33144 29252 33204
rect 31300 31488 31306 31540
rect 31358 31528 31364 31540
rect 31358 31500 31606 31528
rect 31358 31488 31364 31500
rect 29784 30844 29900 30868
rect 29784 30756 29796 30844
rect 29880 30756 29900 30844
rect 29784 30742 29900 30756
rect 28470 30086 28528 30146
rect 28588 30086 28594 30146
rect 31266 28536 31318 28542
rect 31318 28495 31541 28525
rect 31266 28478 31318 28484
rect 29766 27842 29882 27860
rect 29766 27754 29784 27842
rect 29868 27754 29882 27842
rect 29766 27734 29882 27754
rect 28342 27110 28536 27170
rect 28596 27110 28602 27170
rect 31282 25492 31288 25544
rect 31340 25532 31346 25544
rect 31340 25504 31482 25532
rect 31340 25492 31346 25504
rect 29790 24850 29906 24876
rect 29790 24762 29802 24850
rect 29886 24762 29906 24850
rect 29790 24750 29906 24762
rect 28188 24106 28532 24166
rect 28592 24106 28598 24166
rect 31200 22502 31206 22554
rect 31258 22543 31264 22554
rect 31258 22513 31423 22543
rect 31258 22502 31264 22513
rect 29782 21858 29898 21884
rect 29782 21770 29798 21858
rect 29882 21770 29898 21858
rect 29782 21758 29898 21770
rect 28056 21104 28538 21164
rect 28598 21104 28604 21164
rect 27663 20935 29930 20965
rect 27577 20849 29550 20891
rect 27509 20779 29244 20813
rect 27446 20719 28957 20748
rect 27390 20662 28664 20690
rect 23741 20562 28357 20593
rect 23674 20500 28058 20528
rect 23593 20437 27772 20467
rect 23502 20394 27468 20402
rect 23502 20384 27546 20394
rect 23502 20366 27458 20384
rect 27432 20324 27458 20366
rect 23405 20287 27168 20321
rect 27442 20318 27458 20324
rect 27534 20318 27546 20384
rect 27442 20300 27546 20318
rect 27134 19840 27168 20287
rect 27742 19878 27772 20437
rect 28030 20398 28058 20500
rect 28030 20384 28140 20398
rect 28030 20324 28052 20384
rect 28036 20318 28052 20324
rect 28128 20318 28140 20384
rect 28036 20304 28140 20318
rect 27742 19866 27854 19878
rect 27134 19832 27260 19840
rect 27134 19799 27164 19832
rect 27138 19758 27164 19799
rect 27240 19758 27260 19832
rect 27742 19803 27764 19866
rect 27750 19800 27764 19803
rect 27840 19800 27854 19866
rect 27750 19784 27854 19800
rect 28326 19862 28357 20562
rect 28636 20410 28664 20662
rect 28636 20392 28740 20410
rect 28636 20326 28648 20392
rect 28714 20326 28740 20392
rect 28636 20316 28740 20326
rect 28928 19868 28957 20719
rect 29210 20416 29244 20779
rect 29210 20398 29322 20416
rect 29210 20390 29232 20398
rect 29218 20332 29232 20390
rect 29298 20332 29322 20398
rect 29218 20322 29322 20332
rect 29508 19878 29550 20849
rect 29900 20388 29930 20935
rect 31393 20603 31423 22513
rect 29824 20372 29930 20388
rect 29824 20306 29836 20372
rect 29902 20341 29930 20372
rect 30192 20573 31423 20603
rect 29902 20306 29928 20341
rect 29824 20294 29928 20306
rect 28326 19850 28436 19862
rect 28326 19791 28350 19850
rect 28332 19784 28350 19791
rect 28426 19784 28436 19850
rect 28332 19768 28436 19784
rect 28928 19852 29032 19868
rect 28928 19786 28942 19852
rect 29008 19786 29032 19852
rect 29508 19856 29646 19878
rect 30192 19862 30222 20573
rect 31454 20544 31482 25504
rect 30494 20516 31482 20544
rect 30494 20412 30522 20516
rect 31511 20475 31541 28495
rect 30418 20396 30522 20412
rect 30418 20330 30428 20396
rect 30494 20330 30522 20396
rect 30418 20318 30522 20330
rect 30792 20445 31541 20475
rect 29508 19815 29546 19856
rect 28928 19774 29032 19786
rect 29512 19790 29546 19815
rect 29612 19790 29646 19856
rect 29512 19772 29646 19790
rect 30114 19846 30222 19862
rect 30792 19856 30822 20445
rect 31008 20398 31112 20410
rect 31578 20398 31606 31500
rect 31008 20332 31026 20398
rect 31092 20370 31606 20398
rect 31092 20332 31112 20370
rect 31008 20316 31112 20332
rect 31641 19857 31670 34501
rect 30114 19780 30130 19846
rect 30196 19811 30222 19846
rect 30716 19840 30822 19856
rect 30196 19780 30218 19811
rect 30114 19768 30218 19780
rect 30716 19774 30728 19840
rect 30794 19823 30822 19840
rect 31296 19838 31670 19857
rect 31296 19828 31318 19838
rect 30794 19774 30820 19823
rect 30716 19762 30820 19774
rect 31302 19772 31318 19828
rect 31384 19828 31670 19838
rect 31384 19772 31406 19828
rect 27138 19744 27260 19758
rect 31302 19756 31406 19772
rect 21996 18533 22002 18585
rect 22202 18533 22208 18585
rect 22328 18537 22334 18589
rect 22534 18537 22540 18589
rect 22616 18490 23588 18626
rect 23724 18490 23730 18626
rect 25048 16872 25100 16878
rect 24312 16849 24422 16860
rect 24312 16771 24329 16849
rect 24407 16771 24422 16849
rect 25048 16814 25100 16820
rect 24312 16758 24422 16771
rect 25049 16597 25099 16814
rect 26745 16597 26754 16602
rect 20148 16556 20200 16562
rect 22567 16547 26754 16597
rect 22567 16479 22617 16547
rect 26745 16542 26754 16547
rect 26814 16542 26823 16602
rect 20200 16429 22617 16479
rect 20148 16346 20200 16352
rect 27390 15762 27494 15780
rect 27390 15702 27408 15762
rect 27468 15702 27494 15762
rect 27390 15688 27494 15702
rect 27848 15751 27978 15772
rect 27848 15673 27869 15751
rect 27947 15673 27978 15751
rect 27848 15660 27978 15673
<< via2 >>
rect 13850 44468 13910 44528
rect 14424 44374 14484 44434
rect 14963 44297 15023 44357
rect 25096 44298 25152 44354
rect 16064 44201 16124 44261
rect 27816 44206 27872 44262
rect 16626 44136 16686 44196
rect 17166 44059 17226 44119
rect 18265 43984 18325 44044
rect 26456 44030 26512 44086
rect 18800 43916 18860 43976
rect 17720 43854 17780 43914
rect 15516 43774 15576 43834
rect 13306 43702 13366 43762
rect 12740 43596 12800 43656
rect 29624 39091 29684 39151
rect 20206 36494 20514 36802
rect 21696 36020 21752 36076
rect 25096 36040 25152 36096
rect 23736 35870 23792 35926
rect 24416 35732 24472 35788
rect 23056 35614 23112 35670
rect 22376 35476 22432 35532
rect 23624 34946 23754 35296
rect 21782 33766 21866 33854
rect 21776 30760 21860 30848
rect 21774 27762 21858 27850
rect 21776 24762 21860 24850
rect 21766 21760 21850 21848
rect 25776 35886 25832 35942
rect 30536 35838 30592 35894
rect 26456 35744 26512 35800
rect 27136 35600 27192 35656
rect 28496 35456 28552 35512
rect 27592 34944 27722 35294
rect 25754 33768 25838 33856
rect 25748 30774 25832 30862
rect 25756 27760 25840 27848
rect 25736 24772 25820 24860
rect 25766 21768 25850 21856
rect 29176 35692 29232 35748
rect 29856 35550 29912 35606
rect 28936 35312 28992 35368
rect 29626 35418 29682 35474
rect 31540 34944 31670 35294
rect 29792 33764 29876 33852
rect 29796 30756 29880 30844
rect 29784 27754 29868 27842
rect 29802 24762 29886 24850
rect 29798 21770 29882 21858
rect 24334 16776 24402 16844
rect 26754 16542 26814 16602
rect 27410 15704 27466 15760
rect 27874 15678 27942 15746
<< metal3 >>
rect 28492 45082 28556 45088
rect 14422 45074 14486 45080
rect 12738 45062 12802 45068
rect 13848 45066 13912 45072
rect 12738 44992 12802 44998
rect 13304 45058 13368 45064
rect 17164 45070 17228 45076
rect 14422 45004 14486 45010
rect 14961 45060 15025 45066
rect 13848 44996 13912 45002
rect 12740 43661 12800 44992
rect 13304 44988 13368 44994
rect 13306 43767 13366 44988
rect 13850 44533 13910 44996
rect 13845 44528 13915 44533
rect 13845 44468 13850 44528
rect 13910 44468 13915 44528
rect 13845 44463 13915 44468
rect 14424 44439 14484 45004
rect 14961 44990 15025 44996
rect 15514 45064 15578 45070
rect 16624 45054 16688 45060
rect 15514 44994 15578 45000
rect 16062 45048 16126 45054
rect 14419 44434 14489 44439
rect 14419 44374 14424 44434
rect 14484 44374 14489 44434
rect 14419 44369 14489 44374
rect 14963 44362 15023 44990
rect 14958 44357 15028 44362
rect 14958 44297 14963 44357
rect 15023 44297 15028 44357
rect 14958 44292 15028 44297
rect 15516 43839 15576 44994
rect 18798 45068 18862 45074
rect 18263 45062 18327 45068
rect 17164 45000 17228 45006
rect 17718 45056 17782 45062
rect 16624 44984 16688 44990
rect 16062 44978 16126 44984
rect 16064 44266 16124 44978
rect 16059 44261 16129 44266
rect 16059 44201 16064 44261
rect 16124 44201 16129 44261
rect 16626 44201 16686 44984
rect 16059 44196 16129 44201
rect 16621 44196 16691 44201
rect 16621 44136 16626 44196
rect 16686 44136 16691 44196
rect 16621 44131 16691 44136
rect 17166 44124 17226 45000
rect 18798 44998 18862 45004
rect 28480 45018 28492 45026
rect 28556 45018 28568 45026
rect 18263 44992 18327 44998
rect 17718 44986 17782 44992
rect 17161 44119 17231 44124
rect 17161 44059 17166 44119
rect 17226 44059 17231 44119
rect 17161 44054 17231 44059
rect 17720 43919 17780 44986
rect 18265 44049 18325 44992
rect 18260 44044 18330 44049
rect 18260 43984 18265 44044
rect 18325 43984 18330 44044
rect 18260 43979 18330 43984
rect 18800 43981 18860 44998
rect 28480 44946 28568 45018
rect 25091 44354 25157 44359
rect 25091 44298 25096 44354
rect 25152 44298 25157 44354
rect 25091 44293 25157 44298
rect 25094 44052 25154 44293
rect 27811 44262 27877 44267
rect 27811 44206 27816 44262
rect 27872 44206 27877 44262
rect 27811 44201 27877 44206
rect 26451 44086 26517 44091
rect 26451 44030 26456 44086
rect 26512 44030 26517 44086
rect 27814 44064 27874 44201
rect 28494 44094 28554 44946
rect 26451 44025 26517 44030
rect 18795 43976 18865 43981
rect 17715 43914 17785 43919
rect 17715 43854 17720 43914
rect 17780 43854 17785 43914
rect 18795 43916 18800 43976
rect 18860 43916 18865 43976
rect 18795 43911 18865 43916
rect 17715 43849 17785 43854
rect 15511 43834 15581 43839
rect 15511 43774 15516 43834
rect 15576 43774 15581 43834
rect 15511 43769 15581 43774
rect 13301 43762 13371 43767
rect 13301 43702 13306 43762
rect 13366 43702 13371 43762
rect 13301 43697 13371 43702
rect 12735 43656 12805 43661
rect 12735 43596 12740 43656
rect 12800 43596 12805 43656
rect 12735 43591 12805 43596
rect 20775 40753 21093 40754
rect 20770 40437 20776 40753
rect 21092 40437 21098 40753
rect 20196 40095 20524 40102
rect 20196 39948 20202 40095
rect 20201 39779 20202 39948
rect 20518 39948 20524 40095
rect 20518 39779 20519 39948
rect 20201 36814 20519 39779
rect 20194 36802 20526 36814
rect 20194 36494 20206 36802
rect 20514 36494 20526 36802
rect 20194 36482 20526 36494
rect 20775 35297 21093 40437
rect 21968 39778 22700 40096
rect 29619 39151 29689 39156
rect 29619 39091 29624 39151
rect 29684 39091 29689 39151
rect 29619 39086 29689 39091
rect 21694 36081 21754 36532
rect 21691 36076 21757 36081
rect 21691 36020 21696 36076
rect 21752 36020 21757 36076
rect 21691 36015 21757 36020
rect 22374 35568 22434 36646
rect 23054 35675 23114 36548
rect 23734 35931 23794 36502
rect 23731 35926 23797 35931
rect 23731 35870 23736 35926
rect 23792 35870 23797 35926
rect 23731 35865 23797 35870
rect 24414 35793 24474 36532
rect 25094 36101 25154 36568
rect 25091 36096 25157 36101
rect 25091 36040 25096 36096
rect 25152 36040 25157 36096
rect 25091 36035 25157 36040
rect 25774 35947 25834 36572
rect 25771 35942 25837 35947
rect 25771 35886 25776 35942
rect 25832 35886 25837 35942
rect 25771 35881 25837 35886
rect 26454 35805 26514 36600
rect 26451 35800 26517 35805
rect 24411 35788 24477 35793
rect 24411 35732 24416 35788
rect 24472 35732 24477 35788
rect 26451 35744 26456 35800
rect 26512 35744 26517 35800
rect 26451 35739 26517 35744
rect 24411 35727 24477 35732
rect 23051 35670 23117 35675
rect 23051 35614 23056 35670
rect 23112 35614 23117 35670
rect 27134 35661 27194 36596
rect 23051 35609 23117 35614
rect 27131 35656 27197 35661
rect 27131 35600 27136 35656
rect 27192 35600 27197 35656
rect 27131 35595 27197 35600
rect 22370 35532 22438 35568
rect 22370 35486 22376 35532
rect 22371 35476 22376 35486
rect 22432 35486 22438 35532
rect 22432 35476 22437 35486
rect 22371 35471 22437 35476
rect 27814 35370 27874 36480
rect 28494 35564 28554 36578
rect 29174 35753 29234 36538
rect 29171 35748 29237 35753
rect 29171 35692 29176 35748
rect 29232 35692 29237 35748
rect 29171 35687 29237 35692
rect 28490 35512 28558 35564
rect 28490 35488 28496 35512
rect 28491 35456 28496 35488
rect 28552 35488 28558 35512
rect 28552 35456 28557 35488
rect 29624 35479 29684 39086
rect 29854 35611 29914 36530
rect 30534 35899 30594 36508
rect 30531 35894 30597 35899
rect 30531 35838 30536 35894
rect 30592 35838 30597 35894
rect 30531 35833 30597 35838
rect 29851 35606 29917 35611
rect 29851 35550 29856 35606
rect 29912 35550 29917 35606
rect 29851 35545 29917 35550
rect 28491 35451 28557 35456
rect 29621 35474 29687 35479
rect 29621 35418 29626 35474
rect 29682 35418 29687 35474
rect 29621 35413 29687 35418
rect 28931 35370 28997 35373
rect 27814 35368 28997 35370
rect 23596 35297 23776 35328
rect 27560 35297 27740 35324
rect 27814 35312 28936 35368
rect 28992 35312 28997 35368
rect 27814 35310 28997 35312
rect 28931 35307 28997 35310
rect 20773 35296 27740 35297
rect 20773 34975 23624 35296
rect 23596 34946 23624 34975
rect 23754 35294 27740 35296
rect 23754 34975 27592 35294
rect 23754 34946 23776 34975
rect 23596 34924 23776 34946
rect 27560 34944 27592 34975
rect 27722 35250 27740 35294
rect 31514 35294 31694 35320
rect 31514 35250 31540 35294
rect 27722 35246 28870 35250
rect 29060 35246 31540 35250
rect 27722 35022 31540 35246
rect 27722 34944 27740 35022
rect 27560 34920 27740 34944
rect 31514 34944 31540 35022
rect 31670 34944 31694 35294
rect 31514 34916 31694 34944
rect 21764 33870 21880 33880
rect 25736 33870 25852 33878
rect 29776 33870 29892 33874
rect 21760 33856 29896 33870
rect 21760 33854 25754 33856
rect 21760 33766 21782 33854
rect 21866 33768 25754 33854
rect 25838 33852 29896 33856
rect 25838 33768 29792 33852
rect 21866 33766 29792 33768
rect 21760 33764 29792 33766
rect 29876 33764 29896 33852
rect 21760 33744 29896 33764
rect 25736 30868 25852 30886
rect 27813 30868 27939 33744
rect 21748 30862 29900 30868
rect 21748 30848 25748 30862
rect 21748 30760 21776 30848
rect 21860 30774 25748 30848
rect 25832 30844 29900 30862
rect 25832 30774 29796 30844
rect 21860 30760 29796 30774
rect 21748 30756 29796 30760
rect 29880 30756 29900 30844
rect 21748 30742 29900 30756
rect 21758 30738 21874 30742
rect 21758 27868 21874 27874
rect 25736 27868 25852 27872
rect 27813 27868 27939 30742
rect 21758 27850 29898 27868
rect 21758 27762 21774 27850
rect 21858 27848 29898 27850
rect 21858 27762 25756 27848
rect 21758 27760 25756 27762
rect 25840 27842 29898 27848
rect 25840 27760 29784 27842
rect 21758 27754 29784 27760
rect 29868 27754 29898 27842
rect 21758 27748 29898 27754
rect 21762 27742 29898 27748
rect 25722 24876 25838 24884
rect 27813 24876 27939 27742
rect 29766 27734 29882 27742
rect 21760 24874 29906 24876
rect 21758 24860 29906 24874
rect 21758 24850 25736 24860
rect 21758 24762 21776 24850
rect 21860 24772 25736 24850
rect 25820 24850 29906 24860
rect 25820 24772 29802 24850
rect 21860 24762 29802 24772
rect 29886 24762 29906 24850
rect 21758 24750 29906 24762
rect 21758 24748 21874 24750
rect 25746 21866 25862 21878
rect 27813 21866 27939 24750
rect 29782 21866 29898 21884
rect 21748 21858 29898 21866
rect 21748 21856 29798 21858
rect 21748 21848 25766 21856
rect 21748 21760 21766 21848
rect 21850 21768 25766 21848
rect 25850 21770 29798 21856
rect 29882 21770 29898 21858
rect 25850 21768 29898 21770
rect 21850 21760 29898 21768
rect 21748 21758 29898 21760
rect 21748 21740 29884 21758
rect 27813 20461 27939 21740
rect 27813 20335 31673 20461
rect 31547 19445 31673 20335
rect 31547 19313 31673 19319
rect 24312 16848 24422 16860
rect 24312 16772 24330 16848
rect 24406 16772 24422 16848
rect 24312 16758 24422 16772
rect 26749 16602 26819 16607
rect 26749 16542 26754 16602
rect 26814 16542 27468 16602
rect 26749 16537 26819 16542
rect 27408 15765 27468 16542
rect 27405 15760 27471 15765
rect 27405 15704 27410 15760
rect 27466 15704 27471 15760
rect 27405 15699 27471 15704
rect 27848 15750 27978 15772
rect 27848 15674 27870 15750
rect 27946 15674 27978 15750
rect 27848 15660 27978 15674
<< via3 >>
rect 12738 44998 12802 45062
rect 13304 44994 13368 45058
rect 13848 45002 13912 45066
rect 14422 45010 14486 45074
rect 14961 44996 15025 45060
rect 15514 45000 15578 45064
rect 16062 44984 16126 45048
rect 16624 44990 16688 45054
rect 17164 45006 17228 45070
rect 17718 44992 17782 45056
rect 18263 44998 18327 45062
rect 18798 45004 18862 45068
rect 28492 45018 28556 45082
rect 20776 40437 21092 40753
rect 20202 39779 20518 40095
rect 31547 19319 31673 19445
rect 24330 16844 24406 16848
rect 24330 16776 24334 16844
rect 24334 16776 24402 16844
rect 24402 16776 24406 16844
rect 24330 16772 24406 16776
rect 27870 15746 27946 15750
rect 27870 15678 27874 15746
rect 27874 15678 27942 15746
rect 27942 15678 27946 15746
rect 27870 15674 27946 15678
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 45063 12818 45152
rect 12737 45062 12818 45063
rect 12737 44998 12738 45062
rect 12802 44998 12818 45062
rect 13310 45059 13370 45152
rect 13862 45067 13922 45152
rect 12737 44997 12818 44998
rect 12758 44952 12818 44997
rect 13303 45058 13370 45059
rect 13303 44994 13304 45058
rect 13368 44994 13370 45058
rect 13847 45066 13922 45067
rect 13847 45002 13848 45066
rect 13912 45002 13922 45066
rect 13847 45001 13922 45002
rect 13303 44993 13370 44994
rect 13310 44952 13370 44993
rect 13862 44952 13922 45001
rect 14414 45075 14474 45152
rect 14414 45074 14487 45075
rect 14414 45010 14422 45074
rect 14486 45010 14487 45074
rect 14966 45061 15026 45152
rect 15518 45065 15578 45152
rect 14414 45009 14487 45010
rect 14960 45060 15026 45061
rect 14414 44952 14474 45009
rect 14960 44996 14961 45060
rect 15025 44996 15026 45060
rect 15513 45064 15579 45065
rect 15513 45000 15514 45064
rect 15578 45000 15579 45064
rect 16070 45049 16130 45152
rect 15513 44999 15579 45000
rect 16061 45048 16130 45049
rect 14960 44995 15026 44996
rect 14966 44952 15026 44995
rect 15518 44952 15578 44999
rect 16061 44984 16062 45048
rect 16126 44984 16130 45048
rect 16061 44983 16130 44984
rect 16070 44952 16130 44983
rect 16622 45055 16682 45152
rect 17174 45071 17234 45152
rect 17163 45070 17234 45071
rect 16622 45054 16689 45055
rect 16622 44990 16624 45054
rect 16688 44990 16689 45054
rect 17163 45006 17164 45070
rect 17228 45006 17234 45070
rect 17726 45057 17786 45152
rect 18278 45063 18338 45152
rect 18830 45069 18890 45152
rect 17163 45005 17234 45006
rect 16622 44989 16689 44990
rect 16622 44952 16682 44989
rect 17174 44952 17234 45005
rect 17717 45056 17786 45057
rect 17717 44992 17718 45056
rect 17782 44992 17786 45056
rect 18262 45062 18338 45063
rect 18262 44998 18263 45062
rect 18327 44998 18338 45062
rect 18797 45068 18890 45069
rect 18797 45004 18798 45068
rect 18862 45004 18890 45068
rect 18797 45003 18890 45004
rect 18262 44997 18338 44998
rect 17717 44991 17786 44992
rect 17726 44952 17786 44991
rect 18278 44952 18338 44997
rect 18830 44952 18890 45003
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 45115 27722 45152
rect 27660 44979 27722 45115
rect 27662 44952 27722 44979
rect 28214 44952 28274 45152
rect 28491 45082 28557 45083
rect 28491 45018 28492 45082
rect 28556 45080 28557 45082
rect 28766 45080 28826 45152
rect 28556 45020 28826 45080
rect 28556 45018 28557 45020
rect 28491 45017 28557 45018
rect 28766 44952 28826 45020
rect 29318 44952 29378 45152
rect 200 1000 600 44152
rect 800 40096 1200 44152
rect 19756 40753 22696 40754
rect 19756 40437 20776 40753
rect 21092 40437 22696 40753
rect 19756 40436 22696 40437
rect 800 39778 1204 40096
rect 19756 40095 22700 40096
rect 19756 39779 20202 40095
rect 20518 39779 22700 40095
rect 19756 39778 22700 39779
rect 800 1000 1200 39778
rect 31546 19445 31674 19446
rect 31546 19319 31547 19445
rect 31673 19319 31674 19445
rect 31546 19318 31674 19319
rect 24329 16848 27949 16849
rect 24329 16772 24330 16848
rect 24406 16772 27949 16848
rect 24329 16771 27949 16772
rect 27871 15772 27949 16771
rect 27848 15751 27978 15772
rect 31547 15751 31673 19318
rect 27848 15750 31673 15751
rect 27848 15674 27870 15750
rect 27946 15674 31673 15750
rect 27848 15673 31673 15674
rect 27848 15660 27978 15673
rect 31547 213 31673 15673
rect 3314 0 3494 200
rect 7178 0 7358 204
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 202
rect 30409 200 31673 213
rect 30362 87 31673 200
rect 30362 0 30542 87
use bit4_encoder  bit4_encoder_0
timestamp 1730842790
transform 0 1 20296 -1 0 44963
box 0 0 9409 11553
use compr  compr_0
timestamp 1730838366
transform 0 1 20398 -1 0 24630
box 1230 -398 4034 3312
use compr  compr_1
timestamp 1730838366
transform 0 1 20408 -1 0 27618
box 1230 -398 4034 3312
use compr  compr_2
timestamp 1730838366
transform 0 1 20408 -1 0 30618
box 1230 -398 4034 3312
use compr  compr_3
timestamp 1730838366
transform 0 1 20408 -1 0 33628
box 1230 -398 4034 3312
use compr  compr_4
timestamp 1730838366
transform 0 1 20408 -1 0 36628
box 1230 -398 4034 3312
use compr  compr_5
timestamp 1730838366
transform 0 1 24384 -1 0 24630
box 1230 -398 4034 3312
use compr  compr_6
timestamp 1730838366
transform 0 1 24384 -1 0 27630
box 1230 -398 4034 3312
use compr  compr_7
timestamp 1730838366
transform 0 1 24384 -1 0 30618
box 1230 -398 4034 3312
use compr  compr_8
timestamp 1730838366
transform 0 1 24384 -1 0 33628
box 1230 -398 4034 3312
use compr  compr_9
timestamp 1730838366
transform 0 1 24384 -1 0 36618
box 1230 -398 4034 3312
use compr  compr_10
timestamp 1730838366
transform 0 1 28390 -1 0 24630
box 1230 -398 4034 3312
use compr  compr_11
timestamp 1730838366
transform 0 1 28390 -1 0 27630
box 1230 -398 4034 3312
use compr  compr_12
timestamp 1730838366
transform 0 1 28390 -1 0 30618
box 1230 -398 4034 3312
use compr  compr_13
timestamp 1730838366
transform 0 1 28400 -1 0 33618
box 1230 -398 4034 3312
use compr  compr_14
timestamp 1730838366
transform 0 1 28390 -1 0 36628
box 1230 -398 4034 3312
use compr  compr_15
timestamp 1730838366
transform 1 0 22252 0 1 15336
box 1230 -398 4034 3312
use pass_gate2  pass_gate2_0
timestamp 1730493024
transform 1 0 25466 0 1 16056
box 1380 -1118 2522 1056
use r2r_dac  r2r_dac_0
timestamp 1730635755
transform 1 0 18960 0 1 20409
box 1000 -5458 3772 -192
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR1
timestamp 1730493024
transform 1 0 31199 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR2
timestamp 1730493024
transform 1 0 29423 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR3
timestamp 1730493024
transform 1 0 30903 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR4
timestamp 1730493024
transform 1 0 31495 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR5
timestamp 1730493024
transform 1 0 29719 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR6
timestamp 1730493024
transform 1 0 27351 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR7
timestamp 1730493024
transform 1 0 30311 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR8
timestamp 1730493024
transform 1 0 28535 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR9
timestamp 1730493024
transform 1 0 30607 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR10
timestamp 1730493024
transform 1 0 30015 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR11
timestamp 1730493024
transform 1 0 27055 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR12
timestamp 1730493024
transform 1 0 28831 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR13
timestamp 1730493024
transform 1 0 27647 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR14
timestamp 1730493024
transform 1 0 27943 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR15
timestamp 1730493024
transform 1 0 29127 0 1 19932
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR16
timestamp 1730493024
transform 1 0 28239 0 1 19932
box -201 -652 201 652
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
