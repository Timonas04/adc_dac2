magic
tech sky130A
magscale 1 2
timestamp 1730635755
<< pwell >>
rect 3422 508 3600 654
rect 3128 -278 3276 -46
<< locali >>
rect 1274 3300 3834 3310
rect 1274 3128 1288 3300
rect 3822 3288 3834 3300
rect 3822 3232 3836 3288
rect 1274 3120 3638 3128
rect 3616 1178 3638 3120
rect 3830 1996 3836 3232
rect 3830 1178 3840 1996
rect 3830 934 3838 1178
rect 3128 652 3252 868
rect 3638 828 3688 886
rect 3830 828 3842 934
rect 3668 820 3842 828
rect 3128 284 3134 652
rect 3264 350 3498 414
rect 3264 304 3280 350
rect 3264 2 3278 304
rect 3264 -10 3532 2
rect 1270 -256 3134 -246
rect 1270 -378 1282 -256
rect 1270 -380 3532 -378
rect 3148 -382 3532 -380
<< viali >>
rect 1288 3232 3822 3300
rect 1288 3128 3830 3232
rect 3638 886 3830 3128
rect 3688 828 3830 886
rect 3134 -10 3264 652
rect 3134 -256 3532 -10
rect 1282 -378 3532 -256
<< metal1 >>
rect 1268 3300 3838 3312
rect 1268 3128 1288 3300
rect 3822 3286 3838 3300
rect 3822 3232 3844 3286
rect 1268 3120 3638 3128
rect 1354 1538 1416 2960
rect 1352 1366 1416 1538
rect 1352 1250 1400 1366
rect 1482 1322 1576 3052
rect 1676 2956 1720 3120
rect 1868 2960 1908 2962
rect 1648 2926 1720 2956
rect 1648 1378 1710 2926
rect 1826 1548 1908 2960
rect 2024 1690 2204 3050
rect 1824 1384 1908 1548
rect 2018 1488 2218 1690
rect 1352 1152 1416 1250
rect 1264 902 1274 1152
rect 1422 902 1432 1152
rect 1352 686 1400 902
rect 1460 732 1594 1322
rect 1824 924 1888 1384
rect 2024 1292 2204 1488
rect 2324 1380 2334 2958
rect 2412 1380 2422 2958
rect 2518 1378 2594 2962
rect 2734 1682 2898 3054
rect 3012 2956 3280 2958
rect 2716 1482 2916 1682
rect 2520 1054 2572 1378
rect 2734 1290 2898 1482
rect 3012 1388 3024 2956
rect 3114 1388 3280 2956
rect 3012 1384 3280 1388
rect 3350 2934 3434 3052
rect 3616 2958 3638 3120
rect 3350 1324 3434 1460
rect 3500 1386 3638 2958
rect 3308 1104 3466 1324
rect 3616 1184 3638 1386
rect 2520 930 3244 1054
rect 3298 952 3308 1104
rect 3466 952 3476 1104
rect 1352 490 1414 686
rect 1354 -100 1414 490
rect 1482 -176 1570 732
rect 1648 228 1716 690
rect 1824 684 1890 924
rect 1980 684 2248 764
rect 1824 498 2248 684
rect 2520 692 2572 930
rect 3162 800 3242 930
rect 3630 886 3638 1184
rect 3830 2162 3844 3232
rect 3830 1962 3842 2162
rect 3630 828 3688 886
rect 3830 874 3844 1962
rect 3830 828 3842 874
rect 3630 820 3842 828
rect 3442 800 3592 802
rect 3162 790 3592 800
rect 3162 782 3628 790
rect 2520 682 2592 692
rect 2662 682 2936 764
rect 3162 732 3874 782
rect 3162 730 3424 732
rect 3604 714 3874 732
rect 1648 -108 1734 228
rect 1848 -96 2248 498
rect 1694 -232 1734 -108
rect 1980 -176 2248 -96
rect 2330 238 2410 682
rect 2520 624 2936 682
rect 3184 680 3364 682
rect 2330 140 2420 238
rect 2330 6 2438 140
rect 2330 -44 2450 6
rect 2330 -50 2460 -44
rect 2330 -100 2360 -50
rect 2412 -124 2460 -50
rect 2522 -96 2936 624
rect 3018 656 3034 678
rect 3098 656 3364 680
rect 3018 652 3364 656
rect 3018 -58 3134 652
rect 3264 506 3364 652
rect 3418 654 3498 682
rect 3418 508 3810 654
rect 3418 506 3498 508
rect 3264 414 3278 506
rect 3264 360 3498 414
rect 3264 352 3440 360
rect 3264 2 3276 352
rect 3532 316 3808 508
rect 3532 290 3812 316
rect 3388 90 3812 290
rect 3532 84 3812 90
rect 3766 82 3812 84
rect 3264 -10 3546 2
rect 3018 -94 3032 -58
rect 2522 -100 2592 -96
rect 2396 -172 2460 -124
rect 2388 -232 2460 -172
rect 2662 -176 2936 -96
rect 3128 -232 3134 -58
rect 1274 -256 3134 -232
rect 1274 -346 1282 -256
rect 1268 -378 1282 -346
rect 3532 -378 3546 -10
rect 1268 -382 3546 -378
rect 1268 -398 3544 -382
<< rmetal1 >>
rect 3350 1460 3434 2934
<< via1 >>
rect 1274 902 1422 1152
rect 2334 1380 2412 2958
rect 3024 1388 3114 2956
rect 3308 952 3466 1104
<< metal2 >>
rect 2334 2958 2412 2968
rect 3024 2956 3114 2966
rect 2412 1878 3024 2410
rect 2334 1370 2412 1380
rect 3024 1378 3114 1388
rect 1274 1152 1422 1162
rect 1272 960 1274 1100
rect 3308 1104 3466 1114
rect 1422 960 3308 1100
rect 3308 942 3466 952
rect 1274 892 1422 902
use sky130_fd_pr__nfet_01v8_64Z3AY  XM1
timestamp 1730493024
transform 1 0 3401 0 1 625
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_3H2EVM  XM3
timestamp 1730493024
transform 1 0 1526 0 1 2167
box -296 -1019 296 1019
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XM4
timestamp 1730493024
transform 1 0 1528 0 1 292
box -296 -610 296 610
use sky130_fd_pr__nfet_01v8_lvt_AHRV9L  XM5
timestamp 1730493024
transform 1 0 2114 0 1 292
box -396 -610 396 610
use sky130_fd_pr__nfet_01v8_lvt_AHRV9L  XM6
timestamp 1730493024
transform 1 0 2800 0 1 292
box -396 -610 396 610
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM7
timestamp 1730493024
transform 1 0 2112 0 1 2167
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_3H2EVM  XM8
timestamp 1730493024
transform 1 0 3384 0 1 2167
box -296 -1019 296 1019
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM9
timestamp 1730493024
transform 1 0 2798 0 1 2167
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_MGSNAN  XM21
timestamp 1730493024
transform 1 0 3823 0 1 408
box -211 -484 211 484
<< labels >>
flabel metal1 3388 90 3588 290 0 FreeSans 256 0 0 0 out
port 0 nsew
flabel metal1 2716 1482 2916 1682 0 FreeSans 256 0 0 0 in+
port 2 nsew
flabel metal1 3626 1964 3826 2164 0 FreeSans 256 0 0 0 vdd
port 1 nsew
flabel metal1 3212 -288 3412 -88 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 2018 1490 2218 1690 0 FreeSans 256 0 0 0 in-
port 3 nsew
<< end >>
