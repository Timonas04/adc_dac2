magic
tech sky130A
magscale 1 2
timestamp 1730493024
<< error_p >>
rect -125 172 -67 178
rect 67 172 125 178
rect -125 138 -113 172
rect 67 138 79 172
rect -125 132 -67 138
rect 67 132 125 138
rect -221 -138 -163 -132
rect -29 -138 29 -132
rect 163 -138 221 -132
rect -221 -172 -209 -138
rect -29 -172 -17 -138
rect 163 -172 175 -138
rect -221 -178 -163 -172
rect -29 -178 29 -172
rect 163 -178 221 -172
<< pwell >>
rect -407 -310 407 310
<< nmos >>
rect -207 -100 -177 100
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
rect 177 -100 207 100
<< ndiff >>
rect -269 88 -207 100
rect -269 -88 -257 88
rect -223 -88 -207 88
rect -269 -100 -207 -88
rect -177 88 -111 100
rect -177 -88 -161 88
rect -127 -88 -111 88
rect -177 -100 -111 -88
rect -81 88 -15 100
rect -81 -88 -65 88
rect -31 -88 -15 88
rect -81 -100 -15 -88
rect 15 88 81 100
rect 15 -88 31 88
rect 65 -88 81 88
rect 15 -100 81 -88
rect 111 88 177 100
rect 111 -88 127 88
rect 161 -88 177 88
rect 111 -100 177 -88
rect 207 88 269 100
rect 207 -88 223 88
rect 257 -88 269 88
rect 207 -100 269 -88
<< ndiffc >>
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
<< psubdiff >>
rect -371 240 -275 274
rect 275 240 371 274
rect -371 178 -337 240
rect 337 178 371 240
rect -371 -240 -337 -178
rect 337 -240 371 -178
rect -371 -274 -275 -240
rect 275 -274 371 -240
<< psubdiffcont >>
rect -275 240 275 274
rect -371 -178 -337 178
rect 337 -178 371 178
rect -275 -274 275 -240
<< poly >>
rect -129 172 -63 188
rect -129 138 -113 172
rect -79 138 -63 172
rect -207 100 -177 126
rect -129 122 -63 138
rect 63 172 129 188
rect 63 138 79 172
rect 113 138 129 172
rect -111 100 -81 122
rect -15 100 15 126
rect 63 122 129 138
rect 81 100 111 122
rect 177 100 207 126
rect -207 -122 -177 -100
rect -225 -138 -159 -122
rect -111 -126 -81 -100
rect -15 -122 15 -100
rect -225 -172 -209 -138
rect -175 -172 -159 -138
rect -225 -188 -159 -172
rect -33 -138 33 -122
rect 81 -126 111 -100
rect 177 -122 207 -100
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
rect 159 -138 225 -122
rect 159 -172 175 -138
rect 209 -172 225 -138
rect 159 -188 225 -172
<< polycont >>
rect -113 138 -79 172
rect 79 138 113 172
rect -209 -172 -175 -138
rect -17 -172 17 -138
rect 175 -172 209 -138
<< locali >>
rect -371 240 -275 274
rect 275 240 371 274
rect -371 178 -337 240
rect 337 178 371 240
rect -129 138 -113 172
rect -79 138 -63 172
rect 63 138 79 172
rect 113 138 129 172
rect -257 88 -223 104
rect -257 -104 -223 -88
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect 223 88 257 104
rect 223 -104 257 -88
rect -225 -172 -209 -138
rect -175 -172 -159 -138
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect 159 -172 175 -138
rect 209 -172 225 -138
rect -371 -240 -337 -178
rect 337 -240 371 -178
rect -371 -274 -275 -240
rect 275 -274 371 -240
<< viali >>
rect -113 138 -79 172
rect 79 138 113 172
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect -209 -172 -175 -138
rect -17 -172 17 -138
rect 175 -172 209 -138
<< metal1 >>
rect -125 172 -67 178
rect -125 138 -113 172
rect -79 138 -67 172
rect -125 132 -67 138
rect 67 172 125 178
rect 67 138 79 172
rect 113 138 125 172
rect 67 132 125 138
rect -263 88 -217 100
rect -263 -88 -257 88
rect -223 -88 -217 88
rect -263 -100 -217 -88
rect -167 88 -121 100
rect -167 -88 -161 88
rect -127 -88 -121 88
rect -167 -100 -121 -88
rect -71 88 -25 100
rect -71 -88 -65 88
rect -31 -88 -25 88
rect -71 -100 -25 -88
rect 25 88 71 100
rect 25 -88 31 88
rect 65 -88 71 88
rect 25 -100 71 -88
rect 121 88 167 100
rect 121 -88 127 88
rect 161 -88 167 88
rect 121 -100 167 -88
rect 217 88 263 100
rect 217 -88 223 88
rect 257 -88 263 88
rect 217 -100 263 -88
rect -221 -138 -163 -132
rect -221 -172 -209 -138
rect -175 -172 -163 -138
rect -221 -178 -163 -172
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
rect 163 -138 221 -132
rect 163 -172 175 -138
rect 209 -172 221 -138
rect 163 -178 221 -172
<< properties >>
string FIXED_BBOX -354 -257 354 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
