MACRO main
  CLASS BLOCK ;
  FOREIGN main ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 210.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 198.800 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 198.800 ;
    END
  END VPWR
  PIN b0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 206.000 55.110 210.000 ;
    END
  END b0
  PIN b1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 206.000 64.770 210.000 ;
    END
  END b1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END clk
  PIN compr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 68.040 90.000 68.640 ;
    END
  END compr
  PIN dac[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 112.240 90.000 112.840 ;
    END
  END dac[0]
  PIN dac[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 78.240 90.000 78.840 ;
    END
  END dac[1]
  PIN dac[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 71.440 90.000 72.040 ;
    END
  END dac[2]
  PIN dac[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 57.840 90.000 58.440 ;
    END
  END dac[3]
  PIN dac[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 61.240 90.000 61.840 ;
    END
  END dac[4]
  PIN dac[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 64.640 90.000 65.240 ;
    END
  END dac[5]
  PIN dac[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 85.040 90.000 85.640 ;
    END
  END dac[6]
  PIN dac[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 108.840 90.000 109.440 ;
    END
  END dac[7]
  PIN dac_coupl
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END dac_coupl
  PIN m0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END m0
  PIN m1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END m1
  PIN reg0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END reg0[0]
  PIN reg0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END reg0[1]
  PIN reg0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END reg0[2]
  PIN reg0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END reg0[3]
  PIN reg0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END reg0[4]
  PIN reg0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END reg0[5]
  PIN reg0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END reg0[6]
  PIN reg0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END reg0[7]
  PIN reg1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END reg1[0]
  PIN reg1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END reg1[1]
  PIN reg1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END reg1[2]
  PIN reg1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END reg1[3]
  PIN reg1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END reg1[4]
  PIN reg1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END reg1[5]
  PIN reg1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END reg1[6]
  PIN reg1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END reg1[7]
  PIN reg2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END reg2[0]
  PIN reg2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END reg2[1]
  PIN reg2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END reg2[2]
  PIN reg2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END reg2[3]
  PIN reg2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END reg2[4]
  PIN reg2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END reg2[5]
  PIN reg2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END reg2[6]
  PIN reg2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END reg2[7]
  PIN reg3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END reg3[0]
  PIN reg3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END reg3[1]
  PIN reg3[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END reg3[2]
  PIN reg3[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END reg3[3]
  PIN reg3[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END reg3[4]
  PIN reg3[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 27.240 90.000 27.840 ;
    END
  END reg3[5]
  PIN reg3[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 51.040 90.000 51.640 ;
    END
  END reg3[6]
  PIN reg3[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 40.840 90.000 41.440 ;
    END
  END reg3[7]
  PIN reg4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END reg4[0]
  PIN reg4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END reg4[1]
  PIN reg4[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END reg4[2]
  PIN reg4[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END reg4[3]
  PIN reg4[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END reg4[4]
  PIN reg4[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END reg4[5]
  PIN reg4[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END reg4[6]
  PIN reg4[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END reg4[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END rst
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END rx
  PIN tx
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END tx
  OBS
      LAYER nwell ;
        RECT 5.330 197.145 84.370 198.750 ;
      LAYER pwell ;
        RECT 5.525 195.945 6.895 196.755 ;
        RECT 6.905 195.945 12.415 196.755 ;
        RECT 12.425 195.945 17.935 196.755 ;
        RECT 18.415 196.030 18.845 196.815 ;
        RECT 18.865 195.945 24.375 196.755 ;
        RECT 24.385 195.945 29.895 196.755 ;
        RECT 29.905 195.945 31.275 196.755 ;
        RECT 31.295 196.030 31.725 196.815 ;
        RECT 31.745 195.945 37.255 196.755 ;
        RECT 37.265 195.945 42.775 196.755 ;
        RECT 42.785 195.945 44.155 196.755 ;
        RECT 44.175 196.030 44.605 196.815 ;
        RECT 44.625 195.945 50.135 196.755 ;
        RECT 50.145 196.625 51.065 196.855 ;
        RECT 50.145 195.945 52.435 196.625 ;
        RECT 52.445 195.945 55.195 196.755 ;
        RECT 55.205 195.945 56.575 196.725 ;
        RECT 57.055 196.030 57.485 196.815 ;
        RECT 57.505 195.945 63.015 196.755 ;
        RECT 63.025 195.945 64.855 196.755 ;
        RECT 64.865 195.945 66.235 196.725 ;
        RECT 66.245 195.945 69.915 196.755 ;
        RECT 69.935 196.030 70.365 196.815 ;
        RECT 70.385 195.945 75.895 196.755 ;
        RECT 75.905 195.945 81.415 196.755 ;
        RECT 81.425 195.945 82.795 196.755 ;
        RECT 82.805 195.945 84.175 196.755 ;
        RECT 5.665 195.735 5.835 195.945 ;
        RECT 7.045 195.735 7.215 195.945 ;
        RECT 12.565 195.735 12.735 195.945 ;
        RECT 18.085 195.895 18.255 195.925 ;
        RECT 18.080 195.785 18.255 195.895 ;
        RECT 18.085 195.735 18.255 195.785 ;
        RECT 19.005 195.755 19.175 195.945 ;
        RECT 23.605 195.735 23.775 195.925 ;
        RECT 24.525 195.755 24.695 195.945 ;
        RECT 29.125 195.735 29.295 195.925 ;
        RECT 30.045 195.755 30.215 195.945 ;
        RECT 30.960 195.785 31.080 195.895 ;
        RECT 31.885 195.735 32.055 195.945 ;
        RECT 35.560 195.735 35.730 195.925 ;
        RECT 36.025 195.735 36.195 195.925 ;
        RECT 37.405 195.755 37.575 195.945 ;
        RECT 38.325 195.735 38.495 195.925 ;
        RECT 42.925 195.755 43.095 195.945 ;
        RECT 44.765 195.755 44.935 195.945 ;
        RECT 45.685 195.735 45.855 195.925 ;
        RECT 49.365 195.735 49.535 195.925 ;
        RECT 52.125 195.755 52.295 195.945 ;
        RECT 52.585 195.755 52.755 195.945 ;
        RECT 55.345 195.755 55.515 195.945 ;
        RECT 56.720 195.785 56.840 195.895 ;
        RECT 57.645 195.735 57.815 195.945 ;
        RECT 59.480 195.785 59.600 195.895 ;
        RECT 63.165 195.755 63.335 195.945 ;
        RECT 65.925 195.755 66.095 195.945 ;
        RECT 66.385 195.755 66.555 195.945 ;
        RECT 66.845 195.735 67.015 195.925 ;
        RECT 67.305 195.735 67.475 195.925 ;
        RECT 70.525 195.755 70.695 195.945 ;
        RECT 72.825 195.735 72.995 195.925 ;
        RECT 76.045 195.755 76.215 195.945 ;
        RECT 78.345 195.735 78.515 195.925 ;
        RECT 81.565 195.755 81.735 195.945 ;
        RECT 82.035 195.780 82.195 195.890 ;
        RECT 83.865 195.735 84.035 195.945 ;
        RECT 5.525 194.925 6.895 195.735 ;
        RECT 6.905 194.925 12.415 195.735 ;
        RECT 12.425 194.925 17.935 195.735 ;
        RECT 17.945 194.925 23.455 195.735 ;
        RECT 23.465 194.925 28.975 195.735 ;
        RECT 28.985 194.925 30.815 195.735 ;
        RECT 31.295 194.865 31.725 195.650 ;
        RECT 31.745 194.925 34.495 195.735 ;
        RECT 34.525 194.825 35.875 195.735 ;
        RECT 35.885 195.055 38.175 195.735 ;
        RECT 38.185 195.055 45.495 195.735 ;
        RECT 37.255 194.825 38.175 195.055 ;
        RECT 41.700 194.835 42.610 195.055 ;
        RECT 44.145 194.825 45.495 195.055 ;
        RECT 45.545 194.925 49.215 195.735 ;
        RECT 49.225 195.055 56.535 195.735 ;
        RECT 52.740 194.835 53.650 195.055 ;
        RECT 55.185 194.825 56.535 195.055 ;
        RECT 57.055 194.865 57.485 195.650 ;
        RECT 57.505 194.925 59.335 195.735 ;
        RECT 59.845 195.055 67.155 195.735 ;
        RECT 59.845 194.825 61.195 195.055 ;
        RECT 62.730 194.835 63.640 195.055 ;
        RECT 67.165 194.925 72.675 195.735 ;
        RECT 72.685 194.925 78.195 195.735 ;
        RECT 78.205 194.925 81.875 195.735 ;
        RECT 82.805 194.925 84.175 195.735 ;
      LAYER nwell ;
        RECT 5.330 191.705 84.370 194.535 ;
      LAYER pwell ;
        RECT 5.525 190.505 6.895 191.315 ;
        RECT 6.905 190.505 12.415 191.315 ;
        RECT 12.425 190.505 17.935 191.315 ;
        RECT 18.415 190.590 18.845 191.375 ;
        RECT 18.865 190.505 24.375 191.315 ;
        RECT 24.385 190.505 29.895 191.315 ;
        RECT 33.880 191.185 34.790 191.405 ;
        RECT 36.325 191.185 37.675 191.415 ;
        RECT 30.365 190.505 37.675 191.185 ;
        RECT 38.185 191.185 39.105 191.415 ;
        RECT 38.185 190.505 40.475 191.185 ;
        RECT 40.485 190.505 41.835 191.415 ;
        RECT 43.235 191.185 44.155 191.415 ;
        RECT 41.865 190.505 44.155 191.185 ;
        RECT 44.175 190.590 44.605 191.375 ;
        RECT 48.140 191.185 49.050 191.405 ;
        RECT 50.585 191.185 51.935 191.415 ;
        RECT 44.625 190.505 51.935 191.185 ;
        RECT 52.925 190.505 54.275 191.415 ;
        RECT 55.225 190.505 56.575 191.415 ;
        RECT 56.585 190.505 57.955 191.315 ;
        RECT 57.985 190.505 59.335 191.415 ;
        RECT 60.715 191.185 61.635 191.415 ;
        RECT 59.345 190.505 61.635 191.185 ;
        RECT 62.605 191.185 63.955 191.415 ;
        RECT 65.490 191.185 66.400 191.405 ;
        RECT 62.605 190.505 69.915 191.185 ;
        RECT 69.935 190.590 70.365 191.375 ;
        RECT 70.385 190.505 75.895 191.315 ;
        RECT 75.905 190.505 81.415 191.315 ;
        RECT 81.425 190.505 82.795 191.315 ;
        RECT 82.805 190.505 84.175 191.315 ;
        RECT 5.665 190.295 5.835 190.505 ;
        RECT 7.045 190.295 7.215 190.505 ;
        RECT 12.565 190.295 12.735 190.505 ;
        RECT 18.085 190.455 18.255 190.485 ;
        RECT 18.080 190.345 18.255 190.455 ;
        RECT 18.085 190.295 18.255 190.345 ;
        RECT 19.005 190.315 19.175 190.505 ;
        RECT 23.605 190.295 23.775 190.485 ;
        RECT 24.525 190.315 24.695 190.505 ;
        RECT 29.125 190.295 29.295 190.485 ;
        RECT 30.040 190.345 30.160 190.455 ;
        RECT 30.505 190.315 30.675 190.505 ;
        RECT 30.960 190.345 31.080 190.455 ;
        RECT 31.885 190.295 32.055 190.485 ;
        RECT 35.105 190.295 35.275 190.485 ;
        RECT 35.570 190.295 35.740 190.485 ;
        RECT 36.945 190.295 37.115 190.485 ;
        RECT 37.860 190.345 37.980 190.455 ;
        RECT 40.165 190.295 40.335 190.505 ;
        RECT 40.630 190.315 40.800 190.505 ;
        RECT 42.005 190.315 42.175 190.505 ;
        RECT 44.765 190.295 44.935 190.505 ;
        RECT 45.225 190.295 45.395 190.485 ;
        RECT 50.745 190.295 50.915 190.485 ;
        RECT 52.135 190.350 52.295 190.460 ;
        RECT 53.960 190.315 54.130 190.505 ;
        RECT 54.435 190.350 54.595 190.460 ;
        RECT 56.260 190.315 56.430 190.505 ;
        RECT 56.725 190.295 56.895 190.505 ;
        RECT 57.645 190.295 57.815 190.485 ;
        RECT 59.020 190.315 59.190 190.505 ;
        RECT 59.485 190.315 59.655 190.505 ;
        RECT 60.865 190.295 61.035 190.485 ;
        RECT 61.795 190.350 61.955 190.460 ;
        RECT 62.705 190.295 62.875 190.485 ;
        RECT 65.925 190.315 66.095 190.485 ;
        RECT 65.930 190.295 66.095 190.315 ;
        RECT 68.225 190.295 68.395 190.485 ;
        RECT 69.605 190.315 69.775 190.505 ;
        RECT 70.525 190.315 70.695 190.505 ;
        RECT 73.745 190.295 73.915 190.485 ;
        RECT 76.045 190.315 76.215 190.505 ;
        RECT 79.265 190.295 79.435 190.485 ;
        RECT 81.565 190.315 81.735 190.505 ;
        RECT 83.865 190.295 84.035 190.505 ;
        RECT 5.525 189.485 6.895 190.295 ;
        RECT 6.905 189.485 12.415 190.295 ;
        RECT 12.425 189.485 17.935 190.295 ;
        RECT 17.945 189.485 23.455 190.295 ;
        RECT 23.465 189.485 28.975 190.295 ;
        RECT 28.985 189.485 30.815 190.295 ;
        RECT 31.295 189.425 31.725 190.210 ;
        RECT 31.745 189.485 33.115 190.295 ;
        RECT 33.125 189.615 35.415 190.295 ;
        RECT 33.125 189.385 34.045 189.615 ;
        RECT 35.425 189.385 36.775 190.295 ;
        RECT 36.805 189.615 40.015 190.295 ;
        RECT 38.880 189.385 40.015 189.615 ;
        RECT 40.040 189.385 41.855 190.295 ;
        RECT 41.865 189.385 45.035 190.295 ;
        RECT 45.085 189.485 50.595 190.295 ;
        RECT 50.605 189.485 54.275 190.295 ;
        RECT 54.295 189.615 57.035 190.295 ;
        RECT 57.055 189.425 57.485 190.210 ;
        RECT 57.505 189.615 60.715 190.295 ;
        RECT 59.580 189.385 60.715 189.615 ;
        RECT 60.740 189.385 62.555 190.295 ;
        RECT 62.565 189.615 65.775 190.295 ;
        RECT 65.930 189.615 67.765 190.295 ;
        RECT 64.640 189.385 65.775 189.615 ;
        RECT 66.835 189.385 67.765 189.615 ;
        RECT 68.085 189.485 73.595 190.295 ;
        RECT 73.605 189.485 79.115 190.295 ;
        RECT 79.125 189.485 82.795 190.295 ;
        RECT 82.805 189.485 84.175 190.295 ;
      LAYER nwell ;
        RECT 5.330 186.265 84.370 189.095 ;
      LAYER pwell ;
        RECT 5.525 185.065 6.895 185.875 ;
        RECT 6.905 185.065 12.415 185.875 ;
        RECT 12.425 185.065 17.935 185.875 ;
        RECT 18.415 185.150 18.845 185.935 ;
        RECT 18.865 185.065 24.375 185.875 ;
        RECT 24.385 185.065 29.895 185.875 ;
        RECT 29.905 185.065 33.575 185.875 ;
        RECT 33.585 185.745 34.505 185.975 ;
        RECT 33.585 185.065 35.875 185.745 ;
        RECT 35.885 185.065 41.395 185.875 ;
        RECT 41.405 185.065 44.155 185.875 ;
        RECT 44.175 185.150 44.605 185.935 ;
        RECT 44.625 185.065 48.295 185.875 ;
        RECT 49.225 185.065 51.040 185.975 ;
        RECT 51.065 185.065 54.275 185.975 ;
        RECT 54.285 185.065 57.035 185.975 ;
        RECT 57.505 185.745 58.425 185.975 ;
        RECT 57.505 185.065 59.795 185.745 ;
        RECT 59.805 185.065 62.555 185.875 ;
        RECT 63.045 185.065 64.395 185.975 ;
        RECT 64.405 185.065 69.915 185.875 ;
        RECT 69.935 185.150 70.365 185.935 ;
        RECT 70.385 185.065 75.895 185.875 ;
        RECT 75.905 185.065 81.415 185.875 ;
        RECT 81.425 185.065 82.795 185.875 ;
        RECT 82.805 185.065 84.175 185.875 ;
        RECT 5.665 184.855 5.835 185.065 ;
        RECT 7.045 184.855 7.215 185.065 ;
        RECT 12.565 184.855 12.735 185.065 ;
        RECT 15.785 184.855 15.955 185.045 ;
        RECT 16.245 184.855 16.415 185.045 ;
        RECT 18.080 184.905 18.200 185.015 ;
        RECT 19.005 184.875 19.175 185.065 ;
        RECT 19.925 184.855 20.095 185.045 ;
        RECT 24.525 184.875 24.695 185.065 ;
        RECT 27.285 184.855 27.455 185.045 ;
        RECT 30.045 184.875 30.215 185.065 ;
        RECT 30.960 184.905 31.080 185.015 ;
        RECT 31.885 184.855 32.055 185.045 ;
        RECT 35.565 184.875 35.735 185.065 ;
        RECT 36.025 184.875 36.195 185.065 ;
        RECT 39.245 184.855 39.415 185.045 ;
        RECT 41.545 184.875 41.715 185.065 ;
        RECT 44.765 184.855 44.935 185.065 ;
        RECT 48.455 185.015 48.615 185.020 ;
        RECT 48.440 184.910 48.615 185.015 ;
        RECT 48.440 184.905 48.560 184.910 ;
        RECT 50.285 184.855 50.455 185.045 ;
        RECT 50.745 184.855 50.915 185.065 ;
        RECT 51.205 184.875 51.375 185.065 ;
        RECT 52.580 184.905 52.700 185.015 ;
        RECT 53.050 184.855 53.220 185.045 ;
        RECT 54.425 184.875 54.595 185.065 ;
        RECT 54.885 184.855 55.055 185.045 ;
        RECT 56.720 184.905 56.840 185.015 ;
        RECT 57.180 184.905 57.300 185.015 ;
        RECT 57.645 184.855 57.815 185.045 ;
        RECT 59.485 184.875 59.655 185.065 ;
        RECT 59.945 184.875 60.115 185.065 ;
        RECT 63.160 185.045 63.330 185.065 ;
        RECT 62.700 184.905 62.820 185.015 ;
        RECT 63.160 184.875 63.335 185.045 ;
        RECT 64.545 184.875 64.715 185.065 ;
        RECT 63.165 184.855 63.335 184.875 ;
        RECT 68.685 184.855 68.855 185.045 ;
        RECT 70.525 184.875 70.695 185.065 ;
        RECT 74.205 184.855 74.375 185.045 ;
        RECT 76.045 184.875 76.215 185.065 ;
        RECT 79.725 184.855 79.895 185.045 ;
        RECT 81.565 184.875 81.735 185.065 ;
        RECT 82.480 184.905 82.600 185.015 ;
        RECT 83.865 184.855 84.035 185.065 ;
        RECT 5.525 184.045 6.895 184.855 ;
        RECT 6.905 184.045 12.415 184.855 ;
        RECT 12.425 184.045 13.795 184.855 ;
        RECT 13.805 184.175 16.095 184.855 ;
        RECT 13.805 183.945 14.725 184.175 ;
        RECT 16.105 184.045 19.775 184.855 ;
        RECT 19.785 184.175 27.095 184.855 ;
        RECT 23.300 183.955 24.210 184.175 ;
        RECT 25.745 183.945 27.095 184.175 ;
        RECT 27.145 184.045 30.815 184.855 ;
        RECT 31.295 183.985 31.725 184.770 ;
        RECT 31.745 184.175 39.055 184.855 ;
        RECT 35.260 183.955 36.170 184.175 ;
        RECT 37.705 183.945 39.055 184.175 ;
        RECT 39.105 184.045 44.615 184.855 ;
        RECT 44.625 184.045 48.295 184.855 ;
        RECT 48.765 183.945 50.580 184.855 ;
        RECT 50.605 184.045 52.435 184.855 ;
        RECT 52.905 183.945 54.735 184.855 ;
        RECT 54.745 184.045 56.575 184.855 ;
        RECT 57.055 183.985 57.485 184.770 ;
        RECT 57.505 184.045 63.015 184.855 ;
        RECT 63.025 184.045 68.535 184.855 ;
        RECT 68.545 184.045 74.055 184.855 ;
        RECT 74.065 184.045 79.575 184.855 ;
        RECT 79.585 184.045 82.335 184.855 ;
        RECT 82.805 184.045 84.175 184.855 ;
      LAYER nwell ;
        RECT 5.330 180.825 84.370 183.655 ;
      LAYER pwell ;
        RECT 5.525 179.625 6.895 180.435 ;
        RECT 6.905 179.625 9.655 180.435 ;
        RECT 9.685 179.625 11.035 180.535 ;
        RECT 11.085 180.305 12.435 180.535 ;
        RECT 13.970 180.305 14.880 180.525 ;
        RECT 11.085 179.625 18.395 180.305 ;
        RECT 18.415 179.710 18.845 180.495 ;
        RECT 19.785 180.305 20.705 180.535 ;
        RECT 19.785 179.625 22.075 180.305 ;
        RECT 22.085 179.625 25.005 180.535 ;
        RECT 25.315 179.625 28.045 180.535 ;
        RECT 28.265 180.445 29.215 180.535 ;
        RECT 28.265 179.625 30.195 180.445 ;
        RECT 30.365 179.625 32.195 180.535 ;
        RECT 32.245 179.625 35.415 180.535 ;
        RECT 35.425 179.625 39.095 180.435 ;
        RECT 39.105 179.625 40.935 180.305 ;
        RECT 40.945 179.625 43.695 180.435 ;
        RECT 44.175 179.710 44.605 180.495 ;
        RECT 44.635 179.625 47.365 180.535 ;
        RECT 47.385 179.625 51.055 180.435 ;
        RECT 51.525 179.625 55.185 180.535 ;
        RECT 55.405 180.445 56.355 180.535 ;
        RECT 55.405 179.625 57.335 180.445 ;
        RECT 57.515 179.625 58.865 180.535 ;
        RECT 59.345 180.335 60.275 180.535 ;
        RECT 61.605 180.335 62.555 180.535 ;
        RECT 59.345 179.855 62.555 180.335 ;
        RECT 59.490 179.655 62.555 179.855 ;
        RECT 5.665 179.415 5.835 179.625 ;
        RECT 7.045 179.415 7.215 179.625 ;
        RECT 9.800 179.435 9.970 179.625 ;
        RECT 12.565 179.415 12.735 179.605 ;
        RECT 16.245 179.435 16.415 179.605 ;
        RECT 16.245 179.415 16.410 179.435 ;
        RECT 16.705 179.415 16.875 179.605 ;
        RECT 18.085 179.435 18.255 179.625 ;
        RECT 19.015 179.470 19.175 179.580 ;
        RECT 21.765 179.435 21.935 179.625 ;
        RECT 22.230 179.575 22.400 179.625 ;
        RECT 22.220 179.465 22.400 179.575 ;
        RECT 22.230 179.435 22.400 179.465 ;
        RECT 25.445 179.415 25.615 179.625 ;
        RECT 30.045 179.605 30.195 179.625 ;
        RECT 25.900 179.465 26.020 179.575 ;
        RECT 26.365 179.415 26.535 179.605 ;
        RECT 29.585 179.415 29.755 179.605 ;
        RECT 30.045 179.435 30.215 179.605 ;
        RECT 31.880 179.570 32.050 179.625 ;
        RECT 31.880 179.460 32.055 179.570 ;
        RECT 31.880 179.435 32.050 179.460 ;
        RECT 32.345 179.435 32.515 179.625 ;
        RECT 32.805 179.415 32.975 179.605 ;
        RECT 35.565 179.435 35.735 179.625 ;
        RECT 36.950 179.415 37.120 179.605 ;
        RECT 37.405 179.435 37.575 179.605 ;
        RECT 37.410 179.415 37.575 179.435 ;
        RECT 39.705 179.415 39.875 179.605 ;
        RECT 40.625 179.435 40.795 179.625 ;
        RECT 41.085 179.435 41.255 179.625 ;
        RECT 43.390 179.415 43.560 179.605 ;
        RECT 43.840 179.465 43.960 179.575 ;
        RECT 44.765 179.435 44.935 179.625 ;
        RECT 47.525 179.435 47.695 179.625 ;
        RECT 49.360 179.415 49.530 179.605 ;
        RECT 49.825 179.415 49.995 179.605 ;
        RECT 51.200 179.465 51.320 179.575 ;
        RECT 53.500 179.465 53.620 179.575 ;
        RECT 5.525 178.605 6.895 179.415 ;
        RECT 6.905 178.605 12.415 179.415 ;
        RECT 12.425 178.605 14.255 179.415 ;
        RECT 14.575 178.735 16.410 179.415 ;
        RECT 14.575 178.505 15.505 178.735 ;
        RECT 16.565 178.605 22.075 179.415 ;
        RECT 22.545 178.735 25.755 179.415 ;
        RECT 22.545 178.505 23.680 178.735 ;
        RECT 26.305 178.505 29.305 179.415 ;
        RECT 29.445 178.605 31.275 179.415 ;
        RECT 31.295 178.545 31.725 179.330 ;
        RECT 32.765 178.505 35.875 179.415 ;
        RECT 35.885 178.505 37.235 179.415 ;
        RECT 37.410 178.735 39.245 179.415 ;
        RECT 39.565 178.735 43.235 179.415 ;
        RECT 38.315 178.505 39.245 178.735 ;
        RECT 42.305 178.505 43.235 178.735 ;
        RECT 43.245 178.505 45.075 179.415 ;
        RECT 45.285 178.505 49.675 179.415 ;
        RECT 49.685 178.505 53.355 179.415 ;
        RECT 53.965 179.385 54.135 179.605 ;
        RECT 54.890 179.435 55.060 179.625 ;
        RECT 57.185 179.605 57.335 179.625 ;
        RECT 57.185 179.435 57.355 179.605 ;
        RECT 57.645 179.435 57.815 179.625 ;
        RECT 59.020 179.465 59.140 179.575 ;
        RECT 59.490 179.435 59.660 179.655 ;
        RECT 61.620 179.625 62.555 179.655 ;
        RECT 62.605 180.305 63.955 180.535 ;
        RECT 65.490 180.305 66.400 180.525 ;
        RECT 62.605 179.625 69.915 180.305 ;
        RECT 69.935 179.710 70.365 180.495 ;
        RECT 70.385 179.625 75.895 180.435 ;
        RECT 75.905 179.625 81.415 180.435 ;
        RECT 81.425 179.625 82.795 180.435 ;
        RECT 82.805 179.625 84.175 180.435 ;
        RECT 56.090 179.385 57.035 179.415 ;
        RECT 53.965 179.185 57.035 179.385 ;
        RECT 57.505 179.385 58.440 179.415 ;
        RECT 60.400 179.385 60.570 179.605 ;
        RECT 60.865 179.415 61.035 179.605 ;
        RECT 63.165 179.415 63.335 179.605 ;
        RECT 69.605 179.435 69.775 179.625 ;
        RECT 70.525 179.415 70.695 179.625 ;
        RECT 76.045 179.415 76.215 179.625 ;
        RECT 81.565 179.415 81.735 179.625 ;
        RECT 83.865 179.415 84.035 179.625 ;
        RECT 53.825 178.705 57.035 179.185 ;
        RECT 53.825 178.505 54.755 178.705 ;
        RECT 56.090 178.505 57.035 178.705 ;
        RECT 57.055 178.545 57.485 179.330 ;
        RECT 57.505 179.185 60.570 179.385 ;
        RECT 57.505 178.705 60.715 179.185 ;
        RECT 60.725 178.735 63.015 179.415 ;
        RECT 63.025 178.735 70.335 179.415 ;
        RECT 57.505 178.505 58.455 178.705 ;
        RECT 59.785 178.505 60.715 178.705 ;
        RECT 62.095 178.505 63.015 178.735 ;
        RECT 66.540 178.515 67.450 178.735 ;
        RECT 68.985 178.505 70.335 178.735 ;
        RECT 70.385 178.605 75.895 179.415 ;
        RECT 75.905 178.605 81.415 179.415 ;
        RECT 81.425 178.605 82.795 179.415 ;
        RECT 82.805 178.605 84.175 179.415 ;
      LAYER nwell ;
        RECT 5.330 175.385 84.370 178.215 ;
      LAYER pwell ;
        RECT 5.525 174.185 6.895 174.995 ;
        RECT 6.905 174.185 10.575 174.995 ;
        RECT 11.085 174.865 12.435 175.095 ;
        RECT 13.970 174.865 14.880 175.085 ;
        RECT 11.085 174.185 18.395 174.865 ;
        RECT 18.415 174.270 18.845 175.055 ;
        RECT 18.865 174.895 19.795 175.095 ;
        RECT 21.125 174.895 22.075 175.095 ;
        RECT 18.865 174.415 22.075 174.895 ;
        RECT 25.600 174.865 26.510 175.085 ;
        RECT 28.045 174.865 29.395 175.095 ;
        RECT 19.010 174.215 22.075 174.415 ;
        RECT 5.665 173.975 5.835 174.185 ;
        RECT 7.045 173.975 7.215 174.185 ;
        RECT 10.720 174.025 10.840 174.135 ;
        RECT 12.560 174.025 12.680 174.135 ;
        RECT 13.025 173.975 13.195 174.165 ;
        RECT 15.785 173.975 15.955 174.165 ;
        RECT 18.085 173.995 18.255 174.185 ;
        RECT 19.010 173.995 19.180 174.215 ;
        RECT 21.140 174.185 22.075 174.215 ;
        RECT 22.085 174.185 29.395 174.865 ;
        RECT 29.905 174.865 30.835 175.095 ;
        RECT 29.905 174.185 32.655 174.865 ;
        RECT 32.665 174.185 38.175 174.995 ;
        RECT 39.235 174.865 40.165 175.095 ;
        RECT 42.750 174.895 43.695 175.095 ;
        RECT 38.330 174.185 40.165 174.865 ;
        RECT 40.945 174.215 43.695 174.895 ;
        RECT 44.175 174.270 44.605 175.055 ;
        RECT 21.305 173.975 21.475 174.165 ;
        RECT 22.225 173.995 22.395 174.185 ;
        RECT 26.825 173.975 26.995 174.165 ;
        RECT 29.580 174.025 29.700 174.135 ;
        RECT 30.515 174.020 30.675 174.130 ;
        RECT 31.885 173.975 32.055 174.165 ;
        RECT 32.345 173.995 32.515 174.185 ;
        RECT 32.805 173.995 32.975 174.185 ;
        RECT 38.330 174.165 38.495 174.185 ;
        RECT 35.565 173.975 35.735 174.165 ;
        RECT 36.950 173.975 37.120 174.165 ;
        RECT 38.325 173.975 38.495 174.165 ;
        RECT 40.620 174.025 40.740 174.135 ;
        RECT 41.090 173.995 41.260 174.215 ;
        RECT 42.750 174.185 43.695 174.215 ;
        RECT 44.625 174.185 47.835 175.095 ;
        RECT 48.305 174.185 49.655 175.095 ;
        RECT 49.685 174.865 50.605 175.095 ;
        RECT 49.685 174.185 51.975 174.865 ;
        RECT 52.045 174.185 53.815 175.095 ;
        RECT 54.745 174.185 58.220 175.095 ;
        RECT 58.425 174.185 62.095 174.995 ;
        RECT 62.125 174.185 63.475 175.095 ;
        RECT 63.485 174.185 64.835 175.095 ;
        RECT 64.865 174.185 68.535 174.995 ;
        RECT 68.545 174.185 69.915 174.995 ;
        RECT 69.935 174.270 70.365 175.055 ;
        RECT 70.385 174.185 75.895 174.995 ;
        RECT 75.905 174.185 81.415 174.995 ;
        RECT 81.425 174.185 82.795 174.995 ;
        RECT 82.805 174.185 84.175 174.995 ;
        RECT 43.845 174.135 44.015 174.165 ;
        RECT 43.840 174.025 44.015 174.135 ;
        RECT 43.845 173.975 44.015 174.025 ;
        RECT 44.765 173.995 44.935 174.185 ;
        RECT 49.370 174.165 49.540 174.185 ;
        RECT 47.980 174.025 48.100 174.135 ;
        RECT 49.365 173.995 49.540 174.165 ;
        RECT 51.665 173.995 51.835 174.185 ;
        RECT 53.500 173.995 53.670 174.185 ;
        RECT 54.890 174.165 55.060 174.185 ;
        RECT 53.975 174.030 54.135 174.140 ;
        RECT 54.885 173.995 55.060 174.165 ;
        RECT 56.720 174.025 56.840 174.135 ;
        RECT 49.365 173.975 49.535 173.995 ;
        RECT 54.885 173.975 55.055 173.995 ;
        RECT 57.645 173.975 57.815 174.165 ;
        RECT 58.565 173.995 58.735 174.185 ;
        RECT 61.325 173.975 61.495 174.165 ;
        RECT 61.795 174.020 61.955 174.130 ;
        RECT 62.710 173.975 62.880 174.165 ;
        RECT 63.160 173.995 63.330 174.185 ;
        RECT 63.630 173.995 63.800 174.185 ;
        RECT 65.005 174.165 65.175 174.185 ;
        RECT 65.000 173.995 65.175 174.165 ;
        RECT 65.000 173.975 65.170 173.995 ;
        RECT 66.390 173.975 66.560 174.165 ;
        RECT 66.845 173.975 67.015 174.165 ;
        RECT 68.685 173.995 68.855 174.185 ;
        RECT 70.525 173.995 70.695 174.185 ;
        RECT 72.365 173.975 72.535 174.165 ;
        RECT 76.045 173.995 76.215 174.185 ;
        RECT 77.885 173.975 78.055 174.165 ;
        RECT 81.565 173.975 81.735 174.185 ;
        RECT 83.865 173.975 84.035 174.185 ;
        RECT 5.525 173.165 6.895 173.975 ;
        RECT 6.905 173.165 12.415 173.975 ;
        RECT 12.885 173.295 15.635 173.975 ;
        RECT 14.705 173.065 15.635 173.295 ;
        RECT 15.645 173.165 21.155 173.975 ;
        RECT 21.165 173.165 26.675 173.975 ;
        RECT 26.685 173.165 30.355 173.975 ;
        RECT 31.295 173.105 31.725 173.890 ;
        RECT 31.745 173.165 35.415 173.975 ;
        RECT 35.425 173.165 36.795 173.975 ;
        RECT 36.805 173.065 38.155 173.975 ;
        RECT 38.185 173.165 43.695 173.975 ;
        RECT 43.705 173.165 49.215 173.975 ;
        RECT 49.225 173.165 54.735 173.975 ;
        RECT 54.745 173.165 56.575 173.975 ;
        RECT 57.055 173.105 57.485 173.890 ;
        RECT 57.505 173.165 60.255 173.975 ;
        RECT 60.275 173.065 61.625 173.975 ;
        RECT 62.565 173.065 63.915 173.975 ;
        RECT 63.965 173.065 65.315 173.975 ;
        RECT 65.325 173.065 66.675 173.975 ;
        RECT 66.705 173.165 72.215 173.975 ;
        RECT 72.225 173.165 77.735 173.975 ;
        RECT 77.745 173.165 81.415 173.975 ;
        RECT 81.425 173.165 82.795 173.975 ;
        RECT 82.805 173.165 84.175 173.975 ;
      LAYER nwell ;
        RECT 5.330 169.945 84.370 172.775 ;
      LAYER pwell ;
        RECT 5.525 168.745 6.895 169.555 ;
        RECT 6.905 168.745 12.415 169.555 ;
        RECT 12.425 168.745 17.935 169.555 ;
        RECT 18.415 168.830 18.845 169.615 ;
        RECT 18.865 168.745 21.615 169.555 ;
        RECT 23.455 169.425 24.375 169.655 ;
        RECT 22.085 168.745 24.375 169.425 ;
        RECT 24.385 169.425 25.305 169.655 ;
        RECT 24.385 168.745 26.675 169.425 ;
        RECT 26.685 168.745 29.435 169.555 ;
        RECT 34.965 169.425 35.885 169.655 ;
        RECT 37.265 169.425 38.185 169.655 ;
        RECT 30.140 168.745 34.955 169.425 ;
        RECT 34.965 168.745 37.255 169.425 ;
        RECT 37.265 168.745 39.555 169.425 ;
        RECT 39.565 168.745 41.380 169.655 ;
        RECT 41.405 168.745 44.155 169.555 ;
        RECT 44.175 168.830 44.605 169.615 ;
        RECT 44.625 168.745 46.455 169.425 ;
        RECT 46.465 168.745 48.295 169.425 ;
        RECT 48.305 168.745 49.675 169.555 ;
        RECT 49.705 168.745 51.055 169.655 ;
        RECT 51.065 168.745 54.275 169.655 ;
        RECT 54.740 168.975 56.575 169.655 ;
        RECT 54.740 168.745 56.430 168.975 ;
        RECT 56.585 168.745 58.415 169.555 ;
        RECT 58.885 169.425 60.020 169.655 ;
        RECT 62.305 169.565 63.255 169.655 ;
        RECT 58.885 168.745 62.095 169.425 ;
        RECT 62.305 168.745 64.235 169.565 ;
        RECT 66.480 169.425 67.615 169.655 ;
        RECT 64.405 168.745 67.615 169.425 ;
        RECT 67.935 169.425 68.865 169.655 ;
        RECT 67.935 168.745 69.770 169.425 ;
        RECT 69.935 168.830 70.365 169.615 ;
        RECT 73.900 169.425 74.810 169.645 ;
        RECT 76.345 169.425 77.695 169.655 ;
        RECT 70.385 168.745 77.695 169.425 ;
        RECT 77.745 168.745 81.415 169.555 ;
        RECT 81.425 168.745 82.795 169.555 ;
        RECT 82.805 168.745 84.175 169.555 ;
        RECT 5.665 168.535 5.835 168.745 ;
        RECT 7.045 168.535 7.215 168.745 ;
        RECT 12.565 168.535 12.735 168.745 ;
        RECT 14.405 168.535 14.575 168.725 ;
        RECT 18.080 168.585 18.200 168.695 ;
        RECT 19.005 168.555 19.175 168.745 ;
        RECT 21.760 168.535 21.930 168.725 ;
        RECT 22.225 168.555 22.395 168.745 ;
        RECT 23.145 168.535 23.315 168.725 ;
        RECT 26.365 168.555 26.535 168.745 ;
        RECT 26.825 168.555 26.995 168.745 ;
        RECT 29.580 168.585 29.700 168.695 ;
        RECT 30.515 168.580 30.675 168.690 ;
        RECT 31.885 168.535 32.055 168.725 ;
        RECT 34.645 168.555 34.815 168.745 ;
        RECT 36.945 168.555 37.115 168.745 ;
        RECT 39.245 168.555 39.415 168.745 ;
        RECT 41.085 168.555 41.255 168.745 ;
        RECT 41.545 168.555 41.715 168.745 ;
        RECT 42.005 168.535 42.175 168.725 ;
        RECT 44.765 168.555 44.935 168.745 ;
        RECT 47.985 168.555 48.155 168.745 ;
        RECT 48.445 168.555 48.615 168.745 ;
        RECT 50.740 168.555 50.910 168.745 ;
        RECT 51.205 168.535 51.375 168.725 ;
        RECT 51.675 168.580 51.835 168.690 ;
        RECT 53.965 168.535 54.135 168.745 ;
        RECT 54.425 168.535 54.595 168.725 ;
        RECT 56.260 168.555 56.430 168.745 ;
        RECT 56.725 168.555 56.895 168.745 ;
        RECT 57.650 168.535 57.820 168.725 ;
        RECT 58.560 168.585 58.680 168.695 ;
        RECT 61.325 168.535 61.495 168.725 ;
        RECT 61.785 168.555 61.955 168.745 ;
        RECT 64.085 168.725 64.235 168.745 ;
        RECT 64.085 168.555 64.255 168.725 ;
        RECT 64.545 168.555 64.715 168.745 ;
        RECT 69.605 168.725 69.770 168.745 ;
        RECT 69.605 168.555 69.775 168.725 ;
        RECT 70.065 168.535 70.235 168.725 ;
        RECT 70.525 168.535 70.695 168.745 ;
        RECT 76.045 168.535 76.215 168.725 ;
        RECT 77.885 168.555 78.055 168.745 ;
        RECT 81.565 168.535 81.735 168.745 ;
        RECT 83.865 168.535 84.035 168.745 ;
        RECT 5.525 167.725 6.895 168.535 ;
        RECT 6.905 167.725 12.415 168.535 ;
        RECT 12.425 167.725 14.255 168.535 ;
        RECT 14.265 167.855 21.575 168.535 ;
        RECT 17.780 167.635 18.690 167.855 ;
        RECT 20.225 167.625 21.575 167.855 ;
        RECT 21.645 167.625 22.995 168.535 ;
        RECT 23.005 167.855 30.315 168.535 ;
        RECT 26.520 167.635 27.430 167.855 ;
        RECT 28.965 167.625 30.315 167.855 ;
        RECT 31.295 167.665 31.725 168.450 ;
        RECT 31.800 167.625 41.820 168.535 ;
        RECT 41.865 167.855 49.175 168.535 ;
        RECT 45.380 167.635 46.290 167.855 ;
        RECT 47.825 167.625 49.175 167.855 ;
        RECT 49.225 167.625 51.515 168.535 ;
        RECT 52.445 167.855 54.275 168.535 ;
        RECT 52.445 167.625 53.790 167.855 ;
        RECT 54.285 167.725 57.035 168.535 ;
        RECT 57.055 167.665 57.485 168.450 ;
        RECT 57.505 167.855 61.175 168.535 ;
        RECT 57.505 167.625 58.430 167.855 ;
        RECT 61.185 167.725 63.015 168.535 ;
        RECT 63.065 167.855 70.375 168.535 ;
        RECT 63.065 167.625 64.415 167.855 ;
        RECT 65.950 167.635 66.860 167.855 ;
        RECT 70.385 167.725 75.895 168.535 ;
        RECT 75.905 167.725 81.415 168.535 ;
        RECT 81.425 167.725 82.795 168.535 ;
        RECT 82.805 167.725 84.175 168.535 ;
      LAYER nwell ;
        RECT 5.330 164.505 84.370 167.335 ;
      LAYER pwell ;
        RECT 5.525 163.305 6.895 164.115 ;
        RECT 6.905 163.305 12.415 164.115 ;
        RECT 12.425 163.305 14.255 164.115 ;
        RECT 14.725 164.015 15.675 164.215 ;
        RECT 17.005 164.015 17.935 164.215 ;
        RECT 14.725 163.535 17.935 164.015 ;
        RECT 14.725 163.335 17.790 163.535 ;
        RECT 18.415 163.390 18.845 164.175 ;
        RECT 14.725 163.305 15.660 163.335 ;
        RECT 5.665 163.095 5.835 163.305 ;
        RECT 7.045 163.095 7.215 163.305 ;
        RECT 12.565 163.095 12.735 163.305 ;
        RECT 14.400 163.145 14.520 163.255 ;
        RECT 16.245 163.115 16.415 163.285 ;
        RECT 17.620 163.115 17.790 163.335 ;
        RECT 18.875 163.305 21.605 164.215 ;
        RECT 21.790 163.305 25.660 164.215 ;
        RECT 25.765 163.305 27.595 164.115 ;
        RECT 28.655 163.985 29.585 164.215 ;
        RECT 27.750 163.305 29.585 163.985 ;
        RECT 29.955 163.305 33.115 164.215 ;
        RECT 36.640 163.985 37.550 164.205 ;
        RECT 39.085 163.985 40.435 164.215 ;
        RECT 33.125 163.305 40.435 163.985 ;
        RECT 40.680 163.305 44.155 164.215 ;
        RECT 44.175 163.390 44.605 164.175 ;
        RECT 44.645 163.305 45.995 164.215 ;
        RECT 46.015 163.305 47.365 164.215 ;
        RECT 49.205 163.985 50.135 164.215 ;
        RECT 47.385 163.305 50.135 163.985 ;
        RECT 50.145 163.305 54.960 163.985 ;
        RECT 55.245 163.305 58.415 164.215 ;
        RECT 58.425 163.305 60.255 164.115 ;
        RECT 60.775 163.305 63.935 164.215 ;
        RECT 63.945 163.985 64.865 164.215 ;
        RECT 63.945 163.305 66.235 163.985 ;
        RECT 66.245 163.305 69.915 164.115 ;
        RECT 69.935 163.390 70.365 164.175 ;
        RECT 70.385 163.305 75.895 164.115 ;
        RECT 75.905 163.305 81.415 164.115 ;
        RECT 81.425 163.305 82.795 164.115 ;
        RECT 82.805 163.305 84.175 164.115 ;
        RECT 18.080 163.145 18.200 163.255 ;
        RECT 19.005 163.115 19.175 163.305 ;
        RECT 21.790 163.285 21.935 163.305 ;
        RECT 16.250 163.095 16.415 163.115 ;
        RECT 21.305 163.095 21.475 163.285 ;
        RECT 21.765 163.115 21.935 163.285 ;
        RECT 25.905 163.115 26.075 163.305 ;
        RECT 27.750 163.285 27.915 163.305 ;
        RECT 26.365 163.095 26.535 163.285 ;
        RECT 26.825 163.095 26.995 163.285 ;
        RECT 27.745 163.115 27.915 163.285 ;
        RECT 29.585 163.095 29.755 163.285 ;
        RECT 30.045 163.115 30.215 163.305 ;
        RECT 31.885 163.095 32.055 163.285 ;
        RECT 33.265 163.115 33.435 163.305 ;
        RECT 37.405 163.095 37.575 163.285 ;
        RECT 42.925 163.095 43.095 163.285 ;
        RECT 43.840 163.115 44.010 163.305 ;
        RECT 44.760 163.115 44.930 163.305 ;
        RECT 46.145 163.115 46.315 163.305 ;
        RECT 47.525 163.115 47.695 163.305 ;
        RECT 48.445 163.095 48.615 163.285 ;
        RECT 50.285 163.115 50.455 163.305 ;
        RECT 54.420 163.145 54.540 163.255 ;
        RECT 50.310 163.095 50.455 163.115 ;
        RECT 54.890 163.095 55.060 163.285 ;
        RECT 55.345 163.115 55.515 163.305 ;
        RECT 57.645 163.095 57.815 163.285 ;
        RECT 58.565 163.115 58.735 163.305 ;
        RECT 60.400 163.145 60.520 163.255 ;
        RECT 60.865 163.095 61.035 163.305 ;
        RECT 65.925 163.095 66.095 163.305 ;
        RECT 66.385 163.115 66.555 163.305 ;
        RECT 70.525 163.115 70.695 163.305 ;
        RECT 71.445 163.095 71.615 163.285 ;
        RECT 76.045 163.115 76.215 163.305 ;
        RECT 76.965 163.095 77.135 163.285 ;
        RECT 81.565 163.115 81.735 163.305 ;
        RECT 82.480 163.145 82.600 163.255 ;
        RECT 83.865 163.095 84.035 163.305 ;
        RECT 5.525 162.285 6.895 163.095 ;
        RECT 6.905 162.285 12.415 163.095 ;
        RECT 12.425 162.285 16.095 163.095 ;
        RECT 16.250 162.415 18.085 163.095 ;
        RECT 17.155 162.185 18.085 162.415 ;
        RECT 18.405 162.415 21.615 163.095 ;
        RECT 21.860 162.415 26.675 163.095 ;
        RECT 18.405 162.185 19.540 162.415 ;
        RECT 26.695 162.185 29.425 163.095 ;
        RECT 29.445 162.285 31.275 163.095 ;
        RECT 31.295 162.225 31.725 163.010 ;
        RECT 31.745 162.285 37.255 163.095 ;
        RECT 37.265 162.285 42.775 163.095 ;
        RECT 42.785 162.285 48.295 163.095 ;
        RECT 48.305 162.285 50.135 163.095 ;
        RECT 50.310 162.185 54.180 163.095 ;
        RECT 54.890 162.865 56.580 163.095 ;
        RECT 54.745 162.185 56.580 162.865 ;
        RECT 57.055 162.225 57.485 163.010 ;
        RECT 57.505 162.415 60.245 163.095 ;
        RECT 60.725 162.415 65.540 163.095 ;
        RECT 65.785 162.285 71.295 163.095 ;
        RECT 71.305 162.285 76.815 163.095 ;
        RECT 76.825 162.285 82.335 163.095 ;
        RECT 82.805 162.285 84.175 163.095 ;
      LAYER nwell ;
        RECT 5.330 159.065 84.370 161.895 ;
      LAYER pwell ;
        RECT 5.525 157.865 6.895 158.675 ;
        RECT 6.905 157.865 12.415 158.675 ;
        RECT 12.425 157.865 17.935 158.675 ;
        RECT 18.415 157.950 18.845 158.735 ;
        RECT 18.865 158.575 19.795 158.775 ;
        RECT 21.125 158.575 22.075 158.775 ;
        RECT 18.865 158.095 22.075 158.575 ;
        RECT 23.135 158.545 24.065 158.775 ;
        RECT 19.010 157.895 22.075 158.095 ;
        RECT 5.665 157.655 5.835 157.865 ;
        RECT 7.045 157.655 7.215 157.865 ;
        RECT 12.565 157.655 12.735 157.865 ;
        RECT 16.240 157.705 16.360 157.815 ;
        RECT 18.080 157.705 18.200 157.815 ;
        RECT 19.010 157.675 19.180 157.895 ;
        RECT 21.140 157.865 22.075 157.895 ;
        RECT 22.230 157.865 24.065 158.545 ;
        RECT 24.995 157.865 28.650 158.775 ;
        RECT 28.985 157.865 31.735 158.775 ;
        RECT 32.665 157.865 35.775 158.775 ;
        RECT 35.885 157.865 38.635 158.675 ;
        RECT 39.105 157.865 40.935 158.545 ;
        RECT 40.945 157.865 43.865 158.775 ;
        RECT 44.175 157.950 44.605 158.735 ;
        RECT 44.625 157.865 45.995 158.675 ;
        RECT 46.315 158.545 47.245 158.775 ;
        RECT 48.790 158.545 50.135 158.775 ;
        RECT 46.315 157.865 48.150 158.545 ;
        RECT 48.305 157.865 50.135 158.545 ;
        RECT 51.085 157.865 52.435 158.775 ;
        RECT 52.445 157.865 55.655 158.775 ;
        RECT 56.120 158.095 57.955 158.775 ;
        RECT 56.120 157.865 57.810 158.095 ;
        RECT 57.965 157.865 59.795 158.675 ;
        RECT 59.845 157.865 63.015 158.775 ;
        RECT 65.765 158.545 66.695 158.775 ;
        RECT 63.025 157.865 66.695 158.545 ;
        RECT 66.705 157.865 69.455 158.675 ;
        RECT 69.935 157.950 70.365 158.735 ;
        RECT 70.385 157.865 75.895 158.675 ;
        RECT 75.905 157.865 81.415 158.675 ;
        RECT 81.425 157.865 82.795 158.675 ;
        RECT 82.805 157.865 84.175 158.675 ;
        RECT 22.230 157.845 22.395 157.865 ;
        RECT 24.995 157.845 25.155 157.865 ;
        RECT 22.225 157.675 22.395 157.845 ;
        RECT 23.605 157.655 23.775 157.845 ;
        RECT 24.075 157.700 24.235 157.810 ;
        RECT 24.520 157.705 24.640 157.815 ;
        RECT 24.985 157.655 25.155 157.845 ;
        RECT 27.745 157.655 27.915 157.845 ;
        RECT 29.125 157.675 29.295 157.865 ;
        RECT 29.580 157.705 29.700 157.815 ;
        RECT 30.040 157.655 30.210 157.845 ;
        RECT 31.895 157.815 32.055 157.820 ;
        RECT 31.880 157.710 32.055 157.815 ;
        RECT 31.880 157.705 32.000 157.710 ;
        RECT 32.345 157.655 32.515 157.845 ;
        RECT 35.565 157.675 35.735 157.865 ;
        RECT 36.025 157.675 36.195 157.865 ;
        RECT 38.780 157.705 38.900 157.815 ;
        RECT 39.705 157.655 39.875 157.845 ;
        RECT 40.625 157.675 40.795 157.865 ;
        RECT 41.090 157.675 41.260 157.865 ;
        RECT 44.765 157.675 44.935 157.865 ;
        RECT 47.985 157.845 48.150 157.865 ;
        RECT 47.065 157.655 47.235 157.845 ;
        RECT 47.985 157.675 48.155 157.845 ;
        RECT 48.445 157.655 48.615 157.865 ;
        RECT 50.295 157.710 50.455 157.820 ;
        RECT 51.205 157.655 51.375 157.845 ;
        RECT 52.120 157.675 52.290 157.865 ;
        RECT 52.585 157.675 52.755 157.865 ;
        RECT 57.640 157.845 57.810 157.865 ;
        RECT 56.720 157.705 56.840 157.815 ;
        RECT 57.640 157.675 57.815 157.845 ;
        RECT 58.105 157.675 58.275 157.865 ;
        RECT 59.945 157.675 60.115 157.865 ;
        RECT 57.645 157.655 57.815 157.675 ;
        RECT 63.165 157.655 63.335 157.865 ;
        RECT 65.000 157.705 65.120 157.815 ;
        RECT 65.465 157.655 65.635 157.845 ;
        RECT 66.845 157.675 67.015 157.865 ;
        RECT 69.600 157.705 69.720 157.815 ;
        RECT 70.525 157.675 70.695 157.865 ;
        RECT 72.825 157.655 72.995 157.845 ;
        RECT 76.045 157.675 76.215 157.865 ;
        RECT 78.345 157.655 78.515 157.845 ;
        RECT 81.565 157.675 81.735 157.865 ;
        RECT 82.035 157.700 82.195 157.810 ;
        RECT 83.865 157.655 84.035 157.865 ;
        RECT 5.525 156.845 6.895 157.655 ;
        RECT 6.905 156.845 12.415 157.655 ;
        RECT 12.425 156.845 16.095 157.655 ;
        RECT 16.605 156.975 23.915 157.655 ;
        RECT 16.605 156.745 17.955 156.975 ;
        RECT 19.490 156.755 20.400 156.975 ;
        RECT 24.845 156.745 27.595 157.655 ;
        RECT 27.605 156.845 29.435 157.655 ;
        RECT 29.925 156.745 31.275 157.655 ;
        RECT 31.295 156.785 31.725 157.570 ;
        RECT 32.205 156.975 39.515 157.655 ;
        RECT 39.565 156.975 46.875 157.655 ;
        RECT 35.720 156.755 36.630 156.975 ;
        RECT 38.165 156.745 39.515 156.975 ;
        RECT 43.080 156.755 43.990 156.975 ;
        RECT 45.525 156.745 46.875 156.975 ;
        RECT 46.925 156.845 48.295 157.655 ;
        RECT 48.305 156.745 51.055 157.655 ;
        RECT 51.065 156.845 56.575 157.655 ;
        RECT 57.055 156.785 57.485 157.570 ;
        RECT 57.505 156.845 63.015 157.655 ;
        RECT 63.025 156.845 64.855 157.655 ;
        RECT 65.325 156.975 72.635 157.655 ;
        RECT 68.840 156.755 69.750 156.975 ;
        RECT 71.285 156.745 72.635 156.975 ;
        RECT 72.685 156.845 78.195 157.655 ;
        RECT 78.205 156.845 81.875 157.655 ;
        RECT 82.805 156.845 84.175 157.655 ;
      LAYER nwell ;
        RECT 5.330 153.625 84.370 156.455 ;
      LAYER pwell ;
        RECT 5.525 152.425 6.895 153.235 ;
        RECT 6.905 152.425 12.415 153.235 ;
        RECT 12.425 152.425 17.935 153.235 ;
        RECT 18.415 152.510 18.845 153.295 ;
        RECT 18.865 152.425 20.215 153.335 ;
        RECT 25.505 153.245 26.455 153.335 ;
        RECT 20.245 152.425 23.915 153.235 ;
        RECT 23.925 152.425 25.295 153.235 ;
        RECT 25.505 152.425 27.435 153.245 ;
        RECT 27.605 152.425 31.275 153.235 ;
        RECT 31.285 152.425 32.655 153.235 ;
        RECT 32.665 153.105 33.595 153.335 ;
        RECT 32.665 152.425 36.335 153.105 ;
        RECT 36.345 152.425 37.715 153.235 ;
        RECT 40.465 153.105 41.395 153.335 ;
        RECT 37.725 152.425 41.395 153.105 ;
        RECT 41.405 152.425 44.155 153.235 ;
        RECT 44.175 152.510 44.605 153.295 ;
        RECT 44.625 152.425 46.455 153.235 ;
        RECT 46.465 153.105 47.390 153.335 ;
        RECT 50.145 153.135 51.095 153.335 ;
        RECT 46.465 152.425 50.135 153.105 ;
        RECT 50.145 152.455 53.815 153.135 ;
        RECT 50.145 152.425 51.095 152.455 ;
        RECT 5.665 152.215 5.835 152.425 ;
        RECT 7.045 152.215 7.215 152.425 ;
        RECT 12.565 152.215 12.735 152.425 ;
        RECT 14.400 152.265 14.520 152.375 ;
        RECT 14.865 152.215 15.035 152.405 ;
        RECT 18.080 152.265 18.200 152.375 ;
        RECT 19.005 152.235 19.175 152.405 ;
        RECT 19.005 152.215 19.170 152.235 ;
        RECT 19.465 152.215 19.635 152.405 ;
        RECT 19.930 152.235 20.100 152.425 ;
        RECT 20.385 152.235 20.555 152.425 ;
        RECT 24.065 152.235 24.235 152.425 ;
        RECT 27.285 152.405 27.435 152.425 ;
        RECT 26.825 152.215 26.995 152.405 ;
        RECT 27.285 152.235 27.455 152.405 ;
        RECT 27.745 152.235 27.915 152.425 ;
        RECT 30.515 152.260 30.675 152.370 ;
        RECT 31.425 152.235 31.595 152.425 ;
        RECT 31.885 152.215 32.055 152.405 ;
        RECT 36.025 152.235 36.195 152.425 ;
        RECT 36.485 152.235 36.655 152.425 ;
        RECT 37.405 152.215 37.575 152.405 ;
        RECT 37.865 152.235 38.035 152.425 ;
        RECT 41.085 152.215 41.255 152.405 ;
        RECT 41.545 152.235 41.715 152.425 ;
        RECT 42.470 152.215 42.640 152.405 ;
        RECT 43.845 152.215 44.015 152.405 ;
        RECT 44.765 152.235 44.935 152.425 ;
        RECT 46.610 152.235 46.780 152.425 ;
        RECT 5.525 151.405 6.895 152.215 ;
        RECT 6.905 151.405 12.415 152.215 ;
        RECT 12.425 151.405 14.255 152.215 ;
        RECT 14.725 151.535 17.015 152.215 ;
        RECT 16.095 151.305 17.015 151.535 ;
        RECT 17.335 151.535 19.170 152.215 ;
        RECT 19.325 151.535 26.635 152.215 ;
        RECT 17.335 151.305 18.265 151.535 ;
        RECT 22.840 151.315 23.750 151.535 ;
        RECT 25.285 151.305 26.635 151.535 ;
        RECT 26.685 151.405 30.355 152.215 ;
        RECT 31.295 151.345 31.725 152.130 ;
        RECT 31.745 151.405 37.255 152.215 ;
        RECT 37.265 151.405 40.935 152.215 ;
        RECT 40.945 151.405 42.315 152.215 ;
        RECT 42.325 151.305 43.675 152.215 ;
        RECT 43.785 151.305 46.785 152.215 ;
        RECT 47.070 152.185 47.240 152.405 ;
        RECT 49.825 152.215 49.995 152.405 ;
        RECT 53.500 152.370 53.670 152.455 ;
        RECT 53.825 152.425 57.035 153.335 ;
        RECT 57.045 152.425 60.155 153.335 ;
        RECT 60.265 152.425 63.375 153.335 ;
        RECT 63.965 152.425 65.315 153.335 ;
        RECT 68.065 153.105 68.995 153.335 ;
        RECT 65.325 152.425 68.995 153.105 ;
        RECT 69.935 152.510 70.365 153.295 ;
        RECT 73.900 153.105 74.810 153.325 ;
        RECT 76.345 153.105 77.695 153.335 ;
        RECT 70.385 152.425 77.695 153.105 ;
        RECT 77.745 152.425 81.415 153.235 ;
        RECT 81.425 152.425 82.795 153.235 ;
        RECT 82.805 152.425 84.175 153.235 ;
        RECT 53.500 152.260 53.675 152.370 ;
        RECT 53.500 152.235 53.670 152.260 ;
        RECT 53.955 152.235 54.125 152.425 ;
        RECT 48.730 152.185 49.675 152.215 ;
        RECT 46.925 151.505 49.675 152.185 ;
        RECT 48.730 151.305 49.675 151.505 ;
        RECT 49.685 151.405 53.355 152.215 ;
        RECT 54.285 152.185 55.240 152.215 ;
        RECT 56.270 152.185 56.440 152.405 ;
        RECT 56.720 152.265 56.840 152.375 ;
        RECT 57.655 152.260 57.815 152.370 ;
        RECT 59.945 152.235 60.115 152.425 ;
        RECT 58.425 152.185 59.380 152.215 ;
        RECT 60.410 152.185 60.580 152.405 ;
        RECT 60.875 152.260 61.035 152.370 ;
        RECT 63.165 152.235 63.335 152.425 ;
        RECT 65.000 152.405 65.170 152.425 ;
        RECT 63.620 152.265 63.740 152.375 ;
        RECT 64.545 152.215 64.715 152.405 ;
        RECT 65.000 152.235 65.175 152.405 ;
        RECT 65.465 152.235 65.635 152.425 ;
        RECT 65.005 152.215 65.175 152.235 ;
        RECT 68.685 152.215 68.855 152.405 ;
        RECT 69.155 152.270 69.315 152.380 ;
        RECT 70.525 152.215 70.695 152.425 ;
        RECT 70.985 152.215 71.155 152.405 ;
        RECT 76.505 152.215 76.675 152.405 ;
        RECT 77.885 152.235 78.055 152.425 ;
        RECT 81.565 152.235 81.735 152.425 ;
        RECT 82.035 152.260 82.195 152.370 ;
        RECT 83.865 152.215 84.035 152.425 ;
        RECT 54.285 151.505 56.565 152.185 ;
        RECT 54.285 151.305 55.240 151.505 ;
        RECT 57.055 151.345 57.485 152.130 ;
        RECT 58.425 151.505 60.705 152.185 ;
        RECT 61.645 151.535 64.855 152.215 ;
        RECT 58.425 151.305 59.380 151.505 ;
        RECT 61.645 151.305 62.780 151.535 ;
        RECT 64.865 151.405 66.695 152.215 ;
        RECT 66.705 151.535 68.995 152.215 ;
        RECT 66.705 151.305 67.625 151.535 ;
        RECT 69.005 151.305 70.820 152.215 ;
        RECT 70.845 151.405 76.355 152.215 ;
        RECT 76.365 151.405 81.875 152.215 ;
        RECT 82.805 151.405 84.175 152.215 ;
      LAYER nwell ;
        RECT 5.330 148.185 84.370 151.015 ;
      LAYER pwell ;
        RECT 5.525 146.985 6.895 147.795 ;
        RECT 6.905 146.985 10.575 147.795 ;
        RECT 14.560 147.665 15.470 147.885 ;
        RECT 17.005 147.665 18.355 147.895 ;
        RECT 11.045 146.985 18.355 147.665 ;
        RECT 18.415 147.070 18.845 147.855 ;
        RECT 18.875 146.985 21.605 147.895 ;
        RECT 21.625 146.985 24.375 147.795 ;
        RECT 24.385 146.985 28.040 147.895 ;
        RECT 28.065 146.985 29.435 147.795 ;
        RECT 29.900 147.215 31.735 147.895 ;
        RECT 29.900 146.985 31.590 147.215 ;
        RECT 32.245 146.985 35.415 147.895 ;
        RECT 35.425 146.985 36.795 147.795 ;
        RECT 36.905 146.985 40.015 147.895 ;
        RECT 40.025 146.985 41.395 147.795 ;
        RECT 43.210 147.695 44.155 147.895 ;
        RECT 41.405 147.015 44.155 147.695 ;
        RECT 44.175 147.070 44.605 147.855 ;
        RECT 5.665 146.775 5.835 146.985 ;
        RECT 7.045 146.775 7.215 146.985 ;
        RECT 10.720 146.825 10.840 146.935 ;
        RECT 11.185 146.795 11.355 146.985 ;
        RECT 5.525 145.965 6.895 146.775 ;
        RECT 6.905 145.965 12.415 146.775 ;
        RECT 12.425 146.745 13.360 146.775 ;
        RECT 15.320 146.745 15.490 146.965 ;
        RECT 15.780 146.825 15.900 146.935 ;
        RECT 18.085 146.775 18.255 146.965 ;
        RECT 18.545 146.775 18.715 146.965 ;
        RECT 19.005 146.795 19.175 146.985 ;
        RECT 21.765 146.795 21.935 146.985 ;
        RECT 24.070 146.775 24.240 146.965 ;
        RECT 24.530 146.795 24.700 146.985 ;
        RECT 27.285 146.775 27.455 146.965 ;
        RECT 28.205 146.795 28.375 146.985 ;
        RECT 30.960 146.825 31.080 146.935 ;
        RECT 31.420 146.795 31.590 146.985 ;
        RECT 31.880 146.825 32.000 146.935 ;
        RECT 32.345 146.795 32.515 146.985 ;
        RECT 35.565 146.795 35.735 146.985 ;
        RECT 36.945 146.795 37.115 146.985 ;
        RECT 38.785 146.775 38.955 146.965 ;
        RECT 39.245 146.775 39.415 146.965 ;
        RECT 40.165 146.795 40.335 146.985 ;
        RECT 41.080 146.825 41.200 146.935 ;
        RECT 41.550 146.795 41.720 147.015 ;
        RECT 43.210 146.985 44.155 147.015 ;
        RECT 44.625 146.985 52.185 147.895 ;
        RECT 52.445 146.985 56.100 147.895 ;
        RECT 56.125 146.985 57.475 147.895 ;
        RECT 57.505 146.985 63.015 147.795 ;
        RECT 63.025 146.985 65.775 147.795 ;
        RECT 65.805 146.985 67.155 147.895 ;
        RECT 67.165 146.985 68.515 147.895 ;
        RECT 68.545 146.985 69.915 147.795 ;
        RECT 69.935 147.070 70.365 147.855 ;
        RECT 70.385 146.985 75.895 147.795 ;
        RECT 75.905 146.985 81.415 147.795 ;
        RECT 81.425 146.985 82.795 147.795 ;
        RECT 82.805 146.985 84.175 147.795 ;
        RECT 43.845 146.775 44.015 146.965 ;
        RECT 44.305 146.775 44.475 146.965 ;
        RECT 44.770 146.795 44.940 146.985 ;
        RECT 49.825 146.775 49.995 146.965 ;
        RECT 51.205 146.795 51.375 146.965 ;
        RECT 52.590 146.795 52.760 146.985 ;
        RECT 51.210 146.775 51.375 146.795 ;
        RECT 53.510 146.775 53.680 146.965 ;
        RECT 57.190 146.795 57.360 146.985 ;
        RECT 57.645 146.965 57.815 146.985 ;
        RECT 63.165 146.965 63.335 146.985 ;
        RECT 57.645 146.795 57.820 146.965 ;
        RECT 57.650 146.775 57.820 146.795 ;
        RECT 63.160 146.795 63.335 146.965 ;
        RECT 63.160 146.775 63.330 146.795 ;
        RECT 63.625 146.775 63.795 146.965 ;
        RECT 66.840 146.795 67.010 146.985 ;
        RECT 67.310 146.965 67.480 146.985 ;
        RECT 67.305 146.795 67.480 146.965 ;
        RECT 68.685 146.795 68.855 146.985 ;
        RECT 70.525 146.795 70.695 146.985 ;
        RECT 67.305 146.775 67.475 146.795 ;
        RECT 74.665 146.775 74.835 146.965 ;
        RECT 76.045 146.795 76.215 146.985 ;
        RECT 80.185 146.775 80.355 146.965 ;
        RECT 81.565 146.795 81.735 146.985 ;
        RECT 83.865 146.775 84.035 146.985 ;
        RECT 12.425 146.545 15.490 146.745 ;
        RECT 12.425 146.065 15.635 146.545 ;
        RECT 12.425 145.865 13.375 146.065 ;
        RECT 14.705 145.865 15.635 146.065 ;
        RECT 16.105 146.095 18.395 146.775 ;
        RECT 16.105 145.865 17.025 146.095 ;
        RECT 18.405 145.965 23.915 146.775 ;
        RECT 23.925 145.865 26.990 146.775 ;
        RECT 27.145 145.965 30.815 146.775 ;
        RECT 31.295 145.905 31.725 146.690 ;
        RECT 31.785 146.095 39.095 146.775 ;
        RECT 31.785 145.865 33.135 146.095 ;
        RECT 34.670 145.875 35.580 146.095 ;
        RECT 39.105 145.965 40.935 146.775 ;
        RECT 41.415 145.865 44.145 146.775 ;
        RECT 44.165 145.965 49.675 146.775 ;
        RECT 49.685 145.965 51.055 146.775 ;
        RECT 51.210 146.095 53.045 146.775 ;
        RECT 52.115 145.865 53.045 146.095 ;
        RECT 53.365 145.865 56.840 146.775 ;
        RECT 57.055 145.905 57.485 146.690 ;
        RECT 57.505 145.865 60.980 146.775 ;
        RECT 61.640 146.545 63.330 146.775 ;
        RECT 61.640 145.865 63.475 146.545 ;
        RECT 63.485 146.095 67.155 146.775 ;
        RECT 67.165 146.095 74.475 146.775 ;
        RECT 66.225 145.865 67.155 146.095 ;
        RECT 70.680 145.875 71.590 146.095 ;
        RECT 73.125 145.865 74.475 146.095 ;
        RECT 74.525 145.965 80.035 146.775 ;
        RECT 80.045 145.965 82.795 146.775 ;
        RECT 82.805 145.965 84.175 146.775 ;
      LAYER nwell ;
        RECT 5.330 142.745 84.370 145.575 ;
      LAYER pwell ;
        RECT 5.525 141.545 6.895 142.355 ;
        RECT 6.905 141.545 12.415 142.355 ;
        RECT 12.425 141.545 17.935 142.355 ;
        RECT 18.415 141.630 18.845 142.415 ;
        RECT 18.865 141.545 20.235 142.355 ;
        RECT 20.265 141.545 21.615 142.455 ;
        RECT 22.555 141.545 25.285 142.455 ;
        RECT 27.960 142.225 28.880 142.455 ;
        RECT 30.035 142.225 30.965 142.455 ;
        RECT 25.415 141.545 28.880 142.225 ;
        RECT 29.130 141.545 30.965 142.225 ;
        RECT 31.295 141.545 32.645 142.455 ;
        RECT 35.405 142.225 36.335 142.455 ;
        RECT 32.665 141.545 36.335 142.225 ;
        RECT 36.345 141.545 41.855 142.355 ;
        RECT 41.865 141.545 43.695 142.355 ;
        RECT 44.175 141.630 44.605 142.415 ;
        RECT 51.745 142.365 52.695 142.455 ;
        RECT 44.625 141.545 50.135 142.355 ;
        RECT 50.765 141.545 52.695 142.365 ;
        RECT 52.905 142.255 53.835 142.455 ;
        RECT 55.170 142.255 56.115 142.455 ;
        RECT 52.905 141.775 56.115 142.255 ;
        RECT 53.045 141.575 56.115 141.775 ;
        RECT 5.665 141.335 5.835 141.545 ;
        RECT 7.045 141.335 7.215 141.545 ;
        RECT 12.565 141.335 12.735 141.545 ;
        RECT 17.165 141.355 17.335 141.525 ;
        RECT 17.625 141.355 17.795 141.525 ;
        RECT 18.080 141.385 18.200 141.495 ;
        RECT 19.005 141.355 19.175 141.545 ;
        RECT 17.165 141.335 17.315 141.355 ;
        RECT 5.525 140.525 6.895 141.335 ;
        RECT 6.905 140.525 12.415 141.335 ;
        RECT 12.425 140.525 15.175 141.335 ;
        RECT 15.385 140.515 17.315 141.335 ;
        RECT 17.630 141.335 17.795 141.355 ;
        RECT 17.630 140.655 19.465 141.335 ;
        RECT 19.930 141.305 20.100 141.525 ;
        RECT 20.380 141.355 20.550 141.545 ;
        RECT 21.775 141.390 21.935 141.500 ;
        RECT 22.685 141.355 22.855 141.545 ;
        RECT 23.605 141.335 23.775 141.525 ;
        RECT 25.445 141.355 25.615 141.545 ;
        RECT 29.130 141.525 29.295 141.545 ;
        RECT 28.665 141.355 28.835 141.525 ;
        RECT 29.125 141.355 29.295 141.525 ;
        RECT 31.425 141.355 31.595 141.545 ;
        RECT 28.815 141.335 28.835 141.355 ;
        RECT 31.885 141.335 32.055 141.525 ;
        RECT 32.805 141.355 32.975 141.545 ;
        RECT 35.565 141.335 35.735 141.525 ;
        RECT 36.035 141.380 36.195 141.490 ;
        RECT 36.485 141.355 36.655 141.545 ;
        RECT 37.860 141.335 38.030 141.525 ;
        RECT 38.325 141.335 38.495 141.525 ;
        RECT 40.160 141.385 40.280 141.495 ;
        RECT 41.540 141.335 41.710 141.525 ;
        RECT 42.005 141.355 42.175 141.545 ;
        RECT 43.385 141.335 43.555 141.525 ;
        RECT 43.840 141.385 43.960 141.495 ;
        RECT 44.765 141.355 44.935 141.545 ;
        RECT 50.765 141.525 50.915 141.545 ;
        RECT 50.280 141.385 50.400 141.495 ;
        RECT 50.745 141.335 50.915 141.525 ;
        RECT 51.215 141.380 51.375 141.490 ;
        RECT 52.125 141.335 52.295 141.525 ;
        RECT 53.045 141.355 53.215 141.575 ;
        RECT 55.170 141.545 56.115 141.575 ;
        RECT 56.125 141.545 59.285 142.455 ;
        RECT 64.415 142.225 67.415 142.455 ;
        RECT 59.345 141.545 64.160 142.225 ;
        RECT 64.415 142.135 68.995 142.225 ;
        RECT 64.405 141.775 68.995 142.135 ;
        RECT 64.405 141.585 65.335 141.775 ;
        RECT 64.415 141.545 65.335 141.585 ;
        RECT 67.425 141.545 68.995 141.775 ;
        RECT 69.935 141.630 70.365 142.415 ;
        RECT 70.385 141.545 71.755 142.325 ;
        RECT 71.765 141.545 77.275 142.355 ;
        RECT 77.285 141.545 82.795 142.355 ;
        RECT 82.805 141.545 84.175 142.355 ;
        RECT 55.345 141.335 55.515 141.525 ;
        RECT 57.645 141.335 57.815 141.525 ;
        RECT 59.025 141.355 59.195 141.545 ;
        RECT 59.485 141.355 59.655 141.545 ;
        RECT 60.405 141.335 60.575 141.525 ;
        RECT 62.245 141.335 62.415 141.525 ;
        RECT 68.685 141.355 68.855 141.545 ;
        RECT 69.155 141.390 69.315 141.500 ;
        RECT 69.605 141.335 69.775 141.525 ;
        RECT 71.445 141.355 71.615 141.545 ;
        RECT 71.905 141.355 72.075 141.545 ;
        RECT 75.125 141.335 75.295 141.525 ;
        RECT 77.425 141.355 77.595 141.545 ;
        RECT 80.645 141.335 80.815 141.525 ;
        RECT 82.480 141.385 82.600 141.495 ;
        RECT 83.865 141.335 84.035 141.545 ;
        RECT 22.505 141.305 23.455 141.335 ;
        RECT 15.385 140.425 16.335 140.515 ;
        RECT 18.535 140.425 19.465 140.655 ;
        RECT 19.785 140.625 23.455 141.305 ;
        RECT 23.465 140.655 28.280 141.335 ;
        RECT 28.815 140.655 31.265 141.335 ;
        RECT 22.505 140.425 23.455 140.625 ;
        RECT 29.305 140.425 31.265 140.655 ;
        RECT 31.295 140.465 31.725 141.250 ;
        RECT 31.745 140.525 33.835 141.335 ;
        RECT 34.505 140.555 35.875 141.335 ;
        RECT 36.825 140.425 38.175 141.335 ;
        RECT 38.185 140.525 40.015 141.335 ;
        RECT 40.505 140.425 41.855 141.335 ;
        RECT 41.865 140.655 43.695 141.335 ;
        RECT 43.745 140.655 51.055 141.335 ;
        RECT 43.745 140.425 45.095 140.655 ;
        RECT 46.630 140.435 47.540 140.655 ;
        RECT 51.985 140.425 55.195 141.335 ;
        RECT 55.205 140.525 57.035 141.335 ;
        RECT 57.055 140.465 57.485 141.250 ;
        RECT 57.505 140.425 60.255 141.335 ;
        RECT 60.265 140.525 62.095 141.335 ;
        RECT 62.105 140.655 69.415 141.335 ;
        RECT 65.620 140.435 66.530 140.655 ;
        RECT 68.065 140.425 69.415 140.655 ;
        RECT 69.465 140.525 74.975 141.335 ;
        RECT 74.985 140.525 80.495 141.335 ;
        RECT 80.505 140.525 82.335 141.335 ;
        RECT 82.805 140.525 84.175 141.335 ;
      LAYER nwell ;
        RECT 5.330 137.305 84.370 140.135 ;
      LAYER pwell ;
        RECT 5.525 136.105 6.895 136.915 ;
        RECT 6.905 136.105 10.575 136.915 ;
        RECT 14.560 136.785 15.470 137.005 ;
        RECT 17.005 136.785 18.355 137.015 ;
        RECT 11.045 136.105 18.355 136.785 ;
        RECT 18.415 136.190 18.845 136.975 ;
        RECT 21.205 136.785 22.555 137.015 ;
        RECT 24.090 136.785 25.000 137.005 ;
        RECT 28.620 136.785 29.540 137.015 ;
        RECT 19.325 136.105 21.155 136.785 ;
        RECT 21.205 136.105 28.515 136.785 ;
        RECT 28.620 136.105 32.085 136.785 ;
        RECT 32.205 136.105 34.035 136.915 ;
        RECT 37.560 136.785 38.470 137.005 ;
        RECT 40.005 136.785 41.355 137.015 ;
        RECT 43.235 136.785 44.155 137.015 ;
        RECT 34.045 136.105 41.355 136.785 ;
        RECT 41.865 136.105 44.155 136.785 ;
        RECT 44.175 136.190 44.605 136.975 ;
        RECT 47.365 136.785 48.295 137.015 ;
        RECT 44.625 136.105 48.295 136.785 ;
        RECT 48.320 136.105 50.135 137.015 ;
        RECT 50.380 136.105 55.195 136.785 ;
        RECT 55.205 136.105 56.575 136.915 ;
        RECT 56.585 136.785 57.720 137.015 ;
        RECT 56.585 136.105 59.795 136.785 ;
        RECT 59.805 136.105 65.315 136.915 ;
        RECT 65.325 136.105 68.995 136.915 ;
        RECT 69.935 136.190 70.365 136.975 ;
        RECT 70.385 136.105 75.895 136.915 ;
        RECT 75.905 136.105 81.415 136.915 ;
        RECT 81.425 136.105 82.795 136.915 ;
        RECT 82.805 136.105 84.175 136.915 ;
        RECT 5.665 135.895 5.835 136.105 ;
        RECT 7.045 135.915 7.215 136.105 ;
        RECT 8.425 135.895 8.595 136.085 ;
        RECT 8.885 135.895 9.055 136.085 ;
        RECT 10.720 135.945 10.840 136.055 ;
        RECT 11.185 135.915 11.355 136.105 ;
        RECT 12.575 135.940 12.735 136.050 ;
        RECT 5.525 135.085 6.895 135.895 ;
        RECT 6.905 135.215 8.735 135.895 ;
        RECT 6.905 134.985 8.250 135.215 ;
        RECT 8.745 135.085 12.415 135.895 ;
        RECT 13.345 135.865 14.280 135.895 ;
        RECT 16.240 135.865 16.410 136.085 ;
        RECT 16.705 135.895 16.875 136.085 ;
        RECT 18.085 135.915 18.255 136.085 ;
        RECT 19.000 135.945 19.120 136.055 ;
        RECT 19.465 135.915 19.635 136.105 ;
        RECT 18.090 135.895 18.255 135.915 ;
        RECT 20.385 135.895 20.555 136.085 ;
        RECT 22.685 135.895 22.855 136.085 ;
        RECT 28.205 135.915 28.375 136.105 ;
        RECT 30.045 135.895 30.215 136.085 ;
        RECT 31.885 135.915 32.055 136.105 ;
        RECT 32.345 135.915 32.515 136.105 ;
        RECT 32.805 135.895 32.975 136.085 ;
        RECT 34.185 135.915 34.355 136.105 ;
        RECT 41.085 135.895 41.255 136.085 ;
        RECT 41.540 135.945 41.660 136.055 ;
        RECT 42.005 135.915 42.175 136.105 ;
        RECT 44.305 135.895 44.475 136.085 ;
        RECT 44.765 135.915 44.935 136.105 ;
        RECT 45.680 135.895 45.850 136.085 ;
        RECT 46.145 135.895 46.315 136.085 ;
        RECT 48.445 135.915 48.615 136.105 ;
        RECT 49.820 135.945 49.940 136.055 ;
        RECT 50.285 135.895 50.455 136.085 ;
        RECT 53.505 135.895 53.675 136.085 ;
        RECT 54.885 135.915 55.055 136.105 ;
        RECT 55.345 135.915 55.515 136.105 ;
        RECT 57.645 135.895 57.815 136.085 ;
        RECT 59.485 135.915 59.655 136.105 ;
        RECT 59.945 135.915 60.115 136.105 ;
        RECT 60.400 135.895 60.570 136.085 ;
        RECT 60.865 135.895 61.035 136.085 ;
        RECT 62.245 135.895 62.415 136.085 ;
        RECT 65.465 135.915 65.635 136.105 ;
        RECT 69.155 135.950 69.315 136.060 ;
        RECT 70.525 135.915 70.695 136.105 ;
        RECT 72.825 135.895 72.995 136.085 ;
        RECT 73.285 135.895 73.455 136.085 ;
        RECT 76.045 135.915 76.215 136.105 ;
        RECT 78.805 135.895 78.975 136.085 ;
        RECT 81.565 135.915 81.735 136.105 ;
        RECT 82.480 135.945 82.600 136.055 ;
        RECT 83.865 135.895 84.035 136.105 ;
        RECT 13.345 135.665 16.410 135.865 ;
        RECT 13.345 135.185 16.555 135.665 ;
        RECT 13.345 134.985 14.295 135.185 ;
        RECT 15.625 134.985 16.555 135.185 ;
        RECT 16.565 135.085 17.935 135.895 ;
        RECT 18.090 135.215 19.925 135.895 ;
        RECT 20.245 135.215 22.535 135.895 ;
        RECT 22.545 135.215 29.855 135.895 ;
        RECT 18.995 134.985 19.925 135.215 ;
        RECT 21.615 134.985 22.535 135.215 ;
        RECT 26.060 134.995 26.970 135.215 ;
        RECT 28.505 134.985 29.855 135.215 ;
        RECT 29.905 135.085 31.275 135.895 ;
        RECT 31.295 135.025 31.725 135.810 ;
        RECT 32.665 135.215 37.480 135.895 ;
        RECT 37.725 135.215 41.395 135.895 ;
        RECT 41.405 135.215 44.615 135.895 ;
        RECT 37.725 134.985 38.655 135.215 ;
        RECT 41.405 134.985 42.540 135.215 ;
        RECT 44.645 134.985 45.995 135.895 ;
        RECT 46.005 135.085 49.675 135.895 ;
        RECT 50.195 134.985 53.355 135.895 ;
        RECT 53.365 135.085 57.035 135.895 ;
        RECT 57.055 135.025 57.485 135.810 ;
        RECT 57.505 135.085 59.335 135.895 ;
        RECT 59.365 134.985 60.715 135.895 ;
        RECT 60.725 135.085 62.095 135.895 ;
        RECT 62.105 135.215 65.775 135.895 ;
        RECT 64.845 134.985 65.775 135.215 ;
        RECT 65.825 135.215 73.135 135.895 ;
        RECT 65.825 134.985 67.175 135.215 ;
        RECT 68.710 134.995 69.620 135.215 ;
        RECT 73.145 135.085 78.655 135.895 ;
        RECT 78.665 135.085 82.335 135.895 ;
        RECT 82.805 135.085 84.175 135.895 ;
      LAYER nwell ;
        RECT 5.330 131.865 84.370 134.695 ;
      LAYER pwell ;
        RECT 5.525 130.665 6.895 131.475 ;
        RECT 6.905 130.665 12.415 131.475 ;
        RECT 12.425 130.665 17.935 131.475 ;
        RECT 18.415 130.750 18.845 131.535 ;
        RECT 18.865 130.665 22.535 131.475 ;
        RECT 23.465 130.665 25.555 131.475 ;
        RECT 26.240 130.665 28.055 131.575 ;
        RECT 28.065 130.665 29.895 131.475 ;
        RECT 33.880 131.345 34.790 131.565 ;
        RECT 36.325 131.345 37.675 131.575 ;
        RECT 30.365 130.665 37.675 131.345 ;
        RECT 37.725 130.665 43.235 131.475 ;
        RECT 44.175 130.750 44.605 131.535 ;
        RECT 44.625 130.665 46.455 131.345 ;
        RECT 46.465 130.665 50.135 131.475 ;
        RECT 52.885 131.345 53.815 131.575 ;
        RECT 50.145 130.665 53.815 131.345 ;
        RECT 53.845 130.665 55.195 131.575 ;
        RECT 55.685 130.665 57.035 131.575 ;
        RECT 57.965 131.345 58.885 131.575 ;
        RECT 57.965 130.665 60.255 131.345 ;
        RECT 60.280 130.665 62.095 131.575 ;
        RECT 63.065 130.665 66.235 131.575 ;
        RECT 66.245 130.665 69.915 131.475 ;
        RECT 69.935 130.750 70.365 131.535 ;
        RECT 70.385 130.665 75.895 131.475 ;
        RECT 75.905 130.665 81.415 131.475 ;
        RECT 81.425 130.665 82.795 131.475 ;
        RECT 82.805 130.665 84.175 131.475 ;
        RECT 5.665 130.455 5.835 130.665 ;
        RECT 7.045 130.455 7.215 130.665 ;
        RECT 12.565 130.455 12.735 130.665 ;
        RECT 18.085 130.615 18.255 130.645 ;
        RECT 18.080 130.505 18.255 130.615 ;
        RECT 18.085 130.455 18.255 130.505 ;
        RECT 19.005 130.475 19.175 130.665 ;
        RECT 5.525 129.645 6.895 130.455 ;
        RECT 6.905 129.645 12.415 130.455 ;
        RECT 12.425 129.645 17.935 130.455 ;
        RECT 17.945 129.645 19.315 130.455 ;
        RECT 19.325 130.425 20.260 130.455 ;
        RECT 22.220 130.425 22.390 130.645 ;
        RECT 22.695 130.615 22.855 130.620 ;
        RECT 22.680 130.510 22.855 130.615 ;
        RECT 22.680 130.505 22.800 130.510 ;
        RECT 23.145 130.455 23.315 130.645 ;
        RECT 23.605 130.475 23.775 130.665 ;
        RECT 26.365 130.475 26.535 130.665 ;
        RECT 26.835 130.500 26.995 130.610 ;
        RECT 27.745 130.455 27.915 130.645 ;
        RECT 28.205 130.475 28.375 130.665 ;
        RECT 30.040 130.505 30.160 130.615 ;
        RECT 30.505 130.475 30.675 130.665 ;
        RECT 31.885 130.455 32.055 130.645 ;
        RECT 33.725 130.455 33.895 130.645 ;
        RECT 37.865 130.475 38.035 130.665 ;
        RECT 38.325 130.455 38.495 130.645 ;
        RECT 39.710 130.455 39.880 130.645 ;
        RECT 40.175 130.500 40.335 130.610 ;
        RECT 41.085 130.455 41.255 130.645 ;
        RECT 43.395 130.510 43.555 130.620 ;
        RECT 44.305 130.455 44.475 130.645 ;
        RECT 46.145 130.475 46.315 130.665 ;
        RECT 46.605 130.475 46.775 130.665 ;
        RECT 47.985 130.455 48.155 130.645 ;
        RECT 49.825 130.455 49.995 130.645 ;
        RECT 50.285 130.475 50.455 130.665 ;
        RECT 54.880 130.475 55.050 130.665 ;
        RECT 55.340 130.505 55.460 130.615 ;
        RECT 56.720 130.475 56.890 130.665 ;
        RECT 57.195 130.510 57.355 130.620 ;
        RECT 57.655 130.500 57.815 130.610 ;
        RECT 58.565 130.455 58.735 130.645 ;
        RECT 59.945 130.475 60.115 130.665 ;
        RECT 60.405 130.475 60.575 130.665 ;
        RECT 62.255 130.510 62.415 130.620 ;
        RECT 63.165 130.475 63.335 130.665 ;
        RECT 65.925 130.455 66.095 130.645 ;
        RECT 66.385 130.475 66.555 130.665 ;
        RECT 70.525 130.475 70.695 130.665 ;
        RECT 71.445 130.455 71.615 130.645 ;
        RECT 76.045 130.475 76.215 130.665 ;
        RECT 76.965 130.455 77.135 130.645 ;
        RECT 81.565 130.475 81.735 130.665 ;
        RECT 82.480 130.505 82.600 130.615 ;
        RECT 83.865 130.455 84.035 130.665 ;
        RECT 19.325 130.225 22.390 130.425 ;
        RECT 19.325 129.745 22.535 130.225 ;
        RECT 23.115 129.775 26.580 130.455 ;
        RECT 27.715 129.775 31.180 130.455 ;
        RECT 19.325 129.545 20.275 129.745 ;
        RECT 21.605 129.545 22.535 129.745 ;
        RECT 25.660 129.545 26.580 129.775 ;
        RECT 30.260 129.545 31.180 129.775 ;
        RECT 31.295 129.585 31.725 130.370 ;
        RECT 31.760 129.545 33.575 130.455 ;
        RECT 33.585 129.645 34.955 130.455 ;
        RECT 35.060 129.775 38.525 130.455 ;
        RECT 35.060 129.545 35.980 129.775 ;
        RECT 38.645 129.545 39.995 130.455 ;
        RECT 40.985 129.545 44.155 130.455 ;
        RECT 44.165 129.775 47.835 130.455 ;
        RECT 46.905 129.545 47.835 129.775 ;
        RECT 47.845 129.645 49.675 130.455 ;
        RECT 49.685 129.775 56.995 130.455 ;
        RECT 53.200 129.555 54.110 129.775 ;
        RECT 55.645 129.545 56.995 129.775 ;
        RECT 57.055 129.585 57.485 130.370 ;
        RECT 58.425 129.775 65.735 130.455 ;
        RECT 61.940 129.555 62.850 129.775 ;
        RECT 64.385 129.545 65.735 129.775 ;
        RECT 65.785 129.645 71.295 130.455 ;
        RECT 71.305 129.645 76.815 130.455 ;
        RECT 76.825 129.645 82.335 130.455 ;
        RECT 82.805 129.645 84.175 130.455 ;
      LAYER nwell ;
        RECT 5.330 126.425 84.370 129.255 ;
      LAYER pwell ;
        RECT 5.525 125.225 6.895 126.035 ;
        RECT 6.905 125.225 12.415 126.035 ;
        RECT 12.425 125.225 17.935 126.035 ;
        RECT 18.415 125.310 18.845 126.095 ;
        RECT 18.905 125.905 20.255 126.135 ;
        RECT 21.790 125.905 22.700 126.125 ;
        RECT 26.535 125.905 27.465 126.135 ;
        RECT 32.040 125.905 32.950 126.125 ;
        RECT 34.485 125.905 35.835 126.135 ;
        RECT 38.635 125.905 39.555 126.135 ;
        RECT 18.905 125.225 26.215 125.905 ;
        RECT 26.535 125.225 28.370 125.905 ;
        RECT 28.525 125.225 35.835 125.905 ;
        RECT 35.970 125.225 39.555 125.905 ;
        RECT 39.660 125.905 40.580 126.135 ;
        RECT 39.660 125.225 43.125 125.905 ;
        RECT 44.175 125.310 44.605 126.095 ;
        RECT 44.625 125.225 45.975 126.135 ;
        RECT 49.520 125.905 50.430 126.125 ;
        RECT 51.965 125.905 53.315 126.135 ;
        RECT 46.005 125.225 53.315 125.905 ;
        RECT 53.365 125.225 57.035 126.035 ;
        RECT 60.245 125.905 61.175 126.135 ;
        RECT 57.505 125.225 61.175 125.905 ;
        RECT 61.185 125.225 66.695 126.035 ;
        RECT 66.705 125.225 69.455 126.035 ;
        RECT 69.935 125.310 70.365 126.095 ;
        RECT 70.385 125.225 75.895 126.035 ;
        RECT 75.905 125.225 81.415 126.035 ;
        RECT 81.425 125.225 82.795 126.035 ;
        RECT 82.805 125.225 84.175 126.035 ;
        RECT 5.665 125.015 5.835 125.225 ;
        RECT 7.045 125.015 7.215 125.225 ;
        RECT 12.565 125.015 12.735 125.225 ;
        RECT 18.085 125.175 18.255 125.205 ;
        RECT 18.080 125.065 18.255 125.175 ;
        RECT 18.085 125.015 18.255 125.065 ;
        RECT 25.905 125.035 26.075 125.225 ;
        RECT 28.205 125.205 28.370 125.225 ;
        RECT 27.745 125.015 27.915 125.205 ;
        RECT 28.205 125.035 28.375 125.205 ;
        RECT 28.665 125.035 28.835 125.225 ;
        RECT 30.965 125.015 31.135 125.205 ;
        RECT 31.895 125.060 32.055 125.170 ;
        RECT 32.805 125.015 32.975 125.205 ;
        RECT 39.240 125.035 39.410 125.225 ;
        RECT 39.700 125.015 39.870 125.205 ;
        RECT 40.165 125.015 40.335 125.205 ;
        RECT 42.925 125.035 43.095 125.225 ;
        RECT 43.395 125.070 43.555 125.180 ;
        RECT 45.690 125.035 45.860 125.225 ;
        RECT 46.145 125.035 46.315 125.225 ;
        RECT 47.525 125.015 47.695 125.205 ;
        RECT 53.045 125.015 53.215 125.205 ;
        RECT 53.505 125.035 53.675 125.225 ;
        RECT 56.720 125.065 56.840 125.175 ;
        RECT 57.180 125.065 57.300 125.175 ;
        RECT 57.645 125.015 57.815 125.225 ;
        RECT 61.325 125.035 61.495 125.225 ;
        RECT 63.165 125.015 63.335 125.205 ;
        RECT 66.845 125.035 67.015 125.225 ;
        RECT 68.685 125.015 68.855 125.205 ;
        RECT 69.600 125.065 69.720 125.175 ;
        RECT 70.525 125.035 70.695 125.225 ;
        RECT 74.205 125.015 74.375 125.205 ;
        RECT 76.045 125.035 76.215 125.225 ;
        RECT 79.725 125.015 79.895 125.205 ;
        RECT 81.565 125.035 81.735 125.225 ;
        RECT 82.480 125.065 82.600 125.175 ;
        RECT 83.865 125.015 84.035 125.225 ;
        RECT 5.525 124.205 6.895 125.015 ;
        RECT 6.905 124.205 12.415 125.015 ;
        RECT 12.425 124.205 17.935 125.015 ;
        RECT 17.945 124.205 20.695 125.015 ;
        RECT 20.745 124.335 28.055 125.015 ;
        RECT 20.745 124.105 22.095 124.335 ;
        RECT 23.630 124.115 24.540 124.335 ;
        RECT 28.065 124.105 31.175 125.015 ;
        RECT 31.295 124.145 31.725 124.930 ;
        RECT 32.775 124.335 36.240 125.015 ;
        RECT 36.430 124.335 40.015 125.015 ;
        RECT 40.025 124.335 47.335 125.015 ;
        RECT 35.320 124.105 36.240 124.335 ;
        RECT 39.095 124.105 40.015 124.335 ;
        RECT 43.540 124.115 44.450 124.335 ;
        RECT 45.985 124.105 47.335 124.335 ;
        RECT 47.385 124.205 52.895 125.015 ;
        RECT 52.905 124.205 56.575 125.015 ;
        RECT 57.055 124.145 57.485 124.930 ;
        RECT 57.505 124.205 63.015 125.015 ;
        RECT 63.025 124.205 68.535 125.015 ;
        RECT 68.545 124.205 74.055 125.015 ;
        RECT 74.065 124.205 79.575 125.015 ;
        RECT 79.585 124.205 82.335 125.015 ;
        RECT 82.805 124.205 84.175 125.015 ;
      LAYER nwell ;
        RECT 5.330 120.985 84.370 123.815 ;
      LAYER pwell ;
        RECT 5.525 119.785 6.895 120.595 ;
        RECT 6.905 119.785 12.415 120.595 ;
        RECT 12.425 119.785 17.935 120.595 ;
        RECT 18.415 119.870 18.845 120.655 ;
        RECT 18.865 119.785 20.235 120.595 ;
        RECT 22.900 120.465 23.820 120.695 ;
        RECT 20.355 119.785 23.820 120.465 ;
        RECT 23.925 119.785 26.675 120.595 ;
        RECT 27.155 119.785 30.815 120.695 ;
        RECT 30.855 119.785 33.575 120.695 ;
        RECT 37.100 120.465 38.010 120.685 ;
        RECT 39.545 120.465 40.895 120.695 ;
        RECT 42.280 120.495 43.235 120.695 ;
        RECT 33.585 119.785 40.895 120.465 ;
        RECT 40.955 119.815 43.235 120.495 ;
        RECT 44.175 119.870 44.605 120.655 ;
        RECT 5.665 119.575 5.835 119.785 ;
        RECT 7.045 119.575 7.215 119.785 ;
        RECT 12.565 119.575 12.735 119.785 ;
        RECT 15.325 119.575 15.495 119.765 ;
        RECT 18.080 119.625 18.200 119.735 ;
        RECT 19.005 119.595 19.175 119.785 ;
        RECT 20.385 119.595 20.555 119.785 ;
        RECT 22.685 119.575 22.855 119.765 ;
        RECT 24.065 119.595 24.235 119.785 ;
        RECT 26.820 119.625 26.940 119.735 ;
        RECT 27.280 119.595 27.450 119.785 ;
        RECT 28.205 119.575 28.375 119.765 ;
        RECT 30.960 119.625 31.080 119.735 ;
        RECT 31.885 119.575 32.055 119.765 ;
        RECT 33.265 119.595 33.435 119.785 ;
        RECT 33.725 119.595 33.895 119.785 ;
        RECT 39.245 119.595 39.415 119.765 ;
        RECT 39.245 119.575 39.410 119.595 ;
        RECT 40.625 119.575 40.795 119.765 ;
        RECT 41.080 119.595 41.250 119.815 ;
        RECT 42.280 119.785 43.235 119.815 ;
        RECT 44.625 119.785 47.365 120.465 ;
        RECT 47.385 119.785 49.215 120.595 ;
        RECT 49.320 120.465 50.240 120.695 ;
        RECT 49.320 119.785 52.785 120.465 ;
        RECT 52.905 119.785 54.735 120.595 ;
        RECT 54.840 120.465 55.760 120.695 ;
        RECT 54.840 119.785 58.305 120.465 ;
        RECT 58.425 119.785 61.900 120.695 ;
        RECT 62.105 119.785 67.615 120.595 ;
        RECT 67.625 119.785 69.455 120.595 ;
        RECT 69.935 119.870 70.365 120.655 ;
        RECT 70.385 119.785 75.895 120.595 ;
        RECT 75.905 119.785 81.415 120.595 ;
        RECT 81.425 119.785 82.795 120.595 ;
        RECT 82.805 119.785 84.175 120.595 ;
        RECT 42.000 119.575 42.170 119.765 ;
        RECT 42.465 119.575 42.635 119.765 ;
        RECT 43.395 119.630 43.555 119.740 ;
        RECT 44.765 119.595 44.935 119.785 ;
        RECT 46.145 119.575 46.315 119.765 ;
        RECT 47.525 119.575 47.695 119.785 ;
        RECT 52.585 119.595 52.755 119.785 ;
        RECT 53.045 119.595 53.215 119.785 ;
        RECT 54.890 119.575 55.060 119.765 ;
        RECT 56.275 119.620 56.435 119.730 ;
        RECT 57.645 119.575 57.815 119.765 ;
        RECT 58.105 119.595 58.275 119.785 ;
        RECT 58.570 119.595 58.740 119.785 ;
        RECT 62.245 119.595 62.415 119.785 ;
        RECT 66.385 119.575 66.555 119.765 ;
        RECT 66.845 119.575 67.015 119.765 ;
        RECT 67.765 119.595 67.935 119.785 ;
        RECT 69.600 119.625 69.720 119.735 ;
        RECT 70.525 119.595 70.695 119.785 ;
        RECT 72.365 119.575 72.535 119.765 ;
        RECT 76.045 119.595 76.215 119.785 ;
        RECT 77.885 119.575 78.055 119.765 ;
        RECT 81.565 119.575 81.735 119.785 ;
        RECT 83.865 119.575 84.035 119.785 ;
        RECT 5.525 118.765 6.895 119.575 ;
        RECT 6.905 118.765 12.415 119.575 ;
        RECT 12.425 118.765 15.175 119.575 ;
        RECT 15.185 118.895 22.495 119.575 ;
        RECT 18.700 118.675 19.610 118.895 ;
        RECT 21.145 118.665 22.495 118.895 ;
        RECT 22.545 118.765 28.055 119.575 ;
        RECT 28.065 118.765 30.815 119.575 ;
        RECT 31.295 118.705 31.725 119.490 ;
        RECT 31.745 118.765 37.255 119.575 ;
        RECT 37.575 118.895 39.410 119.575 ;
        RECT 37.575 118.665 38.505 118.895 ;
        RECT 39.575 118.665 40.925 119.575 ;
        RECT 40.965 118.665 42.315 119.575 ;
        RECT 42.325 118.765 45.995 119.575 ;
        RECT 46.005 118.765 47.375 119.575 ;
        RECT 47.385 118.895 54.695 119.575 ;
        RECT 50.900 118.675 51.810 118.895 ;
        RECT 53.345 118.665 54.695 118.895 ;
        RECT 54.745 118.665 56.095 119.575 ;
        RECT 57.055 118.705 57.485 119.490 ;
        RECT 57.505 118.765 59.335 119.575 ;
        RECT 59.385 118.895 66.695 119.575 ;
        RECT 59.385 118.665 60.735 118.895 ;
        RECT 62.270 118.675 63.180 118.895 ;
        RECT 66.705 118.765 72.215 119.575 ;
        RECT 72.225 118.765 77.735 119.575 ;
        RECT 77.745 118.765 81.415 119.575 ;
        RECT 81.425 118.765 82.795 119.575 ;
        RECT 82.805 118.765 84.175 119.575 ;
      LAYER nwell ;
        RECT 5.330 115.545 84.370 118.375 ;
      LAYER pwell ;
        RECT 5.525 114.345 6.895 115.155 ;
        RECT 6.905 114.345 8.275 115.155 ;
        RECT 8.325 115.025 9.675 115.255 ;
        RECT 11.210 115.025 12.120 115.245 ;
        RECT 8.325 114.345 15.635 115.025 ;
        RECT 15.645 114.345 18.395 115.255 ;
        RECT 18.415 114.430 18.845 115.215 ;
        RECT 22.380 115.025 23.290 115.245 ;
        RECT 24.825 115.025 26.175 115.255 ;
        RECT 18.865 114.345 26.175 115.025 ;
        RECT 26.320 115.025 27.240 115.255 ;
        RECT 30.460 115.025 31.380 115.255 ;
        RECT 26.320 114.345 29.785 115.025 ;
        RECT 30.460 114.345 33.925 115.025 ;
        RECT 34.045 114.345 39.555 115.155 ;
        RECT 39.565 114.345 43.235 115.155 ;
        RECT 44.175 114.430 44.605 115.215 ;
        RECT 48.140 115.025 49.050 115.245 ;
        RECT 50.585 115.025 51.935 115.255 ;
        RECT 55.960 115.025 56.870 115.245 ;
        RECT 58.405 115.025 59.755 115.255 ;
        RECT 44.625 114.345 51.935 115.025 ;
        RECT 52.445 114.345 59.755 115.025 ;
        RECT 59.900 115.025 60.820 115.255 ;
        RECT 59.900 114.345 63.365 115.025 ;
        RECT 63.485 114.345 66.695 115.255 ;
        RECT 66.705 114.345 69.455 115.155 ;
        RECT 69.935 114.430 70.365 115.215 ;
        RECT 70.385 114.345 75.895 115.155 ;
        RECT 75.905 114.345 81.415 115.155 ;
        RECT 81.425 114.345 82.795 115.155 ;
        RECT 82.805 114.345 84.175 115.155 ;
        RECT 5.665 114.135 5.835 114.345 ;
        RECT 7.045 114.135 7.215 114.345 ;
        RECT 8.885 114.135 9.055 114.325 ;
        RECT 14.405 114.135 14.575 114.325 ;
        RECT 15.325 114.155 15.495 114.345 ;
        RECT 15.785 114.155 15.955 114.345 ;
        RECT 16.245 114.135 16.415 114.325 ;
        RECT 19.005 114.155 19.175 114.345 ;
        RECT 19.925 114.135 20.095 114.325 ;
        RECT 23.605 114.135 23.775 114.325 ;
        RECT 24.070 114.135 24.240 114.325 ;
        RECT 25.445 114.135 25.615 114.325 ;
        RECT 28.210 114.135 28.380 114.325 ;
        RECT 29.585 114.155 29.755 114.345 ;
        RECT 30.040 114.185 30.160 114.295 ;
        RECT 31.880 114.185 32.000 114.295 ;
        RECT 33.270 114.135 33.440 114.325 ;
        RECT 33.725 114.135 33.895 114.345 ;
        RECT 34.185 114.155 34.355 114.345 ;
        RECT 37.400 114.135 37.570 114.325 ;
        RECT 39.705 114.155 39.875 114.345 ;
        RECT 42.005 114.135 42.175 114.325 ;
        RECT 42.465 114.135 42.635 114.325 ;
        RECT 43.395 114.190 43.555 114.300 ;
        RECT 44.765 114.155 44.935 114.345 ;
        RECT 49.825 114.135 49.995 114.325 ;
        RECT 52.120 114.185 52.240 114.295 ;
        RECT 52.585 114.155 52.755 114.345 ;
        RECT 55.345 114.135 55.515 114.325 ;
        RECT 57.640 114.185 57.760 114.295 ;
        RECT 59.030 114.135 59.200 114.325 ;
        RECT 59.485 114.135 59.655 114.325 ;
        RECT 60.870 114.135 61.040 114.325 ;
        RECT 62.245 114.135 62.415 114.325 ;
        RECT 63.165 114.155 63.335 114.345 ;
        RECT 63.625 114.155 63.795 114.345 ;
        RECT 64.080 114.185 64.200 114.295 ;
        RECT 64.545 114.135 64.715 114.325 ;
        RECT 66.845 114.155 67.015 114.345 ;
        RECT 67.305 114.135 67.475 114.325 ;
        RECT 69.600 114.185 69.720 114.295 ;
        RECT 70.525 114.155 70.695 114.345 ;
        RECT 72.825 114.135 72.995 114.325 ;
        RECT 76.045 114.155 76.215 114.345 ;
        RECT 78.345 114.135 78.515 114.325 ;
        RECT 81.105 114.135 81.275 114.325 ;
        RECT 81.565 114.155 81.735 114.345 ;
        RECT 83.865 114.135 84.035 114.345 ;
        RECT 5.525 113.325 6.895 114.135 ;
        RECT 6.905 113.455 8.735 114.135 ;
        RECT 8.745 113.325 14.255 114.135 ;
        RECT 14.265 113.325 16.095 114.135 ;
        RECT 16.120 113.225 17.935 114.135 ;
        RECT 17.945 113.455 20.235 114.135 ;
        RECT 20.340 113.455 23.805 114.135 ;
        RECT 17.945 113.225 18.865 113.455 ;
        RECT 20.340 113.225 21.260 113.455 ;
        RECT 23.925 113.225 25.275 114.135 ;
        RECT 25.305 113.325 28.055 114.135 ;
        RECT 28.065 113.225 30.985 114.135 ;
        RECT 31.295 113.265 31.725 114.050 ;
        RECT 32.205 113.225 33.555 114.135 ;
        RECT 33.695 113.455 37.160 114.135 ;
        RECT 36.240 113.225 37.160 113.455 ;
        RECT 37.285 113.225 38.635 114.135 ;
        RECT 38.740 113.455 42.205 114.135 ;
        RECT 42.325 113.455 49.635 114.135 ;
        RECT 38.740 113.225 39.660 113.455 ;
        RECT 45.840 113.235 46.750 113.455 ;
        RECT 48.285 113.225 49.635 113.455 ;
        RECT 49.685 113.325 55.195 114.135 ;
        RECT 55.205 113.325 57.035 114.135 ;
        RECT 57.055 113.265 57.485 114.050 ;
        RECT 57.965 113.225 59.315 114.135 ;
        RECT 59.345 113.325 60.715 114.135 ;
        RECT 60.725 113.225 62.075 114.135 ;
        RECT 62.105 113.325 63.935 114.135 ;
        RECT 64.405 113.455 67.155 114.135 ;
        RECT 66.225 113.225 67.155 113.455 ;
        RECT 67.165 113.325 72.675 114.135 ;
        RECT 72.685 113.325 78.195 114.135 ;
        RECT 78.205 113.325 80.955 114.135 ;
        RECT 80.965 113.455 82.795 114.135 ;
        RECT 81.450 113.225 82.795 113.455 ;
        RECT 82.805 113.325 84.175 114.135 ;
      LAYER nwell ;
        RECT 5.330 110.105 84.370 112.935 ;
      LAYER pwell ;
        RECT 5.525 108.905 6.895 109.715 ;
        RECT 7.565 109.585 11.495 109.815 ;
        RECT 7.080 108.905 11.495 109.585 ;
        RECT 11.600 109.585 12.520 109.815 ;
        RECT 11.600 108.905 15.065 109.585 ;
        RECT 15.185 108.905 17.935 109.715 ;
        RECT 18.415 108.990 18.845 109.775 ;
        RECT 18.865 108.905 24.375 109.715 ;
        RECT 24.385 108.905 26.215 109.715 ;
        RECT 30.200 109.585 31.110 109.805 ;
        RECT 32.645 109.585 33.995 109.815 ;
        RECT 26.685 108.905 33.995 109.585 ;
        RECT 34.055 108.905 36.785 109.815 ;
        RECT 40.320 109.585 41.230 109.805 ;
        RECT 42.765 109.585 44.115 109.815 ;
        RECT 36.805 108.905 44.115 109.585 ;
        RECT 44.175 108.990 44.605 109.775 ;
        RECT 44.625 108.905 47.375 109.715 ;
        RECT 47.385 109.615 48.315 109.815 ;
        RECT 49.645 109.615 50.595 109.815 ;
        RECT 47.385 109.135 50.595 109.615 ;
        RECT 54.120 109.585 55.030 109.805 ;
        RECT 56.565 109.585 57.915 109.815 ;
        RECT 47.530 108.935 50.595 109.135 ;
        RECT 5.665 108.695 5.835 108.905 ;
        RECT 7.080 108.885 7.190 108.905 ;
        RECT 7.020 108.715 7.215 108.885 ;
        RECT 7.045 108.695 7.215 108.715 ;
        RECT 8.430 108.695 8.600 108.885 ;
        RECT 10.265 108.695 10.435 108.885 ;
        RECT 13.945 108.695 14.115 108.885 ;
        RECT 14.865 108.715 15.035 108.905 ;
        RECT 15.325 108.715 15.495 108.905 ;
        RECT 18.080 108.745 18.200 108.855 ;
        RECT 19.005 108.715 19.175 108.905 ;
        RECT 21.310 108.695 21.480 108.885 ;
        RECT 22.695 108.740 22.855 108.850 ;
        RECT 23.605 108.695 23.775 108.885 ;
        RECT 24.525 108.715 24.695 108.905 ;
        RECT 26.360 108.745 26.480 108.855 ;
        RECT 26.825 108.715 26.995 108.905 ;
        RECT 30.960 108.745 31.080 108.855 ;
        RECT 5.525 107.885 6.895 108.695 ;
        RECT 6.905 107.885 8.275 108.695 ;
        RECT 8.285 107.785 10.115 108.695 ;
        RECT 10.235 108.015 13.700 108.695 ;
        RECT 13.805 108.015 21.115 108.695 ;
        RECT 12.780 107.785 13.700 108.015 ;
        RECT 17.320 107.795 18.230 108.015 ;
        RECT 19.765 107.785 21.115 108.015 ;
        RECT 21.165 107.785 22.515 108.695 ;
        RECT 23.465 108.015 30.775 108.695 ;
        RECT 31.880 108.665 32.050 108.885 ;
        RECT 34.185 108.855 34.355 108.905 ;
        RECT 36.945 108.885 37.115 108.905 ;
        RECT 34.180 108.745 34.355 108.855 ;
        RECT 34.185 108.715 34.355 108.745 ;
        RECT 34.645 108.715 34.815 108.885 ;
        RECT 36.945 108.715 37.120 108.885 ;
        RECT 34.650 108.695 34.815 108.715 ;
        RECT 36.950 108.695 37.120 108.715 ;
        RECT 38.785 108.695 38.955 108.885 ;
        RECT 40.165 108.695 40.335 108.885 ;
        RECT 44.765 108.715 44.935 108.905 ;
        RECT 45.685 108.695 45.855 108.885 ;
        RECT 47.530 108.855 47.700 108.935 ;
        RECT 49.660 108.905 50.595 108.935 ;
        RECT 50.605 108.905 57.915 109.585 ;
        RECT 57.965 108.905 59.315 109.815 ;
        RECT 59.345 108.905 60.715 109.715 ;
        RECT 60.735 108.905 62.085 109.815 ;
        RECT 62.145 109.585 63.495 109.815 ;
        RECT 65.030 109.585 65.940 109.805 ;
        RECT 62.145 108.905 69.455 109.585 ;
        RECT 69.935 108.990 70.365 109.775 ;
        RECT 70.385 108.905 75.895 109.715 ;
        RECT 75.905 108.905 79.575 109.715 ;
        RECT 79.585 108.905 80.955 109.685 ;
        RECT 81.450 109.585 82.795 109.815 ;
        RECT 80.965 108.905 82.795 109.585 ;
        RECT 82.805 108.905 84.175 109.715 ;
        RECT 47.520 108.745 47.700 108.855 ;
        RECT 47.530 108.715 47.700 108.745 ;
        RECT 47.990 108.695 48.160 108.885 ;
        RECT 50.745 108.715 50.915 108.905 ;
        RECT 52.125 108.695 52.295 108.885 ;
        RECT 53.960 108.745 54.080 108.855 ;
        RECT 56.725 108.695 56.895 108.885 ;
        RECT 57.645 108.695 57.815 108.885 ;
        RECT 58.110 108.715 58.280 108.905 ;
        RECT 59.485 108.715 59.655 108.905 ;
        RECT 61.335 108.740 61.495 108.850 ;
        RECT 61.785 108.715 61.955 108.905 ;
        RECT 65.465 108.695 65.635 108.885 ;
        RECT 65.925 108.695 66.095 108.885 ;
        RECT 68.225 108.695 68.395 108.885 ;
        RECT 69.145 108.715 69.315 108.905 ;
        RECT 69.600 108.745 69.720 108.855 ;
        RECT 70.525 108.715 70.695 108.905 ;
        RECT 71.905 108.695 72.075 108.885 ;
        RECT 76.045 108.715 76.215 108.905 ;
        RECT 79.725 108.715 79.895 108.905 ;
        RECT 81.105 108.715 81.275 108.905 ;
        RECT 82.485 108.695 82.655 108.885 ;
        RECT 83.865 108.695 84.035 108.905 ;
        RECT 33.080 108.665 34.035 108.695 ;
        RECT 26.980 107.795 27.890 108.015 ;
        RECT 29.425 107.785 30.775 108.015 ;
        RECT 31.295 107.825 31.725 108.610 ;
        RECT 31.755 107.985 34.035 108.665 ;
        RECT 34.650 108.015 36.485 108.695 ;
        RECT 33.080 107.785 34.035 107.985 ;
        RECT 35.555 107.785 36.485 108.015 ;
        RECT 36.805 107.785 38.635 108.695 ;
        RECT 38.655 107.785 40.005 108.695 ;
        RECT 40.025 107.885 45.535 108.695 ;
        RECT 45.545 107.885 47.375 108.695 ;
        RECT 47.845 108.015 51.940 108.695 ;
        RECT 48.330 107.785 51.940 108.015 ;
        RECT 51.985 107.885 53.815 108.695 ;
        RECT 54.285 107.785 57.035 108.695 ;
        RECT 57.055 107.825 57.485 108.610 ;
        RECT 57.505 108.015 61.175 108.695 ;
        RECT 60.245 107.785 61.175 108.015 ;
        RECT 62.200 108.015 65.665 108.695 ;
        RECT 62.200 107.785 63.120 108.015 ;
        RECT 65.785 107.785 68.075 108.695 ;
        RECT 68.085 107.885 71.755 108.695 ;
        RECT 71.765 108.015 79.075 108.695 ;
        RECT 75.280 107.795 76.190 108.015 ;
        RECT 77.725 107.785 79.075 108.015 ;
        RECT 79.220 108.015 82.685 108.695 ;
        RECT 79.220 107.785 80.140 108.015 ;
        RECT 82.805 107.885 84.175 108.695 ;
      LAYER nwell ;
        RECT 5.330 104.665 84.370 107.495 ;
      LAYER pwell ;
        RECT 5.525 103.465 6.895 104.275 ;
        RECT 10.420 104.145 11.330 104.365 ;
        RECT 12.865 104.145 14.215 104.375 ;
        RECT 6.905 103.465 14.215 104.145 ;
        RECT 14.265 103.465 16.095 104.375 ;
        RECT 16.415 104.145 17.345 104.375 ;
        RECT 16.415 103.465 18.250 104.145 ;
        RECT 18.415 103.550 18.845 104.335 ;
        RECT 21.155 104.175 22.510 104.375 ;
        RECT 19.830 104.145 22.510 104.175 ;
        RECT 23.005 104.175 23.960 104.375 ;
        RECT 19.830 103.495 22.995 104.145 ;
        RECT 21.155 103.465 22.995 103.495 ;
        RECT 23.005 103.495 25.285 104.175 ;
        RECT 23.005 103.465 23.960 103.495 ;
        RECT 5.665 103.255 5.835 103.465 ;
        RECT 7.045 103.415 7.215 103.465 ;
        RECT 7.040 103.305 7.215 103.415 ;
        RECT 7.045 103.275 7.215 103.305 ;
        RECT 7.510 103.255 7.680 103.445 ;
        RECT 12.565 103.255 12.735 103.445 ;
        RECT 13.035 103.300 13.195 103.410 ;
        RECT 13.940 103.255 14.110 103.445 ;
        RECT 14.410 103.275 14.580 103.465 ;
        RECT 18.085 103.445 18.250 103.465 ;
        RECT 15.335 103.255 15.505 103.445 ;
        RECT 16.700 103.305 16.820 103.415 ;
        RECT 18.085 103.275 18.255 103.445 ;
        RECT 18.540 103.255 18.710 103.445 ;
        RECT 19.005 103.255 19.175 103.445 ;
        RECT 22.685 103.275 22.855 103.465 ;
        RECT 23.605 103.255 23.775 103.445 ;
        RECT 24.065 103.255 24.235 103.445 ;
        RECT 24.990 103.275 25.160 103.495 ;
        RECT 25.305 103.465 27.135 104.275 ;
        RECT 27.625 103.465 28.975 104.375 ;
        RECT 28.985 104.175 29.930 104.375 ;
        RECT 31.265 104.175 32.195 104.375 ;
        RECT 28.985 103.695 32.195 104.175 ;
        RECT 32.300 104.145 33.220 104.375 ;
        RECT 37.025 104.285 37.975 104.375 ;
        RECT 28.985 103.495 32.055 103.695 ;
        RECT 28.985 103.465 29.930 103.495 ;
        RECT 25.445 103.275 25.615 103.465 ;
        RECT 27.280 103.305 27.400 103.415 ;
        RECT 27.740 103.275 27.910 103.465 ;
        RECT 31.885 103.275 32.055 103.495 ;
        RECT 32.300 103.465 35.765 104.145 ;
        RECT 36.045 103.465 37.975 104.285 ;
        RECT 38.185 103.465 41.855 104.275 ;
        RECT 43.235 104.145 44.155 104.375 ;
        RECT 41.865 103.465 44.155 104.145 ;
        RECT 44.175 103.550 44.605 104.335 ;
        RECT 44.625 103.465 53.730 104.145 ;
        RECT 53.825 103.465 57.495 104.275 ;
        RECT 58.435 103.465 59.785 104.375 ;
        RECT 59.805 103.465 61.175 104.275 ;
        RECT 61.185 104.175 62.135 104.375 ;
        RECT 63.465 104.175 64.395 104.375 ;
        RECT 65.740 104.175 66.695 104.375 ;
        RECT 61.185 103.695 64.395 104.175 ;
        RECT 61.185 103.495 64.250 103.695 ;
        RECT 64.415 103.495 66.695 104.175 ;
        RECT 61.185 103.465 62.120 103.495 ;
        RECT 35.565 103.445 35.735 103.465 ;
        RECT 36.045 103.445 36.195 103.465 ;
        RECT 34.185 103.255 34.355 103.445 ;
        RECT 35.560 103.275 35.735 103.445 ;
        RECT 35.560 103.255 35.730 103.275 ;
        RECT 36.025 103.255 36.195 103.445 ;
        RECT 38.325 103.275 38.495 103.465 ;
        RECT 42.005 103.275 42.175 103.465 ;
        RECT 43.395 103.300 43.555 103.410 ;
        RECT 44.765 103.275 44.935 103.465 ;
        RECT 47.525 103.255 47.695 103.445 ;
        RECT 47.980 103.305 48.100 103.415 ;
        RECT 48.445 103.255 48.615 103.445 ;
        RECT 50.745 103.255 50.915 103.445 ;
        RECT 53.965 103.275 54.135 103.465 ;
        RECT 54.425 103.255 54.595 103.445 ;
        RECT 57.650 103.255 57.820 103.445 ;
        RECT 58.565 103.275 58.735 103.465 ;
        RECT 59.485 103.255 59.655 103.445 ;
        RECT 59.945 103.275 60.115 103.465 ;
        RECT 64.080 103.275 64.250 103.495 ;
        RECT 64.540 103.275 64.710 103.495 ;
        RECT 65.740 103.465 66.695 103.495 ;
        RECT 66.705 103.465 68.895 104.375 ;
        RECT 69.935 103.550 70.365 104.335 ;
        RECT 70.385 103.695 72.220 104.375 ;
        RECT 70.530 103.465 72.220 103.695 ;
        RECT 72.685 103.465 74.055 104.275 ;
        RECT 74.065 104.145 74.995 104.375 ;
        RECT 74.065 103.465 77.965 104.145 ;
        RECT 78.205 103.465 79.575 104.275 ;
        RECT 79.585 103.465 80.955 104.245 ;
        RECT 80.965 103.465 82.795 104.275 ;
        RECT 82.805 103.465 84.175 104.275 ;
        RECT 65.000 103.305 65.120 103.415 ;
        RECT 65.470 103.255 65.640 103.445 ;
        RECT 66.850 103.275 67.020 103.465 ;
        RECT 69.155 103.310 69.315 103.420 ;
        RECT 70.530 103.275 70.700 103.465 ;
        RECT 70.980 103.255 71.150 103.445 ;
        RECT 72.825 103.255 72.995 103.465 ;
        RECT 73.285 103.255 73.455 103.445 ;
        RECT 74.480 103.275 74.650 103.465 ;
        RECT 76.965 103.255 77.135 103.445 ;
        RECT 78.345 103.275 78.515 103.465 ;
        RECT 79.725 103.275 79.895 103.465 ;
        RECT 81.105 103.275 81.275 103.465 ;
        RECT 81.565 103.255 81.735 103.445 ;
        RECT 82.035 103.300 82.195 103.410 ;
        RECT 83.865 103.255 84.035 103.465 ;
        RECT 5.525 102.445 6.895 103.255 ;
        RECT 7.365 102.345 11.035 103.255 ;
        RECT 11.045 102.575 12.875 103.255 ;
        RECT 11.045 102.345 12.390 102.575 ;
        RECT 13.825 102.345 15.175 103.255 ;
        RECT 15.185 102.475 16.555 103.255 ;
        RECT 17.025 102.345 18.855 103.255 ;
        RECT 18.865 102.445 20.235 103.255 ;
        RECT 20.340 102.575 23.805 103.255 ;
        RECT 23.925 102.575 31.235 103.255 ;
        RECT 20.340 102.345 21.260 102.575 ;
        RECT 27.440 102.355 28.350 102.575 ;
        RECT 29.885 102.345 31.235 102.575 ;
        RECT 31.295 102.385 31.725 103.170 ;
        RECT 31.755 102.345 34.485 103.255 ;
        RECT 34.525 102.345 35.875 103.255 ;
        RECT 35.885 102.575 43.195 103.255 ;
        RECT 39.400 102.355 40.310 102.575 ;
        RECT 41.845 102.345 43.195 102.575 ;
        RECT 44.260 102.575 47.725 103.255 ;
        RECT 48.305 102.575 50.595 103.255 ;
        RECT 50.715 102.575 54.180 103.255 ;
        RECT 44.260 102.345 45.180 102.575 ;
        RECT 49.675 102.345 50.595 102.575 ;
        RECT 53.260 102.345 54.180 102.575 ;
        RECT 54.285 102.445 57.035 103.255 ;
        RECT 57.055 102.385 57.485 103.170 ;
        RECT 57.505 102.345 59.335 103.255 ;
        RECT 59.345 102.445 64.855 103.255 ;
        RECT 65.325 102.575 67.600 103.255 ;
        RECT 66.230 102.345 67.600 102.575 ;
        RECT 67.820 102.345 71.295 103.255 ;
        RECT 71.305 102.575 73.135 103.255 ;
        RECT 71.305 102.345 72.650 102.575 ;
        RECT 73.145 102.445 76.815 103.255 ;
        RECT 76.825 102.445 78.195 103.255 ;
        RECT 78.300 102.575 81.765 103.255 ;
        RECT 78.300 102.345 79.220 102.575 ;
        RECT 82.805 102.445 84.175 103.255 ;
      LAYER nwell ;
        RECT 5.330 99.225 84.370 102.055 ;
      LAYER pwell ;
        RECT 5.525 98.025 6.895 98.835 ;
        RECT 6.905 98.025 8.735 98.705 ;
        RECT 9.685 98.025 11.035 98.935 ;
        RECT 13.700 98.705 14.620 98.935 ;
        RECT 11.155 98.025 14.620 98.705 ;
        RECT 15.285 98.025 18.395 98.935 ;
        RECT 18.415 98.110 18.845 98.895 ;
        RECT 22.380 98.705 23.290 98.925 ;
        RECT 24.825 98.705 26.175 98.935 ;
        RECT 18.865 98.025 26.175 98.705 ;
        RECT 26.225 98.025 29.895 98.835 ;
        RECT 30.365 98.025 31.715 98.935 ;
        RECT 32.205 98.025 35.415 98.935 ;
        RECT 35.425 98.025 38.925 98.935 ;
        RECT 39.105 98.025 42.775 98.835 ;
        RECT 42.795 98.025 44.145 98.935 ;
        RECT 44.175 98.110 44.605 98.895 ;
        RECT 45.585 98.705 46.935 98.935 ;
        RECT 48.470 98.705 49.380 98.925 ;
        RECT 52.905 98.705 53.835 98.935 ;
        RECT 57.530 98.705 58.875 98.935 ;
        RECT 45.585 98.025 52.895 98.705 ;
        RECT 52.905 98.025 56.805 98.705 ;
        RECT 57.045 98.025 58.875 98.705 ;
        RECT 58.885 98.025 60.235 98.935 ;
        RECT 60.265 98.025 63.935 98.835 ;
        RECT 64.865 98.025 66.215 98.935 ;
        RECT 66.245 98.025 69.455 98.935 ;
        RECT 69.935 98.110 70.365 98.895 ;
        RECT 70.385 98.025 72.215 98.835 ;
        RECT 76.200 98.705 77.110 98.925 ;
        RECT 78.645 98.705 79.995 98.935 ;
        RECT 72.685 98.025 79.995 98.705 ;
        RECT 80.045 98.025 82.795 98.835 ;
        RECT 82.805 98.025 84.175 98.835 ;
        RECT 5.665 97.815 5.835 98.025 ;
        RECT 7.045 97.815 7.215 98.025 ;
        RECT 8.895 97.870 9.055 97.980 ;
        RECT 9.800 97.835 9.970 98.025 ;
        RECT 11.185 97.835 11.355 98.025 ;
        RECT 14.860 97.865 14.980 97.975 ;
        RECT 15.325 97.835 15.495 98.025 ;
        RECT 17.625 97.815 17.795 98.005 ;
        RECT 18.080 97.815 18.250 98.005 ;
        RECT 19.005 97.835 19.175 98.025 ;
        RECT 19.465 97.815 19.635 98.005 ;
        RECT 24.985 97.815 25.155 98.005 ;
        RECT 26.365 97.835 26.535 98.025 ;
        RECT 30.040 97.865 30.160 97.975 ;
        RECT 30.515 97.860 30.675 97.970 ;
        RECT 31.430 97.835 31.600 98.025 ;
        RECT 31.885 97.975 32.055 98.005 ;
        RECT 31.880 97.865 32.055 97.975 ;
        RECT 31.885 97.815 32.055 97.865 ;
        RECT 32.335 97.835 32.505 98.025 ;
        RECT 38.790 98.005 38.925 98.025 ;
        RECT 34.640 97.865 34.760 97.975 ;
        RECT 35.380 97.815 35.550 98.005 ;
        RECT 38.790 97.835 38.960 98.005 ;
        RECT 39.245 97.815 39.415 98.025 ;
        RECT 43.845 97.835 44.015 98.025 ;
        RECT 44.775 97.870 44.935 97.980 ;
        RECT 49.360 97.815 49.530 98.005 ;
        RECT 49.825 97.815 49.995 98.005 ;
        RECT 52.585 97.835 52.755 98.025 ;
        RECT 53.320 97.835 53.490 98.025 ;
        RECT 57.185 97.835 57.355 98.025 ;
        RECT 57.920 97.815 58.090 98.005 ;
        RECT 59.030 97.835 59.200 98.025 ;
        RECT 60.405 97.835 60.575 98.025 ;
        RECT 61.785 97.815 61.955 98.005 ;
        RECT 63.620 97.865 63.740 97.975 ;
        RECT 64.095 97.870 64.255 97.980 ;
        RECT 65.930 97.835 66.100 98.025 ;
        RECT 69.145 98.005 69.315 98.025 ;
        RECT 66.845 97.815 67.015 98.005 ;
        RECT 69.140 97.835 69.315 98.005 ;
        RECT 69.600 97.865 69.720 97.975 ;
        RECT 70.525 97.835 70.695 98.025 ;
        RECT 69.140 97.815 69.310 97.835 ;
        RECT 5.525 97.005 6.895 97.815 ;
        RECT 6.905 97.135 14.215 97.815 ;
        RECT 10.420 96.915 11.330 97.135 ;
        RECT 12.865 96.905 14.215 97.135 ;
        RECT 14.265 97.135 17.935 97.815 ;
        RECT 14.265 96.905 15.195 97.135 ;
        RECT 17.965 96.905 19.315 97.815 ;
        RECT 19.325 97.005 24.835 97.815 ;
        RECT 24.845 97.005 30.355 97.815 ;
        RECT 31.295 96.945 31.725 97.730 ;
        RECT 31.745 97.005 34.495 97.815 ;
        RECT 34.965 97.135 38.865 97.815 ;
        RECT 39.105 97.135 46.415 97.815 ;
        RECT 34.965 96.905 35.895 97.135 ;
        RECT 42.620 96.915 43.530 97.135 ;
        RECT 45.065 96.905 46.415 97.135 ;
        RECT 46.560 96.905 49.675 97.815 ;
        RECT 49.685 97.135 56.995 97.815 ;
        RECT 53.200 96.915 54.110 97.135 ;
        RECT 55.645 96.905 56.995 97.135 ;
        RECT 57.055 96.945 57.485 97.730 ;
        RECT 57.505 97.135 61.405 97.815 ;
        RECT 57.505 96.905 58.435 97.135 ;
        RECT 61.645 97.005 63.475 97.815 ;
        RECT 64.075 96.905 67.075 97.815 ;
        RECT 67.245 96.905 69.455 97.815 ;
        RECT 69.465 97.785 70.420 97.815 ;
        RECT 71.450 97.785 71.620 98.005 ;
        RECT 71.910 97.815 72.080 98.005 ;
        RECT 72.360 97.865 72.480 97.975 ;
        RECT 72.825 97.835 72.995 98.025 ;
        RECT 74.200 97.865 74.320 97.975 ;
        RECT 74.940 97.815 75.110 98.005 ;
        RECT 78.805 97.815 78.975 98.005 ;
        RECT 80.185 97.835 80.355 98.025 ;
        RECT 82.480 97.865 82.600 97.975 ;
        RECT 83.865 97.815 84.035 98.025 ;
        RECT 69.465 97.105 71.745 97.785 ;
        RECT 71.765 97.135 74.040 97.815 ;
        RECT 69.465 96.905 70.420 97.105 ;
        RECT 72.670 96.905 74.040 97.135 ;
        RECT 74.525 97.135 78.425 97.815 ;
        RECT 74.525 96.905 75.455 97.135 ;
        RECT 78.665 97.005 82.335 97.815 ;
        RECT 82.805 97.005 84.175 97.815 ;
      LAYER nwell ;
        RECT 5.330 93.785 84.370 96.615 ;
      LAYER pwell ;
        RECT 5.525 92.585 6.895 93.395 ;
        RECT 6.905 92.585 10.575 93.395 ;
        RECT 10.585 92.585 12.415 93.495 ;
        RECT 12.520 93.265 13.440 93.495 ;
        RECT 12.520 92.585 15.985 93.265 ;
        RECT 16.105 92.585 17.935 93.395 ;
        RECT 18.415 92.670 18.845 93.455 ;
        RECT 18.865 92.585 24.375 93.395 ;
        RECT 24.385 92.585 26.215 93.395 ;
        RECT 29.740 93.265 30.650 93.485 ;
        RECT 32.185 93.265 33.535 93.495 ;
        RECT 26.225 92.585 33.535 93.265 ;
        RECT 33.680 93.265 34.600 93.495 ;
        RECT 33.680 92.585 37.145 93.265 ;
        RECT 37.265 92.585 40.015 93.395 ;
        RECT 40.025 93.265 40.955 93.495 ;
        RECT 40.025 92.585 43.925 93.265 ;
        RECT 44.175 92.670 44.605 93.455 ;
        RECT 44.625 93.265 45.555 93.495 ;
        RECT 44.625 92.585 48.525 93.265 ;
        RECT 48.765 92.585 52.435 93.395 ;
        RECT 52.445 92.585 53.815 93.395 ;
        RECT 56.480 93.265 57.400 93.495 ;
        RECT 53.935 92.585 57.400 93.265 ;
        RECT 57.505 92.585 59.335 93.395 ;
        RECT 59.345 93.265 60.265 93.495 ;
        RECT 59.345 92.585 61.635 93.265 ;
        RECT 61.645 92.585 62.995 93.495 ;
        RECT 63.025 92.585 65.775 93.395 ;
        RECT 67.580 93.295 68.535 93.495 ;
        RECT 66.255 92.615 68.535 93.295 ;
        RECT 5.665 92.375 5.835 92.585 ;
        RECT 7.045 92.375 7.215 92.585 ;
        RECT 8.700 92.375 8.870 92.565 ;
        RECT 10.730 92.395 10.900 92.585 ;
        RECT 12.560 92.425 12.680 92.535 ;
        RECT 5.525 91.565 6.895 92.375 ;
        RECT 6.905 91.565 8.275 92.375 ;
        RECT 8.285 91.695 12.185 92.375 ;
        RECT 13.025 92.345 13.195 92.565 ;
        RECT 15.785 92.375 15.955 92.585 ;
        RECT 16.245 92.395 16.415 92.585 ;
        RECT 18.080 92.425 18.200 92.535 ;
        RECT 18.545 92.375 18.715 92.565 ;
        RECT 19.005 92.395 19.175 92.585 ;
        RECT 24.525 92.395 24.695 92.585 ;
        RECT 26.365 92.395 26.535 92.585 ;
        RECT 27.560 92.375 27.730 92.565 ;
        RECT 31.880 92.425 32.000 92.535 ;
        RECT 32.620 92.375 32.790 92.565 ;
        RECT 36.485 92.375 36.655 92.565 ;
        RECT 36.945 92.395 37.115 92.585 ;
        RECT 37.405 92.395 37.575 92.585 ;
        RECT 38.785 92.375 38.955 92.565 ;
        RECT 40.440 92.395 40.610 92.585 ;
        RECT 44.305 92.375 44.475 92.565 ;
        RECT 45.040 92.395 45.210 92.585 ;
        RECT 47.060 92.425 47.180 92.535 ;
        RECT 48.905 92.395 49.075 92.585 ;
        RECT 52.585 92.395 52.755 92.585 ;
        RECT 53.965 92.395 54.135 92.585 ;
        RECT 54.425 92.375 54.595 92.565 ;
        RECT 54.885 92.375 55.055 92.565 ;
        RECT 56.720 92.425 56.840 92.535 ;
        RECT 57.645 92.395 57.815 92.585 ;
        RECT 61.325 92.565 61.495 92.585 ;
        RECT 60.405 92.375 60.575 92.565 ;
        RECT 60.860 92.425 60.980 92.535 ;
        RECT 61.315 92.395 61.495 92.565 ;
        RECT 61.790 92.395 61.960 92.585 ;
        RECT 63.165 92.395 63.335 92.585 ;
        RECT 61.315 92.375 61.485 92.395 ;
        RECT 64.545 92.375 64.715 92.565 ;
        RECT 65.920 92.425 66.040 92.535 ;
        RECT 14.225 92.345 15.605 92.375 ;
        RECT 8.285 91.465 9.215 91.695 ;
        RECT 12.900 91.665 15.605 92.345 ;
        RECT 14.225 91.465 15.605 91.665 ;
        RECT 15.645 91.565 18.395 92.375 ;
        RECT 18.405 91.695 26.135 92.375 ;
        RECT 21.920 91.475 22.830 91.695 ;
        RECT 24.365 91.465 26.135 91.695 ;
        RECT 27.145 91.695 31.045 92.375 ;
        RECT 27.145 91.465 28.075 91.695 ;
        RECT 31.295 91.505 31.725 92.290 ;
        RECT 32.205 91.695 36.105 92.375 ;
        RECT 36.345 91.695 38.635 92.375 ;
        RECT 32.205 91.465 33.135 91.695 ;
        RECT 37.715 91.465 38.635 91.695 ;
        RECT 38.645 91.565 44.155 92.375 ;
        RECT 44.165 91.565 46.915 92.375 ;
        RECT 47.425 91.695 54.735 92.375 ;
        RECT 47.425 91.465 48.775 91.695 ;
        RECT 50.310 91.475 51.220 91.695 ;
        RECT 54.745 91.565 56.575 92.375 ;
        RECT 57.055 91.505 57.485 92.290 ;
        RECT 57.505 91.465 60.715 92.375 ;
        RECT 61.185 91.465 64.395 92.375 ;
        RECT 64.405 91.565 66.235 92.375 ;
        RECT 66.380 92.345 66.550 92.615 ;
        RECT 67.580 92.585 68.535 92.615 ;
        RECT 68.545 92.585 69.915 93.395 ;
        RECT 69.935 92.670 70.365 93.455 ;
        RECT 74.505 93.265 75.435 93.495 ;
        RECT 71.535 92.585 75.435 93.265 ;
        RECT 75.445 92.585 80.955 93.395 ;
        RECT 80.965 92.585 82.795 93.395 ;
        RECT 82.805 92.585 84.175 93.395 ;
        RECT 68.685 92.395 68.855 92.585 ;
        RECT 70.535 92.430 70.695 92.540 ;
        RECT 70.995 92.420 71.155 92.530 ;
        RECT 68.690 92.375 68.855 92.395 ;
        RECT 71.905 92.375 72.075 92.565 ;
        RECT 74.850 92.395 75.020 92.585 ;
        RECT 75.125 92.375 75.295 92.565 ;
        RECT 75.585 92.395 75.755 92.585 ;
        RECT 80.645 92.375 80.815 92.565 ;
        RECT 81.105 92.395 81.275 92.585 ;
        RECT 82.480 92.425 82.600 92.535 ;
        RECT 83.865 92.375 84.035 92.585 ;
        RECT 67.580 92.345 68.535 92.375 ;
        RECT 66.255 91.665 68.535 92.345 ;
        RECT 68.690 91.695 70.525 92.375 ;
        RECT 67.580 91.465 68.535 91.665 ;
        RECT 69.595 91.465 70.525 91.695 ;
        RECT 71.765 91.465 74.975 92.375 ;
        RECT 74.985 91.565 80.495 92.375 ;
        RECT 80.505 91.565 82.335 92.375 ;
        RECT 82.805 91.565 84.175 92.375 ;
      LAYER nwell ;
        RECT 5.330 88.345 84.370 91.175 ;
      LAYER pwell ;
        RECT 5.525 87.145 6.895 87.955 ;
        RECT 10.420 87.825 11.330 88.045 ;
        RECT 12.865 87.825 14.635 88.055 ;
        RECT 17.015 87.825 17.935 88.055 ;
        RECT 6.905 87.145 14.635 87.825 ;
        RECT 15.645 87.145 17.935 87.825 ;
        RECT 18.415 87.230 18.845 88.015 ;
        RECT 19.325 87.825 20.255 88.055 ;
        RECT 19.325 87.145 23.225 87.825 ;
        RECT 23.465 87.145 28.975 87.955 ;
        RECT 28.985 87.145 32.655 87.955 ;
        RECT 35.320 87.825 36.240 88.055 ;
        RECT 32.775 87.145 36.240 87.825 ;
        RECT 36.345 87.145 38.175 87.955 ;
        RECT 41.365 87.855 42.315 88.055 ;
        RECT 38.645 87.175 42.315 87.855 ;
        RECT 5.665 86.935 5.835 87.145 ;
        RECT 7.045 86.935 7.215 87.145 ;
        RECT 8.880 86.985 9.000 87.095 ;
        RECT 5.525 86.125 6.895 86.935 ;
        RECT 6.905 86.125 8.735 86.935 ;
        RECT 9.205 86.905 10.160 86.935 ;
        RECT 11.190 86.905 11.360 87.125 ;
        RECT 11.645 86.935 11.815 87.125 ;
        RECT 14.875 86.990 15.035 87.100 ;
        RECT 15.785 86.955 15.955 87.145 ;
        RECT 19.005 87.095 19.175 87.125 ;
        RECT 18.080 86.985 18.200 87.095 ;
        RECT 19.000 86.985 19.175 87.095 ;
        RECT 19.005 86.935 19.175 86.985 ;
        RECT 19.740 86.955 19.910 87.145 ;
        RECT 21.305 86.935 21.475 87.125 ;
        RECT 23.605 86.955 23.775 87.145 ;
        RECT 24.065 86.935 24.235 87.125 ;
        RECT 29.125 86.955 29.295 87.145 ;
        RECT 32.160 86.935 32.330 87.125 ;
        RECT 32.805 86.955 32.975 87.145 ;
        RECT 36.025 86.935 36.195 87.125 ;
        RECT 36.485 86.955 36.655 87.145 ;
        RECT 37.870 86.935 38.040 87.125 ;
        RECT 38.320 86.985 38.440 87.095 ;
        RECT 38.790 86.955 38.960 87.175 ;
        RECT 41.365 87.145 42.315 87.175 ;
        RECT 42.325 87.145 44.155 87.955 ;
        RECT 44.175 87.230 44.605 88.015 ;
        RECT 44.625 87.145 50.135 87.955 ;
        RECT 50.145 87.145 55.655 87.955 ;
        RECT 55.665 87.145 59.335 87.955 ;
        RECT 59.445 87.145 61.635 88.055 ;
        RECT 61.645 87.145 63.475 87.955 ;
        RECT 64.855 87.825 65.775 88.055 ;
        RECT 63.485 87.145 65.775 87.825 ;
        RECT 65.785 87.145 69.455 87.955 ;
        RECT 69.935 87.230 70.365 88.015 ;
        RECT 70.385 87.145 72.595 88.055 ;
        RECT 72.695 87.145 74.045 88.055 ;
        RECT 74.065 87.145 77.735 87.955 ;
        RECT 77.745 87.145 79.115 87.955 ;
        RECT 79.220 87.825 80.140 88.055 ;
        RECT 79.220 87.145 82.685 87.825 ;
        RECT 82.805 87.145 84.175 87.955 ;
        RECT 42.465 86.955 42.635 87.145 ;
        RECT 9.205 86.225 11.485 86.905 ;
        RECT 11.505 86.255 18.815 86.935 ;
        RECT 18.865 86.255 21.155 86.935 ;
        RECT 9.205 86.025 10.160 86.225 ;
        RECT 15.020 86.035 15.930 86.255 ;
        RECT 17.465 86.025 18.815 86.255 ;
        RECT 20.235 86.025 21.155 86.255 ;
        RECT 21.165 86.125 23.915 86.935 ;
        RECT 23.925 86.255 31.235 86.935 ;
        RECT 27.440 86.035 28.350 86.255 ;
        RECT 29.885 86.025 31.235 86.255 ;
        RECT 31.295 86.065 31.725 86.850 ;
        RECT 31.745 86.255 35.645 86.935 ;
        RECT 31.745 86.025 32.675 86.255 ;
        RECT 35.885 86.125 37.715 86.935 ;
        RECT 37.725 86.025 41.200 86.935 ;
        RECT 41.405 86.905 42.340 86.935 ;
        RECT 44.300 86.905 44.470 87.125 ;
        RECT 44.765 86.955 44.935 87.145 ;
        RECT 47.065 86.935 47.235 87.125 ;
        RECT 47.525 86.935 47.695 87.125 ;
        RECT 49.365 86.935 49.535 87.125 ;
        RECT 50.285 86.955 50.455 87.145 ;
        RECT 55.805 86.955 55.975 87.145 ;
        RECT 56.720 86.985 56.840 87.095 ;
        RECT 57.650 86.935 57.820 87.125 ;
        RECT 61.320 87.090 61.490 87.145 ;
        RECT 61.320 86.980 61.495 87.090 ;
        RECT 61.320 86.955 61.490 86.980 ;
        RECT 61.785 86.955 61.955 87.145 ;
        RECT 62.245 86.935 62.415 87.125 ;
        RECT 63.625 86.955 63.795 87.145 ;
        RECT 65.010 86.935 65.180 87.125 ;
        RECT 65.925 86.955 66.095 87.145 ;
        RECT 66.845 86.935 67.015 87.125 ;
        RECT 69.600 86.985 69.720 87.095 ;
        RECT 70.065 86.935 70.235 87.125 ;
        RECT 70.530 86.955 70.700 87.145 ;
        RECT 73.280 86.985 73.400 87.095 ;
        RECT 73.745 86.935 73.915 87.145 ;
        RECT 74.205 86.955 74.375 87.145 ;
        RECT 77.885 86.955 78.055 87.145 ;
        RECT 81.105 86.935 81.275 87.125 ;
        RECT 82.485 86.955 82.655 87.145 ;
        RECT 83.865 86.935 84.035 87.145 ;
        RECT 41.405 86.705 44.470 86.905 ;
        RECT 41.405 86.225 44.615 86.705 ;
        RECT 41.405 86.025 42.355 86.225 ;
        RECT 43.685 86.025 44.615 86.225 ;
        RECT 44.625 86.255 47.375 86.935 ;
        RECT 44.625 86.025 45.555 86.255 ;
        RECT 47.385 86.125 49.215 86.935 ;
        RECT 49.225 86.255 56.535 86.935 ;
        RECT 52.740 86.035 53.650 86.255 ;
        RECT 55.185 86.025 56.535 86.255 ;
        RECT 57.055 86.065 57.485 86.850 ;
        RECT 57.505 86.025 61.175 86.935 ;
        RECT 62.105 86.255 64.855 86.935 ;
        RECT 63.925 86.025 64.855 86.255 ;
        RECT 64.865 86.025 66.695 86.935 ;
        RECT 66.705 86.125 69.455 86.935 ;
        RECT 69.925 86.025 73.135 86.935 ;
        RECT 73.605 86.255 80.915 86.935 ;
        RECT 80.965 86.255 82.795 86.935 ;
        RECT 77.120 86.035 78.030 86.255 ;
        RECT 79.565 86.025 80.915 86.255 ;
        RECT 81.450 86.025 82.795 86.255 ;
        RECT 82.805 86.125 84.175 86.935 ;
      LAYER nwell ;
        RECT 5.330 82.905 84.370 85.735 ;
      LAYER pwell ;
        RECT 5.525 81.705 6.895 82.515 ;
        RECT 6.905 81.705 10.575 82.515 ;
        RECT 10.585 81.705 11.955 82.515 ;
        RECT 13.015 82.385 13.945 82.615 ;
        RECT 12.110 81.705 13.945 82.385 ;
        RECT 14.465 82.525 15.415 82.615 ;
        RECT 14.465 81.705 16.395 82.525 ;
        RECT 17.035 81.705 18.385 82.615 ;
        RECT 18.415 81.790 18.845 82.575 ;
        RECT 23.300 82.385 24.210 82.605 ;
        RECT 25.745 82.385 27.515 82.615 ;
        RECT 19.785 81.705 27.515 82.385 ;
        RECT 27.605 81.705 31.275 82.515 ;
        RECT 32.300 82.385 33.220 82.615 ;
        RECT 35.885 82.415 36.815 82.615 ;
        RECT 38.145 82.415 39.095 82.615 ;
        RECT 32.300 81.705 35.765 82.385 ;
        RECT 35.885 81.935 39.095 82.415 ;
        RECT 36.030 81.735 39.095 81.935 ;
        RECT 5.665 81.495 5.835 81.705 ;
        RECT 7.045 81.495 7.215 81.705 ;
        RECT 10.725 81.515 10.895 81.705 ;
        RECT 12.110 81.685 12.275 81.705 ;
        RECT 16.245 81.685 16.395 81.705 ;
        RECT 12.105 81.515 12.275 81.685 ;
        RECT 12.565 81.495 12.735 81.685 ;
        RECT 16.245 81.515 16.415 81.685 ;
        RECT 16.700 81.545 16.820 81.655 ;
        RECT 17.165 81.515 17.335 81.705 ;
        RECT 18.085 81.495 18.255 81.685 ;
        RECT 19.015 81.550 19.175 81.660 ;
        RECT 19.925 81.655 20.095 81.705 ;
        RECT 19.920 81.545 20.095 81.655 ;
        RECT 19.925 81.515 20.095 81.545 ;
        RECT 20.660 81.495 20.830 81.685 ;
        RECT 24.525 81.495 24.695 81.685 ;
        RECT 27.745 81.515 27.915 81.705 ;
        RECT 30.045 81.495 30.215 81.685 ;
        RECT 31.435 81.550 31.595 81.660 ;
        RECT 31.885 81.495 32.055 81.685 ;
        RECT 35.565 81.515 35.735 81.705 ;
        RECT 36.030 81.515 36.200 81.735 ;
        RECT 38.160 81.705 39.095 81.735 ;
        RECT 40.025 82.385 40.955 82.615 ;
        RECT 40.025 81.705 42.775 82.385 ;
        RECT 42.785 81.705 44.155 82.515 ;
        RECT 44.175 81.790 44.605 82.575 ;
        RECT 44.625 82.385 45.555 82.615 ;
        RECT 52.740 82.385 53.650 82.605 ;
        RECT 55.185 82.385 56.535 82.615 ;
        RECT 44.625 81.705 48.525 82.385 ;
        RECT 49.225 81.705 56.535 82.385 ;
        RECT 56.585 81.705 59.795 82.615 ;
        RECT 60.115 82.385 61.045 82.615 ;
        RECT 60.115 81.705 61.950 82.385 ;
        RECT 62.105 81.705 63.455 82.615 ;
        RECT 63.485 81.705 64.855 82.515 ;
        RECT 64.865 81.705 66.695 82.615 ;
        RECT 68.675 82.385 69.605 82.615 ;
        RECT 67.770 81.705 69.605 82.385 ;
        RECT 69.935 81.790 70.365 82.575 ;
        RECT 70.535 81.705 74.190 82.615 ;
        RECT 75.445 82.385 76.375 82.615 ;
        RECT 75.445 81.705 79.345 82.385 ;
        RECT 79.585 81.705 80.955 82.485 ;
        RECT 80.965 81.705 82.795 82.515 ;
        RECT 82.805 81.705 84.175 82.515 ;
        RECT 39.255 81.550 39.415 81.660 ;
        RECT 5.525 80.685 6.895 81.495 ;
        RECT 6.905 80.685 12.415 81.495 ;
        RECT 12.425 80.685 17.935 81.495 ;
        RECT 17.945 80.685 19.775 81.495 ;
        RECT 20.245 80.815 24.145 81.495 ;
        RECT 20.245 80.585 21.175 80.815 ;
        RECT 24.385 80.685 29.895 81.495 ;
        RECT 29.905 80.685 31.275 81.495 ;
        RECT 31.295 80.625 31.725 81.410 ;
        RECT 31.745 80.815 39.055 81.495 ;
        RECT 35.260 80.595 36.170 80.815 ;
        RECT 37.705 80.585 39.055 80.815 ;
        RECT 39.105 81.465 40.050 81.495 ;
        RECT 41.540 81.465 41.710 81.685 ;
        RECT 42.000 81.545 42.120 81.655 ;
        RECT 42.465 81.495 42.635 81.705 ;
        RECT 42.925 81.515 43.095 81.705 ;
        RECT 45.040 81.515 45.210 81.705 ;
        RECT 48.900 81.545 49.020 81.655 ;
        RECT 49.365 81.515 49.535 81.705 ;
        RECT 53.045 81.495 53.215 81.685 ;
        RECT 53.505 81.495 53.675 81.685 ;
        RECT 56.715 81.515 56.885 81.705 ;
        RECT 61.785 81.685 61.950 81.705 ;
        RECT 57.655 81.540 57.815 81.650 ;
        RECT 39.105 80.785 41.855 81.465 ;
        RECT 42.325 80.815 49.635 81.495 ;
        RECT 39.105 80.585 40.050 80.785 ;
        RECT 45.840 80.595 46.750 80.815 ;
        RECT 48.285 80.585 49.635 80.815 ;
        RECT 49.780 80.815 53.245 81.495 ;
        RECT 49.780 80.585 50.700 80.815 ;
        RECT 53.365 80.685 57.035 81.495 ;
        RECT 58.570 81.465 58.740 81.685 ;
        RECT 61.785 81.515 61.955 81.685 ;
        RECT 63.170 81.515 63.340 81.705 ;
        RECT 63.625 81.515 63.795 81.705 ;
        RECT 64.085 81.495 64.255 81.685 ;
        RECT 64.545 81.495 64.715 81.685 ;
        RECT 65.010 81.515 65.180 81.705 ;
        RECT 67.770 81.685 67.935 81.705 ;
        RECT 70.535 81.685 70.695 81.705 ;
        RECT 66.855 81.550 67.015 81.660 ;
        RECT 67.765 81.515 67.935 81.685 ;
        RECT 69.145 81.495 69.315 81.685 ;
        RECT 69.605 81.495 69.775 81.685 ;
        RECT 70.525 81.515 70.695 81.685 ;
        RECT 74.675 81.550 74.835 81.660 ;
        RECT 75.125 81.495 75.295 81.685 ;
        RECT 75.860 81.515 76.030 81.705 ;
        RECT 77.885 81.495 78.055 81.685 ;
        RECT 79.725 81.515 79.895 81.705 ;
        RECT 81.105 81.515 81.275 81.705 ;
        RECT 82.485 81.495 82.655 81.685 ;
        RECT 83.865 81.495 84.035 81.705 ;
        RECT 60.700 81.465 61.635 81.495 ;
        RECT 57.055 80.625 57.485 81.410 ;
        RECT 58.570 81.265 61.635 81.465 ;
        RECT 58.425 80.785 61.635 81.265 ;
        RECT 58.425 80.585 59.355 80.785 ;
        RECT 60.685 80.585 61.635 80.785 ;
        RECT 61.645 80.815 64.395 81.495 ;
        RECT 61.645 80.585 62.575 80.815 ;
        RECT 64.405 80.685 67.155 81.495 ;
        RECT 67.165 80.815 69.455 81.495 ;
        RECT 67.165 80.585 68.085 80.815 ;
        RECT 69.465 80.685 74.975 81.495 ;
        RECT 74.985 80.685 77.735 81.495 ;
        RECT 77.745 80.715 79.115 81.495 ;
        RECT 79.220 80.815 82.685 81.495 ;
        RECT 79.220 80.585 80.140 80.815 ;
        RECT 82.805 80.685 84.175 81.495 ;
      LAYER nwell ;
        RECT 5.330 77.465 84.370 80.295 ;
      LAYER pwell ;
        RECT 9.405 77.085 10.355 77.175 ;
        RECT 5.525 76.265 6.895 77.075 ;
        RECT 6.905 76.265 8.735 77.075 ;
        RECT 9.405 76.265 11.335 77.085 ;
        RECT 11.505 76.265 12.855 77.175 ;
        RECT 12.885 76.265 14.235 77.175 ;
        RECT 15.185 76.975 16.115 77.175 ;
        RECT 17.450 76.975 18.395 77.175 ;
        RECT 15.185 76.495 18.395 76.975 ;
        RECT 15.325 76.295 18.395 76.495 ;
        RECT 18.415 76.350 18.845 77.135 ;
        RECT 5.665 76.055 5.835 76.265 ;
        RECT 7.045 76.075 7.215 76.265 ;
        RECT 11.185 76.245 11.335 76.265 ;
        RECT 7.965 76.055 8.135 76.245 ;
        RECT 8.880 76.105 9.000 76.215 ;
        RECT 11.185 76.075 11.355 76.245 ;
        RECT 12.570 76.075 12.740 76.265 ;
        RECT 13.030 76.075 13.200 76.265 ;
        RECT 14.415 76.110 14.575 76.220 ;
        RECT 15.325 76.055 15.495 76.295 ;
        RECT 17.450 76.265 18.395 76.295 ;
        RECT 18.865 76.265 20.235 77.075 ;
        RECT 20.245 76.945 21.175 77.175 ;
        RECT 20.245 76.265 24.145 76.945 ;
        RECT 24.385 76.265 29.895 77.075 ;
        RECT 34.025 76.945 34.955 77.175 ;
        RECT 31.055 76.265 34.955 76.945 ;
        RECT 34.965 76.265 36.795 77.075 ;
        RECT 36.900 76.945 37.820 77.175 ;
        RECT 43.140 76.945 44.060 77.175 ;
        RECT 36.900 76.265 40.365 76.945 ;
        RECT 40.595 76.265 44.060 76.945 ;
        RECT 44.175 76.350 44.605 77.135 ;
        RECT 44.625 76.945 45.545 77.175 ;
        RECT 46.925 76.945 47.855 77.175 ;
        RECT 44.625 76.265 46.915 76.945 ;
        RECT 46.925 76.265 50.825 76.945 ;
        RECT 51.065 76.265 56.575 77.075 ;
        RECT 59.240 76.945 60.160 77.175 ;
        RECT 61.635 76.945 62.555 77.175 ;
        RECT 56.695 76.265 60.160 76.945 ;
        RECT 60.265 76.265 62.555 76.945 ;
        RECT 62.565 76.265 65.315 77.075 ;
        RECT 65.935 76.265 69.590 77.175 ;
        RECT 69.935 76.350 70.365 77.135 ;
        RECT 70.385 76.265 73.595 77.175 ;
        RECT 77.120 76.945 78.030 77.165 ;
        RECT 79.565 76.945 80.915 77.175 ;
        RECT 81.450 76.945 82.795 77.175 ;
        RECT 73.605 76.265 80.915 76.945 ;
        RECT 80.965 76.265 82.795 76.945 ;
        RECT 82.805 76.265 84.175 77.075 ;
        RECT 5.525 75.245 6.895 76.055 ;
        RECT 7.825 75.375 15.135 76.055 ;
        RECT 11.340 75.155 12.250 75.375 ;
        RECT 13.785 75.145 15.135 75.375 ;
        RECT 15.185 75.245 17.015 76.055 ;
        RECT 17.165 76.025 17.335 76.245 ;
        RECT 19.005 76.075 19.175 76.265 ;
        RECT 20.380 76.105 20.500 76.215 ;
        RECT 20.660 76.075 20.830 76.265 ;
        RECT 20.845 76.055 21.015 76.245 ;
        RECT 24.525 76.075 24.695 76.265 ;
        RECT 28.665 76.055 28.835 76.245 ;
        RECT 30.055 76.110 30.215 76.220 ;
        RECT 31.885 76.055 32.055 76.245 ;
        RECT 34.370 76.075 34.540 76.265 ;
        RECT 35.105 76.075 35.275 76.265 ;
        RECT 39.240 76.105 39.360 76.215 ;
        RECT 40.165 76.075 40.335 76.265 ;
        RECT 40.625 76.075 40.795 76.265 ;
        RECT 46.605 76.055 46.775 76.265 ;
        RECT 47.065 76.055 47.235 76.245 ;
        RECT 47.340 76.075 47.510 76.265 ;
        RECT 51.205 76.075 51.375 76.265 ;
        RECT 56.725 76.055 56.895 76.265 ;
        RECT 57.645 76.055 57.815 76.245 ;
        RECT 60.405 76.075 60.575 76.265 ;
        RECT 60.870 76.055 61.040 76.245 ;
        RECT 62.705 76.075 62.875 76.265 ;
        RECT 65.935 76.245 66.095 76.265 ;
        RECT 64.095 76.100 64.255 76.210 ;
        RECT 65.460 76.105 65.580 76.215 ;
        RECT 65.925 76.075 66.095 76.245 ;
        RECT 67.305 76.055 67.475 76.245 ;
        RECT 70.065 76.055 70.235 76.245 ;
        RECT 70.525 76.055 70.695 76.265 ;
        RECT 73.745 76.075 73.915 76.265 ;
        RECT 74.205 76.055 74.375 76.245 ;
        RECT 75.860 76.055 76.030 76.245 ;
        RECT 79.725 76.055 79.895 76.245 ;
        RECT 81.105 76.055 81.275 76.265 ;
        RECT 83.865 76.055 84.035 76.265 ;
        RECT 19.290 76.025 20.235 76.055 ;
        RECT 17.165 75.825 20.235 76.025 ;
        RECT 17.025 75.345 20.235 75.825 ;
        RECT 20.705 75.375 28.435 76.055 ;
        RECT 17.025 75.145 17.955 75.345 ;
        RECT 19.290 75.145 20.235 75.345 ;
        RECT 24.220 75.155 25.130 75.375 ;
        RECT 26.665 75.145 28.435 75.375 ;
        RECT 28.525 75.245 31.275 76.055 ;
        RECT 31.295 75.185 31.725 75.970 ;
        RECT 31.745 75.375 39.055 76.055 ;
        RECT 35.260 75.155 36.170 75.375 ;
        RECT 37.705 75.145 39.055 75.375 ;
        RECT 39.605 75.375 46.915 76.055 ;
        RECT 39.605 75.145 40.955 75.375 ;
        RECT 42.490 75.155 43.400 75.375 ;
        RECT 46.925 75.245 49.675 76.055 ;
        RECT 49.725 75.375 57.035 76.055 ;
        RECT 49.725 75.145 51.075 75.375 ;
        RECT 52.610 75.155 53.520 75.375 ;
        RECT 57.055 75.185 57.485 75.970 ;
        RECT 57.585 75.145 60.585 76.055 ;
        RECT 60.725 75.145 63.645 76.055 ;
        RECT 64.875 75.145 67.605 76.055 ;
        RECT 67.635 75.145 70.365 76.055 ;
        RECT 70.385 75.245 74.055 76.055 ;
        RECT 74.065 75.245 75.435 76.055 ;
        RECT 75.445 75.375 79.345 76.055 ;
        RECT 75.445 75.145 76.375 75.375 ;
        RECT 79.585 75.275 80.955 76.055 ;
        RECT 80.965 75.245 82.795 76.055 ;
        RECT 82.805 75.245 84.175 76.055 ;
      LAYER nwell ;
        RECT 5.330 72.025 84.370 74.855 ;
      LAYER pwell ;
        RECT 5.525 70.825 6.895 71.635 ;
        RECT 6.905 70.825 8.735 71.635 ;
        RECT 9.055 71.505 9.985 71.735 ;
        RECT 11.505 71.535 12.435 71.735 ;
        RECT 13.765 71.535 14.715 71.735 ;
        RECT 9.055 70.825 10.890 71.505 ;
        RECT 11.505 71.055 14.715 71.535 ;
        RECT 15.185 71.535 16.115 71.735 ;
        RECT 17.450 71.535 18.395 71.735 ;
        RECT 15.185 71.055 18.395 71.535 ;
        RECT 5.665 70.615 5.835 70.825 ;
        RECT 7.045 70.775 7.215 70.825 ;
        RECT 10.725 70.805 10.890 70.825 ;
        RECT 11.650 70.855 14.715 71.055 ;
        RECT 7.040 70.665 7.215 70.775 ;
        RECT 7.045 70.635 7.215 70.665 ;
        RECT 7.780 70.615 7.950 70.805 ;
        RECT 10.725 70.635 10.895 70.805 ;
        RECT 11.180 70.665 11.300 70.775 ;
        RECT 11.650 70.635 11.820 70.855 ;
        RECT 13.780 70.825 14.715 70.855 ;
        RECT 15.325 70.855 18.395 71.055 ;
        RECT 18.415 70.910 18.845 71.695 ;
        RECT 11.920 70.615 12.090 70.805 ;
        RECT 14.860 70.665 14.980 70.775 ;
        RECT 15.325 70.635 15.495 70.855 ;
        RECT 17.450 70.825 18.395 70.855 ;
        RECT 18.865 70.825 20.695 71.635 ;
        RECT 24.680 71.505 25.590 71.725 ;
        RECT 27.125 71.505 28.895 71.735 ;
        RECT 21.165 70.825 28.895 71.505 ;
        RECT 28.985 70.825 32.655 71.635 ;
        RECT 34.505 71.505 35.435 71.735 ;
        RECT 38.645 71.505 39.575 71.735 ;
        RECT 33.130 70.825 34.495 71.505 ;
        RECT 34.505 70.825 38.405 71.505 ;
        RECT 38.645 70.825 42.545 71.505 ;
        RECT 42.785 70.825 44.155 71.635 ;
        RECT 44.175 70.910 44.605 71.695 ;
        RECT 44.625 71.505 45.555 71.735 ;
        RECT 49.265 71.505 50.615 71.735 ;
        RECT 52.150 71.505 53.060 71.725 ;
        RECT 59.240 71.505 60.160 71.735 ;
        RECT 44.625 70.825 48.525 71.505 ;
        RECT 49.265 70.825 56.575 71.505 ;
        RECT 56.695 70.825 60.160 71.505 ;
        RECT 60.265 70.825 63.475 71.735 ;
        RECT 64.625 71.645 65.575 71.735 ;
        RECT 63.645 70.825 65.575 71.645 ;
        RECT 65.785 70.825 67.135 71.735 ;
        RECT 68.110 71.505 69.455 71.735 ;
        RECT 67.625 70.825 69.455 71.505 ;
        RECT 69.935 70.910 70.365 71.695 ;
        RECT 70.385 70.825 73.135 71.635 ;
        RECT 77.120 71.505 78.030 71.725 ;
        RECT 79.565 71.505 80.915 71.735 ;
        RECT 81.450 71.505 82.795 71.735 ;
        RECT 73.605 70.825 80.915 71.505 ;
        RECT 80.965 70.825 82.795 71.505 ;
        RECT 82.805 70.825 84.175 71.635 ;
        RECT 15.795 70.660 15.955 70.770 ;
        RECT 19.005 70.635 19.175 70.825 ;
        RECT 20.110 70.615 20.280 70.805 ;
        RECT 20.845 70.775 21.015 70.805 ;
        RECT 20.840 70.665 21.015 70.775 ;
        RECT 20.845 70.615 21.015 70.665 ;
        RECT 21.305 70.635 21.475 70.825 ;
        RECT 25.905 70.615 26.075 70.805 ;
        RECT 29.125 70.635 29.295 70.825 ;
        RECT 31.895 70.660 32.055 70.770 ;
        RECT 32.805 70.615 32.975 70.805 ;
        RECT 34.920 70.635 35.090 70.825 ;
        RECT 37.865 70.615 38.035 70.805 ;
        RECT 39.060 70.635 39.230 70.825 ;
        RECT 40.625 70.615 40.795 70.805 ;
        RECT 42.925 70.635 43.095 70.825 ;
        RECT 45.040 70.635 45.210 70.825 ;
        RECT 48.260 70.615 48.430 70.805 ;
        RECT 48.900 70.665 49.020 70.775 ;
        RECT 55.345 70.615 55.515 70.805 ;
        RECT 55.805 70.615 55.975 70.805 ;
        RECT 56.265 70.635 56.435 70.825 ;
        RECT 56.725 70.635 56.895 70.825 ;
        RECT 57.645 70.635 57.815 70.805 ;
        RECT 60.405 70.635 60.575 70.825 ;
        RECT 63.645 70.805 63.795 70.825 ;
        RECT 61.790 70.615 61.960 70.805 ;
        RECT 63.170 70.615 63.340 70.805 ;
        RECT 63.625 70.635 63.795 70.805 ;
        RECT 64.540 70.615 64.710 70.805 ;
        RECT 65.015 70.660 65.175 70.770 ;
        RECT 65.925 70.615 66.095 70.805 ;
        RECT 66.850 70.635 67.020 70.825 ;
        RECT 67.300 70.665 67.420 70.775 ;
        RECT 67.765 70.635 67.935 70.825 ;
        RECT 69.600 70.665 69.720 70.775 ;
        RECT 70.525 70.635 70.695 70.825 ;
        RECT 72.360 70.615 72.530 70.805 ;
        RECT 72.825 70.615 72.995 70.805 ;
        RECT 73.280 70.665 73.400 70.775 ;
        RECT 73.745 70.635 73.915 70.825 ;
        RECT 74.660 70.665 74.780 70.775 ;
        RECT 75.400 70.615 75.570 70.805 ;
        RECT 81.105 70.635 81.275 70.825 ;
        RECT 82.485 70.615 82.655 70.805 ;
        RECT 83.865 70.615 84.035 70.825 ;
        RECT 5.525 69.805 6.895 70.615 ;
        RECT 7.365 69.935 11.265 70.615 ;
        RECT 11.505 69.935 15.405 70.615 ;
        RECT 16.795 69.935 20.695 70.615 ;
        RECT 20.705 69.935 25.520 70.615 ;
        RECT 7.365 69.705 8.295 69.935 ;
        RECT 11.505 69.705 12.435 69.935 ;
        RECT 19.765 69.705 20.695 69.935 ;
        RECT 25.765 69.805 31.275 70.615 ;
        RECT 31.295 69.745 31.725 70.530 ;
        RECT 32.665 69.935 37.480 70.615 ;
        RECT 37.725 69.805 40.475 70.615 ;
        RECT 40.485 69.935 47.795 70.615 ;
        RECT 44.000 69.715 44.910 69.935 ;
        RECT 46.445 69.705 47.795 69.935 ;
        RECT 47.845 69.935 51.745 70.615 ;
        RECT 52.080 69.935 55.545 70.615 ;
        RECT 47.845 69.705 48.775 69.935 ;
        RECT 52.080 69.705 53.000 69.935 ;
        RECT 55.665 69.805 57.035 70.615 ;
        RECT 57.055 69.745 57.485 70.530 ;
        RECT 57.910 69.935 60.335 70.615 ;
        RECT 60.725 69.705 62.075 70.615 ;
        RECT 62.105 69.705 63.455 70.615 ;
        RECT 63.505 69.705 64.855 70.615 ;
        RECT 65.785 69.705 68.995 70.615 ;
        RECT 69.200 69.705 72.675 70.615 ;
        RECT 72.685 69.805 74.515 70.615 ;
        RECT 74.985 69.935 78.885 70.615 ;
        RECT 79.220 69.935 82.685 70.615 ;
        RECT 74.985 69.705 75.915 69.935 ;
        RECT 79.220 69.705 80.140 69.935 ;
        RECT 82.805 69.805 84.175 70.615 ;
      LAYER nwell ;
        RECT 5.330 66.585 84.370 69.415 ;
      LAYER pwell ;
        RECT 5.525 65.385 6.895 66.195 ;
        RECT 10.420 66.065 11.330 66.285 ;
        RECT 12.865 66.065 14.635 66.295 ;
        RECT 6.905 65.385 14.635 66.065 ;
        RECT 14.725 65.385 18.395 66.195 ;
        RECT 18.415 65.470 18.845 66.255 ;
        RECT 22.380 66.065 23.290 66.285 ;
        RECT 24.825 66.065 26.595 66.295 ;
        RECT 18.865 65.385 26.595 66.065 ;
        RECT 26.685 65.385 28.515 66.195 ;
        RECT 28.525 66.065 29.455 66.295 ;
        RECT 36.180 66.065 37.090 66.285 ;
        RECT 38.625 66.065 39.975 66.295 ;
        RECT 28.525 65.385 32.425 66.065 ;
        RECT 32.665 65.385 39.975 66.065 ;
        RECT 40.025 66.065 40.955 66.295 ;
        RECT 40.025 65.385 43.925 66.065 ;
        RECT 44.175 65.470 44.605 66.255 ;
        RECT 44.720 66.065 45.640 66.295 ;
        RECT 44.720 65.385 48.185 66.065 ;
        RECT 48.305 65.385 51.975 66.195 ;
        RECT 60.620 66.065 61.540 66.295 ;
        RECT 52.905 65.385 57.720 66.065 ;
        RECT 58.075 65.385 61.540 66.065 ;
        RECT 61.845 66.205 62.795 66.295 ;
        RECT 61.845 65.385 63.775 66.205 ;
        RECT 63.955 65.385 65.305 66.295 ;
        RECT 65.345 65.385 66.695 66.295 ;
        RECT 68.040 66.095 68.995 66.295 ;
        RECT 66.715 65.415 68.995 66.095 ;
        RECT 69.935 65.470 70.365 66.255 ;
        RECT 5.665 65.175 5.835 65.385 ;
        RECT 7.045 65.195 7.215 65.385 ;
        RECT 8.425 65.175 8.595 65.365 ;
        RECT 8.895 65.220 9.055 65.330 ;
        RECT 9.805 65.175 9.975 65.365 ;
        RECT 14.865 65.195 15.035 65.385 ;
        RECT 19.005 65.195 19.175 65.385 ;
        RECT 21.030 65.175 21.200 65.365 ;
        RECT 21.765 65.175 21.935 65.365 ;
        RECT 26.825 65.195 26.995 65.385 ;
        RECT 27.285 65.175 27.455 65.365 ;
        RECT 28.940 65.195 29.110 65.385 ;
        RECT 30.960 65.225 31.080 65.335 ;
        RECT 31.880 65.225 32.000 65.335 ;
        RECT 32.805 65.195 32.975 65.385 ;
        RECT 35.565 65.175 35.735 65.365 ;
        RECT 38.795 65.175 38.965 65.365 ;
        RECT 39.245 65.175 39.415 65.365 ;
        RECT 40.440 65.195 40.610 65.385 ;
        RECT 43.845 65.175 44.015 65.365 ;
        RECT 44.315 65.220 44.475 65.330 ;
        RECT 45.500 65.175 45.670 65.365 ;
        RECT 47.985 65.195 48.155 65.385 ;
        RECT 48.445 65.195 48.615 65.385 ;
        RECT 52.135 65.230 52.295 65.340 ;
        RECT 53.045 65.195 53.215 65.385 ;
        RECT 56.265 65.175 56.435 65.365 ;
        RECT 56.720 65.225 56.840 65.335 ;
        RECT 57.920 65.175 58.090 65.365 ;
        RECT 58.105 65.195 58.275 65.385 ;
        RECT 63.625 65.365 63.775 65.385 ;
        RECT 65.005 65.365 65.175 65.385 ;
        RECT 61.785 65.175 61.955 65.365 ;
        RECT 63.625 65.195 63.795 65.365 ;
        RECT 64.540 65.225 64.660 65.335 ;
        RECT 65.000 65.195 65.175 65.365 ;
        RECT 65.460 65.195 65.630 65.385 ;
        RECT 66.840 65.195 67.010 65.415 ;
        RECT 68.040 65.385 68.995 65.415 ;
        RECT 71.305 65.385 74.515 66.295 ;
        RECT 74.525 65.385 77.275 66.195 ;
        RECT 77.285 66.065 78.630 66.295 ;
        RECT 79.220 66.065 80.140 66.295 ;
        RECT 77.285 65.385 79.115 66.065 ;
        RECT 79.220 65.385 82.685 66.065 ;
        RECT 82.805 65.385 84.175 66.195 ;
        RECT 70.520 65.340 70.690 65.365 ;
        RECT 69.155 65.230 69.315 65.340 ;
        RECT 70.520 65.230 70.695 65.340 ;
        RECT 5.525 64.365 6.895 65.175 ;
        RECT 6.905 64.495 8.735 65.175 ;
        RECT 9.665 64.495 17.395 65.175 ;
        RECT 17.715 64.495 21.615 65.175 ;
        RECT 6.905 64.265 8.250 64.495 ;
        RECT 13.180 64.275 14.090 64.495 ;
        RECT 15.625 64.265 17.395 64.495 ;
        RECT 20.685 64.265 21.615 64.495 ;
        RECT 21.625 64.365 27.135 65.175 ;
        RECT 27.145 64.365 30.815 65.175 ;
        RECT 31.295 64.305 31.725 65.090 ;
        RECT 32.300 64.495 35.765 65.175 ;
        RECT 32.300 64.265 33.220 64.495 ;
        RECT 35.885 64.265 39.095 65.175 ;
        RECT 39.105 64.365 40.475 65.175 ;
        RECT 40.580 64.495 44.045 65.175 ;
        RECT 45.085 64.495 48.985 65.175 ;
        RECT 49.265 64.495 56.575 65.175 ;
        RECT 40.580 64.265 41.500 64.495 ;
        RECT 45.085 64.265 46.015 64.495 ;
        RECT 49.265 64.265 50.615 64.495 ;
        RECT 52.150 64.275 53.060 64.495 ;
        RECT 57.055 64.305 57.485 65.090 ;
        RECT 57.505 64.495 61.405 65.175 ;
        RECT 57.505 64.265 58.435 64.495 ;
        RECT 61.645 64.365 64.395 65.175 ;
        RECT 65.000 65.145 65.170 65.195 ;
        RECT 70.520 65.175 70.690 65.230 ;
        RECT 70.985 65.175 71.155 65.365 ;
        RECT 71.445 65.195 71.615 65.385 ;
        RECT 74.205 65.175 74.375 65.365 ;
        RECT 74.665 65.195 74.835 65.385 ;
        RECT 78.805 65.195 78.975 65.385 ;
        RECT 82.485 65.175 82.655 65.385 ;
        RECT 83.865 65.175 84.035 65.385 ;
        RECT 66.200 65.145 67.155 65.175 ;
        RECT 64.875 64.465 67.155 65.145 ;
        RECT 66.200 64.265 67.155 64.465 ;
        RECT 67.360 64.265 70.835 65.175 ;
        RECT 70.845 64.265 74.055 65.175 ;
        RECT 74.065 64.495 81.375 65.175 ;
        RECT 77.580 64.275 78.490 64.495 ;
        RECT 80.025 64.265 81.375 64.495 ;
        RECT 81.425 64.395 82.795 65.175 ;
        RECT 82.805 64.365 84.175 65.175 ;
      LAYER nwell ;
        RECT 5.330 61.145 84.370 63.975 ;
      LAYER pwell ;
        RECT 5.525 59.945 6.895 60.755 ;
        RECT 6.905 60.625 8.250 60.855 ;
        RECT 8.745 60.625 10.090 60.855 ;
        RECT 6.905 59.945 8.735 60.625 ;
        RECT 8.745 59.945 10.575 60.625 ;
        RECT 10.585 59.945 11.955 60.755 ;
        RECT 11.965 60.625 13.310 60.855 ;
        RECT 11.965 59.945 13.795 60.625 ;
        RECT 13.805 59.945 17.475 60.755 ;
        RECT 18.415 60.030 18.845 60.815 ;
        RECT 18.865 59.945 22.340 60.855 ;
        RECT 23.595 60.625 24.525 60.855 ;
        RECT 22.690 59.945 24.525 60.625 ;
        RECT 24.845 59.945 26.675 60.755 ;
        RECT 30.200 60.625 31.110 60.845 ;
        RECT 32.645 60.625 33.995 60.855 ;
        RECT 26.685 59.945 33.995 60.625 ;
        RECT 34.045 59.945 36.795 60.755 ;
        RECT 36.805 60.625 37.735 60.855 ;
        RECT 36.805 59.945 40.705 60.625 ;
        RECT 41.415 59.945 44.155 60.625 ;
        RECT 44.175 60.030 44.605 60.815 ;
        RECT 48.140 60.625 49.050 60.845 ;
        RECT 50.585 60.625 51.935 60.855 ;
        RECT 44.625 59.945 51.935 60.625 ;
        RECT 52.080 60.625 53.000 60.855 ;
        RECT 58.320 60.625 59.240 60.855 ;
        RECT 52.080 59.945 55.545 60.625 ;
        RECT 55.775 59.945 59.240 60.625 ;
        RECT 59.345 59.945 61.175 60.855 ;
        RECT 68.675 60.625 69.605 60.855 ;
        RECT 62.105 59.945 66.920 60.625 ;
        RECT 67.770 59.945 69.605 60.625 ;
        RECT 69.935 60.030 70.365 60.815 ;
        RECT 70.385 59.945 72.215 60.755 ;
        RECT 74.880 60.625 75.800 60.855 ;
        RECT 72.335 59.945 75.800 60.625 ;
        RECT 75.905 60.625 76.835 60.855 ;
        RECT 81.450 60.625 82.795 60.855 ;
        RECT 75.905 59.945 79.805 60.625 ;
        RECT 80.965 59.945 82.795 60.625 ;
        RECT 82.805 59.945 84.175 60.755 ;
        RECT 5.665 59.735 5.835 59.945 ;
        RECT 7.045 59.735 7.215 59.925 ;
        RECT 8.425 59.755 8.595 59.945 ;
        RECT 10.265 59.755 10.435 59.945 ;
        RECT 8.430 59.735 8.595 59.755 ;
        RECT 10.725 59.735 10.895 59.945 ;
        RECT 13.485 59.755 13.655 59.945 ;
        RECT 13.945 59.755 14.115 59.945 ;
        RECT 16.270 59.755 16.440 59.925 ;
        RECT 16.270 59.735 16.380 59.755 ;
        RECT 16.705 59.735 16.875 59.925 ;
        RECT 17.635 59.790 17.795 59.900 ;
        RECT 19.010 59.755 19.180 59.945 ;
        RECT 22.690 59.925 22.855 59.945 ;
        RECT 22.685 59.755 22.855 59.925 ;
        RECT 24.065 59.735 24.235 59.925 ;
        RECT 24.985 59.755 25.155 59.945 ;
        RECT 26.825 59.755 26.995 59.945 ;
        RECT 31.885 59.735 32.055 59.925 ;
        RECT 34.185 59.755 34.355 59.945 ;
        RECT 34.645 59.735 34.815 59.925 ;
        RECT 37.220 59.755 37.390 59.945 ;
        RECT 41.080 59.785 41.200 59.895 ;
        RECT 42.005 59.735 42.175 59.925 ;
        RECT 43.845 59.755 44.015 59.945 ;
        RECT 44.765 59.755 44.935 59.945 ;
        RECT 47.250 59.735 47.420 59.925 ;
        RECT 47.985 59.735 48.155 59.925 ;
        RECT 55.345 59.755 55.515 59.945 ;
        RECT 55.805 59.755 55.975 59.945 ;
        RECT 56.725 59.735 56.895 59.925 ;
        RECT 60.405 59.735 60.575 59.925 ;
        RECT 60.860 59.755 61.030 59.945 ;
        RECT 62.245 59.925 62.415 59.945 ;
        RECT 67.770 59.925 67.935 59.945 ;
        RECT 61.335 59.790 61.495 59.900 ;
        RECT 61.790 59.735 61.960 59.925 ;
        RECT 62.245 59.755 62.420 59.925 ;
        RECT 67.300 59.785 67.420 59.895 ;
        RECT 67.765 59.755 67.935 59.925 ;
        RECT 70.525 59.755 70.695 59.945 ;
        RECT 72.365 59.755 72.535 59.945 ;
        RECT 62.250 59.735 62.420 59.755 ;
        RECT 73.280 59.735 73.450 59.925 ;
        RECT 74.675 59.780 74.835 59.890 ;
        RECT 75.860 59.735 76.030 59.925 ;
        RECT 76.320 59.755 76.490 59.945 ;
        RECT 80.195 59.790 80.355 59.900 ;
        RECT 80.645 59.735 80.815 59.925 ;
        RECT 81.105 59.735 81.275 59.945 ;
        RECT 83.865 59.735 84.035 59.945 ;
        RECT 5.525 58.925 6.895 59.735 ;
        RECT 6.905 58.925 8.275 59.735 ;
        RECT 8.430 59.055 10.265 59.735 ;
        RECT 9.335 58.825 10.265 59.055 ;
        RECT 10.585 58.925 11.955 59.735 ;
        RECT 11.965 59.055 16.380 59.735 ;
        RECT 16.565 59.055 23.875 59.735 ;
        RECT 23.925 59.055 31.235 59.735 ;
        RECT 11.965 58.825 15.895 59.055 ;
        RECT 20.080 58.835 20.990 59.055 ;
        RECT 22.525 58.825 23.875 59.055 ;
        RECT 27.440 58.835 28.350 59.055 ;
        RECT 29.885 58.825 31.235 59.055 ;
        RECT 31.295 58.865 31.725 59.650 ;
        RECT 31.745 58.925 34.495 59.735 ;
        RECT 34.505 59.055 41.815 59.735 ;
        RECT 38.020 58.835 38.930 59.055 ;
        RECT 40.465 58.825 41.815 59.055 ;
        RECT 41.865 58.925 43.695 59.735 ;
        RECT 43.935 59.055 47.835 59.735 ;
        RECT 46.905 58.825 47.835 59.055 ;
        RECT 47.845 58.925 49.675 59.735 ;
        RECT 49.725 59.055 57.035 59.735 ;
        RECT 49.725 58.825 51.075 59.055 ;
        RECT 52.610 58.835 53.520 59.055 ;
        RECT 57.055 58.865 57.485 59.650 ;
        RECT 57.505 58.825 60.715 59.735 ;
        RECT 60.725 58.825 62.075 59.735 ;
        RECT 62.105 58.825 73.115 59.735 ;
        RECT 73.165 58.825 74.515 59.735 ;
        RECT 75.445 59.055 79.345 59.735 ;
        RECT 75.445 58.825 76.375 59.055 ;
        RECT 79.585 58.955 80.955 59.735 ;
        RECT 80.965 59.055 82.795 59.735 ;
        RECT 81.450 58.825 82.795 59.055 ;
        RECT 82.805 58.925 84.175 59.735 ;
      LAYER nwell ;
        RECT 5.330 55.705 84.370 58.535 ;
      LAYER pwell ;
        RECT 5.525 54.505 6.895 55.315 ;
        RECT 6.905 55.185 8.250 55.415 ;
        RECT 12.260 55.185 13.170 55.405 ;
        RECT 14.705 55.185 16.055 55.415 ;
        RECT 6.905 54.505 8.735 55.185 ;
        RECT 8.745 54.505 16.055 55.185 ;
        RECT 16.105 54.505 17.935 55.315 ;
        RECT 18.415 54.590 18.845 55.375 ;
        RECT 19.915 55.185 20.845 55.415 ;
        RECT 19.010 54.505 20.845 55.185 ;
        RECT 21.820 54.505 25.295 55.415 ;
        RECT 25.305 54.505 27.135 55.315 ;
        RECT 30.660 55.185 31.570 55.405 ;
        RECT 33.105 55.185 34.455 55.415 ;
        RECT 27.145 54.505 34.455 55.185 ;
        RECT 34.505 55.185 35.435 55.415 ;
        RECT 42.305 55.185 43.235 55.415 ;
        RECT 34.505 54.505 38.405 55.185 ;
        RECT 39.335 54.505 43.235 55.185 ;
        RECT 44.175 54.590 44.605 55.375 ;
        RECT 44.625 54.505 48.295 55.315 ;
        RECT 48.305 55.185 49.235 55.415 ;
        RECT 48.305 54.505 52.205 55.185 ;
        RECT 52.445 54.505 57.955 55.315 ;
        RECT 57.965 54.505 61.175 55.415 ;
        RECT 61.205 54.505 62.555 55.415 ;
        RECT 62.565 54.505 65.485 55.415 ;
        RECT 65.935 54.505 69.590 55.415 ;
        RECT 69.935 54.590 70.365 55.375 ;
        RECT 70.385 54.505 73.595 55.415 ;
        RECT 77.580 55.185 78.490 55.405 ;
        RECT 80.025 55.185 81.375 55.415 ;
        RECT 74.065 54.505 81.375 55.185 ;
        RECT 81.425 54.505 82.795 55.285 ;
        RECT 82.805 54.505 84.175 55.315 ;
        RECT 5.665 54.295 5.835 54.505 ;
        RECT 8.425 54.485 8.595 54.505 ;
        RECT 7.045 54.295 7.215 54.485 ;
        RECT 8.425 54.315 8.600 54.485 ;
        RECT 8.885 54.315 9.055 54.505 ;
        RECT 8.430 54.295 8.600 54.315 ;
        RECT 12.110 54.295 12.280 54.485 ;
        RECT 16.245 54.315 16.415 54.505 ;
        RECT 19.010 54.485 19.175 54.505 ;
        RECT 18.080 54.345 18.200 54.455 ;
        RECT 18.555 54.295 18.725 54.485 ;
        RECT 19.005 54.315 19.175 54.485 ;
        RECT 21.300 54.345 21.420 54.455 ;
        RECT 22.220 54.295 22.390 54.485 ;
        RECT 22.685 54.295 22.855 54.485 ;
        RECT 24.980 54.315 25.150 54.505 ;
        RECT 25.445 54.315 25.615 54.505 ;
        RECT 27.285 54.315 27.455 54.505 ;
        RECT 30.045 54.295 30.215 54.485 ;
        RECT 32.160 54.295 32.330 54.485 ;
        RECT 34.920 54.315 35.090 54.505 ;
        RECT 38.780 54.345 38.900 54.455 ;
        RECT 39.245 54.295 39.415 54.485 ;
        RECT 39.695 54.295 39.865 54.485 ;
        RECT 42.650 54.315 42.820 54.505 ;
        RECT 42.925 54.295 43.095 54.485 ;
        RECT 43.395 54.350 43.555 54.460 ;
        RECT 44.765 54.315 44.935 54.505 ;
        RECT 45.040 54.295 45.210 54.485 ;
        RECT 48.720 54.315 48.890 54.505 ;
        RECT 52.125 54.295 52.295 54.485 ;
        RECT 52.585 54.455 52.755 54.505 ;
        RECT 52.580 54.345 52.755 54.455 ;
        RECT 52.585 54.315 52.755 54.345 ;
        RECT 56.265 54.295 56.435 54.485 ;
        RECT 56.720 54.345 56.840 54.455 ;
        RECT 57.645 54.295 57.815 54.485 ;
        RECT 60.865 54.315 61.035 54.505 ;
        RECT 61.320 54.315 61.490 54.505 ;
        RECT 62.710 54.485 62.880 54.505 ;
        RECT 65.935 54.485 66.095 54.505 ;
        RECT 62.700 54.315 62.880 54.485 ;
        RECT 62.700 54.295 62.870 54.315 ;
        RECT 64.540 54.295 64.710 54.485 ;
        RECT 65.015 54.340 65.175 54.450 ;
        RECT 65.925 54.315 66.095 54.485 ;
        RECT 69.140 54.295 69.310 54.485 ;
        RECT 70.525 54.315 70.695 54.505 ;
        RECT 71.905 54.315 72.075 54.485 ;
        RECT 72.360 54.345 72.480 54.455 ;
        RECT 71.905 54.295 71.925 54.315 ;
        RECT 72.825 54.295 72.995 54.485 ;
        RECT 73.740 54.345 73.860 54.455 ;
        RECT 74.205 54.315 74.375 54.505 ;
        RECT 80.195 54.340 80.355 54.450 ;
        RECT 81.105 54.295 81.275 54.485 ;
        RECT 82.485 54.315 82.655 54.505 ;
        RECT 83.865 54.295 84.035 54.505 ;
        RECT 5.525 53.485 6.895 54.295 ;
        RECT 6.905 53.485 8.275 54.295 ;
        RECT 8.285 53.385 11.760 54.295 ;
        RECT 11.965 53.385 15.440 54.295 ;
        RECT 15.645 53.385 18.855 54.295 ;
        RECT 19.060 53.385 22.535 54.295 ;
        RECT 22.545 53.615 29.855 54.295 ;
        RECT 26.060 53.395 26.970 53.615 ;
        RECT 28.505 53.385 29.855 53.615 ;
        RECT 29.905 53.485 31.275 54.295 ;
        RECT 31.295 53.425 31.725 54.210 ;
        RECT 31.745 53.615 35.645 54.295 ;
        RECT 35.980 53.615 39.445 54.295 ;
        RECT 31.745 53.385 32.675 53.615 ;
        RECT 35.980 53.385 36.900 53.615 ;
        RECT 39.565 53.385 42.775 54.295 ;
        RECT 42.785 53.485 44.615 54.295 ;
        RECT 44.625 53.615 48.525 54.295 ;
        RECT 48.860 53.615 52.325 54.295 ;
        RECT 53.000 53.615 56.465 54.295 ;
        RECT 44.625 53.385 45.555 53.615 ;
        RECT 48.860 53.385 49.780 53.615 ;
        RECT 53.000 53.385 53.920 53.615 ;
        RECT 57.055 53.425 57.485 54.210 ;
        RECT 57.615 53.615 61.080 54.295 ;
        RECT 60.160 53.385 61.080 53.615 ;
        RECT 61.185 53.385 63.015 54.295 ;
        RECT 63.025 53.385 64.855 54.295 ;
        RECT 65.870 53.615 69.455 54.295 ;
        RECT 68.535 53.385 69.455 53.615 ;
        RECT 69.475 53.615 71.925 54.295 ;
        RECT 72.685 53.615 79.995 54.295 ;
        RECT 80.965 53.615 82.795 54.295 ;
        RECT 69.475 53.385 71.435 53.615 ;
        RECT 76.200 53.395 77.110 53.615 ;
        RECT 78.645 53.385 79.995 53.615 ;
        RECT 81.450 53.385 82.795 53.615 ;
        RECT 82.805 53.485 84.175 54.295 ;
      LAYER nwell ;
        RECT 5.330 50.265 84.370 53.095 ;
      LAYER pwell ;
        RECT 5.525 49.065 6.895 49.875 ;
        RECT 7.955 49.745 8.885 49.975 ;
        RECT 12.720 49.745 13.630 49.965 ;
        RECT 15.165 49.745 16.515 49.975 ;
        RECT 7.050 49.065 8.885 49.745 ;
        RECT 9.205 49.065 16.515 49.745 ;
        RECT 16.565 49.065 18.395 49.875 ;
        RECT 18.415 49.150 18.845 49.935 ;
        RECT 18.865 49.065 23.680 49.745 ;
        RECT 23.925 49.065 27.135 49.975 ;
        RECT 27.145 49.065 32.655 49.875 ;
        RECT 32.665 49.065 38.175 49.875 ;
        RECT 38.185 49.065 40.935 49.875 ;
        RECT 40.945 49.065 44.155 49.975 ;
        RECT 44.175 49.150 44.605 49.935 ;
        RECT 49.060 49.745 49.970 49.965 ;
        RECT 51.505 49.745 52.855 49.975 ;
        RECT 45.545 49.065 52.855 49.745 ;
        RECT 52.945 49.745 54.295 49.975 ;
        RECT 55.830 49.745 56.740 49.965 ;
        RECT 60.305 49.745 61.655 49.975 ;
        RECT 63.190 49.745 64.100 49.965 ;
        RECT 52.945 49.065 60.255 49.745 ;
        RECT 60.305 49.065 67.615 49.745 ;
        RECT 67.645 49.065 68.995 49.975 ;
        RECT 69.935 49.150 70.365 49.935 ;
        RECT 70.480 49.745 71.400 49.975 ;
        RECT 74.525 49.745 75.455 49.975 ;
        RECT 78.760 49.745 79.680 49.975 ;
        RECT 70.480 49.065 73.945 49.745 ;
        RECT 74.525 49.065 78.425 49.745 ;
        RECT 78.760 49.065 82.225 49.745 ;
        RECT 82.805 49.065 84.175 49.875 ;
        RECT 5.665 48.855 5.835 49.065 ;
        RECT 7.050 49.045 7.215 49.065 ;
        RECT 7.045 48.875 7.215 49.045 ;
        RECT 8.425 48.855 8.595 49.045 ;
        RECT 9.345 48.875 9.515 49.065 ;
        RECT 10.265 48.855 10.435 49.045 ;
        RECT 10.725 48.855 10.895 49.045 ;
        RECT 16.240 48.905 16.360 49.015 ;
        RECT 16.705 48.875 16.875 49.065 ;
        RECT 19.005 48.875 19.175 49.065 ;
        RECT 16.710 48.855 16.875 48.875 ;
        RECT 23.605 48.855 23.775 49.045 ;
        RECT 24.065 48.875 24.235 49.045 ;
        RECT 24.070 48.855 24.235 48.875 ;
        RECT 26.365 48.855 26.535 49.045 ;
        RECT 26.835 48.875 27.005 49.065 ;
        RECT 27.285 48.875 27.455 49.065 ;
        RECT 30.965 48.875 31.135 49.045 ;
        RECT 31.880 48.905 32.000 49.015 ;
        RECT 32.335 48.855 32.505 49.045 ;
        RECT 32.805 48.875 32.975 49.065 ;
        RECT 35.560 48.905 35.680 49.015 ;
        RECT 36.025 48.855 36.195 49.045 ;
        RECT 38.325 48.875 38.495 49.065 ;
        RECT 41.075 48.875 41.245 49.065 ;
        RECT 43.385 48.855 43.555 49.045 ;
        RECT 44.775 48.910 44.935 49.020 ;
        RECT 45.685 48.875 45.855 49.065 ;
        RECT 51.020 48.855 51.190 49.045 ;
        RECT 54.885 48.855 55.055 49.045 ;
        RECT 56.720 48.905 56.840 49.015 ;
        RECT 57.645 48.855 57.815 49.045 ;
        RECT 59.945 48.875 60.115 49.065 ;
        RECT 63.165 48.855 63.335 49.045 ;
        RECT 67.305 48.875 67.475 49.065 ;
        RECT 67.760 48.875 67.930 49.065 ;
        RECT 68.685 48.855 68.855 49.045 ;
        RECT 69.155 48.910 69.315 49.020 ;
        RECT 70.525 48.855 70.695 49.045 ;
        RECT 71.905 48.855 72.075 49.045 ;
        RECT 73.745 48.875 73.915 49.065 ;
        RECT 74.200 48.905 74.320 49.015 ;
        RECT 74.940 48.875 75.110 49.065 ;
        RECT 77.425 48.855 77.595 49.045 ;
        RECT 81.100 48.905 81.220 49.015 ;
        RECT 82.025 48.875 82.195 49.065 ;
        RECT 82.485 49.015 82.655 49.045 ;
        RECT 82.480 48.905 82.655 49.015 ;
        RECT 82.485 48.855 82.655 48.905 ;
        RECT 83.865 48.855 84.035 49.065 ;
        RECT 5.525 48.045 6.895 48.855 ;
        RECT 6.905 48.175 8.735 48.855 ;
        RECT 8.745 48.175 10.575 48.855 ;
        RECT 6.905 47.945 8.250 48.175 ;
        RECT 8.745 47.945 10.090 48.175 ;
        RECT 10.585 48.045 16.095 48.855 ;
        RECT 16.710 48.175 18.545 48.855 ;
        RECT 19.100 48.175 23.915 48.855 ;
        RECT 24.070 48.175 25.905 48.855 ;
        RECT 17.615 47.945 18.545 48.175 ;
        RECT 24.975 47.945 25.905 48.175 ;
        RECT 26.225 48.045 28.055 48.855 ;
        RECT 28.445 48.175 30.870 48.855 ;
        RECT 31.295 47.985 31.725 48.770 ;
        RECT 32.205 47.945 35.415 48.855 ;
        RECT 35.885 48.175 43.195 48.855 ;
        RECT 43.245 48.175 50.555 48.855 ;
        RECT 39.400 47.955 40.310 48.175 ;
        RECT 41.845 47.945 43.195 48.175 ;
        RECT 46.760 47.955 47.670 48.175 ;
        RECT 49.205 47.945 50.555 48.175 ;
        RECT 50.605 48.175 54.505 48.855 ;
        RECT 50.605 47.945 51.535 48.175 ;
        RECT 54.745 48.045 56.575 48.855 ;
        RECT 57.055 47.985 57.485 48.770 ;
        RECT 57.505 48.045 63.015 48.855 ;
        RECT 63.025 48.045 68.535 48.855 ;
        RECT 68.545 48.045 70.375 48.855 ;
        RECT 70.395 47.945 71.745 48.855 ;
        RECT 71.765 48.045 77.275 48.855 ;
        RECT 77.285 48.045 80.955 48.855 ;
        RECT 81.425 48.075 82.795 48.855 ;
        RECT 82.805 48.045 84.175 48.855 ;
      LAYER nwell ;
        RECT 5.330 44.825 84.370 47.655 ;
      LAYER pwell ;
        RECT 5.525 43.625 6.895 44.435 ;
        RECT 6.905 44.305 8.250 44.535 ;
        RECT 6.905 43.625 8.735 44.305 ;
        RECT 9.860 43.625 13.335 44.535 ;
        RECT 13.345 44.305 14.690 44.535 ;
        RECT 13.345 43.625 15.175 44.305 ;
        RECT 15.185 43.625 17.935 44.435 ;
        RECT 18.415 43.710 18.845 44.495 ;
        RECT 19.520 43.625 22.995 44.535 ;
        RECT 26.520 44.305 27.430 44.525 ;
        RECT 28.965 44.305 30.315 44.535 ;
        RECT 33.880 44.305 34.790 44.525 ;
        RECT 36.325 44.305 37.675 44.535 ;
        RECT 23.005 43.625 30.315 44.305 ;
        RECT 30.365 43.625 37.675 44.305 ;
        RECT 37.725 44.305 38.655 44.535 ;
        RECT 37.725 43.625 41.625 44.305 ;
        RECT 41.865 43.625 43.695 44.435 ;
        RECT 44.175 43.710 44.605 44.495 ;
        RECT 44.720 44.305 45.640 44.535 ;
        RECT 49.645 44.335 51.055 44.535 ;
        RECT 44.720 43.625 48.185 44.305 ;
        RECT 48.320 43.655 51.055 44.335 ;
        RECT 5.665 43.415 5.835 43.625 ;
        RECT 7.045 43.415 7.215 43.605 ;
        RECT 8.425 43.435 8.595 43.625 ;
        RECT 8.895 43.470 9.055 43.580 ;
        RECT 8.430 43.415 8.595 43.435 ;
        RECT 10.725 43.415 10.895 43.605 ;
        RECT 13.020 43.435 13.190 43.625 ;
        RECT 14.865 43.435 15.035 43.625 ;
        RECT 15.325 43.435 15.495 43.625 ;
        RECT 18.085 43.575 18.255 43.605 ;
        RECT 18.080 43.465 18.255 43.575 ;
        RECT 19.000 43.465 19.120 43.575 ;
        RECT 18.085 43.435 18.255 43.465 ;
        RECT 22.680 43.435 22.850 43.625 ;
        RECT 23.145 43.435 23.315 43.625 ;
        RECT 18.090 43.415 18.255 43.435 ;
        RECT 23.600 43.415 23.770 43.605 ;
        RECT 24.065 43.415 24.235 43.605 ;
        RECT 30.505 43.435 30.675 43.625 ;
        RECT 31.885 43.415 32.055 43.605 ;
        RECT 38.140 43.435 38.310 43.625 ;
        RECT 40.165 43.415 40.335 43.605 ;
        RECT 40.625 43.415 40.795 43.605 ;
        RECT 42.005 43.435 42.175 43.625 ;
        RECT 43.390 43.415 43.560 43.605 ;
        RECT 43.840 43.465 43.960 43.575 ;
        RECT 47.065 43.415 47.235 43.605 ;
        RECT 47.985 43.435 48.155 43.625 ;
        RECT 48.445 43.435 48.615 43.655 ;
        RECT 49.660 43.625 51.055 43.655 ;
        RECT 51.065 43.625 52.895 44.305 ;
        RECT 52.905 43.625 54.275 44.435 ;
        RECT 54.285 43.625 57.495 44.535 ;
        RECT 58.165 44.305 62.095 44.535 ;
        RECT 57.680 43.625 62.095 44.305 ;
        RECT 62.105 43.625 65.315 44.535 ;
        RECT 65.635 44.305 66.565 44.535 ;
        RECT 65.635 43.625 67.470 44.305 ;
        RECT 67.625 43.625 69.455 44.435 ;
        RECT 69.935 43.710 70.365 44.495 ;
        RECT 70.580 43.625 74.055 44.535 ;
        RECT 74.065 43.625 79.575 44.435 ;
        RECT 79.585 43.625 82.335 44.435 ;
        RECT 82.805 43.625 84.175 44.435 ;
        RECT 48.905 43.415 49.075 43.605 ;
        RECT 51.205 43.435 51.375 43.625 ;
        RECT 51.675 43.460 51.835 43.570 ;
        RECT 53.045 43.435 53.215 43.625 ;
        RECT 54.420 43.415 54.590 43.605 ;
        RECT 54.885 43.415 55.055 43.605 ;
        RECT 56.720 43.465 56.840 43.575 ;
        RECT 57.185 43.435 57.355 43.625 ;
        RECT 57.680 43.605 57.790 43.625 ;
        RECT 57.620 43.435 57.815 43.605 ;
        RECT 60.865 43.435 61.035 43.605 ;
        RECT 57.645 43.415 57.815 43.435 ;
        RECT 61.325 43.415 61.495 43.605 ;
        RECT 62.245 43.435 62.415 43.625 ;
        RECT 67.305 43.605 67.470 43.625 ;
        RECT 66.385 43.415 66.555 43.605 ;
        RECT 67.305 43.435 67.475 43.605 ;
        RECT 67.765 43.435 67.935 43.625 ;
        RECT 73.740 43.605 73.910 43.625 ;
        RECT 69.600 43.465 69.720 43.575 ;
        RECT 73.740 43.435 73.915 43.605 ;
        RECT 74.205 43.435 74.375 43.625 ;
        RECT 73.745 43.415 73.915 43.435 ;
        RECT 79.265 43.415 79.435 43.605 ;
        RECT 79.725 43.435 79.895 43.625 ;
        RECT 81.105 43.415 81.275 43.605 ;
        RECT 82.480 43.465 82.600 43.575 ;
        RECT 83.865 43.415 84.035 43.625 ;
        RECT 5.525 42.605 6.895 43.415 ;
        RECT 6.905 42.605 8.275 43.415 ;
        RECT 8.430 42.735 10.265 43.415 ;
        RECT 10.585 42.735 17.895 43.415 ;
        RECT 18.090 42.735 19.925 43.415 ;
        RECT 9.335 42.505 10.265 42.735 ;
        RECT 14.100 42.515 15.010 42.735 ;
        RECT 16.545 42.505 17.895 42.735 ;
        RECT 18.995 42.505 19.925 42.735 ;
        RECT 20.440 42.505 23.915 43.415 ;
        RECT 23.925 42.735 31.235 43.415 ;
        RECT 27.440 42.515 28.350 42.735 ;
        RECT 29.885 42.505 31.235 42.735 ;
        RECT 31.295 42.545 31.725 43.330 ;
        RECT 31.745 42.735 36.560 43.415 ;
        RECT 36.900 42.735 40.365 43.415 ;
        RECT 40.485 42.735 43.225 43.415 ;
        RECT 36.900 42.505 37.820 42.735 ;
        RECT 43.250 42.505 46.835 43.415 ;
        RECT 46.925 42.605 48.755 43.415 ;
        RECT 48.765 42.605 50.855 43.415 ;
        RECT 52.545 42.505 54.735 43.415 ;
        RECT 54.745 42.605 56.575 43.415 ;
        RECT 57.055 42.545 57.485 43.330 ;
        RECT 57.505 42.605 59.335 43.415 ;
        RECT 59.345 42.735 60.710 43.415 ;
        RECT 61.185 42.735 66.000 43.415 ;
        RECT 66.245 42.735 73.555 43.415 ;
        RECT 69.760 42.515 70.670 42.735 ;
        RECT 72.205 42.505 73.555 42.735 ;
        RECT 73.605 42.605 79.115 43.415 ;
        RECT 79.125 42.605 80.955 43.415 ;
        RECT 80.965 42.735 82.795 43.415 ;
        RECT 81.450 42.505 82.795 42.735 ;
        RECT 82.805 42.605 84.175 43.415 ;
      LAYER nwell ;
        RECT 5.330 39.385 84.370 42.215 ;
      LAYER pwell ;
        RECT 5.525 38.185 6.895 38.995 ;
        RECT 10.420 38.865 11.330 39.085 ;
        RECT 12.865 38.865 14.215 39.095 ;
        RECT 6.905 38.185 14.215 38.865 ;
        RECT 14.265 38.865 15.610 39.095 ;
        RECT 14.265 38.185 16.095 38.865 ;
        RECT 16.105 38.185 17.935 38.995 ;
        RECT 18.415 38.270 18.845 39.055 ;
        RECT 18.865 38.185 22.075 39.095 ;
        RECT 22.100 38.865 23.470 39.095 ;
        RECT 22.100 38.185 24.375 38.865 ;
        RECT 24.395 38.185 25.745 39.095 ;
        RECT 25.765 38.185 31.275 38.995 ;
        RECT 31.745 38.865 32.675 39.095 ;
        RECT 40.320 38.865 41.230 39.085 ;
        RECT 42.765 38.865 44.115 39.095 ;
        RECT 31.745 38.185 35.645 38.865 ;
        RECT 36.805 38.185 44.115 38.865 ;
        RECT 44.175 38.270 44.605 39.055 ;
        RECT 44.635 38.185 45.985 39.095 ;
        RECT 49.520 38.865 50.430 39.085 ;
        RECT 51.965 38.865 53.315 39.095 ;
        RECT 57.800 38.865 58.710 39.085 ;
        RECT 60.245 38.865 61.595 39.095 ;
        RECT 46.005 38.185 53.315 38.865 ;
        RECT 54.285 38.185 61.595 38.865 ;
        RECT 62.760 38.185 66.235 39.095 ;
        RECT 67.295 38.865 68.225 39.095 ;
        RECT 66.390 38.185 68.225 38.865 ;
        RECT 68.545 38.185 69.915 38.995 ;
        RECT 69.935 38.270 70.365 39.055 ;
        RECT 73.900 38.865 74.810 39.085 ;
        RECT 76.345 38.865 77.695 39.095 ;
        RECT 70.385 38.185 77.695 38.865 ;
        RECT 77.745 38.185 81.415 38.995 ;
        RECT 81.425 38.185 82.795 38.995 ;
        RECT 82.805 38.185 84.175 38.995 ;
        RECT 5.665 37.975 5.835 38.185 ;
        RECT 7.045 37.995 7.215 38.185 ;
        RECT 7.970 37.975 8.140 38.165 ;
        RECT 13.485 37.995 13.655 38.165 ;
        RECT 13.485 37.975 13.650 37.995 ;
        RECT 13.945 37.975 14.115 38.165 ;
        RECT 15.785 37.995 15.955 38.185 ;
        RECT 16.245 37.995 16.415 38.185 ;
        RECT 17.165 37.975 17.335 38.165 ;
        RECT 18.080 38.025 18.200 38.135 ;
        RECT 20.840 38.025 20.960 38.135 ;
        RECT 21.310 37.975 21.480 38.165 ;
        RECT 21.775 37.995 21.945 38.185 ;
        RECT 22.685 37.975 22.855 38.165 ;
        RECT 24.060 37.995 24.230 38.185 ;
        RECT 24.525 37.995 24.695 38.185 ;
        RECT 25.905 37.995 26.075 38.185 ;
        RECT 25.905 37.975 26.055 37.995 ;
        RECT 26.365 37.975 26.535 38.165 ;
        RECT 30.045 37.975 30.215 38.165 ;
        RECT 31.420 38.025 31.540 38.135 ;
        RECT 31.885 37.975 32.055 38.165 ;
        RECT 32.160 37.995 32.330 38.185 ;
        RECT 33.715 37.975 33.885 38.165 ;
        RECT 36.035 38.030 36.195 38.140 ;
        RECT 36.945 37.975 37.115 38.185 ;
        RECT 39.700 38.025 39.820 38.135 ;
        RECT 40.440 37.975 40.610 38.165 ;
        RECT 44.765 37.995 44.935 38.185 ;
        RECT 46.145 37.995 46.315 38.185 ;
        RECT 5.525 37.165 6.895 37.975 ;
        RECT 7.825 37.065 11.300 37.975 ;
        RECT 11.815 37.295 13.650 37.975 ;
        RECT 11.815 37.065 12.745 37.295 ;
        RECT 13.805 37.065 17.015 37.975 ;
        RECT 17.025 37.165 20.695 37.975 ;
        RECT 21.165 37.065 22.515 37.975 ;
        RECT 22.545 37.165 23.915 37.975 ;
        RECT 24.125 37.155 26.055 37.975 ;
        RECT 26.225 37.165 29.895 37.975 ;
        RECT 29.905 37.165 31.275 37.975 ;
        RECT 24.125 37.065 25.075 37.155 ;
        RECT 31.295 37.105 31.725 37.890 ;
        RECT 31.745 37.165 33.575 37.975 ;
        RECT 33.585 37.065 36.795 37.975 ;
        RECT 36.805 37.165 39.555 37.975 ;
        RECT 40.025 37.295 43.925 37.975 ;
        RECT 44.165 37.945 45.560 37.975 ;
        RECT 46.605 37.945 46.775 38.165 ;
        RECT 47.060 38.025 47.180 38.135 ;
        RECT 48.445 37.975 48.615 38.165 ;
        RECT 53.505 37.975 53.675 38.165 ;
        RECT 53.965 37.995 54.135 38.165 ;
        RECT 54.425 37.995 54.595 38.185 ;
        RECT 56.720 38.025 56.840 38.135 ;
        RECT 53.995 37.975 54.135 37.995 ;
        RECT 57.650 37.975 57.820 38.165 ;
        RECT 61.320 38.025 61.440 38.135 ;
        RECT 61.785 37.995 61.955 38.165 ;
        RECT 61.790 37.975 61.955 37.995 ;
        RECT 64.090 37.975 64.260 38.165 ;
        RECT 65.920 37.995 66.090 38.185 ;
        RECT 66.390 38.165 66.555 38.185 ;
        RECT 66.385 37.995 66.555 38.165 ;
        RECT 66.405 37.975 66.555 37.995 ;
        RECT 68.685 37.975 68.855 38.185 ;
        RECT 70.525 37.995 70.695 38.185 ;
        RECT 75.580 37.975 75.750 38.165 ;
        RECT 76.955 37.975 77.125 38.165 ;
        RECT 77.425 37.975 77.595 38.165 ;
        RECT 77.885 37.995 78.055 38.185 ;
        RECT 81.565 37.995 81.735 38.185 ;
        RECT 83.865 37.975 84.035 38.185 ;
        RECT 40.025 37.065 40.955 37.295 ;
        RECT 44.165 37.265 46.900 37.945 ;
        RECT 44.165 37.065 45.575 37.265 ;
        RECT 47.395 37.065 48.745 37.975 ;
        RECT 49.000 37.295 53.815 37.975 ;
        RECT 53.995 37.155 56.565 37.975 ;
        RECT 54.975 37.065 56.565 37.155 ;
        RECT 57.055 37.105 57.485 37.890 ;
        RECT 57.505 37.065 60.980 37.975 ;
        RECT 61.790 37.295 63.625 37.975 ;
        RECT 62.695 37.065 63.625 37.295 ;
        RECT 63.945 37.065 66.135 37.975 ;
        RECT 66.405 37.155 68.335 37.975 ;
        RECT 68.545 37.165 72.215 37.975 ;
        RECT 67.385 37.065 68.335 37.155 ;
        RECT 72.420 37.065 75.895 37.975 ;
        RECT 75.905 37.195 77.275 37.975 ;
        RECT 77.285 37.165 82.795 37.975 ;
        RECT 82.805 37.165 84.175 37.975 ;
      LAYER nwell ;
        RECT 5.330 33.945 84.370 36.775 ;
      LAYER pwell ;
        RECT 5.525 32.745 6.895 33.555 ;
        RECT 6.905 32.745 9.655 33.555 ;
        RECT 13.640 33.425 14.550 33.645 ;
        RECT 16.085 33.425 17.435 33.655 ;
        RECT 10.125 32.745 17.435 33.425 ;
        RECT 18.415 32.830 18.845 33.615 ;
        RECT 19.175 33.425 20.105 33.655 ;
        RECT 19.175 32.745 21.010 33.425 ;
        RECT 22.280 32.745 25.755 33.655 ;
        RECT 25.865 32.745 28.055 33.655 ;
        RECT 28.065 32.745 29.895 33.555 ;
        RECT 29.945 33.425 31.295 33.655 ;
        RECT 32.830 33.425 33.740 33.645 ;
        RECT 29.945 32.745 37.255 33.425 ;
        RECT 37.265 32.745 40.740 33.655 ;
        RECT 40.945 32.745 43.695 33.555 ;
        RECT 44.175 32.830 44.605 33.615 ;
        RECT 44.625 32.745 47.375 33.555 ;
        RECT 47.385 33.425 48.315 33.655 ;
        RECT 51.620 33.425 52.540 33.655 ;
        RECT 47.385 32.745 51.285 33.425 ;
        RECT 51.620 32.745 55.085 33.425 ;
        RECT 55.205 32.745 57.035 33.425 ;
        RECT 57.045 32.745 62.555 33.555 ;
        RECT 62.565 32.745 66.235 33.555 ;
        RECT 66.245 32.745 67.615 33.555 ;
        RECT 68.675 33.425 69.605 33.655 ;
        RECT 67.770 32.745 69.605 33.425 ;
        RECT 69.935 32.830 70.365 33.615 ;
        RECT 71.500 32.745 74.975 33.655 ;
        RECT 78.500 33.425 79.410 33.645 ;
        RECT 80.945 33.425 82.295 33.655 ;
        RECT 74.985 32.745 82.295 33.425 ;
        RECT 82.805 32.745 84.175 33.555 ;
        RECT 5.665 32.535 5.835 32.745 ;
        RECT 7.045 32.535 7.215 32.745 ;
        RECT 9.800 32.585 9.920 32.695 ;
        RECT 10.265 32.555 10.435 32.745 ;
        RECT 20.845 32.725 21.010 32.745 ;
        RECT 12.575 32.580 12.735 32.690 ;
        RECT 13.490 32.535 13.660 32.725 ;
        RECT 17.165 32.535 17.335 32.725 ;
        RECT 17.635 32.590 17.795 32.700 ;
        RECT 19.005 32.535 19.175 32.725 ;
        RECT 20.845 32.555 21.015 32.725 ;
        RECT 21.315 32.590 21.475 32.700 ;
        RECT 20.850 32.535 21.015 32.555 ;
        RECT 23.145 32.535 23.315 32.725 ;
        RECT 25.440 32.555 25.610 32.745 ;
        RECT 27.740 32.555 27.910 32.745 ;
        RECT 28.205 32.555 28.375 32.745 ;
        RECT 30.515 32.580 30.675 32.690 ;
        RECT 31.885 32.535 32.055 32.725 ;
        RECT 35.105 32.555 35.275 32.725 ;
        RECT 36.945 32.555 37.115 32.745 ;
        RECT 37.410 32.725 37.580 32.745 ;
        RECT 37.405 32.555 37.580 32.725 ;
        RECT 41.085 32.555 41.255 32.745 ;
        RECT 44.765 32.725 44.935 32.745 ;
        RECT 35.110 32.535 35.275 32.555 ;
        RECT 37.405 32.535 37.575 32.555 ;
        RECT 42.925 32.535 43.095 32.725 ;
        RECT 43.840 32.585 43.960 32.695 ;
        RECT 44.765 32.555 44.940 32.725 ;
        RECT 47.800 32.555 47.970 32.745 ;
        RECT 44.770 32.535 44.940 32.555 ;
        RECT 48.445 32.535 48.615 32.725 ;
        RECT 49.825 32.535 49.995 32.725 ;
        RECT 54.885 32.555 55.055 32.745 ;
        RECT 55.345 32.555 55.515 32.745 ;
        RECT 57.185 32.555 57.355 32.745 ;
        RECT 57.645 32.535 57.815 32.725 ;
        RECT 61.320 32.585 61.440 32.695 ;
        RECT 62.705 32.555 62.875 32.745 ;
        RECT 64.085 32.555 64.255 32.725 ;
        RECT 64.085 32.535 64.225 32.555 ;
        RECT 64.550 32.535 64.720 32.725 ;
        RECT 66.385 32.555 66.555 32.745 ;
        RECT 67.770 32.725 67.935 32.745 ;
        RECT 66.845 32.535 67.015 32.725 ;
        RECT 67.765 32.555 67.935 32.725 ;
        RECT 68.680 32.585 68.800 32.695 ;
        RECT 69.145 32.555 69.315 32.725 ;
        RECT 70.535 32.590 70.695 32.700 ;
        RECT 69.150 32.535 69.315 32.555 ;
        RECT 74.205 32.535 74.375 32.725 ;
        RECT 74.660 32.690 74.830 32.745 ;
        RECT 74.660 32.580 74.835 32.690 ;
        RECT 74.660 32.555 74.830 32.580 ;
        RECT 75.125 32.555 75.295 32.745 ;
        RECT 75.585 32.535 75.755 32.725 ;
        RECT 82.480 32.585 82.600 32.695 ;
        RECT 83.865 32.535 84.035 32.745 ;
        RECT 5.525 31.725 6.895 32.535 ;
        RECT 6.905 31.725 12.415 32.535 ;
        RECT 13.345 31.625 16.820 32.535 ;
        RECT 17.025 31.855 18.855 32.535 ;
        RECT 17.510 31.625 18.855 31.855 ;
        RECT 18.865 31.725 20.695 32.535 ;
        RECT 20.850 31.855 22.685 32.535 ;
        RECT 23.005 31.855 30.315 32.535 ;
        RECT 21.755 31.625 22.685 31.855 ;
        RECT 26.520 31.635 27.430 31.855 ;
        RECT 28.965 31.625 30.315 31.855 ;
        RECT 31.295 31.665 31.725 32.450 ;
        RECT 31.745 31.625 34.955 32.535 ;
        RECT 35.110 31.855 36.945 32.535 ;
        RECT 36.015 31.625 36.945 31.855 ;
        RECT 37.265 31.725 42.775 32.535 ;
        RECT 42.785 31.725 44.615 32.535 ;
        RECT 44.630 31.625 48.215 32.535 ;
        RECT 48.305 31.725 49.675 32.535 ;
        RECT 49.685 31.855 56.995 32.535 ;
        RECT 53.200 31.635 54.110 31.855 ;
        RECT 55.645 31.625 56.995 31.855 ;
        RECT 57.055 31.665 57.485 32.450 ;
        RECT 57.505 31.725 61.175 32.535 ;
        RECT 61.655 31.715 64.225 32.535 ;
        RECT 61.655 31.625 63.245 31.715 ;
        RECT 64.405 31.625 66.595 32.535 ;
        RECT 66.705 31.725 68.535 32.535 ;
        RECT 69.150 31.855 70.985 32.535 ;
        RECT 70.055 31.625 70.985 31.855 ;
        RECT 71.305 31.625 74.515 32.535 ;
        RECT 75.445 31.855 82.755 32.535 ;
        RECT 78.960 31.635 79.870 31.855 ;
        RECT 81.405 31.625 82.755 31.855 ;
        RECT 82.805 31.725 84.175 32.535 ;
      LAYER nwell ;
        RECT 5.330 28.505 84.370 31.335 ;
      LAYER pwell ;
        RECT 5.525 27.305 6.895 28.115 ;
        RECT 6.905 27.985 8.250 28.215 ;
        RECT 9.515 27.985 10.445 28.215 ;
        RECT 6.905 27.305 8.735 27.985 ;
        RECT 9.515 27.305 11.350 27.985 ;
        RECT 11.505 27.305 13.335 28.115 ;
        RECT 13.805 27.305 17.280 28.215 ;
        RECT 18.415 27.390 18.845 28.175 ;
        RECT 18.865 27.305 24.375 28.115 ;
        RECT 24.385 27.305 29.895 28.115 ;
        RECT 29.905 27.305 35.415 28.115 ;
        RECT 37.395 27.985 38.325 28.215 ;
        RECT 36.490 27.305 38.325 27.985 ;
        RECT 38.645 27.305 40.475 28.115 ;
        RECT 40.945 27.305 44.155 28.215 ;
        RECT 44.175 27.390 44.605 28.175 ;
        RECT 44.625 27.305 45.995 28.115 ;
        RECT 46.200 27.305 49.675 28.215 ;
        RECT 49.995 27.985 50.925 28.215 ;
        RECT 55.500 27.985 56.410 28.205 ;
        RECT 57.945 27.985 59.295 28.215 ;
        RECT 49.995 27.305 51.830 27.985 ;
        RECT 51.985 27.305 59.295 27.985 ;
        RECT 59.655 27.985 60.585 28.215 ;
        RECT 65.160 27.985 66.070 28.205 ;
        RECT 67.605 27.985 68.955 28.215 ;
        RECT 59.655 27.305 61.490 27.985 ;
        RECT 61.645 27.305 68.955 27.985 ;
        RECT 69.935 27.390 70.365 28.175 ;
        RECT 71.895 27.985 72.825 28.215 ;
        RECT 70.990 27.305 72.825 27.985 ;
        RECT 73.145 27.305 78.655 28.115 ;
        RECT 78.665 27.305 80.495 28.115 ;
        RECT 81.450 27.985 82.795 28.215 ;
        RECT 80.965 27.305 82.795 27.985 ;
        RECT 82.805 27.305 84.175 28.115 ;
        RECT 5.665 27.095 5.835 27.305 ;
        RECT 7.040 27.145 7.160 27.255 ;
        RECT 7.510 27.095 7.680 27.285 ;
        RECT 8.425 27.115 8.595 27.305 ;
        RECT 11.185 27.285 11.350 27.305 ;
        RECT 8.880 27.145 9.000 27.255 ;
        RECT 11.185 27.095 11.355 27.285 ;
        RECT 11.645 27.115 11.815 27.305 ;
        RECT 13.480 27.145 13.600 27.255 ;
        RECT 13.950 27.115 14.120 27.305 ;
        RECT 17.635 27.150 17.795 27.260 ;
        RECT 19.005 27.115 19.175 27.305 ;
        RECT 20.385 27.115 20.555 27.285 ;
        RECT 20.840 27.145 20.960 27.255 ;
        RECT 20.385 27.095 20.550 27.115 ;
        RECT 21.310 27.095 21.480 27.285 ;
        RECT 24.525 27.115 24.695 27.305 ;
        RECT 24.980 27.145 25.100 27.255 ;
        RECT 28.660 27.095 28.830 27.285 ;
        RECT 29.125 27.115 29.295 27.285 ;
        RECT 30.045 27.115 30.215 27.305 ;
        RECT 36.490 27.285 36.655 27.305 ;
        RECT 29.130 27.095 29.295 27.115 ;
        RECT 31.885 27.095 32.055 27.285 ;
        RECT 34.645 27.095 34.815 27.285 ;
        RECT 35.575 27.150 35.735 27.260 ;
        RECT 36.485 27.115 36.655 27.285 ;
        RECT 38.785 27.115 38.955 27.305 ;
        RECT 40.620 27.145 40.740 27.255 ;
        RECT 41.085 27.115 41.255 27.305 ;
        RECT 42.005 27.095 42.175 27.285 ;
        RECT 43.385 27.095 43.555 27.285 ;
        RECT 44.765 27.115 44.935 27.305 ;
        RECT 49.360 27.115 49.530 27.305 ;
        RECT 51.665 27.285 51.830 27.305 ;
        RECT 50.740 27.145 50.860 27.255 ;
        RECT 51.210 27.095 51.380 27.285 ;
        RECT 51.665 27.115 51.835 27.285 ;
        RECT 52.125 27.115 52.295 27.305 ;
        RECT 61.325 27.285 61.490 27.305 ;
        RECT 56.725 27.115 56.895 27.285 ;
        RECT 57.655 27.140 57.815 27.250 ;
        RECT 56.725 27.095 56.890 27.115 ;
        RECT 61.325 27.095 61.495 27.285 ;
        RECT 61.785 27.115 61.955 27.305 ;
        RECT 70.990 27.285 71.155 27.305 ;
        RECT 65.000 27.095 65.170 27.285 ;
        RECT 65.465 27.095 65.635 27.285 ;
        RECT 67.300 27.145 67.420 27.255 ;
        RECT 67.765 27.095 67.935 27.285 ;
        RECT 69.155 27.150 69.315 27.260 ;
        RECT 70.520 27.145 70.640 27.255 ;
        RECT 70.985 27.115 71.155 27.285 ;
        RECT 73.285 27.115 73.455 27.305 ;
        RECT 77.885 27.095 78.055 27.285 ;
        RECT 78.345 27.095 78.515 27.285 ;
        RECT 78.805 27.115 78.975 27.305 ;
        RECT 80.640 27.145 80.760 27.255 ;
        RECT 81.105 27.115 81.275 27.305 ;
        RECT 82.035 27.140 82.195 27.250 ;
        RECT 83.865 27.095 84.035 27.305 ;
        RECT 5.525 26.285 6.895 27.095 ;
        RECT 7.365 26.185 10.840 27.095 ;
        RECT 11.045 26.415 18.355 27.095 ;
        RECT 14.560 26.195 15.470 26.415 ;
        RECT 17.005 26.185 18.355 26.415 ;
        RECT 18.715 26.415 20.550 27.095 ;
        RECT 18.715 26.185 19.645 26.415 ;
        RECT 21.165 26.185 24.640 27.095 ;
        RECT 25.500 26.185 28.975 27.095 ;
        RECT 29.130 26.415 30.965 27.095 ;
        RECT 30.035 26.185 30.965 26.415 ;
        RECT 31.295 26.225 31.725 27.010 ;
        RECT 31.745 26.285 34.495 27.095 ;
        RECT 34.505 26.415 41.815 27.095 ;
        RECT 38.020 26.195 38.930 26.415 ;
        RECT 40.465 26.185 41.815 26.415 ;
        RECT 41.865 26.285 43.235 27.095 ;
        RECT 43.245 26.415 50.555 27.095 ;
        RECT 46.760 26.195 47.670 26.415 ;
        RECT 49.205 26.185 50.555 26.415 ;
        RECT 51.065 26.185 54.540 27.095 ;
        RECT 55.055 26.415 56.890 27.095 ;
        RECT 55.055 26.185 55.985 26.415 ;
        RECT 57.055 26.225 57.485 27.010 ;
        RECT 58.425 26.185 61.635 27.095 ;
        RECT 61.840 26.185 65.315 27.095 ;
        RECT 65.325 26.285 67.155 27.095 ;
        RECT 67.625 26.415 74.935 27.095 ;
        RECT 71.140 26.195 72.050 26.415 ;
        RECT 73.585 26.185 74.935 26.415 ;
        RECT 74.985 26.185 78.195 27.095 ;
        RECT 78.205 26.285 81.875 27.095 ;
        RECT 82.805 26.285 84.175 27.095 ;
      LAYER nwell ;
        RECT 5.330 23.065 84.370 25.895 ;
      LAYER pwell ;
        RECT 5.525 21.865 6.895 22.675 ;
        RECT 10.420 22.545 11.330 22.765 ;
        RECT 12.865 22.545 14.215 22.775 ;
        RECT 6.905 21.865 14.215 22.545 ;
        RECT 14.265 21.865 17.475 22.775 ;
        RECT 18.415 21.950 18.845 22.735 ;
        RECT 18.865 21.865 20.235 22.675 ;
        RECT 23.760 22.545 24.670 22.765 ;
        RECT 26.205 22.545 27.555 22.775 ;
        RECT 31.120 22.545 32.030 22.765 ;
        RECT 33.565 22.545 34.915 22.775 ;
        RECT 20.245 21.865 27.555 22.545 ;
        RECT 27.605 21.865 34.915 22.545 ;
        RECT 35.885 21.865 39.360 22.775 ;
        RECT 39.565 21.865 41.395 22.675 ;
        RECT 42.915 22.545 43.845 22.775 ;
        RECT 42.010 21.865 43.845 22.545 ;
        RECT 44.175 21.950 44.605 22.735 ;
        RECT 44.625 21.865 48.100 22.775 ;
        RECT 48.305 21.865 50.135 22.675 ;
        RECT 50.145 22.545 51.490 22.775 ;
        RECT 50.145 21.865 51.975 22.545 ;
        RECT 51.985 21.865 57.495 22.675 ;
        RECT 57.505 21.865 63.015 22.675 ;
        RECT 63.025 21.865 66.695 22.675 ;
        RECT 68.675 22.545 69.605 22.775 ;
        RECT 67.770 21.865 69.605 22.545 ;
        RECT 69.935 21.950 70.365 22.735 ;
        RECT 70.385 21.865 73.860 22.775 ;
        RECT 74.065 21.865 75.435 22.675 ;
        RECT 78.960 22.545 79.870 22.765 ;
        RECT 81.405 22.545 82.755 22.775 ;
        RECT 75.445 21.865 82.755 22.545 ;
        RECT 82.805 21.865 84.175 22.675 ;
        RECT 5.665 21.655 5.835 21.865 ;
        RECT 7.045 21.675 7.215 21.865 ;
        RECT 8.425 21.655 8.595 21.845 ;
        RECT 8.885 21.655 9.055 21.845 ;
        RECT 11.645 21.655 11.815 21.845 ;
        RECT 13.485 21.655 13.655 21.845 ;
        RECT 13.955 21.700 14.115 21.810 ;
        RECT 14.405 21.675 14.575 21.865 ;
        RECT 14.865 21.655 15.035 21.845 ;
        RECT 17.635 21.710 17.795 21.820 ;
        RECT 18.085 21.655 18.255 21.845 ;
        RECT 19.005 21.675 19.175 21.865 ;
        RECT 19.935 21.700 20.095 21.810 ;
        RECT 20.385 21.675 20.555 21.865 ;
        RECT 20.845 21.675 21.015 21.845 ;
        RECT 20.850 21.655 21.015 21.675 ;
        RECT 23.145 21.655 23.315 21.845 ;
        RECT 27.745 21.675 27.915 21.865 ;
        RECT 28.665 21.655 28.835 21.845 ;
        RECT 31.885 21.655 32.055 21.845 ;
        RECT 33.725 21.655 33.895 21.845 ;
        RECT 35.115 21.710 35.275 21.820 ;
        RECT 36.030 21.675 36.200 21.865 ;
        RECT 36.945 21.655 37.115 21.845 ;
        RECT 38.325 21.655 38.495 21.845 ;
        RECT 39.705 21.675 39.875 21.865 ;
        RECT 42.010 21.845 42.175 21.865 ;
        RECT 41.545 21.815 41.715 21.845 ;
        RECT 41.540 21.705 41.715 21.815 ;
        RECT 41.545 21.655 41.715 21.705 ;
        RECT 42.005 21.675 42.175 21.845 ;
        RECT 44.770 21.675 44.940 21.865 ;
        RECT 47.065 21.655 47.235 21.845 ;
        RECT 48.445 21.675 48.615 21.865 ;
        RECT 50.740 21.705 50.860 21.815 ;
        RECT 51.210 21.655 51.380 21.845 ;
        RECT 51.665 21.675 51.835 21.865 ;
        RECT 52.125 21.675 52.295 21.865 ;
        RECT 56.725 21.675 56.895 21.845 ;
        RECT 57.645 21.675 57.815 21.865 ;
        RECT 56.725 21.655 56.890 21.675 ;
        RECT 60.405 21.655 60.575 21.845 ;
        RECT 60.870 21.655 61.040 21.845 ;
        RECT 63.165 21.675 63.335 21.865 ;
        RECT 67.770 21.845 67.935 21.865 ;
        RECT 66.385 21.675 66.555 21.845 ;
        RECT 66.385 21.655 66.550 21.675 ;
        RECT 66.845 21.655 67.015 21.845 ;
        RECT 67.765 21.675 67.935 21.845 ;
        RECT 68.680 21.705 68.800 21.815 ;
        RECT 70.530 21.675 70.700 21.865 ;
        RECT 71.905 21.655 72.075 21.845 ;
        RECT 74.205 21.675 74.375 21.865 ;
        RECT 75.585 21.845 75.755 21.865 ;
        RECT 75.580 21.675 75.755 21.845 ;
        RECT 75.580 21.655 75.750 21.675 ;
        RECT 76.045 21.655 76.215 21.845 ;
        RECT 77.425 21.655 77.595 21.845 ;
        RECT 79.265 21.655 79.435 21.845 ;
        RECT 82.485 21.655 82.655 21.845 ;
        RECT 83.865 21.655 84.035 21.865 ;
        RECT 5.525 20.845 6.895 21.655 ;
        RECT 6.905 20.975 8.735 21.655 ;
        RECT 6.905 20.745 8.250 20.975 ;
        RECT 8.745 20.845 10.115 21.655 ;
        RECT 10.125 20.975 11.955 21.655 ;
        RECT 11.965 20.975 13.795 21.655 ;
        RECT 10.125 20.745 11.470 20.975 ;
        RECT 11.965 20.745 13.310 20.975 ;
        RECT 14.725 20.745 17.935 21.655 ;
        RECT 17.945 20.975 19.775 21.655 ;
        RECT 20.850 20.975 22.685 21.655 ;
        RECT 18.430 20.745 19.775 20.975 ;
        RECT 21.755 20.745 22.685 20.975 ;
        RECT 23.005 20.845 28.515 21.655 ;
        RECT 28.525 20.845 31.275 21.655 ;
        RECT 31.295 20.785 31.725 21.570 ;
        RECT 31.745 20.845 33.575 21.655 ;
        RECT 33.585 20.745 36.795 21.655 ;
        RECT 36.805 20.845 38.175 21.655 ;
        RECT 38.185 20.745 41.395 21.655 ;
        RECT 41.405 20.845 46.915 21.655 ;
        RECT 46.925 20.845 50.595 21.655 ;
        RECT 51.065 20.745 54.540 21.655 ;
        RECT 55.055 20.975 56.890 21.655 ;
        RECT 55.055 20.745 55.985 20.975 ;
        RECT 57.055 20.785 57.485 21.570 ;
        RECT 57.505 20.745 60.715 21.655 ;
        RECT 60.725 20.745 64.200 21.655 ;
        RECT 64.715 20.975 66.550 21.655 ;
        RECT 64.715 20.745 65.645 20.975 ;
        RECT 66.705 20.845 68.535 21.655 ;
        RECT 69.005 20.745 72.215 21.655 ;
        RECT 72.420 20.745 75.895 21.655 ;
        RECT 75.905 20.845 77.275 21.655 ;
        RECT 77.285 20.975 79.115 21.655 ;
        RECT 79.125 20.975 80.955 21.655 ;
        RECT 77.770 20.745 79.115 20.975 ;
        RECT 79.610 20.745 80.955 20.975 ;
        RECT 80.965 20.975 82.795 21.655 ;
        RECT 80.965 20.745 82.310 20.975 ;
        RECT 82.805 20.845 84.175 21.655 ;
      LAYER nwell ;
        RECT 5.330 17.625 84.370 20.455 ;
      LAYER pwell ;
        RECT 5.525 16.425 6.895 17.235 ;
        RECT 7.365 16.425 10.840 17.335 ;
        RECT 11.965 17.105 13.310 17.335 ;
        RECT 11.965 16.425 13.795 17.105 ;
        RECT 13.805 16.425 17.280 17.335 ;
        RECT 18.415 16.510 18.845 17.295 ;
        RECT 19.520 16.425 22.995 17.335 ;
        RECT 23.200 16.425 26.675 17.335 ;
        RECT 30.200 17.105 31.110 17.325 ;
        RECT 32.645 17.105 33.995 17.335 ;
        RECT 26.685 16.425 33.995 17.105 ;
        RECT 34.965 16.425 38.440 17.335 ;
        RECT 38.645 16.425 40.475 17.235 ;
        RECT 40.485 16.425 43.960 17.335 ;
        RECT 44.175 16.510 44.605 17.295 ;
        RECT 44.625 16.425 46.455 17.235 ;
        RECT 46.925 16.425 50.400 17.335 ;
        RECT 54.120 17.105 55.030 17.325 ;
        RECT 56.565 17.105 57.915 17.335 ;
        RECT 61.480 17.105 62.390 17.325 ;
        RECT 63.925 17.105 65.275 17.335 ;
        RECT 50.605 16.425 57.915 17.105 ;
        RECT 57.965 16.425 65.275 17.105 ;
        RECT 65.325 16.425 68.800 17.335 ;
        RECT 69.935 16.510 70.365 17.295 ;
        RECT 71.040 16.425 74.515 17.335 ;
        RECT 74.720 16.425 78.195 17.335 ;
        RECT 78.690 17.105 80.035 17.335 ;
        RECT 80.530 17.105 81.875 17.335 ;
        RECT 78.205 16.425 80.035 17.105 ;
        RECT 80.045 16.425 81.875 17.105 ;
        RECT 82.805 16.425 84.175 17.235 ;
        RECT 5.665 16.215 5.835 16.425 ;
        RECT 7.040 16.370 7.160 16.375 ;
        RECT 7.040 16.265 7.215 16.370 ;
        RECT 7.055 16.260 7.215 16.265 ;
        RECT 7.510 16.235 7.680 16.425 ;
        RECT 7.965 16.235 8.135 16.405 ;
        RECT 7.970 16.215 8.135 16.235 ;
        RECT 10.265 16.215 10.435 16.405 ;
        RECT 11.195 16.270 11.355 16.380 ;
        RECT 11.645 16.215 11.815 16.405 ;
        RECT 13.485 16.235 13.655 16.425 ;
        RECT 13.950 16.235 14.120 16.425 ;
        RECT 17.635 16.270 17.795 16.380 ;
        RECT 19.005 16.375 19.175 16.405 ;
        RECT 19.000 16.265 19.175 16.375 ;
        RECT 19.005 16.235 19.175 16.265 ;
        RECT 19.010 16.215 19.175 16.235 ;
        RECT 21.305 16.215 21.475 16.405 ;
        RECT 22.680 16.235 22.850 16.425 ;
        RECT 26.360 16.235 26.530 16.425 ;
        RECT 26.825 16.235 26.995 16.425 ;
        RECT 30.505 16.235 30.675 16.405 ;
        RECT 30.960 16.265 31.080 16.375 ;
        RECT 31.880 16.265 32.000 16.375 ;
        RECT 34.195 16.270 34.355 16.380 ;
        RECT 35.110 16.235 35.280 16.425 ;
        RECT 38.785 16.235 38.955 16.425 ;
        RECT 30.505 16.215 30.670 16.235 ;
        RECT 39.245 16.215 39.415 16.405 ;
        RECT 39.700 16.265 39.820 16.375 ;
        RECT 40.165 16.215 40.335 16.405 ;
        RECT 40.630 16.235 40.800 16.425 ;
        RECT 44.765 16.235 44.935 16.425 ;
        RECT 46.600 16.265 46.720 16.375 ;
        RECT 47.070 16.235 47.240 16.425 ;
        RECT 47.525 16.215 47.695 16.405 ;
        RECT 50.745 16.235 50.915 16.425 ;
        RECT 56.725 16.235 56.895 16.405 ;
        RECT 58.105 16.235 58.275 16.425 ;
        RECT 56.725 16.215 56.890 16.235 ;
        RECT 60.405 16.215 60.575 16.405 ;
        RECT 60.865 16.215 61.035 16.405 ;
        RECT 62.245 16.215 62.415 16.405 ;
        RECT 65.470 16.235 65.640 16.425 ;
        RECT 69.155 16.270 69.315 16.380 ;
        RECT 69.605 16.235 69.775 16.405 ;
        RECT 70.520 16.265 70.640 16.375 ;
        RECT 69.610 16.215 69.775 16.235 ;
        RECT 71.905 16.215 72.075 16.405 ;
        RECT 73.285 16.215 73.455 16.405 ;
        RECT 74.200 16.235 74.370 16.425 ;
        RECT 77.880 16.235 78.050 16.425 ;
        RECT 78.345 16.235 78.515 16.425 ;
        RECT 80.185 16.235 80.355 16.425 ;
        RECT 80.645 16.215 80.815 16.405 ;
        RECT 82.035 16.270 82.195 16.380 ;
        RECT 82.480 16.265 82.600 16.375 ;
        RECT 83.865 16.215 84.035 16.425 ;
        RECT 5.525 15.405 6.895 16.215 ;
        RECT 7.970 15.535 9.805 16.215 ;
        RECT 8.875 15.305 9.805 15.535 ;
        RECT 10.125 15.405 11.495 16.215 ;
        RECT 11.505 15.535 18.815 16.215 ;
        RECT 19.010 15.535 20.845 16.215 ;
        RECT 21.165 15.535 28.475 16.215 ;
        RECT 15.020 15.315 15.930 15.535 ;
        RECT 17.465 15.305 18.815 15.535 ;
        RECT 19.915 15.305 20.845 15.535 ;
        RECT 24.680 15.315 25.590 15.535 ;
        RECT 27.125 15.305 28.475 15.535 ;
        RECT 28.835 15.535 30.670 16.215 ;
        RECT 28.835 15.305 29.765 15.535 ;
        RECT 31.295 15.345 31.725 16.130 ;
        RECT 32.245 15.535 39.555 16.215 ;
        RECT 40.025 15.535 47.335 16.215 ;
        RECT 47.385 15.535 54.695 16.215 ;
        RECT 32.245 15.305 33.595 15.535 ;
        RECT 35.130 15.315 36.040 15.535 ;
        RECT 43.540 15.315 44.450 15.535 ;
        RECT 45.985 15.305 47.335 15.535 ;
        RECT 50.900 15.315 51.810 15.535 ;
        RECT 53.345 15.305 54.695 15.535 ;
        RECT 55.055 15.535 56.890 16.215 ;
        RECT 55.055 15.305 55.985 15.535 ;
        RECT 57.055 15.345 57.485 16.130 ;
        RECT 57.505 15.305 60.715 16.215 ;
        RECT 60.725 15.405 62.095 16.215 ;
        RECT 62.105 15.535 69.415 16.215 ;
        RECT 69.610 15.535 71.445 16.215 ;
        RECT 65.620 15.315 66.530 15.535 ;
        RECT 68.065 15.305 69.415 15.535 ;
        RECT 70.515 15.305 71.445 15.535 ;
        RECT 71.765 15.405 73.135 16.215 ;
        RECT 73.145 15.535 80.455 16.215 ;
        RECT 80.505 15.535 82.335 16.215 ;
        RECT 76.660 15.315 77.570 15.535 ;
        RECT 79.105 15.305 80.455 15.535 ;
        RECT 80.990 15.305 82.335 15.535 ;
        RECT 82.805 15.405 84.175 16.215 ;
      LAYER nwell ;
        RECT 5.330 12.185 84.370 15.015 ;
      LAYER pwell ;
        RECT 5.525 10.985 6.895 11.795 ;
        RECT 10.420 11.665 11.330 11.885 ;
        RECT 12.865 11.665 14.215 11.895 ;
        RECT 6.905 10.985 14.215 11.665 ;
        RECT 15.495 11.665 16.425 11.895 ;
        RECT 15.495 10.985 17.330 11.665 ;
        RECT 18.415 11.070 18.845 11.855 ;
        RECT 19.785 11.665 21.130 11.895 ;
        RECT 22.085 11.665 23.430 11.895 ;
        RECT 23.925 11.665 25.270 11.895 ;
        RECT 25.765 11.665 27.110 11.895 ;
        RECT 27.605 11.665 28.950 11.895 ;
        RECT 29.445 11.665 30.790 11.895 ;
        RECT 19.785 10.985 21.615 11.665 ;
        RECT 22.085 10.985 23.915 11.665 ;
        RECT 23.925 10.985 25.755 11.665 ;
        RECT 25.765 10.985 27.595 11.665 ;
        RECT 27.605 10.985 29.435 11.665 ;
        RECT 29.445 10.985 31.275 11.665 ;
        RECT 31.295 11.070 31.725 11.855 ;
        RECT 32.665 10.985 35.875 11.895 ;
        RECT 36.935 11.665 37.865 11.895 ;
        RECT 36.030 10.985 37.865 11.665 ;
        RECT 38.185 11.665 39.530 11.895 ;
        RECT 40.510 11.665 41.855 11.895 ;
        RECT 42.915 11.665 43.845 11.895 ;
        RECT 38.185 10.985 40.015 11.665 ;
        RECT 40.025 10.985 41.855 11.665 ;
        RECT 42.010 10.985 43.845 11.665 ;
        RECT 44.175 11.070 44.605 11.855 ;
        RECT 45.545 11.665 46.890 11.895 ;
        RECT 45.545 10.985 47.375 11.665 ;
        RECT 47.385 10.985 48.755 11.795 ;
        RECT 48.765 11.665 50.110 11.895 ;
        RECT 48.765 10.985 50.595 11.665 ;
        RECT 50.605 10.985 51.975 11.795 ;
        RECT 52.470 11.665 53.815 11.895 ;
        RECT 51.985 10.985 53.815 11.665 ;
        RECT 53.825 10.985 55.195 11.795 ;
        RECT 55.205 11.665 56.550 11.895 ;
        RECT 55.205 10.985 57.035 11.665 ;
        RECT 57.055 11.070 57.485 11.855 ;
        RECT 58.425 11.665 59.770 11.895 ;
        RECT 58.425 10.985 60.255 11.665 ;
        RECT 60.265 10.985 61.635 11.795 ;
        RECT 61.645 11.665 62.990 11.895 ;
        RECT 61.645 10.985 63.475 11.665 ;
        RECT 63.485 10.985 64.855 11.795 ;
        RECT 65.350 11.665 66.695 11.895 ;
        RECT 64.865 10.985 66.695 11.665 ;
        RECT 66.705 10.985 68.075 11.795 ;
        RECT 68.085 11.665 69.430 11.895 ;
        RECT 68.085 10.985 69.915 11.665 ;
        RECT 69.935 11.070 70.365 11.855 ;
        RECT 71.435 11.665 72.365 11.895 ;
        RECT 73.735 11.665 74.665 11.895 ;
        RECT 78.960 11.665 79.870 11.885 ;
        RECT 81.405 11.665 82.755 11.895 ;
        RECT 70.530 10.985 72.365 11.665 ;
        RECT 72.830 10.985 74.665 11.665 ;
        RECT 75.445 10.985 82.755 11.665 ;
        RECT 82.805 10.985 84.175 11.795 ;
        RECT 5.665 10.795 5.835 10.985 ;
        RECT 7.045 10.795 7.215 10.985 ;
        RECT 17.165 10.965 17.330 10.985 ;
        RECT 14.415 10.830 14.575 10.940 ;
        RECT 17.165 10.795 17.335 10.965 ;
        RECT 17.635 10.830 17.795 10.940 ;
        RECT 19.015 10.830 19.175 10.940 ;
        RECT 21.305 10.795 21.475 10.985 ;
        RECT 21.760 10.825 21.880 10.935 ;
        RECT 23.605 10.795 23.775 10.985 ;
        RECT 25.445 10.795 25.615 10.985 ;
        RECT 27.285 10.795 27.455 10.985 ;
        RECT 29.125 10.795 29.295 10.985 ;
        RECT 30.965 10.795 31.135 10.985 ;
        RECT 31.895 10.830 32.055 10.940 ;
        RECT 32.805 10.795 32.975 10.985 ;
        RECT 36.030 10.965 36.195 10.985 ;
        RECT 36.025 10.795 36.195 10.965 ;
        RECT 39.705 10.795 39.875 10.985 ;
        RECT 40.165 10.795 40.335 10.985 ;
        RECT 42.010 10.965 42.175 10.985 ;
        RECT 42.005 10.795 42.175 10.965 ;
        RECT 44.775 10.830 44.935 10.940 ;
        RECT 47.065 10.795 47.235 10.985 ;
        RECT 47.525 10.795 47.695 10.985 ;
        RECT 50.285 10.795 50.455 10.985 ;
        RECT 50.745 10.795 50.915 10.985 ;
        RECT 52.125 10.795 52.295 10.985 ;
        RECT 53.965 10.795 54.135 10.985 ;
        RECT 56.725 10.795 56.895 10.985 ;
        RECT 57.655 10.830 57.815 10.940 ;
        RECT 59.945 10.795 60.115 10.985 ;
        RECT 60.405 10.795 60.575 10.985 ;
        RECT 63.165 10.795 63.335 10.985 ;
        RECT 63.625 10.795 63.795 10.985 ;
        RECT 65.005 10.795 65.175 10.985 ;
        RECT 66.845 10.795 67.015 10.985 ;
        RECT 69.605 10.795 69.775 10.985 ;
        RECT 70.530 10.965 70.695 10.985 ;
        RECT 72.830 10.965 72.995 10.985 ;
        RECT 70.525 10.795 70.695 10.965 ;
        RECT 72.825 10.795 72.995 10.965 ;
        RECT 75.120 10.825 75.240 10.935 ;
        RECT 75.585 10.795 75.755 10.985 ;
        RECT 83.865 10.795 84.035 10.985 ;
      LAYER li1 ;
        RECT 5.520 198.475 84.180 198.645 ;
        RECT 5.605 197.385 6.815 198.475 ;
        RECT 6.985 198.040 12.330 198.475 ;
        RECT 12.505 198.040 17.850 198.475 ;
        RECT 5.605 196.675 6.125 197.215 ;
        RECT 6.295 196.845 6.815 197.385 ;
        RECT 5.605 195.925 6.815 196.675 ;
        RECT 8.570 196.470 8.910 197.300 ;
        RECT 10.390 196.790 10.740 198.040 ;
        RECT 14.090 196.470 14.430 197.300 ;
        RECT 15.910 196.790 16.260 198.040 ;
        RECT 18.485 197.310 18.775 198.475 ;
        RECT 18.945 198.040 24.290 198.475 ;
        RECT 24.465 198.040 29.810 198.475 ;
        RECT 6.985 195.925 12.330 196.470 ;
        RECT 12.505 195.925 17.850 196.470 ;
        RECT 18.485 195.925 18.775 196.650 ;
        RECT 20.530 196.470 20.870 197.300 ;
        RECT 22.350 196.790 22.700 198.040 ;
        RECT 26.050 196.470 26.390 197.300 ;
        RECT 27.870 196.790 28.220 198.040 ;
        RECT 29.985 197.385 31.195 198.475 ;
        RECT 29.985 196.675 30.505 197.215 ;
        RECT 30.675 196.845 31.195 197.385 ;
        RECT 31.365 197.310 31.655 198.475 ;
        RECT 31.825 198.040 37.170 198.475 ;
        RECT 37.345 198.040 42.690 198.475 ;
        RECT 18.945 195.925 24.290 196.470 ;
        RECT 24.465 195.925 29.810 196.470 ;
        RECT 29.985 195.925 31.195 196.675 ;
        RECT 31.365 195.925 31.655 196.650 ;
        RECT 33.410 196.470 33.750 197.300 ;
        RECT 35.230 196.790 35.580 198.040 ;
        RECT 38.930 196.470 39.270 197.300 ;
        RECT 40.750 196.790 41.100 198.040 ;
        RECT 42.865 197.385 44.075 198.475 ;
        RECT 42.865 196.675 43.385 197.215 ;
        RECT 43.555 196.845 44.075 197.385 ;
        RECT 44.245 197.310 44.535 198.475 ;
        RECT 44.705 198.040 50.050 198.475 ;
        RECT 31.825 195.925 37.170 196.470 ;
        RECT 37.345 195.925 42.690 196.470 ;
        RECT 42.865 195.925 44.075 196.675 ;
        RECT 44.245 195.925 44.535 196.650 ;
        RECT 46.290 196.470 46.630 197.300 ;
        RECT 48.110 196.790 48.460 198.040 ;
        RECT 50.225 197.605 50.500 198.305 ;
        RECT 50.670 197.930 50.925 198.475 ;
        RECT 51.095 197.965 51.575 198.305 ;
        RECT 51.750 197.920 52.355 198.475 ;
        RECT 51.740 197.820 52.355 197.920 ;
        RECT 51.740 197.795 51.925 197.820 ;
        RECT 50.225 196.575 50.395 197.605 ;
        RECT 50.670 197.475 51.425 197.725 ;
        RECT 51.595 197.550 51.925 197.795 ;
        RECT 50.670 197.440 51.440 197.475 ;
        RECT 50.670 197.430 51.455 197.440 ;
        RECT 50.565 197.415 51.460 197.430 ;
        RECT 50.565 197.400 51.480 197.415 ;
        RECT 50.565 197.390 51.500 197.400 ;
        RECT 50.565 197.380 51.525 197.390 ;
        RECT 50.565 197.350 51.595 197.380 ;
        RECT 50.565 197.320 51.615 197.350 ;
        RECT 50.565 197.290 51.635 197.320 ;
        RECT 50.565 197.265 51.665 197.290 ;
        RECT 50.565 197.230 51.700 197.265 ;
        RECT 50.565 197.225 51.730 197.230 ;
        RECT 50.565 196.830 50.795 197.225 ;
        RECT 51.340 197.220 51.730 197.225 ;
        RECT 51.365 197.210 51.730 197.220 ;
        RECT 51.380 197.205 51.730 197.210 ;
        RECT 51.395 197.200 51.730 197.205 ;
        RECT 52.095 197.200 52.355 197.650 ;
        RECT 52.525 197.385 55.115 198.475 ;
        RECT 51.395 197.195 52.355 197.200 ;
        RECT 51.405 197.185 52.355 197.195 ;
        RECT 51.415 197.180 52.355 197.185 ;
        RECT 51.425 197.170 52.355 197.180 ;
        RECT 51.430 197.160 52.355 197.170 ;
        RECT 51.435 197.155 52.355 197.160 ;
        RECT 51.445 197.140 52.355 197.155 ;
        RECT 51.450 197.125 52.355 197.140 ;
        RECT 51.460 197.100 52.355 197.125 ;
        RECT 50.965 196.630 51.295 197.055 ;
        RECT 44.705 195.925 50.050 196.470 ;
        RECT 50.225 196.095 50.485 196.575 ;
        RECT 50.655 195.925 50.905 196.465 ;
        RECT 51.075 196.145 51.295 196.630 ;
        RECT 51.465 197.030 52.355 197.100 ;
        RECT 51.465 196.305 51.635 197.030 ;
        RECT 51.805 196.475 52.355 196.860 ;
        RECT 52.525 196.695 53.735 197.215 ;
        RECT 53.905 196.865 55.115 197.385 ;
        RECT 55.375 197.545 55.545 198.305 ;
        RECT 55.725 197.715 56.055 198.475 ;
        RECT 55.375 197.375 56.040 197.545 ;
        RECT 56.225 197.400 56.495 198.305 ;
        RECT 55.870 197.230 56.040 197.375 ;
        RECT 55.305 196.825 55.635 197.195 ;
        RECT 55.870 196.900 56.155 197.230 ;
        RECT 51.465 196.135 52.355 196.305 ;
        RECT 52.525 195.925 55.115 196.695 ;
        RECT 55.870 196.645 56.040 196.900 ;
        RECT 55.375 196.475 56.040 196.645 ;
        RECT 56.325 196.600 56.495 197.400 ;
        RECT 57.125 197.310 57.415 198.475 ;
        RECT 57.585 198.040 62.930 198.475 ;
        RECT 55.375 196.095 55.545 196.475 ;
        RECT 55.725 195.925 56.055 196.305 ;
        RECT 56.235 196.095 56.495 196.600 ;
        RECT 57.125 195.925 57.415 196.650 ;
        RECT 59.170 196.470 59.510 197.300 ;
        RECT 60.990 196.790 61.340 198.040 ;
        RECT 63.105 197.385 64.775 198.475 ;
        RECT 63.105 196.695 63.855 197.215 ;
        RECT 64.025 196.865 64.775 197.385 ;
        RECT 64.945 197.400 65.215 198.305 ;
        RECT 65.385 197.715 65.715 198.475 ;
        RECT 65.895 197.545 66.065 198.305 ;
        RECT 57.585 195.925 62.930 196.470 ;
        RECT 63.105 195.925 64.775 196.695 ;
        RECT 64.945 196.600 65.115 197.400 ;
        RECT 65.400 197.375 66.065 197.545 ;
        RECT 66.325 197.385 69.835 198.475 ;
        RECT 65.400 197.230 65.570 197.375 ;
        RECT 65.285 196.900 65.570 197.230 ;
        RECT 65.400 196.645 65.570 196.900 ;
        RECT 65.805 196.825 66.135 197.195 ;
        RECT 66.325 196.695 67.975 197.215 ;
        RECT 68.145 196.865 69.835 197.385 ;
        RECT 70.005 197.310 70.295 198.475 ;
        RECT 70.465 198.040 75.810 198.475 ;
        RECT 75.985 198.040 81.330 198.475 ;
        RECT 64.945 196.095 65.205 196.600 ;
        RECT 65.400 196.475 66.065 196.645 ;
        RECT 65.385 195.925 65.715 196.305 ;
        RECT 65.895 196.095 66.065 196.475 ;
        RECT 66.325 195.925 69.835 196.695 ;
        RECT 70.005 195.925 70.295 196.650 ;
        RECT 72.050 196.470 72.390 197.300 ;
        RECT 73.870 196.790 74.220 198.040 ;
        RECT 77.570 196.470 77.910 197.300 ;
        RECT 79.390 196.790 79.740 198.040 ;
        RECT 81.505 197.385 82.715 198.475 ;
        RECT 81.505 196.675 82.025 197.215 ;
        RECT 82.195 196.845 82.715 197.385 ;
        RECT 82.885 197.385 84.095 198.475 ;
        RECT 82.885 196.845 83.405 197.385 ;
        RECT 83.575 196.675 84.095 197.215 ;
        RECT 70.465 195.925 75.810 196.470 ;
        RECT 75.985 195.925 81.330 196.470 ;
        RECT 81.505 195.925 82.715 196.675 ;
        RECT 82.885 195.925 84.095 196.675 ;
        RECT 5.520 195.755 84.180 195.925 ;
        RECT 5.605 195.005 6.815 195.755 ;
        RECT 6.985 195.210 12.330 195.755 ;
        RECT 12.505 195.210 17.850 195.755 ;
        RECT 18.025 195.210 23.370 195.755 ;
        RECT 23.545 195.210 28.890 195.755 ;
        RECT 5.605 194.465 6.125 195.005 ;
        RECT 6.295 194.295 6.815 194.835 ;
        RECT 8.570 194.380 8.910 195.210 ;
        RECT 5.605 193.205 6.815 194.295 ;
        RECT 10.390 193.640 10.740 194.890 ;
        RECT 14.090 194.380 14.430 195.210 ;
        RECT 15.910 193.640 16.260 194.890 ;
        RECT 19.610 194.380 19.950 195.210 ;
        RECT 21.430 193.640 21.780 194.890 ;
        RECT 25.130 194.380 25.470 195.210 ;
        RECT 29.065 194.985 30.735 195.755 ;
        RECT 31.365 195.030 31.655 195.755 ;
        RECT 31.825 194.985 34.415 195.755 ;
        RECT 26.950 193.640 27.300 194.890 ;
        RECT 29.065 194.465 29.815 194.985 ;
        RECT 29.985 194.295 30.735 194.815 ;
        RECT 31.825 194.465 33.035 194.985 ;
        RECT 34.595 194.945 34.865 195.755 ;
        RECT 35.035 194.945 35.365 195.585 ;
        RECT 35.535 194.945 35.775 195.755 ;
        RECT 35.965 195.375 36.855 195.545 ;
        RECT 6.985 193.205 12.330 193.640 ;
        RECT 12.505 193.205 17.850 193.640 ;
        RECT 18.025 193.205 23.370 193.640 ;
        RECT 23.545 193.205 28.890 193.640 ;
        RECT 29.065 193.205 30.735 194.295 ;
        RECT 31.365 193.205 31.655 194.370 ;
        RECT 33.205 194.295 34.415 194.815 ;
        RECT 34.585 194.515 34.935 194.765 ;
        RECT 35.105 194.345 35.275 194.945 ;
        RECT 35.965 194.820 36.515 195.205 ;
        RECT 35.445 194.515 35.795 194.765 ;
        RECT 36.685 194.650 36.855 195.375 ;
        RECT 35.965 194.580 36.855 194.650 ;
        RECT 37.025 195.050 37.245 195.535 ;
        RECT 37.415 195.215 37.665 195.755 ;
        RECT 37.835 195.105 38.095 195.585 ;
        RECT 37.025 194.625 37.355 195.050 ;
        RECT 35.965 194.555 36.860 194.580 ;
        RECT 35.965 194.540 36.870 194.555 ;
        RECT 35.965 194.525 36.875 194.540 ;
        RECT 35.965 194.520 36.885 194.525 ;
        RECT 35.965 194.510 36.890 194.520 ;
        RECT 35.965 194.500 36.895 194.510 ;
        RECT 35.965 194.495 36.905 194.500 ;
        RECT 35.965 194.485 36.915 194.495 ;
        RECT 35.965 194.480 36.925 194.485 ;
        RECT 31.825 193.205 34.415 194.295 ;
        RECT 34.595 193.205 34.925 194.345 ;
        RECT 35.105 194.175 35.785 194.345 ;
        RECT 35.455 193.390 35.785 194.175 ;
        RECT 35.965 194.030 36.225 194.480 ;
        RECT 36.590 194.475 36.925 194.480 ;
        RECT 36.590 194.470 36.940 194.475 ;
        RECT 36.590 194.460 36.955 194.470 ;
        RECT 36.590 194.455 36.980 194.460 ;
        RECT 37.525 194.455 37.755 194.850 ;
        RECT 36.590 194.450 37.755 194.455 ;
        RECT 36.620 194.415 37.755 194.450 ;
        RECT 36.655 194.390 37.755 194.415 ;
        RECT 36.685 194.360 37.755 194.390 ;
        RECT 36.705 194.330 37.755 194.360 ;
        RECT 36.725 194.300 37.755 194.330 ;
        RECT 36.795 194.290 37.755 194.300 ;
        RECT 36.820 194.280 37.755 194.290 ;
        RECT 36.840 194.265 37.755 194.280 ;
        RECT 36.860 194.250 37.755 194.265 ;
        RECT 36.865 194.240 37.650 194.250 ;
        RECT 36.880 194.205 37.650 194.240 ;
        RECT 36.395 193.885 36.725 194.130 ;
        RECT 36.895 193.955 37.650 194.205 ;
        RECT 37.925 194.075 38.095 195.105 ;
        RECT 38.355 195.205 38.525 195.495 ;
        RECT 38.695 195.375 39.025 195.755 ;
        RECT 38.355 195.035 39.020 195.205 ;
        RECT 38.270 194.215 38.620 194.865 ;
        RECT 36.395 193.860 36.580 193.885 ;
        RECT 35.965 193.760 36.580 193.860 ;
        RECT 35.965 193.205 36.570 193.760 ;
        RECT 36.745 193.375 37.225 193.715 ;
        RECT 37.395 193.205 37.650 193.750 ;
        RECT 37.820 193.375 38.095 194.075 ;
        RECT 38.790 194.045 39.020 195.035 ;
        RECT 38.355 193.875 39.020 194.045 ;
        RECT 38.355 193.375 38.525 193.875 ;
        RECT 38.695 193.205 39.025 193.705 ;
        RECT 39.195 193.375 39.380 195.495 ;
        RECT 39.635 195.295 39.885 195.755 ;
        RECT 40.055 195.305 40.390 195.475 ;
        RECT 40.585 195.305 41.260 195.475 ;
        RECT 40.055 195.165 40.225 195.305 ;
        RECT 39.550 194.175 39.830 195.125 ;
        RECT 40.000 195.035 40.225 195.165 ;
        RECT 40.000 193.930 40.170 195.035 ;
        RECT 40.395 194.885 40.920 195.105 ;
        RECT 40.340 194.120 40.580 194.715 ;
        RECT 40.750 194.185 40.920 194.885 ;
        RECT 41.090 194.525 41.260 195.305 ;
        RECT 41.580 195.255 41.950 195.755 ;
        RECT 42.130 195.305 42.535 195.475 ;
        RECT 42.705 195.305 43.490 195.475 ;
        RECT 42.130 195.075 42.300 195.305 ;
        RECT 41.470 194.775 42.300 195.075 ;
        RECT 42.685 194.805 43.150 195.135 ;
        RECT 41.470 194.745 41.670 194.775 ;
        RECT 41.790 194.525 41.960 194.595 ;
        RECT 41.090 194.355 41.960 194.525 ;
        RECT 41.450 194.265 41.960 194.355 ;
        RECT 40.000 193.800 40.305 193.930 ;
        RECT 40.750 193.820 41.280 194.185 ;
        RECT 39.620 193.205 39.885 193.665 ;
        RECT 40.055 193.375 40.305 193.800 ;
        RECT 41.450 193.650 41.620 194.265 ;
        RECT 40.515 193.480 41.620 193.650 ;
        RECT 41.790 193.205 41.960 194.005 ;
        RECT 42.130 193.705 42.300 194.775 ;
        RECT 42.470 193.875 42.660 194.595 ;
        RECT 42.830 193.845 43.150 194.805 ;
        RECT 43.320 194.845 43.490 195.305 ;
        RECT 43.765 195.225 43.975 195.755 ;
        RECT 44.235 195.015 44.565 195.540 ;
        RECT 44.735 195.145 44.905 195.755 ;
        RECT 45.075 195.100 45.405 195.535 ;
        RECT 45.075 195.015 45.455 195.100 ;
        RECT 44.365 194.845 44.565 195.015 ;
        RECT 45.230 194.975 45.455 195.015 ;
        RECT 43.320 194.515 44.195 194.845 ;
        RECT 44.365 194.515 45.115 194.845 ;
        RECT 42.130 193.375 42.380 193.705 ;
        RECT 43.320 193.675 43.490 194.515 ;
        RECT 44.365 194.310 44.555 194.515 ;
        RECT 45.285 194.395 45.455 194.975 ;
        RECT 45.625 194.985 49.135 195.755 ;
        RECT 49.395 195.205 49.565 195.495 ;
        RECT 49.735 195.375 50.065 195.755 ;
        RECT 49.395 195.035 50.060 195.205 ;
        RECT 45.625 194.465 47.275 194.985 ;
        RECT 45.240 194.345 45.455 194.395 ;
        RECT 43.660 193.935 44.555 194.310 ;
        RECT 45.065 194.265 45.455 194.345 ;
        RECT 47.445 194.295 49.135 194.815 ;
        RECT 42.605 193.505 43.490 193.675 ;
        RECT 43.670 193.205 43.985 193.705 ;
        RECT 44.215 193.375 44.555 193.935 ;
        RECT 44.725 193.205 44.895 194.215 ;
        RECT 45.065 193.420 45.395 194.265 ;
        RECT 45.625 193.205 49.135 194.295 ;
        RECT 49.310 194.215 49.660 194.865 ;
        RECT 49.830 194.045 50.060 195.035 ;
        RECT 49.395 193.875 50.060 194.045 ;
        RECT 49.395 193.375 49.565 193.875 ;
        RECT 49.735 193.205 50.065 193.705 ;
        RECT 50.235 193.375 50.420 195.495 ;
        RECT 50.675 195.295 50.925 195.755 ;
        RECT 51.095 195.305 51.430 195.475 ;
        RECT 51.625 195.305 52.300 195.475 ;
        RECT 51.095 195.165 51.265 195.305 ;
        RECT 50.590 194.175 50.870 195.125 ;
        RECT 51.040 195.035 51.265 195.165 ;
        RECT 51.040 193.930 51.210 195.035 ;
        RECT 51.435 194.885 51.960 195.105 ;
        RECT 51.380 194.120 51.620 194.715 ;
        RECT 51.790 194.185 51.960 194.885 ;
        RECT 52.130 194.525 52.300 195.305 ;
        RECT 52.620 195.255 52.990 195.755 ;
        RECT 53.170 195.305 53.575 195.475 ;
        RECT 53.745 195.305 54.530 195.475 ;
        RECT 53.170 195.075 53.340 195.305 ;
        RECT 52.510 194.775 53.340 195.075 ;
        RECT 53.725 194.805 54.190 195.135 ;
        RECT 52.510 194.745 52.710 194.775 ;
        RECT 52.830 194.525 53.000 194.595 ;
        RECT 52.130 194.355 53.000 194.525 ;
        RECT 52.490 194.265 53.000 194.355 ;
        RECT 51.040 193.800 51.345 193.930 ;
        RECT 51.790 193.820 52.320 194.185 ;
        RECT 50.660 193.205 50.925 193.665 ;
        RECT 51.095 193.375 51.345 193.800 ;
        RECT 52.490 193.650 52.660 194.265 ;
        RECT 51.555 193.480 52.660 193.650 ;
        RECT 52.830 193.205 53.000 194.005 ;
        RECT 53.170 193.705 53.340 194.775 ;
        RECT 53.510 193.875 53.700 194.595 ;
        RECT 53.870 193.845 54.190 194.805 ;
        RECT 54.360 194.845 54.530 195.305 ;
        RECT 54.805 195.225 55.015 195.755 ;
        RECT 55.275 195.015 55.605 195.540 ;
        RECT 55.775 195.145 55.945 195.755 ;
        RECT 56.115 195.100 56.445 195.535 ;
        RECT 56.115 195.015 56.495 195.100 ;
        RECT 57.125 195.030 57.415 195.755 ;
        RECT 55.405 194.845 55.605 195.015 ;
        RECT 56.270 194.975 56.495 195.015 ;
        RECT 54.360 194.515 55.235 194.845 ;
        RECT 55.405 194.515 56.155 194.845 ;
        RECT 53.170 193.375 53.420 193.705 ;
        RECT 54.360 193.675 54.530 194.515 ;
        RECT 55.405 194.310 55.595 194.515 ;
        RECT 56.325 194.395 56.495 194.975 ;
        RECT 57.585 194.985 59.255 195.755 ;
        RECT 59.935 195.100 60.265 195.535 ;
        RECT 60.435 195.145 60.605 195.755 ;
        RECT 59.885 195.015 60.265 195.100 ;
        RECT 60.775 195.015 61.105 195.540 ;
        RECT 61.365 195.225 61.575 195.755 ;
        RECT 61.850 195.305 62.635 195.475 ;
        RECT 62.805 195.305 63.210 195.475 ;
        RECT 57.585 194.465 58.335 194.985 ;
        RECT 59.885 194.975 60.110 195.015 ;
        RECT 56.280 194.345 56.495 194.395 ;
        RECT 54.700 193.935 55.595 194.310 ;
        RECT 56.105 194.265 56.495 194.345 ;
        RECT 53.645 193.505 54.530 193.675 ;
        RECT 54.710 193.205 55.025 193.705 ;
        RECT 55.255 193.375 55.595 193.935 ;
        RECT 55.765 193.205 55.935 194.215 ;
        RECT 56.105 193.420 56.435 194.265 ;
        RECT 57.125 193.205 57.415 194.370 ;
        RECT 58.505 194.295 59.255 194.815 ;
        RECT 57.585 193.205 59.255 194.295 ;
        RECT 59.885 194.395 60.055 194.975 ;
        RECT 60.775 194.845 60.975 195.015 ;
        RECT 61.850 194.845 62.020 195.305 ;
        RECT 60.225 194.515 60.975 194.845 ;
        RECT 61.145 194.515 62.020 194.845 ;
        RECT 59.885 194.345 60.100 194.395 ;
        RECT 59.885 194.265 60.275 194.345 ;
        RECT 59.945 193.420 60.275 194.265 ;
        RECT 60.785 194.310 60.975 194.515 ;
        RECT 60.445 193.205 60.615 194.215 ;
        RECT 60.785 193.935 61.680 194.310 ;
        RECT 60.785 193.375 61.125 193.935 ;
        RECT 61.355 193.205 61.670 193.705 ;
        RECT 61.850 193.675 62.020 194.515 ;
        RECT 62.190 194.805 62.655 195.135 ;
        RECT 63.040 195.075 63.210 195.305 ;
        RECT 63.390 195.255 63.760 195.755 ;
        RECT 64.080 195.305 64.755 195.475 ;
        RECT 64.950 195.305 65.285 195.475 ;
        RECT 62.190 193.845 62.510 194.805 ;
        RECT 63.040 194.775 63.870 195.075 ;
        RECT 62.680 193.875 62.870 194.595 ;
        RECT 63.040 193.705 63.210 194.775 ;
        RECT 63.670 194.745 63.870 194.775 ;
        RECT 63.380 194.525 63.550 194.595 ;
        RECT 64.080 194.525 64.250 195.305 ;
        RECT 65.115 195.165 65.285 195.305 ;
        RECT 65.455 195.295 65.705 195.755 ;
        RECT 63.380 194.355 64.250 194.525 ;
        RECT 64.420 194.885 64.945 195.105 ;
        RECT 65.115 195.035 65.340 195.165 ;
        RECT 63.380 194.265 63.890 194.355 ;
        RECT 61.850 193.505 62.735 193.675 ;
        RECT 62.960 193.375 63.210 193.705 ;
        RECT 63.380 193.205 63.550 194.005 ;
        RECT 63.720 193.650 63.890 194.265 ;
        RECT 64.420 194.185 64.590 194.885 ;
        RECT 64.060 193.820 64.590 194.185 ;
        RECT 64.760 194.120 65.000 194.715 ;
        RECT 65.170 193.930 65.340 195.035 ;
        RECT 65.510 194.175 65.790 195.125 ;
        RECT 65.035 193.800 65.340 193.930 ;
        RECT 63.720 193.480 64.825 193.650 ;
        RECT 65.035 193.375 65.285 193.800 ;
        RECT 65.455 193.205 65.720 193.665 ;
        RECT 65.960 193.375 66.145 195.495 ;
        RECT 66.315 195.375 66.645 195.755 ;
        RECT 66.815 195.205 66.985 195.495 ;
        RECT 67.245 195.210 72.590 195.755 ;
        RECT 72.765 195.210 78.110 195.755 ;
        RECT 66.320 195.035 66.985 195.205 ;
        RECT 66.320 194.045 66.550 195.035 ;
        RECT 66.720 194.215 67.070 194.865 ;
        RECT 68.830 194.380 69.170 195.210 ;
        RECT 66.320 193.875 66.985 194.045 ;
        RECT 66.315 193.205 66.645 193.705 ;
        RECT 66.815 193.375 66.985 193.875 ;
        RECT 70.650 193.640 71.000 194.890 ;
        RECT 74.350 194.380 74.690 195.210 ;
        RECT 78.285 194.985 81.795 195.755 ;
        RECT 82.885 195.005 84.095 195.755 ;
        RECT 76.170 193.640 76.520 194.890 ;
        RECT 78.285 194.465 79.935 194.985 ;
        RECT 80.105 194.295 81.795 194.815 ;
        RECT 67.245 193.205 72.590 193.640 ;
        RECT 72.765 193.205 78.110 193.640 ;
        RECT 78.285 193.205 81.795 194.295 ;
        RECT 82.885 194.295 83.405 194.835 ;
        RECT 83.575 194.465 84.095 195.005 ;
        RECT 82.885 193.205 84.095 194.295 ;
        RECT 5.520 193.035 84.180 193.205 ;
        RECT 5.605 191.945 6.815 193.035 ;
        RECT 6.985 192.600 12.330 193.035 ;
        RECT 12.505 192.600 17.850 193.035 ;
        RECT 5.605 191.235 6.125 191.775 ;
        RECT 6.295 191.405 6.815 191.945 ;
        RECT 5.605 190.485 6.815 191.235 ;
        RECT 8.570 191.030 8.910 191.860 ;
        RECT 10.390 191.350 10.740 192.600 ;
        RECT 14.090 191.030 14.430 191.860 ;
        RECT 15.910 191.350 16.260 192.600 ;
        RECT 18.485 191.870 18.775 193.035 ;
        RECT 18.945 192.600 24.290 193.035 ;
        RECT 24.465 192.600 29.810 193.035 ;
        RECT 6.985 190.485 12.330 191.030 ;
        RECT 12.505 190.485 17.850 191.030 ;
        RECT 18.485 190.485 18.775 191.210 ;
        RECT 20.530 191.030 20.870 191.860 ;
        RECT 22.350 191.350 22.700 192.600 ;
        RECT 26.050 191.030 26.390 191.860 ;
        RECT 27.870 191.350 28.220 192.600 ;
        RECT 30.535 192.365 30.705 192.865 ;
        RECT 30.875 192.535 31.205 193.035 ;
        RECT 30.535 192.195 31.200 192.365 ;
        RECT 30.450 191.375 30.800 192.025 ;
        RECT 30.970 191.205 31.200 192.195 ;
        RECT 30.535 191.035 31.200 191.205 ;
        RECT 18.945 190.485 24.290 191.030 ;
        RECT 24.465 190.485 29.810 191.030 ;
        RECT 30.535 190.745 30.705 191.035 ;
        RECT 30.875 190.485 31.205 190.865 ;
        RECT 31.375 190.745 31.560 192.865 ;
        RECT 31.800 192.575 32.065 193.035 ;
        RECT 32.235 192.440 32.485 192.865 ;
        RECT 32.695 192.590 33.800 192.760 ;
        RECT 32.180 192.310 32.485 192.440 ;
        RECT 31.730 191.115 32.010 192.065 ;
        RECT 32.180 191.205 32.350 192.310 ;
        RECT 32.520 191.525 32.760 192.120 ;
        RECT 32.930 192.055 33.460 192.420 ;
        RECT 32.930 191.355 33.100 192.055 ;
        RECT 33.630 191.975 33.800 192.590 ;
        RECT 33.970 192.235 34.140 193.035 ;
        RECT 34.310 192.535 34.560 192.865 ;
        RECT 34.785 192.565 35.670 192.735 ;
        RECT 33.630 191.885 34.140 191.975 ;
        RECT 32.180 191.075 32.405 191.205 ;
        RECT 32.575 191.135 33.100 191.355 ;
        RECT 33.270 191.715 34.140 191.885 ;
        RECT 31.815 190.485 32.065 190.945 ;
        RECT 32.235 190.935 32.405 191.075 ;
        RECT 33.270 190.935 33.440 191.715 ;
        RECT 33.970 191.645 34.140 191.715 ;
        RECT 33.650 191.465 33.850 191.495 ;
        RECT 34.310 191.465 34.480 192.535 ;
        RECT 34.650 191.645 34.840 192.365 ;
        RECT 33.650 191.165 34.480 191.465 ;
        RECT 35.010 191.435 35.330 192.395 ;
        RECT 32.235 190.765 32.570 190.935 ;
        RECT 32.765 190.765 33.440 190.935 ;
        RECT 33.760 190.485 34.130 190.985 ;
        RECT 34.310 190.935 34.480 191.165 ;
        RECT 34.865 191.105 35.330 191.435 ;
        RECT 35.500 191.725 35.670 192.565 ;
        RECT 35.850 192.535 36.165 193.035 ;
        RECT 36.395 192.305 36.735 192.865 ;
        RECT 35.840 191.930 36.735 192.305 ;
        RECT 36.905 192.025 37.075 193.035 ;
        RECT 36.545 191.725 36.735 191.930 ;
        RECT 37.245 191.975 37.575 192.820 ;
        RECT 38.265 192.165 38.540 192.865 ;
        RECT 38.710 192.490 38.965 193.035 ;
        RECT 39.135 192.525 39.615 192.865 ;
        RECT 39.790 192.480 40.395 193.035 ;
        RECT 39.780 192.380 40.395 192.480 ;
        RECT 39.780 192.355 39.965 192.380 ;
        RECT 37.245 191.895 37.635 191.975 ;
        RECT 37.420 191.845 37.635 191.895 ;
        RECT 35.500 191.395 36.375 191.725 ;
        RECT 36.545 191.395 37.295 191.725 ;
        RECT 35.500 190.935 35.670 191.395 ;
        RECT 36.545 191.225 36.745 191.395 ;
        RECT 37.465 191.265 37.635 191.845 ;
        RECT 37.410 191.225 37.635 191.265 ;
        RECT 34.310 190.765 34.715 190.935 ;
        RECT 34.885 190.765 35.670 190.935 ;
        RECT 35.945 190.485 36.155 191.015 ;
        RECT 36.415 190.700 36.745 191.225 ;
        RECT 37.255 191.140 37.635 191.225 ;
        RECT 36.915 190.485 37.085 191.095 ;
        RECT 37.255 190.705 37.585 191.140 ;
        RECT 38.265 191.135 38.435 192.165 ;
        RECT 38.710 192.035 39.465 192.285 ;
        RECT 39.635 192.110 39.965 192.355 ;
        RECT 38.710 192.000 39.480 192.035 ;
        RECT 38.710 191.990 39.495 192.000 ;
        RECT 38.605 191.975 39.500 191.990 ;
        RECT 38.605 191.960 39.520 191.975 ;
        RECT 38.605 191.950 39.540 191.960 ;
        RECT 38.605 191.940 39.565 191.950 ;
        RECT 38.605 191.910 39.635 191.940 ;
        RECT 38.605 191.880 39.655 191.910 ;
        RECT 38.605 191.850 39.675 191.880 ;
        RECT 38.605 191.825 39.705 191.850 ;
        RECT 38.605 191.790 39.740 191.825 ;
        RECT 38.605 191.785 39.770 191.790 ;
        RECT 38.605 191.390 38.835 191.785 ;
        RECT 39.380 191.780 39.770 191.785 ;
        RECT 39.405 191.770 39.770 191.780 ;
        RECT 39.420 191.765 39.770 191.770 ;
        RECT 39.435 191.760 39.770 191.765 ;
        RECT 40.135 191.760 40.395 192.210 ;
        RECT 40.575 192.065 40.905 192.850 ;
        RECT 40.575 191.895 41.255 192.065 ;
        RECT 41.435 191.895 41.765 193.035 ;
        RECT 41.945 192.480 42.550 193.035 ;
        RECT 42.725 192.525 43.205 192.865 ;
        RECT 43.375 192.490 43.630 193.035 ;
        RECT 41.945 192.380 42.560 192.480 ;
        RECT 42.375 192.355 42.560 192.380 ;
        RECT 39.435 191.755 40.395 191.760 ;
        RECT 39.445 191.745 40.395 191.755 ;
        RECT 39.455 191.740 40.395 191.745 ;
        RECT 39.465 191.730 40.395 191.740 ;
        RECT 39.470 191.720 40.395 191.730 ;
        RECT 39.475 191.715 40.395 191.720 ;
        RECT 39.485 191.700 40.395 191.715 ;
        RECT 39.490 191.685 40.395 191.700 ;
        RECT 39.500 191.660 40.395 191.685 ;
        RECT 39.005 191.190 39.335 191.615 ;
        RECT 38.265 190.655 38.525 191.135 ;
        RECT 38.695 190.485 38.945 191.025 ;
        RECT 39.115 190.705 39.335 191.190 ;
        RECT 39.505 191.590 40.395 191.660 ;
        RECT 39.505 190.865 39.675 191.590 ;
        RECT 40.565 191.475 40.915 191.725 ;
        RECT 39.845 191.035 40.395 191.420 ;
        RECT 41.085 191.295 41.255 191.895 ;
        RECT 41.945 191.760 42.205 192.210 ;
        RECT 42.375 192.110 42.705 192.355 ;
        RECT 42.875 192.035 43.630 192.285 ;
        RECT 43.800 192.165 44.075 192.865 ;
        RECT 42.860 192.000 43.630 192.035 ;
        RECT 42.845 191.990 43.630 192.000 ;
        RECT 42.840 191.975 43.735 191.990 ;
        RECT 42.820 191.960 43.735 191.975 ;
        RECT 42.800 191.950 43.735 191.960 ;
        RECT 42.775 191.940 43.735 191.950 ;
        RECT 42.705 191.910 43.735 191.940 ;
        RECT 42.685 191.880 43.735 191.910 ;
        RECT 42.665 191.850 43.735 191.880 ;
        RECT 42.635 191.825 43.735 191.850 ;
        RECT 42.600 191.790 43.735 191.825 ;
        RECT 42.570 191.785 43.735 191.790 ;
        RECT 42.570 191.780 42.960 191.785 ;
        RECT 42.570 191.770 42.935 191.780 ;
        RECT 42.570 191.765 42.920 191.770 ;
        RECT 42.570 191.760 42.905 191.765 ;
        RECT 41.945 191.755 42.905 191.760 ;
        RECT 41.945 191.745 42.895 191.755 ;
        RECT 41.945 191.740 42.885 191.745 ;
        RECT 41.945 191.730 42.875 191.740 ;
        RECT 41.425 191.475 41.775 191.725 ;
        RECT 41.945 191.720 42.870 191.730 ;
        RECT 41.945 191.715 42.865 191.720 ;
        RECT 41.945 191.700 42.855 191.715 ;
        RECT 41.945 191.685 42.850 191.700 ;
        RECT 41.945 191.660 42.840 191.685 ;
        RECT 41.945 191.590 42.835 191.660 ;
        RECT 39.505 190.695 40.395 190.865 ;
        RECT 40.585 190.485 40.825 191.295 ;
        RECT 40.995 190.655 41.325 191.295 ;
        RECT 41.495 190.485 41.765 191.295 ;
        RECT 41.945 191.035 42.495 191.420 ;
        RECT 42.665 190.865 42.835 191.590 ;
        RECT 41.945 190.695 42.835 190.865 ;
        RECT 43.005 191.190 43.335 191.615 ;
        RECT 43.505 191.390 43.735 191.785 ;
        RECT 43.005 190.705 43.225 191.190 ;
        RECT 43.905 191.135 44.075 192.165 ;
        RECT 44.245 191.870 44.535 193.035 ;
        RECT 44.795 192.365 44.965 192.865 ;
        RECT 45.135 192.535 45.465 193.035 ;
        RECT 44.795 192.195 45.460 192.365 ;
        RECT 44.710 191.375 45.060 192.025 ;
        RECT 43.395 190.485 43.645 191.025 ;
        RECT 43.815 190.655 44.075 191.135 ;
        RECT 44.245 190.485 44.535 191.210 ;
        RECT 45.230 191.205 45.460 192.195 ;
        RECT 44.795 191.035 45.460 191.205 ;
        RECT 44.795 190.745 44.965 191.035 ;
        RECT 45.135 190.485 45.465 190.865 ;
        RECT 45.635 190.745 45.820 192.865 ;
        RECT 46.060 192.575 46.325 193.035 ;
        RECT 46.495 192.440 46.745 192.865 ;
        RECT 46.955 192.590 48.060 192.760 ;
        RECT 46.440 192.310 46.745 192.440 ;
        RECT 45.990 191.115 46.270 192.065 ;
        RECT 46.440 191.205 46.610 192.310 ;
        RECT 46.780 191.525 47.020 192.120 ;
        RECT 47.190 192.055 47.720 192.420 ;
        RECT 47.190 191.355 47.360 192.055 ;
        RECT 47.890 191.975 48.060 192.590 ;
        RECT 48.230 192.235 48.400 193.035 ;
        RECT 48.570 192.535 48.820 192.865 ;
        RECT 49.045 192.565 49.930 192.735 ;
        RECT 47.890 191.885 48.400 191.975 ;
        RECT 46.440 191.075 46.665 191.205 ;
        RECT 46.835 191.135 47.360 191.355 ;
        RECT 47.530 191.715 48.400 191.885 ;
        RECT 46.075 190.485 46.325 190.945 ;
        RECT 46.495 190.935 46.665 191.075 ;
        RECT 47.530 190.935 47.700 191.715 ;
        RECT 48.230 191.645 48.400 191.715 ;
        RECT 47.910 191.465 48.110 191.495 ;
        RECT 48.570 191.465 48.740 192.535 ;
        RECT 48.910 191.645 49.100 192.365 ;
        RECT 47.910 191.165 48.740 191.465 ;
        RECT 49.270 191.435 49.590 192.395 ;
        RECT 46.495 190.765 46.830 190.935 ;
        RECT 47.025 190.765 47.700 190.935 ;
        RECT 48.020 190.485 48.390 190.985 ;
        RECT 48.570 190.935 48.740 191.165 ;
        RECT 49.125 191.105 49.590 191.435 ;
        RECT 49.760 191.725 49.930 192.565 ;
        RECT 50.110 192.535 50.425 193.035 ;
        RECT 50.655 192.305 50.995 192.865 ;
        RECT 50.100 191.930 50.995 192.305 ;
        RECT 51.165 192.025 51.335 193.035 ;
        RECT 50.805 191.725 50.995 191.930 ;
        RECT 51.505 191.975 51.835 192.820 ;
        RECT 51.505 191.895 51.895 191.975 ;
        RECT 52.995 191.895 53.325 193.035 ;
        RECT 53.855 192.065 54.185 192.850 ;
        RECT 53.505 191.895 54.185 192.065 ;
        RECT 55.295 191.895 55.625 193.035 ;
        RECT 56.155 192.065 56.485 192.850 ;
        RECT 55.805 191.895 56.485 192.065 ;
        RECT 56.665 191.945 57.875 193.035 ;
        RECT 51.680 191.845 51.895 191.895 ;
        RECT 49.760 191.395 50.635 191.725 ;
        RECT 50.805 191.395 51.555 191.725 ;
        RECT 49.760 190.935 49.930 191.395 ;
        RECT 50.805 191.225 51.005 191.395 ;
        RECT 51.725 191.265 51.895 191.845 ;
        RECT 52.985 191.475 53.335 191.725 ;
        RECT 53.505 191.295 53.675 191.895 ;
        RECT 53.845 191.475 54.195 191.725 ;
        RECT 55.285 191.475 55.635 191.725 ;
        RECT 55.805 191.295 55.975 191.895 ;
        RECT 56.145 191.475 56.495 191.725 ;
        RECT 51.670 191.225 51.895 191.265 ;
        RECT 48.570 190.765 48.975 190.935 ;
        RECT 49.145 190.765 49.930 190.935 ;
        RECT 50.205 190.485 50.415 191.015 ;
        RECT 50.675 190.700 51.005 191.225 ;
        RECT 51.515 191.140 51.895 191.225 ;
        RECT 51.175 190.485 51.345 191.095 ;
        RECT 51.515 190.705 51.845 191.140 ;
        RECT 52.995 190.485 53.265 191.295 ;
        RECT 53.435 190.655 53.765 191.295 ;
        RECT 53.935 190.485 54.175 191.295 ;
        RECT 55.295 190.485 55.565 191.295 ;
        RECT 55.735 190.655 56.065 191.295 ;
        RECT 56.235 190.485 56.475 191.295 ;
        RECT 56.665 191.235 57.185 191.775 ;
        RECT 57.355 191.405 57.875 191.945 ;
        RECT 58.055 191.895 58.385 193.035 ;
        RECT 58.915 192.065 59.245 192.850 ;
        RECT 59.425 192.480 60.030 193.035 ;
        RECT 60.205 192.525 60.685 192.865 ;
        RECT 60.855 192.490 61.110 193.035 ;
        RECT 59.425 192.380 60.040 192.480 ;
        RECT 59.855 192.355 60.040 192.380 ;
        RECT 58.565 191.895 59.245 192.065 ;
        RECT 58.045 191.475 58.395 191.725 ;
        RECT 58.565 191.295 58.735 191.895 ;
        RECT 59.425 191.760 59.685 192.210 ;
        RECT 59.855 192.110 60.185 192.355 ;
        RECT 60.355 192.035 61.110 192.285 ;
        RECT 61.280 192.165 61.555 192.865 ;
        RECT 60.340 192.000 61.110 192.035 ;
        RECT 60.325 191.990 61.110 192.000 ;
        RECT 60.320 191.975 61.215 191.990 ;
        RECT 60.300 191.960 61.215 191.975 ;
        RECT 60.280 191.950 61.215 191.960 ;
        RECT 60.255 191.940 61.215 191.950 ;
        RECT 60.185 191.910 61.215 191.940 ;
        RECT 60.165 191.880 61.215 191.910 ;
        RECT 60.145 191.850 61.215 191.880 ;
        RECT 60.115 191.825 61.215 191.850 ;
        RECT 60.080 191.790 61.215 191.825 ;
        RECT 60.050 191.785 61.215 191.790 ;
        RECT 60.050 191.780 60.440 191.785 ;
        RECT 60.050 191.770 60.415 191.780 ;
        RECT 60.050 191.765 60.400 191.770 ;
        RECT 60.050 191.760 60.385 191.765 ;
        RECT 59.425 191.755 60.385 191.760 ;
        RECT 59.425 191.745 60.375 191.755 ;
        RECT 59.425 191.740 60.365 191.745 ;
        RECT 59.425 191.730 60.355 191.740 ;
        RECT 58.905 191.475 59.255 191.725 ;
        RECT 59.425 191.720 60.350 191.730 ;
        RECT 59.425 191.715 60.345 191.720 ;
        RECT 59.425 191.700 60.335 191.715 ;
        RECT 59.425 191.685 60.330 191.700 ;
        RECT 59.425 191.660 60.320 191.685 ;
        RECT 59.425 191.590 60.315 191.660 ;
        RECT 56.665 190.485 57.875 191.235 ;
        RECT 58.055 190.485 58.325 191.295 ;
        RECT 58.495 190.655 58.825 191.295 ;
        RECT 58.995 190.485 59.235 191.295 ;
        RECT 59.425 191.035 59.975 191.420 ;
        RECT 60.145 190.865 60.315 191.590 ;
        RECT 59.425 190.695 60.315 190.865 ;
        RECT 60.485 191.190 60.815 191.615 ;
        RECT 60.985 191.390 61.215 191.785 ;
        RECT 60.485 190.705 60.705 191.190 ;
        RECT 61.385 191.135 61.555 192.165 ;
        RECT 62.705 191.975 63.035 192.820 ;
        RECT 63.205 192.025 63.375 193.035 ;
        RECT 63.545 192.305 63.885 192.865 ;
        RECT 64.115 192.535 64.430 193.035 ;
        RECT 64.610 192.565 65.495 192.735 ;
        RECT 62.645 191.895 63.035 191.975 ;
        RECT 63.545 191.930 64.440 192.305 ;
        RECT 62.645 191.845 62.860 191.895 ;
        RECT 62.645 191.265 62.815 191.845 ;
        RECT 63.545 191.725 63.735 191.930 ;
        RECT 64.610 191.725 64.780 192.565 ;
        RECT 65.720 192.535 65.970 192.865 ;
        RECT 62.985 191.395 63.735 191.725 ;
        RECT 63.905 191.395 64.780 191.725 ;
        RECT 62.645 191.225 62.870 191.265 ;
        RECT 63.535 191.225 63.735 191.395 ;
        RECT 62.645 191.140 63.025 191.225 ;
        RECT 60.875 190.485 61.125 191.025 ;
        RECT 61.295 190.655 61.555 191.135 ;
        RECT 62.695 190.705 63.025 191.140 ;
        RECT 63.195 190.485 63.365 191.095 ;
        RECT 63.535 190.700 63.865 191.225 ;
        RECT 64.125 190.485 64.335 191.015 ;
        RECT 64.610 190.935 64.780 191.395 ;
        RECT 64.950 191.435 65.270 192.395 ;
        RECT 65.440 191.645 65.630 192.365 ;
        RECT 65.800 191.465 65.970 192.535 ;
        RECT 66.140 192.235 66.310 193.035 ;
        RECT 66.480 192.590 67.585 192.760 ;
        RECT 66.480 191.975 66.650 192.590 ;
        RECT 67.795 192.440 68.045 192.865 ;
        RECT 68.215 192.575 68.480 193.035 ;
        RECT 66.820 192.055 67.350 192.420 ;
        RECT 67.795 192.310 68.100 192.440 ;
        RECT 66.140 191.885 66.650 191.975 ;
        RECT 66.140 191.715 67.010 191.885 ;
        RECT 66.140 191.645 66.310 191.715 ;
        RECT 66.430 191.465 66.630 191.495 ;
        RECT 64.950 191.105 65.415 191.435 ;
        RECT 65.800 191.165 66.630 191.465 ;
        RECT 65.800 190.935 65.970 191.165 ;
        RECT 64.610 190.765 65.395 190.935 ;
        RECT 65.565 190.765 65.970 190.935 ;
        RECT 66.150 190.485 66.520 190.985 ;
        RECT 66.840 190.935 67.010 191.715 ;
        RECT 67.180 191.355 67.350 192.055 ;
        RECT 67.520 191.525 67.760 192.120 ;
        RECT 67.180 191.135 67.705 191.355 ;
        RECT 67.930 191.205 68.100 192.310 ;
        RECT 67.875 191.075 68.100 191.205 ;
        RECT 68.270 191.115 68.550 192.065 ;
        RECT 67.875 190.935 68.045 191.075 ;
        RECT 66.840 190.765 67.515 190.935 ;
        RECT 67.710 190.765 68.045 190.935 ;
        RECT 68.215 190.485 68.465 190.945 ;
        RECT 68.720 190.745 68.905 192.865 ;
        RECT 69.075 192.535 69.405 193.035 ;
        RECT 69.575 192.365 69.745 192.865 ;
        RECT 69.080 192.195 69.745 192.365 ;
        RECT 69.080 191.205 69.310 192.195 ;
        RECT 69.480 191.375 69.830 192.025 ;
        RECT 70.005 191.870 70.295 193.035 ;
        RECT 70.465 192.600 75.810 193.035 ;
        RECT 75.985 192.600 81.330 193.035 ;
        RECT 69.080 191.035 69.745 191.205 ;
        RECT 69.075 190.485 69.405 190.865 ;
        RECT 69.575 190.745 69.745 191.035 ;
        RECT 70.005 190.485 70.295 191.210 ;
        RECT 72.050 191.030 72.390 191.860 ;
        RECT 73.870 191.350 74.220 192.600 ;
        RECT 77.570 191.030 77.910 191.860 ;
        RECT 79.390 191.350 79.740 192.600 ;
        RECT 81.505 191.945 82.715 193.035 ;
        RECT 81.505 191.235 82.025 191.775 ;
        RECT 82.195 191.405 82.715 191.945 ;
        RECT 82.885 191.945 84.095 193.035 ;
        RECT 82.885 191.405 83.405 191.945 ;
        RECT 83.575 191.235 84.095 191.775 ;
        RECT 70.465 190.485 75.810 191.030 ;
        RECT 75.985 190.485 81.330 191.030 ;
        RECT 81.505 190.485 82.715 191.235 ;
        RECT 82.885 190.485 84.095 191.235 ;
        RECT 5.520 190.315 84.180 190.485 ;
        RECT 5.605 189.565 6.815 190.315 ;
        RECT 6.985 189.770 12.330 190.315 ;
        RECT 12.505 189.770 17.850 190.315 ;
        RECT 18.025 189.770 23.370 190.315 ;
        RECT 23.545 189.770 28.890 190.315 ;
        RECT 5.605 189.025 6.125 189.565 ;
        RECT 6.295 188.855 6.815 189.395 ;
        RECT 8.570 188.940 8.910 189.770 ;
        RECT 5.605 187.765 6.815 188.855 ;
        RECT 10.390 188.200 10.740 189.450 ;
        RECT 14.090 188.940 14.430 189.770 ;
        RECT 15.910 188.200 16.260 189.450 ;
        RECT 19.610 188.940 19.950 189.770 ;
        RECT 21.430 188.200 21.780 189.450 ;
        RECT 25.130 188.940 25.470 189.770 ;
        RECT 29.065 189.545 30.735 190.315 ;
        RECT 31.365 189.590 31.655 190.315 ;
        RECT 31.825 189.565 33.035 190.315 ;
        RECT 33.205 189.665 33.465 190.145 ;
        RECT 33.635 189.775 33.885 190.315 ;
        RECT 26.950 188.200 27.300 189.450 ;
        RECT 29.065 189.025 29.815 189.545 ;
        RECT 29.985 188.855 30.735 189.375 ;
        RECT 31.825 189.025 32.345 189.565 ;
        RECT 6.985 187.765 12.330 188.200 ;
        RECT 12.505 187.765 17.850 188.200 ;
        RECT 18.025 187.765 23.370 188.200 ;
        RECT 23.545 187.765 28.890 188.200 ;
        RECT 29.065 187.765 30.735 188.855 ;
        RECT 31.365 187.765 31.655 188.930 ;
        RECT 32.515 188.855 33.035 189.395 ;
        RECT 31.825 187.765 33.035 188.855 ;
        RECT 33.205 188.635 33.375 189.665 ;
        RECT 34.055 189.610 34.275 190.095 ;
        RECT 33.545 189.015 33.775 189.410 ;
        RECT 33.945 189.185 34.275 189.610 ;
        RECT 34.445 189.935 35.335 190.105 ;
        RECT 34.445 189.210 34.615 189.935 ;
        RECT 34.785 189.380 35.335 189.765 ;
        RECT 35.525 189.505 35.765 190.315 ;
        RECT 35.935 189.505 36.265 190.145 ;
        RECT 36.435 189.505 36.705 190.315 ;
        RECT 36.970 189.815 37.465 190.145 ;
        RECT 34.445 189.140 35.335 189.210 ;
        RECT 34.440 189.115 35.335 189.140 ;
        RECT 34.430 189.100 35.335 189.115 ;
        RECT 34.425 189.085 35.335 189.100 ;
        RECT 34.415 189.080 35.335 189.085 ;
        RECT 34.410 189.070 35.335 189.080 ;
        RECT 35.505 189.075 35.855 189.325 ;
        RECT 34.405 189.060 35.335 189.070 ;
        RECT 34.395 189.055 35.335 189.060 ;
        RECT 34.385 189.045 35.335 189.055 ;
        RECT 34.375 189.040 35.335 189.045 ;
        RECT 34.375 189.035 34.710 189.040 ;
        RECT 34.360 189.030 34.710 189.035 ;
        RECT 34.345 189.020 34.710 189.030 ;
        RECT 34.320 189.015 34.710 189.020 ;
        RECT 33.545 189.010 34.710 189.015 ;
        RECT 33.545 188.975 34.680 189.010 ;
        RECT 33.545 188.950 34.645 188.975 ;
        RECT 33.545 188.920 34.615 188.950 ;
        RECT 33.545 188.890 34.595 188.920 ;
        RECT 33.545 188.860 34.575 188.890 ;
        RECT 33.545 188.850 34.505 188.860 ;
        RECT 33.545 188.840 34.480 188.850 ;
        RECT 33.545 188.825 34.460 188.840 ;
        RECT 33.545 188.810 34.440 188.825 ;
        RECT 33.650 188.800 34.435 188.810 ;
        RECT 33.650 188.765 34.420 188.800 ;
        RECT 33.205 187.935 33.480 188.635 ;
        RECT 33.650 188.515 34.405 188.765 ;
        RECT 34.575 188.445 34.905 188.690 ;
        RECT 35.075 188.590 35.335 189.040 ;
        RECT 36.025 188.905 36.195 189.505 ;
        RECT 36.365 189.075 36.715 189.325 ;
        RECT 35.515 188.735 36.195 188.905 ;
        RECT 34.720 188.420 34.905 188.445 ;
        RECT 34.720 188.320 35.335 188.420 ;
        RECT 33.650 187.765 33.905 188.310 ;
        RECT 34.075 187.935 34.555 188.275 ;
        RECT 34.730 187.765 35.335 188.320 ;
        RECT 35.515 187.950 35.845 188.735 ;
        RECT 36.375 187.765 36.705 188.905 ;
        RECT 36.885 188.325 37.125 189.635 ;
        RECT 37.295 188.905 37.465 189.815 ;
        RECT 37.685 189.075 38.035 190.040 ;
        RECT 38.215 189.075 38.515 190.045 ;
        RECT 38.695 189.075 38.975 190.045 ;
        RECT 39.155 189.515 39.425 190.315 ;
        RECT 39.595 189.595 39.935 190.105 ;
        RECT 40.130 189.925 40.460 190.315 ;
        RECT 40.630 189.755 40.855 190.135 ;
        RECT 39.170 189.075 39.500 189.325 ;
        RECT 39.170 188.905 39.485 189.075 ;
        RECT 37.295 188.735 39.485 188.905 ;
        RECT 36.890 187.765 37.225 188.145 ;
        RECT 37.395 187.935 37.645 188.735 ;
        RECT 37.865 187.765 38.195 188.485 ;
        RECT 38.380 187.935 38.630 188.735 ;
        RECT 39.095 187.765 39.425 188.565 ;
        RECT 39.675 188.195 39.935 189.595 ;
        RECT 40.115 189.075 40.355 189.725 ;
        RECT 40.525 189.575 40.855 189.755 ;
        RECT 40.525 188.905 40.700 189.575 ;
        RECT 41.055 189.405 41.285 190.025 ;
        RECT 41.465 189.585 41.765 190.315 ;
        RECT 41.945 189.480 42.235 190.315 ;
        RECT 42.405 189.915 43.360 190.085 ;
        RECT 43.775 189.925 44.105 190.315 ;
        RECT 40.870 189.075 41.285 189.405 ;
        RECT 41.465 189.075 41.760 189.405 ;
        RECT 42.405 189.035 42.575 189.915 ;
        RECT 44.275 189.745 44.445 190.065 ;
        RECT 44.615 189.925 44.945 190.315 ;
        RECT 45.165 189.770 50.510 190.315 ;
        RECT 42.745 189.575 44.995 189.745 ;
        RECT 42.745 189.075 42.975 189.575 ;
        RECT 43.145 189.155 43.520 189.325 ;
        RECT 39.595 187.935 39.935 188.195 ;
        RECT 40.115 188.715 40.700 188.905 ;
        RECT 40.115 187.945 40.390 188.715 ;
        RECT 40.870 188.545 41.765 188.875 ;
        RECT 40.560 188.375 41.765 188.545 ;
        RECT 40.560 187.945 40.890 188.375 ;
        RECT 41.060 187.765 41.255 188.205 ;
        RECT 41.435 187.945 41.765 188.375 ;
        RECT 41.945 188.865 42.575 189.035 ;
        RECT 43.350 188.955 43.520 189.155 ;
        RECT 43.690 189.125 44.240 189.325 ;
        RECT 44.410 188.955 44.655 189.405 ;
        RECT 41.945 187.935 42.265 188.865 ;
        RECT 43.350 188.785 44.655 188.955 ;
        RECT 44.825 188.615 44.995 189.575 ;
        RECT 46.750 188.940 47.090 189.770 ;
        RECT 50.685 189.545 54.195 190.315 ;
        RECT 54.425 189.835 54.705 190.315 ;
        RECT 54.875 189.665 55.135 190.055 ;
        RECT 55.310 189.835 55.565 190.315 ;
        RECT 55.735 189.665 56.030 190.055 ;
        RECT 56.210 189.835 56.485 190.315 ;
        RECT 56.655 189.815 56.955 190.145 ;
        RECT 42.445 188.445 43.685 188.615 ;
        RECT 42.445 187.935 42.845 188.445 ;
        RECT 43.015 187.765 43.185 188.275 ;
        RECT 43.355 187.935 43.685 188.445 ;
        RECT 43.855 187.765 44.025 188.615 ;
        RECT 44.615 187.935 44.995 188.615 ;
        RECT 48.570 188.200 48.920 189.450 ;
        RECT 50.685 189.025 52.335 189.545 ;
        RECT 54.380 189.495 56.030 189.665 ;
        RECT 52.505 188.855 54.195 189.375 ;
        RECT 45.165 187.765 50.510 188.200 ;
        RECT 50.685 187.765 54.195 188.855 ;
        RECT 54.380 188.985 54.785 189.495 ;
        RECT 54.955 189.155 56.095 189.325 ;
        RECT 54.380 188.815 55.135 188.985 ;
        RECT 54.420 187.765 54.705 188.635 ;
        RECT 54.875 188.565 55.135 188.815 ;
        RECT 55.925 188.905 56.095 189.155 ;
        RECT 56.265 189.075 56.615 189.645 ;
        RECT 56.785 188.905 56.955 189.815 ;
        RECT 57.125 189.590 57.415 190.315 ;
        RECT 57.670 189.815 58.165 190.145 ;
        RECT 55.925 188.735 56.955 188.905 ;
        RECT 54.875 188.395 55.995 188.565 ;
        RECT 54.875 187.935 55.135 188.395 ;
        RECT 55.310 187.765 55.565 188.225 ;
        RECT 55.735 187.935 55.995 188.395 ;
        RECT 56.165 187.765 56.475 188.565 ;
        RECT 56.645 187.935 56.955 188.735 ;
        RECT 57.125 187.765 57.415 188.930 ;
        RECT 57.585 188.325 57.825 189.635 ;
        RECT 57.995 188.905 58.165 189.815 ;
        RECT 58.385 189.075 58.735 190.040 ;
        RECT 58.915 189.075 59.215 190.045 ;
        RECT 59.395 189.075 59.675 190.045 ;
        RECT 59.855 189.515 60.125 190.315 ;
        RECT 60.295 189.595 60.635 190.105 ;
        RECT 60.830 189.925 61.160 190.315 ;
        RECT 61.330 189.755 61.555 190.135 ;
        RECT 59.870 189.075 60.200 189.325 ;
        RECT 59.870 188.905 60.185 189.075 ;
        RECT 57.995 188.735 60.185 188.905 ;
        RECT 57.590 187.765 57.925 188.145 ;
        RECT 58.095 187.935 58.345 188.735 ;
        RECT 58.565 187.765 58.895 188.485 ;
        RECT 59.080 187.935 59.330 188.735 ;
        RECT 59.795 187.765 60.125 188.565 ;
        RECT 60.375 188.195 60.635 189.595 ;
        RECT 60.815 189.075 61.055 189.725 ;
        RECT 61.225 189.575 61.555 189.755 ;
        RECT 61.225 188.905 61.400 189.575 ;
        RECT 61.755 189.405 61.985 190.025 ;
        RECT 62.165 189.585 62.465 190.315 ;
        RECT 62.730 189.815 63.225 190.145 ;
        RECT 61.570 189.075 61.985 189.405 ;
        RECT 62.165 189.075 62.460 189.405 ;
        RECT 60.295 187.935 60.635 188.195 ;
        RECT 60.815 188.715 61.400 188.905 ;
        RECT 60.815 187.945 61.090 188.715 ;
        RECT 61.570 188.545 62.465 188.875 ;
        RECT 61.260 188.375 62.465 188.545 ;
        RECT 61.260 187.945 61.590 188.375 ;
        RECT 61.760 187.765 61.955 188.205 ;
        RECT 62.135 187.945 62.465 188.375 ;
        RECT 62.645 188.325 62.885 189.635 ;
        RECT 63.055 188.905 63.225 189.815 ;
        RECT 63.445 189.075 63.795 190.040 ;
        RECT 63.975 189.075 64.275 190.045 ;
        RECT 64.455 189.075 64.735 190.045 ;
        RECT 64.915 189.515 65.185 190.315 ;
        RECT 65.355 189.595 65.695 190.105 ;
        RECT 66.030 189.805 66.270 190.315 ;
        RECT 66.450 189.805 66.730 190.135 ;
        RECT 66.960 189.805 67.175 190.315 ;
        RECT 64.930 189.075 65.260 189.325 ;
        RECT 64.930 188.905 65.245 189.075 ;
        RECT 63.055 188.735 65.245 188.905 ;
        RECT 62.650 187.765 62.985 188.145 ;
        RECT 63.155 187.935 63.405 188.735 ;
        RECT 63.625 187.765 63.955 188.485 ;
        RECT 64.140 187.935 64.390 188.735 ;
        RECT 64.855 187.765 65.185 188.565 ;
        RECT 65.435 188.195 65.695 189.595 ;
        RECT 65.925 189.075 66.280 189.635 ;
        RECT 66.450 188.905 66.620 189.805 ;
        RECT 66.790 189.075 67.055 189.635 ;
        RECT 67.345 189.575 67.960 190.145 ;
        RECT 68.165 189.770 73.510 190.315 ;
        RECT 73.685 189.770 79.030 190.315 ;
        RECT 67.305 188.905 67.475 189.405 ;
        RECT 66.050 188.735 67.475 188.905 ;
        RECT 66.050 188.560 66.440 188.735 ;
        RECT 65.355 187.935 65.695 188.195 ;
        RECT 66.925 187.765 67.255 188.565 ;
        RECT 67.645 188.555 67.960 189.575 ;
        RECT 69.750 188.940 70.090 189.770 ;
        RECT 67.425 187.935 67.960 188.555 ;
        RECT 71.570 188.200 71.920 189.450 ;
        RECT 75.270 188.940 75.610 189.770 ;
        RECT 79.205 189.545 82.715 190.315 ;
        RECT 82.885 189.565 84.095 190.315 ;
        RECT 77.090 188.200 77.440 189.450 ;
        RECT 79.205 189.025 80.855 189.545 ;
        RECT 81.025 188.855 82.715 189.375 ;
        RECT 68.165 187.765 73.510 188.200 ;
        RECT 73.685 187.765 79.030 188.200 ;
        RECT 79.205 187.765 82.715 188.855 ;
        RECT 82.885 188.855 83.405 189.395 ;
        RECT 83.575 189.025 84.095 189.565 ;
        RECT 82.885 187.765 84.095 188.855 ;
        RECT 5.520 187.595 84.180 187.765 ;
        RECT 5.605 186.505 6.815 187.595 ;
        RECT 6.985 187.160 12.330 187.595 ;
        RECT 12.505 187.160 17.850 187.595 ;
        RECT 5.605 185.795 6.125 186.335 ;
        RECT 6.295 185.965 6.815 186.505 ;
        RECT 5.605 185.045 6.815 185.795 ;
        RECT 8.570 185.590 8.910 186.420 ;
        RECT 10.390 185.910 10.740 187.160 ;
        RECT 14.090 185.590 14.430 186.420 ;
        RECT 15.910 185.910 16.260 187.160 ;
        RECT 18.485 186.430 18.775 187.595 ;
        RECT 18.945 187.160 24.290 187.595 ;
        RECT 24.465 187.160 29.810 187.595 ;
        RECT 6.985 185.045 12.330 185.590 ;
        RECT 12.505 185.045 17.850 185.590 ;
        RECT 18.485 185.045 18.775 185.770 ;
        RECT 20.530 185.590 20.870 186.420 ;
        RECT 22.350 185.910 22.700 187.160 ;
        RECT 26.050 185.590 26.390 186.420 ;
        RECT 27.870 185.910 28.220 187.160 ;
        RECT 29.985 186.505 33.495 187.595 ;
        RECT 29.985 185.815 31.635 186.335 ;
        RECT 31.805 185.985 33.495 186.505 ;
        RECT 33.665 186.725 33.940 187.425 ;
        RECT 34.110 187.050 34.365 187.595 ;
        RECT 34.535 187.085 35.015 187.425 ;
        RECT 35.190 187.040 35.795 187.595 ;
        RECT 35.965 187.160 41.310 187.595 ;
        RECT 35.180 186.940 35.795 187.040 ;
        RECT 35.180 186.915 35.365 186.940 ;
        RECT 18.945 185.045 24.290 185.590 ;
        RECT 24.465 185.045 29.810 185.590 ;
        RECT 29.985 185.045 33.495 185.815 ;
        RECT 33.665 185.695 33.835 186.725 ;
        RECT 34.110 186.595 34.865 186.845 ;
        RECT 35.035 186.670 35.365 186.915 ;
        RECT 34.110 186.560 34.880 186.595 ;
        RECT 34.110 186.550 34.895 186.560 ;
        RECT 34.005 186.535 34.900 186.550 ;
        RECT 34.005 186.520 34.920 186.535 ;
        RECT 34.005 186.510 34.940 186.520 ;
        RECT 34.005 186.500 34.965 186.510 ;
        RECT 34.005 186.470 35.035 186.500 ;
        RECT 34.005 186.440 35.055 186.470 ;
        RECT 34.005 186.410 35.075 186.440 ;
        RECT 34.005 186.385 35.105 186.410 ;
        RECT 34.005 186.350 35.140 186.385 ;
        RECT 34.005 186.345 35.170 186.350 ;
        RECT 34.005 185.950 34.235 186.345 ;
        RECT 34.780 186.340 35.170 186.345 ;
        RECT 34.805 186.330 35.170 186.340 ;
        RECT 34.820 186.325 35.170 186.330 ;
        RECT 34.835 186.320 35.170 186.325 ;
        RECT 35.535 186.320 35.795 186.770 ;
        RECT 34.835 186.315 35.795 186.320 ;
        RECT 34.845 186.305 35.795 186.315 ;
        RECT 34.855 186.300 35.795 186.305 ;
        RECT 34.865 186.290 35.795 186.300 ;
        RECT 34.870 186.280 35.795 186.290 ;
        RECT 34.875 186.275 35.795 186.280 ;
        RECT 34.885 186.260 35.795 186.275 ;
        RECT 34.890 186.245 35.795 186.260 ;
        RECT 34.900 186.220 35.795 186.245 ;
        RECT 34.405 185.750 34.735 186.175 ;
        RECT 33.665 185.215 33.925 185.695 ;
        RECT 34.095 185.045 34.345 185.585 ;
        RECT 34.515 185.265 34.735 185.750 ;
        RECT 34.905 186.150 35.795 186.220 ;
        RECT 34.905 185.425 35.075 186.150 ;
        RECT 35.245 185.595 35.795 185.980 ;
        RECT 37.550 185.590 37.890 186.420 ;
        RECT 39.370 185.910 39.720 187.160 ;
        RECT 41.485 186.505 44.075 187.595 ;
        RECT 41.485 185.815 42.695 186.335 ;
        RECT 42.865 185.985 44.075 186.505 ;
        RECT 44.245 186.430 44.535 187.595 ;
        RECT 44.705 186.505 48.215 187.595 ;
        RECT 44.705 185.815 46.355 186.335 ;
        RECT 46.525 185.985 48.215 186.505 ;
        RECT 49.315 186.985 49.645 187.415 ;
        RECT 49.825 187.155 50.020 187.595 ;
        RECT 50.190 186.985 50.520 187.415 ;
        RECT 49.315 186.815 50.520 186.985 ;
        RECT 49.315 186.485 50.210 186.815 ;
        RECT 50.690 186.645 50.965 187.415 ;
        RECT 50.380 186.455 50.965 186.645 ;
        RECT 49.320 185.955 49.615 186.285 ;
        RECT 49.795 185.955 50.210 186.285 ;
        RECT 34.905 185.255 35.795 185.425 ;
        RECT 35.965 185.045 41.310 185.590 ;
        RECT 41.485 185.045 44.075 185.815 ;
        RECT 44.245 185.045 44.535 185.770 ;
        RECT 44.705 185.045 48.215 185.815 ;
        RECT 49.315 185.045 49.615 185.775 ;
        RECT 49.795 185.335 50.025 185.955 ;
        RECT 50.380 185.785 50.555 186.455 ;
        RECT 50.225 185.605 50.555 185.785 ;
        RECT 50.725 185.635 50.965 186.285 ;
        RECT 50.225 185.225 50.450 185.605 ;
        RECT 50.620 185.045 50.950 185.435 ;
        RECT 51.145 185.325 51.425 187.425 ;
        RECT 51.615 186.835 52.400 187.595 ;
        RECT 52.795 186.765 53.180 187.425 ;
        RECT 52.795 186.665 53.205 186.765 ;
        RECT 51.595 186.455 53.205 186.665 ;
        RECT 53.505 186.575 53.705 187.365 ;
        RECT 51.595 185.855 51.870 186.455 ;
        RECT 53.375 186.405 53.705 186.575 ;
        RECT 53.875 186.415 54.195 187.595 ;
        RECT 53.375 186.285 53.555 186.405 ;
        RECT 52.040 186.035 52.395 186.285 ;
        RECT 52.590 186.235 53.055 186.285 ;
        RECT 52.585 186.065 53.055 186.235 ;
        RECT 52.590 186.035 53.055 186.065 ;
        RECT 53.225 186.035 53.555 186.285 ;
        RECT 53.730 186.035 54.195 186.235 ;
        RECT 54.365 185.990 54.645 187.425 ;
        RECT 54.815 186.820 55.525 187.595 ;
        RECT 55.695 186.650 56.025 187.425 ;
        RECT 54.875 186.435 56.025 186.650 ;
        RECT 51.595 185.675 52.845 185.855 ;
        RECT 52.480 185.605 52.845 185.675 ;
        RECT 53.015 185.655 54.195 185.825 ;
        RECT 51.655 185.045 51.825 185.505 ;
        RECT 53.015 185.435 53.345 185.655 ;
        RECT 52.095 185.255 53.345 185.435 ;
        RECT 53.515 185.045 53.685 185.485 ;
        RECT 53.855 185.240 54.195 185.655 ;
        RECT 54.365 185.215 54.705 185.990 ;
        RECT 54.875 185.865 55.160 186.435 ;
        RECT 55.345 186.035 55.815 186.265 ;
        RECT 56.220 186.235 56.435 187.350 ;
        RECT 56.615 186.875 56.945 187.595 ;
        RECT 57.585 186.725 57.860 187.425 ;
        RECT 58.030 187.050 58.285 187.595 ;
        RECT 58.455 187.085 58.935 187.425 ;
        RECT 59.110 187.040 59.715 187.595 ;
        RECT 59.100 186.940 59.715 187.040 ;
        RECT 59.100 186.915 59.285 186.940 ;
        RECT 56.725 186.235 56.955 186.575 ;
        RECT 55.985 186.055 56.435 186.235 ;
        RECT 55.985 186.035 56.315 186.055 ;
        RECT 56.625 186.035 56.955 186.235 ;
        RECT 54.875 185.675 55.585 185.865 ;
        RECT 55.285 185.535 55.585 185.675 ;
        RECT 55.775 185.675 56.955 185.865 ;
        RECT 55.775 185.595 56.105 185.675 ;
        RECT 55.285 185.525 55.600 185.535 ;
        RECT 55.285 185.515 55.610 185.525 ;
        RECT 55.285 185.510 55.620 185.515 ;
        RECT 54.875 185.045 55.045 185.505 ;
        RECT 55.285 185.500 55.625 185.510 ;
        RECT 55.285 185.495 55.630 185.500 ;
        RECT 55.285 185.485 55.635 185.495 ;
        RECT 55.285 185.480 55.640 185.485 ;
        RECT 55.285 185.215 55.645 185.480 ;
        RECT 56.275 185.045 56.445 185.505 ;
        RECT 56.615 185.215 56.955 185.675 ;
        RECT 57.585 185.695 57.755 186.725 ;
        RECT 58.030 186.595 58.785 186.845 ;
        RECT 58.955 186.670 59.285 186.915 ;
        RECT 58.030 186.560 58.800 186.595 ;
        RECT 58.030 186.550 58.815 186.560 ;
        RECT 57.925 186.535 58.820 186.550 ;
        RECT 57.925 186.520 58.840 186.535 ;
        RECT 57.925 186.510 58.860 186.520 ;
        RECT 57.925 186.500 58.885 186.510 ;
        RECT 57.925 186.470 58.955 186.500 ;
        RECT 57.925 186.440 58.975 186.470 ;
        RECT 57.925 186.410 58.995 186.440 ;
        RECT 57.925 186.385 59.025 186.410 ;
        RECT 57.925 186.350 59.060 186.385 ;
        RECT 57.925 186.345 59.090 186.350 ;
        RECT 57.925 185.950 58.155 186.345 ;
        RECT 58.700 186.340 59.090 186.345 ;
        RECT 58.725 186.330 59.090 186.340 ;
        RECT 58.740 186.325 59.090 186.330 ;
        RECT 58.755 186.320 59.090 186.325 ;
        RECT 59.455 186.320 59.715 186.770 ;
        RECT 59.885 186.505 62.475 187.595 ;
        RECT 58.755 186.315 59.715 186.320 ;
        RECT 58.765 186.305 59.715 186.315 ;
        RECT 58.775 186.300 59.715 186.305 ;
        RECT 58.785 186.290 59.715 186.300 ;
        RECT 58.790 186.280 59.715 186.290 ;
        RECT 58.795 186.275 59.715 186.280 ;
        RECT 58.805 186.260 59.715 186.275 ;
        RECT 58.810 186.245 59.715 186.260 ;
        RECT 58.820 186.220 59.715 186.245 ;
        RECT 58.325 185.750 58.655 186.175 ;
        RECT 57.585 185.215 57.845 185.695 ;
        RECT 58.015 185.045 58.265 185.585 ;
        RECT 58.435 185.265 58.655 185.750 ;
        RECT 58.825 186.150 59.715 186.220 ;
        RECT 58.825 185.425 58.995 186.150 ;
        RECT 59.165 185.595 59.715 185.980 ;
        RECT 59.885 185.815 61.095 186.335 ;
        RECT 61.265 185.985 62.475 186.505 ;
        RECT 63.105 186.455 63.385 187.595 ;
        RECT 63.555 186.445 63.885 187.425 ;
        RECT 64.055 186.455 64.315 187.595 ;
        RECT 64.485 187.160 69.830 187.595 ;
        RECT 63.115 186.015 63.450 186.285 ;
        RECT 63.620 185.845 63.790 186.445 ;
        RECT 63.960 186.035 64.295 186.285 ;
        RECT 58.825 185.255 59.715 185.425 ;
        RECT 59.885 185.045 62.475 185.815 ;
        RECT 63.105 185.045 63.415 185.845 ;
        RECT 63.620 185.215 64.315 185.845 ;
        RECT 66.070 185.590 66.410 186.420 ;
        RECT 67.890 185.910 68.240 187.160 ;
        RECT 70.005 186.430 70.295 187.595 ;
        RECT 70.465 187.160 75.810 187.595 ;
        RECT 75.985 187.160 81.330 187.595 ;
        RECT 64.485 185.045 69.830 185.590 ;
        RECT 70.005 185.045 70.295 185.770 ;
        RECT 72.050 185.590 72.390 186.420 ;
        RECT 73.870 185.910 74.220 187.160 ;
        RECT 77.570 185.590 77.910 186.420 ;
        RECT 79.390 185.910 79.740 187.160 ;
        RECT 81.505 186.505 82.715 187.595 ;
        RECT 81.505 185.795 82.025 186.335 ;
        RECT 82.195 185.965 82.715 186.505 ;
        RECT 82.885 186.505 84.095 187.595 ;
        RECT 82.885 185.965 83.405 186.505 ;
        RECT 83.575 185.795 84.095 186.335 ;
        RECT 70.465 185.045 75.810 185.590 ;
        RECT 75.985 185.045 81.330 185.590 ;
        RECT 81.505 185.045 82.715 185.795 ;
        RECT 82.885 185.045 84.095 185.795 ;
        RECT 5.520 184.875 84.180 185.045 ;
        RECT 5.605 184.125 6.815 184.875 ;
        RECT 6.985 184.330 12.330 184.875 ;
        RECT 5.605 183.585 6.125 184.125 ;
        RECT 6.295 183.415 6.815 183.955 ;
        RECT 8.570 183.500 8.910 184.330 ;
        RECT 12.505 184.125 13.715 184.875 ;
        RECT 13.885 184.225 14.145 184.705 ;
        RECT 14.315 184.335 14.565 184.875 ;
        RECT 5.605 182.325 6.815 183.415 ;
        RECT 10.390 182.760 10.740 184.010 ;
        RECT 12.505 183.585 13.025 184.125 ;
        RECT 13.195 183.415 13.715 183.955 ;
        RECT 6.985 182.325 12.330 182.760 ;
        RECT 12.505 182.325 13.715 183.415 ;
        RECT 13.885 183.195 14.055 184.225 ;
        RECT 14.735 184.170 14.955 184.655 ;
        RECT 14.225 183.575 14.455 183.970 ;
        RECT 14.625 183.745 14.955 184.170 ;
        RECT 15.125 184.495 16.015 184.665 ;
        RECT 15.125 183.770 15.295 184.495 ;
        RECT 15.465 183.940 16.015 184.325 ;
        RECT 16.185 184.105 19.695 184.875 ;
        RECT 19.955 184.325 20.125 184.615 ;
        RECT 20.295 184.495 20.625 184.875 ;
        RECT 19.955 184.155 20.620 184.325 ;
        RECT 15.125 183.700 16.015 183.770 ;
        RECT 15.120 183.675 16.015 183.700 ;
        RECT 15.110 183.660 16.015 183.675 ;
        RECT 15.105 183.645 16.015 183.660 ;
        RECT 15.095 183.640 16.015 183.645 ;
        RECT 15.090 183.630 16.015 183.640 ;
        RECT 15.085 183.620 16.015 183.630 ;
        RECT 15.075 183.615 16.015 183.620 ;
        RECT 15.065 183.605 16.015 183.615 ;
        RECT 15.055 183.600 16.015 183.605 ;
        RECT 15.055 183.595 15.390 183.600 ;
        RECT 15.040 183.590 15.390 183.595 ;
        RECT 15.025 183.580 15.390 183.590 ;
        RECT 15.000 183.575 15.390 183.580 ;
        RECT 14.225 183.570 15.390 183.575 ;
        RECT 14.225 183.535 15.360 183.570 ;
        RECT 14.225 183.510 15.325 183.535 ;
        RECT 14.225 183.480 15.295 183.510 ;
        RECT 14.225 183.450 15.275 183.480 ;
        RECT 14.225 183.420 15.255 183.450 ;
        RECT 14.225 183.410 15.185 183.420 ;
        RECT 14.225 183.400 15.160 183.410 ;
        RECT 14.225 183.385 15.140 183.400 ;
        RECT 14.225 183.370 15.120 183.385 ;
        RECT 14.330 183.360 15.115 183.370 ;
        RECT 14.330 183.325 15.100 183.360 ;
        RECT 13.885 182.495 14.160 183.195 ;
        RECT 14.330 183.075 15.085 183.325 ;
        RECT 15.255 183.005 15.585 183.250 ;
        RECT 15.755 183.150 16.015 183.600 ;
        RECT 16.185 183.585 17.835 184.105 ;
        RECT 18.005 183.415 19.695 183.935 ;
        RECT 15.400 182.980 15.585 183.005 ;
        RECT 15.400 182.880 16.015 182.980 ;
        RECT 14.330 182.325 14.585 182.870 ;
        RECT 14.755 182.495 15.235 182.835 ;
        RECT 15.410 182.325 16.015 182.880 ;
        RECT 16.185 182.325 19.695 183.415 ;
        RECT 19.870 183.335 20.220 183.985 ;
        RECT 20.390 183.165 20.620 184.155 ;
        RECT 19.955 182.995 20.620 183.165 ;
        RECT 19.955 182.495 20.125 182.995 ;
        RECT 20.295 182.325 20.625 182.825 ;
        RECT 20.795 182.495 20.980 184.615 ;
        RECT 21.235 184.415 21.485 184.875 ;
        RECT 21.655 184.425 21.990 184.595 ;
        RECT 22.185 184.425 22.860 184.595 ;
        RECT 21.655 184.285 21.825 184.425 ;
        RECT 21.150 183.295 21.430 184.245 ;
        RECT 21.600 184.155 21.825 184.285 ;
        RECT 21.600 183.050 21.770 184.155 ;
        RECT 21.995 184.005 22.520 184.225 ;
        RECT 21.940 183.240 22.180 183.835 ;
        RECT 22.350 183.305 22.520 184.005 ;
        RECT 22.690 183.645 22.860 184.425 ;
        RECT 23.180 184.375 23.550 184.875 ;
        RECT 23.730 184.425 24.135 184.595 ;
        RECT 24.305 184.425 25.090 184.595 ;
        RECT 23.730 184.195 23.900 184.425 ;
        RECT 23.070 183.895 23.900 184.195 ;
        RECT 24.285 183.925 24.750 184.255 ;
        RECT 23.070 183.865 23.270 183.895 ;
        RECT 23.390 183.645 23.560 183.715 ;
        RECT 22.690 183.475 23.560 183.645 ;
        RECT 23.050 183.385 23.560 183.475 ;
        RECT 21.600 182.920 21.905 183.050 ;
        RECT 22.350 182.940 22.880 183.305 ;
        RECT 21.220 182.325 21.485 182.785 ;
        RECT 21.655 182.495 21.905 182.920 ;
        RECT 23.050 182.770 23.220 183.385 ;
        RECT 22.115 182.600 23.220 182.770 ;
        RECT 23.390 182.325 23.560 183.125 ;
        RECT 23.730 182.825 23.900 183.895 ;
        RECT 24.070 182.995 24.260 183.715 ;
        RECT 24.430 182.965 24.750 183.925 ;
        RECT 24.920 183.965 25.090 184.425 ;
        RECT 25.365 184.345 25.575 184.875 ;
        RECT 25.835 184.135 26.165 184.660 ;
        RECT 26.335 184.265 26.505 184.875 ;
        RECT 26.675 184.220 27.005 184.655 ;
        RECT 26.675 184.135 27.055 184.220 ;
        RECT 25.965 183.965 26.165 184.135 ;
        RECT 26.830 184.095 27.055 184.135 ;
        RECT 24.920 183.635 25.795 183.965 ;
        RECT 25.965 183.635 26.715 183.965 ;
        RECT 23.730 182.495 23.980 182.825 ;
        RECT 24.920 182.795 25.090 183.635 ;
        RECT 25.965 183.430 26.155 183.635 ;
        RECT 26.885 183.515 27.055 184.095 ;
        RECT 27.225 184.105 30.735 184.875 ;
        RECT 31.365 184.150 31.655 184.875 ;
        RECT 31.915 184.325 32.085 184.615 ;
        RECT 32.255 184.495 32.585 184.875 ;
        RECT 31.915 184.155 32.580 184.325 ;
        RECT 27.225 183.585 28.875 184.105 ;
        RECT 26.840 183.465 27.055 183.515 ;
        RECT 25.260 183.055 26.155 183.430 ;
        RECT 26.665 183.385 27.055 183.465 ;
        RECT 29.045 183.415 30.735 183.935 ;
        RECT 24.205 182.625 25.090 182.795 ;
        RECT 25.270 182.325 25.585 182.825 ;
        RECT 25.815 182.495 26.155 183.055 ;
        RECT 26.325 182.325 26.495 183.335 ;
        RECT 26.665 182.540 26.995 183.385 ;
        RECT 27.225 182.325 30.735 183.415 ;
        RECT 31.365 182.325 31.655 183.490 ;
        RECT 31.830 183.335 32.180 183.985 ;
        RECT 32.350 183.165 32.580 184.155 ;
        RECT 31.915 182.995 32.580 183.165 ;
        RECT 31.915 182.495 32.085 182.995 ;
        RECT 32.255 182.325 32.585 182.825 ;
        RECT 32.755 182.495 32.940 184.615 ;
        RECT 33.195 184.415 33.445 184.875 ;
        RECT 33.615 184.425 33.950 184.595 ;
        RECT 34.145 184.425 34.820 184.595 ;
        RECT 33.615 184.285 33.785 184.425 ;
        RECT 33.110 183.295 33.390 184.245 ;
        RECT 33.560 184.155 33.785 184.285 ;
        RECT 33.560 183.050 33.730 184.155 ;
        RECT 33.955 184.005 34.480 184.225 ;
        RECT 33.900 183.240 34.140 183.835 ;
        RECT 34.310 183.305 34.480 184.005 ;
        RECT 34.650 183.645 34.820 184.425 ;
        RECT 35.140 184.375 35.510 184.875 ;
        RECT 35.690 184.425 36.095 184.595 ;
        RECT 36.265 184.425 37.050 184.595 ;
        RECT 35.690 184.195 35.860 184.425 ;
        RECT 35.030 183.895 35.860 184.195 ;
        RECT 36.245 183.925 36.710 184.255 ;
        RECT 35.030 183.865 35.230 183.895 ;
        RECT 35.350 183.645 35.520 183.715 ;
        RECT 34.650 183.475 35.520 183.645 ;
        RECT 35.010 183.385 35.520 183.475 ;
        RECT 33.560 182.920 33.865 183.050 ;
        RECT 34.310 182.940 34.840 183.305 ;
        RECT 33.180 182.325 33.445 182.785 ;
        RECT 33.615 182.495 33.865 182.920 ;
        RECT 35.010 182.770 35.180 183.385 ;
        RECT 34.075 182.600 35.180 182.770 ;
        RECT 35.350 182.325 35.520 183.125 ;
        RECT 35.690 182.825 35.860 183.895 ;
        RECT 36.030 182.995 36.220 183.715 ;
        RECT 36.390 182.965 36.710 183.925 ;
        RECT 36.880 183.965 37.050 184.425 ;
        RECT 37.325 184.345 37.535 184.875 ;
        RECT 37.795 184.135 38.125 184.660 ;
        RECT 38.295 184.265 38.465 184.875 ;
        RECT 38.635 184.220 38.965 184.655 ;
        RECT 39.185 184.330 44.530 184.875 ;
        RECT 38.635 184.135 39.015 184.220 ;
        RECT 37.925 183.965 38.125 184.135 ;
        RECT 38.790 184.095 39.015 184.135 ;
        RECT 36.880 183.635 37.755 183.965 ;
        RECT 37.925 183.635 38.675 183.965 ;
        RECT 35.690 182.495 35.940 182.825 ;
        RECT 36.880 182.795 37.050 183.635 ;
        RECT 37.925 183.430 38.115 183.635 ;
        RECT 38.845 183.515 39.015 184.095 ;
        RECT 38.800 183.465 39.015 183.515 ;
        RECT 40.770 183.500 41.110 184.330 ;
        RECT 44.705 184.105 48.215 184.875 ;
        RECT 48.855 184.145 49.155 184.875 ;
        RECT 37.220 183.055 38.115 183.430 ;
        RECT 38.625 183.385 39.015 183.465 ;
        RECT 36.165 182.625 37.050 182.795 ;
        RECT 37.230 182.325 37.545 182.825 ;
        RECT 37.775 182.495 38.115 183.055 ;
        RECT 38.285 182.325 38.455 183.335 ;
        RECT 38.625 182.540 38.955 183.385 ;
        RECT 42.590 182.760 42.940 184.010 ;
        RECT 44.705 183.585 46.355 184.105 ;
        RECT 49.335 183.965 49.565 184.585 ;
        RECT 49.765 184.315 49.990 184.695 ;
        RECT 50.160 184.485 50.490 184.875 ;
        RECT 49.765 184.135 50.095 184.315 ;
        RECT 46.525 183.415 48.215 183.935 ;
        RECT 48.860 183.635 49.155 183.965 ;
        RECT 49.335 183.635 49.750 183.965 ;
        RECT 49.920 183.465 50.095 184.135 ;
        RECT 50.265 183.635 50.505 184.285 ;
        RECT 50.685 184.105 52.355 184.875 ;
        RECT 52.990 184.345 53.280 184.695 ;
        RECT 53.475 184.515 53.805 184.875 ;
        RECT 53.975 184.345 54.205 184.650 ;
        RECT 52.990 184.175 54.205 184.345 ;
        RECT 50.685 183.585 51.435 184.105 ;
        RECT 54.395 184.005 54.565 184.570 ;
        RECT 39.185 182.325 44.530 182.760 ;
        RECT 44.705 182.325 48.215 183.415 ;
        RECT 48.855 183.105 49.750 183.435 ;
        RECT 49.920 183.275 50.505 183.465 ;
        RECT 51.605 183.415 52.355 183.935 ;
        RECT 53.050 183.855 53.310 183.965 ;
        RECT 53.045 183.685 53.310 183.855 ;
        RECT 53.050 183.635 53.310 183.685 ;
        RECT 53.490 183.635 53.875 183.965 ;
        RECT 54.045 183.835 54.565 184.005 ;
        RECT 54.825 184.105 56.495 184.875 ;
        RECT 57.125 184.150 57.415 184.875 ;
        RECT 57.585 184.330 62.930 184.875 ;
        RECT 63.105 184.330 68.450 184.875 ;
        RECT 68.625 184.330 73.970 184.875 ;
        RECT 74.145 184.330 79.490 184.875 ;
        RECT 48.855 182.935 50.060 183.105 ;
        RECT 48.855 182.505 49.185 182.935 ;
        RECT 49.365 182.325 49.560 182.765 ;
        RECT 49.730 182.505 50.060 182.935 ;
        RECT 50.230 182.505 50.505 183.275 ;
        RECT 50.685 182.325 52.355 183.415 ;
        RECT 52.990 182.325 53.310 183.465 ;
        RECT 53.490 182.585 53.685 183.635 ;
        RECT 54.045 183.455 54.215 183.835 ;
        RECT 53.865 183.175 54.215 183.455 ;
        RECT 54.405 183.305 54.650 183.665 ;
        RECT 54.825 183.585 55.575 184.105 ;
        RECT 55.745 183.415 56.495 183.935 ;
        RECT 59.170 183.500 59.510 184.330 ;
        RECT 53.865 182.495 54.195 183.175 ;
        RECT 54.395 182.325 54.650 183.125 ;
        RECT 54.825 182.325 56.495 183.415 ;
        RECT 57.125 182.325 57.415 183.490 ;
        RECT 60.990 182.760 61.340 184.010 ;
        RECT 64.690 183.500 65.030 184.330 ;
        RECT 66.510 182.760 66.860 184.010 ;
        RECT 70.210 183.500 70.550 184.330 ;
        RECT 72.030 182.760 72.380 184.010 ;
        RECT 75.730 183.500 76.070 184.330 ;
        RECT 79.665 184.105 82.255 184.875 ;
        RECT 82.885 184.125 84.095 184.875 ;
        RECT 77.550 182.760 77.900 184.010 ;
        RECT 79.665 183.585 80.875 184.105 ;
        RECT 81.045 183.415 82.255 183.935 ;
        RECT 57.585 182.325 62.930 182.760 ;
        RECT 63.105 182.325 68.450 182.760 ;
        RECT 68.625 182.325 73.970 182.760 ;
        RECT 74.145 182.325 79.490 182.760 ;
        RECT 79.665 182.325 82.255 183.415 ;
        RECT 82.885 183.415 83.405 183.955 ;
        RECT 83.575 183.585 84.095 184.125 ;
        RECT 82.885 182.325 84.095 183.415 ;
        RECT 5.520 182.155 84.180 182.325 ;
        RECT 5.605 181.065 6.815 182.155 ;
        RECT 6.985 181.065 9.575 182.155 ;
        RECT 5.605 180.355 6.125 180.895 ;
        RECT 6.295 180.525 6.815 181.065 ;
        RECT 6.985 180.375 8.195 180.895 ;
        RECT 8.365 180.545 9.575 181.065 ;
        RECT 9.745 181.015 10.025 182.155 ;
        RECT 10.195 181.005 10.525 181.985 ;
        RECT 10.695 181.015 10.955 182.155 ;
        RECT 11.185 181.095 11.515 181.940 ;
        RECT 11.685 181.145 11.855 182.155 ;
        RECT 12.025 181.425 12.365 181.985 ;
        RECT 12.595 181.655 12.910 182.155 ;
        RECT 13.090 181.685 13.975 181.855 ;
        RECT 11.125 181.015 11.515 181.095 ;
        RECT 12.025 181.050 12.920 181.425 ;
        RECT 9.755 180.575 10.090 180.845 ;
        RECT 10.260 180.405 10.430 181.005 ;
        RECT 11.125 180.965 11.340 181.015 ;
        RECT 10.600 180.595 10.935 180.845 ;
        RECT 5.605 179.605 6.815 180.355 ;
        RECT 6.985 179.605 9.575 180.375 ;
        RECT 9.745 179.605 10.055 180.405 ;
        RECT 10.260 179.775 10.955 180.405 ;
        RECT 11.125 180.385 11.295 180.965 ;
        RECT 12.025 180.845 12.215 181.050 ;
        RECT 13.090 180.845 13.260 181.685 ;
        RECT 14.200 181.655 14.450 181.985 ;
        RECT 11.465 180.515 12.215 180.845 ;
        RECT 12.385 180.515 13.260 180.845 ;
        RECT 11.125 180.345 11.350 180.385 ;
        RECT 12.015 180.345 12.215 180.515 ;
        RECT 11.125 180.260 11.505 180.345 ;
        RECT 11.175 179.825 11.505 180.260 ;
        RECT 11.675 179.605 11.845 180.215 ;
        RECT 12.015 179.820 12.345 180.345 ;
        RECT 12.605 179.605 12.815 180.135 ;
        RECT 13.090 180.055 13.260 180.515 ;
        RECT 13.430 180.555 13.750 181.515 ;
        RECT 13.920 180.765 14.110 181.485 ;
        RECT 14.280 180.585 14.450 181.655 ;
        RECT 14.620 181.355 14.790 182.155 ;
        RECT 14.960 181.710 16.065 181.880 ;
        RECT 14.960 181.095 15.130 181.710 ;
        RECT 16.275 181.560 16.525 181.985 ;
        RECT 16.695 181.695 16.960 182.155 ;
        RECT 15.300 181.175 15.830 181.540 ;
        RECT 16.275 181.430 16.580 181.560 ;
        RECT 14.620 181.005 15.130 181.095 ;
        RECT 14.620 180.835 15.490 181.005 ;
        RECT 14.620 180.765 14.790 180.835 ;
        RECT 14.910 180.585 15.110 180.615 ;
        RECT 13.430 180.225 13.895 180.555 ;
        RECT 14.280 180.285 15.110 180.585 ;
        RECT 14.280 180.055 14.450 180.285 ;
        RECT 13.090 179.885 13.875 180.055 ;
        RECT 14.045 179.885 14.450 180.055 ;
        RECT 14.630 179.605 15.000 180.105 ;
        RECT 15.320 180.055 15.490 180.835 ;
        RECT 15.660 180.475 15.830 181.175 ;
        RECT 16.000 180.645 16.240 181.240 ;
        RECT 15.660 180.255 16.185 180.475 ;
        RECT 16.410 180.325 16.580 181.430 ;
        RECT 16.355 180.195 16.580 180.325 ;
        RECT 16.750 180.235 17.030 181.185 ;
        RECT 16.355 180.055 16.525 180.195 ;
        RECT 15.320 179.885 15.995 180.055 ;
        RECT 16.190 179.885 16.525 180.055 ;
        RECT 16.695 179.605 16.945 180.065 ;
        RECT 17.200 179.865 17.385 181.985 ;
        RECT 17.555 181.655 17.885 182.155 ;
        RECT 18.055 181.485 18.225 181.985 ;
        RECT 17.560 181.315 18.225 181.485 ;
        RECT 17.560 180.325 17.790 181.315 ;
        RECT 17.960 180.495 18.310 181.145 ;
        RECT 18.485 180.990 18.775 182.155 ;
        RECT 19.865 181.285 20.140 181.985 ;
        RECT 20.310 181.610 20.565 182.155 ;
        RECT 20.735 181.645 21.215 181.985 ;
        RECT 21.390 181.600 21.995 182.155 ;
        RECT 21.380 181.500 21.995 181.600 ;
        RECT 21.380 181.475 21.565 181.500 ;
        RECT 17.560 180.155 18.225 180.325 ;
        RECT 17.555 179.605 17.885 179.985 ;
        RECT 18.055 179.865 18.225 180.155 ;
        RECT 18.485 179.605 18.775 180.330 ;
        RECT 19.865 180.255 20.035 181.285 ;
        RECT 20.310 181.155 21.065 181.405 ;
        RECT 21.235 181.230 21.565 181.475 ;
        RECT 20.310 181.120 21.080 181.155 ;
        RECT 20.310 181.110 21.095 181.120 ;
        RECT 20.205 181.095 21.100 181.110 ;
        RECT 20.205 181.080 21.120 181.095 ;
        RECT 20.205 181.070 21.140 181.080 ;
        RECT 20.205 181.060 21.165 181.070 ;
        RECT 20.205 181.030 21.235 181.060 ;
        RECT 20.205 181.000 21.255 181.030 ;
        RECT 20.205 180.970 21.275 181.000 ;
        RECT 20.205 180.945 21.305 180.970 ;
        RECT 20.205 180.910 21.340 180.945 ;
        RECT 20.205 180.905 21.370 180.910 ;
        RECT 20.205 180.510 20.435 180.905 ;
        RECT 20.980 180.900 21.370 180.905 ;
        RECT 21.005 180.890 21.370 180.900 ;
        RECT 21.020 180.885 21.370 180.890 ;
        RECT 21.035 180.880 21.370 180.885 ;
        RECT 21.735 180.880 21.995 181.330 ;
        RECT 21.035 180.875 21.995 180.880 ;
        RECT 21.045 180.865 21.995 180.875 ;
        RECT 21.055 180.860 21.995 180.865 ;
        RECT 21.065 180.850 21.995 180.860 ;
        RECT 21.070 180.840 21.995 180.850 ;
        RECT 21.075 180.835 21.995 180.840 ;
        RECT 21.085 180.820 21.995 180.835 ;
        RECT 21.090 180.805 21.995 180.820 ;
        RECT 21.100 180.780 21.995 180.805 ;
        RECT 20.605 180.310 20.935 180.735 ;
        RECT 19.865 179.775 20.125 180.255 ;
        RECT 20.295 179.605 20.545 180.145 ;
        RECT 20.715 179.825 20.935 180.310 ;
        RECT 21.105 180.710 21.995 180.780 ;
        RECT 22.175 181.095 22.505 181.945 ;
        RECT 21.105 179.985 21.275 180.710 ;
        RECT 21.445 180.155 21.995 180.540 ;
        RECT 22.175 180.330 22.365 181.095 ;
        RECT 22.675 181.015 22.925 182.155 ;
        RECT 23.115 181.515 23.365 181.935 ;
        RECT 23.595 181.685 23.925 182.155 ;
        RECT 24.155 181.515 24.405 181.935 ;
        RECT 23.115 181.345 24.405 181.515 ;
        RECT 24.585 181.515 24.915 181.945 ;
        RECT 24.585 181.345 25.040 181.515 ;
        RECT 23.105 180.845 23.320 181.175 ;
        RECT 22.535 180.515 22.845 180.845 ;
        RECT 23.015 180.515 23.320 180.845 ;
        RECT 23.495 180.515 23.780 181.175 ;
        RECT 23.975 180.515 24.240 181.175 ;
        RECT 24.455 180.515 24.700 181.175 ;
        RECT 22.675 180.345 22.845 180.515 ;
        RECT 24.870 180.345 25.040 181.345 ;
        RECT 21.105 179.815 21.995 179.985 ;
        RECT 22.175 179.820 22.505 180.330 ;
        RECT 22.675 180.175 25.040 180.345 ;
        RECT 22.675 179.605 23.005 180.005 ;
        RECT 24.055 179.835 24.385 180.175 ;
        RECT 24.555 179.605 24.885 180.005 ;
        RECT 25.395 179.785 25.655 181.975 ;
        RECT 25.825 181.425 26.165 182.155 ;
        RECT 26.345 181.245 26.615 181.975 ;
        RECT 25.845 181.025 26.615 181.245 ;
        RECT 26.795 181.265 27.025 181.975 ;
        RECT 27.195 181.445 27.525 182.155 ;
        RECT 27.695 181.265 27.955 181.975 ;
        RECT 26.795 181.025 27.955 181.265 ;
        RECT 28.145 181.435 28.605 181.985 ;
        RECT 28.795 181.435 29.125 182.155 ;
        RECT 25.845 180.355 26.135 181.025 ;
        RECT 26.315 180.535 26.780 180.845 ;
        RECT 26.960 180.535 27.485 180.845 ;
        RECT 25.845 180.155 27.075 180.355 ;
        RECT 25.915 179.605 26.585 179.975 ;
        RECT 26.765 179.785 27.075 180.155 ;
        RECT 27.255 179.895 27.485 180.535 ;
        RECT 27.665 180.515 27.965 180.845 ;
        RECT 27.665 179.605 27.955 180.335 ;
        RECT 28.145 180.065 28.395 181.435 ;
        RECT 29.325 181.265 29.625 181.815 ;
        RECT 29.795 181.485 30.075 182.155 ;
        RECT 28.685 181.095 29.625 181.265 ;
        RECT 28.685 180.845 28.855 181.095 ;
        RECT 29.995 180.845 30.260 181.205 ;
        RECT 30.455 181.185 30.785 181.985 ;
        RECT 30.955 181.355 31.185 182.155 ;
        RECT 31.355 181.185 31.685 181.985 ;
        RECT 30.455 181.015 31.685 181.185 ;
        RECT 31.855 181.015 32.110 182.155 ;
        RECT 32.285 181.305 32.665 181.985 ;
        RECT 33.255 181.305 33.425 182.155 ;
        RECT 33.595 181.475 33.925 181.985 ;
        RECT 34.095 181.645 34.265 182.155 ;
        RECT 34.435 181.475 34.835 181.985 ;
        RECT 33.595 181.305 34.835 181.475 ;
        RECT 28.565 180.515 28.855 180.845 ;
        RECT 29.025 180.595 29.365 180.845 ;
        RECT 29.585 180.595 30.260 180.845 ;
        RECT 30.445 180.515 30.755 180.845 ;
        RECT 28.685 180.425 28.855 180.515 ;
        RECT 28.685 180.235 30.075 180.425 ;
        RECT 28.145 179.775 28.705 180.065 ;
        RECT 28.875 179.605 29.125 180.065 ;
        RECT 29.745 179.875 30.075 180.235 ;
        RECT 30.455 180.115 30.785 180.345 ;
        RECT 30.960 180.285 31.335 180.845 ;
        RECT 31.505 180.115 31.685 181.015 ;
        RECT 31.870 180.265 32.090 180.845 ;
        RECT 32.285 180.345 32.455 181.305 ;
        RECT 32.625 180.965 33.930 181.135 ;
        RECT 35.015 181.055 35.335 181.985 ;
        RECT 35.505 181.065 39.015 182.155 ;
        RECT 39.190 181.730 39.525 182.155 ;
        RECT 39.695 181.550 39.880 181.955 ;
        RECT 32.625 180.515 32.870 180.965 ;
        RECT 33.040 180.595 33.590 180.795 ;
        RECT 33.760 180.765 33.930 180.965 ;
        RECT 34.705 180.885 35.335 181.055 ;
        RECT 33.760 180.595 34.135 180.765 ;
        RECT 34.305 180.345 34.535 180.845 ;
        RECT 32.285 180.175 34.535 180.345 ;
        RECT 30.455 179.775 31.685 180.115 ;
        RECT 31.855 179.605 32.110 180.095 ;
        RECT 32.335 179.605 32.665 179.995 ;
        RECT 32.835 179.855 33.005 180.175 ;
        RECT 34.705 180.005 34.875 180.885 ;
        RECT 33.175 179.605 33.505 179.995 ;
        RECT 33.920 179.835 34.875 180.005 ;
        RECT 35.045 179.605 35.335 180.440 ;
        RECT 35.505 180.375 37.155 180.895 ;
        RECT 37.325 180.545 39.015 181.065 ;
        RECT 39.215 181.375 39.880 181.550 ;
        RECT 40.085 181.375 40.415 182.155 ;
        RECT 35.505 179.605 39.015 180.375 ;
        RECT 39.215 180.345 39.555 181.375 ;
        RECT 40.585 181.185 40.855 181.955 ;
        RECT 39.725 181.015 40.855 181.185 ;
        RECT 41.025 181.065 43.615 182.155 ;
        RECT 39.725 180.515 39.975 181.015 ;
        RECT 39.215 180.175 39.900 180.345 ;
        RECT 40.155 180.265 40.515 180.845 ;
        RECT 39.190 179.605 39.525 180.005 ;
        RECT 39.695 179.775 39.900 180.175 ;
        RECT 40.685 180.105 40.855 181.015 ;
        RECT 40.110 179.605 40.385 180.085 ;
        RECT 40.595 179.775 40.855 180.105 ;
        RECT 41.025 180.375 42.235 180.895 ;
        RECT 42.405 180.545 43.615 181.065 ;
        RECT 44.245 180.990 44.535 182.155 ;
        RECT 41.025 179.605 43.615 180.375 ;
        RECT 44.245 179.605 44.535 180.330 ;
        RECT 44.715 179.785 44.975 181.975 ;
        RECT 45.145 181.425 45.485 182.155 ;
        RECT 45.665 181.245 45.935 181.975 ;
        RECT 45.165 181.025 45.935 181.245 ;
        RECT 46.115 181.265 46.345 181.975 ;
        RECT 46.515 181.445 46.845 182.155 ;
        RECT 47.015 181.265 47.275 181.975 ;
        RECT 46.115 181.025 47.275 181.265 ;
        RECT 47.465 181.065 50.975 182.155 ;
        RECT 45.165 180.355 45.455 181.025 ;
        RECT 45.635 180.535 46.100 180.845 ;
        RECT 46.280 180.535 46.805 180.845 ;
        RECT 45.165 180.155 46.395 180.355 ;
        RECT 45.235 179.605 45.905 179.975 ;
        RECT 46.085 179.785 46.395 180.155 ;
        RECT 46.575 179.895 46.805 180.535 ;
        RECT 46.985 180.515 47.285 180.845 ;
        RECT 47.465 180.375 49.115 180.895 ;
        RECT 49.285 180.545 50.975 181.065 ;
        RECT 51.605 181.185 51.895 181.985 ;
        RECT 52.065 181.355 52.300 182.155 ;
        RECT 52.485 181.815 54.020 181.985 ;
        RECT 52.485 181.185 52.815 181.815 ;
        RECT 51.605 181.015 52.815 181.185 ;
        RECT 51.605 180.515 51.850 180.845 ;
        RECT 46.985 179.605 47.275 180.335 ;
        RECT 47.465 179.605 50.975 180.375 ;
        RECT 52.020 180.345 52.190 181.015 ;
        RECT 52.985 180.845 53.220 181.590 ;
        RECT 52.360 180.515 52.760 180.845 ;
        RECT 52.930 180.515 53.220 180.845 ;
        RECT 53.410 180.845 53.680 181.590 ;
        RECT 53.850 181.185 54.020 181.815 ;
        RECT 54.190 181.355 54.595 182.155 ;
        RECT 53.850 181.015 54.595 181.185 ;
        RECT 53.410 180.515 53.750 180.845 ;
        RECT 53.920 180.515 54.255 180.845 ;
        RECT 54.425 180.515 54.595 181.015 ;
        RECT 54.765 180.590 55.115 181.985 ;
        RECT 51.605 179.775 52.190 180.345 ;
        RECT 52.440 180.175 53.835 180.345 ;
        RECT 52.440 179.830 52.770 180.175 ;
        RECT 52.985 179.605 53.360 180.005 ;
        RECT 53.540 179.830 53.835 180.175 ;
        RECT 54.005 179.605 54.675 180.345 ;
        RECT 54.845 179.775 55.115 180.590 ;
        RECT 55.285 181.435 55.745 181.985 ;
        RECT 55.935 181.435 56.265 182.155 ;
        RECT 55.285 180.065 55.535 181.435 ;
        RECT 56.465 181.265 56.765 181.815 ;
        RECT 56.935 181.485 57.215 182.155 ;
        RECT 55.825 181.095 56.765 181.265 ;
        RECT 55.825 180.845 55.995 181.095 ;
        RECT 57.135 180.845 57.400 181.205 ;
        RECT 57.625 181.015 57.855 182.155 ;
        RECT 58.025 181.005 58.355 181.985 ;
        RECT 58.525 181.015 58.735 182.155 ;
        RECT 59.425 181.645 59.685 182.155 ;
        RECT 55.705 180.515 55.995 180.845 ;
        RECT 56.165 180.595 56.505 180.845 ;
        RECT 56.725 180.595 57.400 180.845 ;
        RECT 57.605 180.595 57.935 180.845 ;
        RECT 55.825 180.425 55.995 180.515 ;
        RECT 55.825 180.235 57.215 180.425 ;
        RECT 55.285 179.775 55.845 180.065 ;
        RECT 56.015 179.605 56.265 180.065 ;
        RECT 56.885 179.875 57.215 180.235 ;
        RECT 57.625 179.605 57.855 180.425 ;
        RECT 58.105 180.405 58.355 181.005 ;
        RECT 59.425 180.595 59.765 181.475 ;
        RECT 59.935 180.765 60.105 181.985 ;
        RECT 60.345 181.650 60.960 182.155 ;
        RECT 60.345 181.115 60.595 181.480 ;
        RECT 60.765 181.475 60.960 181.650 ;
        RECT 61.130 181.645 61.605 181.985 ;
        RECT 61.775 181.610 61.990 182.155 ;
        RECT 60.765 181.285 61.095 181.475 ;
        RECT 61.315 181.115 62.030 181.410 ;
        RECT 62.200 181.285 62.475 181.985 ;
        RECT 60.345 180.945 62.135 181.115 ;
        RECT 59.935 180.515 60.730 180.765 ;
        RECT 59.935 180.425 60.185 180.515 ;
        RECT 58.025 179.775 58.355 180.405 ;
        RECT 58.525 179.605 58.735 180.425 ;
        RECT 59.425 179.605 59.685 180.425 ;
        RECT 59.855 180.005 60.185 180.425 ;
        RECT 60.900 180.090 61.155 180.945 ;
        RECT 60.365 179.825 61.155 180.090 ;
        RECT 61.325 180.245 61.735 180.765 ;
        RECT 61.905 180.515 62.135 180.945 ;
        RECT 62.305 180.255 62.475 181.285 ;
        RECT 62.705 181.095 63.035 181.940 ;
        RECT 63.205 181.145 63.375 182.155 ;
        RECT 63.545 181.425 63.885 181.985 ;
        RECT 64.115 181.655 64.430 182.155 ;
        RECT 64.610 181.685 65.495 181.855 ;
        RECT 62.645 181.015 63.035 181.095 ;
        RECT 63.545 181.050 64.440 181.425 ;
        RECT 62.645 180.965 62.860 181.015 ;
        RECT 62.645 180.385 62.815 180.965 ;
        RECT 63.545 180.845 63.735 181.050 ;
        RECT 64.610 180.845 64.780 181.685 ;
        RECT 65.720 181.655 65.970 181.985 ;
        RECT 62.985 180.515 63.735 180.845 ;
        RECT 63.905 180.515 64.780 180.845 ;
        RECT 62.645 180.345 62.870 180.385 ;
        RECT 63.535 180.345 63.735 180.515 ;
        RECT 62.645 180.260 63.025 180.345 ;
        RECT 61.325 179.825 61.525 180.245 ;
        RECT 61.715 179.605 62.045 180.065 ;
        RECT 62.215 179.775 62.475 180.255 ;
        RECT 62.695 179.825 63.025 180.260 ;
        RECT 63.195 179.605 63.365 180.215 ;
        RECT 63.535 179.820 63.865 180.345 ;
        RECT 64.125 179.605 64.335 180.135 ;
        RECT 64.610 180.055 64.780 180.515 ;
        RECT 64.950 180.555 65.270 181.515 ;
        RECT 65.440 180.765 65.630 181.485 ;
        RECT 65.800 180.585 65.970 181.655 ;
        RECT 66.140 181.355 66.310 182.155 ;
        RECT 66.480 181.710 67.585 181.880 ;
        RECT 66.480 181.095 66.650 181.710 ;
        RECT 67.795 181.560 68.045 181.985 ;
        RECT 68.215 181.695 68.480 182.155 ;
        RECT 66.820 181.175 67.350 181.540 ;
        RECT 67.795 181.430 68.100 181.560 ;
        RECT 66.140 181.005 66.650 181.095 ;
        RECT 66.140 180.835 67.010 181.005 ;
        RECT 66.140 180.765 66.310 180.835 ;
        RECT 66.430 180.585 66.630 180.615 ;
        RECT 64.950 180.225 65.415 180.555 ;
        RECT 65.800 180.285 66.630 180.585 ;
        RECT 65.800 180.055 65.970 180.285 ;
        RECT 64.610 179.885 65.395 180.055 ;
        RECT 65.565 179.885 65.970 180.055 ;
        RECT 66.150 179.605 66.520 180.105 ;
        RECT 66.840 180.055 67.010 180.835 ;
        RECT 67.180 180.475 67.350 181.175 ;
        RECT 67.520 180.645 67.760 181.240 ;
        RECT 67.180 180.255 67.705 180.475 ;
        RECT 67.930 180.325 68.100 181.430 ;
        RECT 67.875 180.195 68.100 180.325 ;
        RECT 68.270 180.235 68.550 181.185 ;
        RECT 67.875 180.055 68.045 180.195 ;
        RECT 66.840 179.885 67.515 180.055 ;
        RECT 67.710 179.885 68.045 180.055 ;
        RECT 68.215 179.605 68.465 180.065 ;
        RECT 68.720 179.865 68.905 181.985 ;
        RECT 69.075 181.655 69.405 182.155 ;
        RECT 69.575 181.485 69.745 181.985 ;
        RECT 69.080 181.315 69.745 181.485 ;
        RECT 69.080 180.325 69.310 181.315 ;
        RECT 69.480 180.495 69.830 181.145 ;
        RECT 70.005 180.990 70.295 182.155 ;
        RECT 70.465 181.720 75.810 182.155 ;
        RECT 75.985 181.720 81.330 182.155 ;
        RECT 69.080 180.155 69.745 180.325 ;
        RECT 69.075 179.605 69.405 179.985 ;
        RECT 69.575 179.865 69.745 180.155 ;
        RECT 70.005 179.605 70.295 180.330 ;
        RECT 72.050 180.150 72.390 180.980 ;
        RECT 73.870 180.470 74.220 181.720 ;
        RECT 77.570 180.150 77.910 180.980 ;
        RECT 79.390 180.470 79.740 181.720 ;
        RECT 81.505 181.065 82.715 182.155 ;
        RECT 81.505 180.355 82.025 180.895 ;
        RECT 82.195 180.525 82.715 181.065 ;
        RECT 82.885 181.065 84.095 182.155 ;
        RECT 82.885 180.525 83.405 181.065 ;
        RECT 83.575 180.355 84.095 180.895 ;
        RECT 70.465 179.605 75.810 180.150 ;
        RECT 75.985 179.605 81.330 180.150 ;
        RECT 81.505 179.605 82.715 180.355 ;
        RECT 82.885 179.605 84.095 180.355 ;
        RECT 5.520 179.435 84.180 179.605 ;
        RECT 5.605 178.685 6.815 179.435 ;
        RECT 6.985 178.890 12.330 179.435 ;
        RECT 5.605 178.145 6.125 178.685 ;
        RECT 6.295 177.975 6.815 178.515 ;
        RECT 8.570 178.060 8.910 178.890 ;
        RECT 12.505 178.665 14.175 179.435 ;
        RECT 14.380 178.695 14.995 179.265 ;
        RECT 15.165 178.925 15.380 179.435 ;
        RECT 15.610 178.925 15.890 179.255 ;
        RECT 16.070 178.925 16.310 179.435 ;
        RECT 5.605 176.885 6.815 177.975 ;
        RECT 10.390 177.320 10.740 178.570 ;
        RECT 12.505 178.145 13.255 178.665 ;
        RECT 13.425 177.975 14.175 178.495 ;
        RECT 6.985 176.885 12.330 177.320 ;
        RECT 12.505 176.885 14.175 177.975 ;
        RECT 14.380 177.675 14.695 178.695 ;
        RECT 14.865 178.025 15.035 178.525 ;
        RECT 15.285 178.195 15.550 178.755 ;
        RECT 15.720 178.025 15.890 178.925 ;
        RECT 16.645 178.890 21.990 179.435 ;
        RECT 16.060 178.195 16.415 178.755 ;
        RECT 18.230 178.060 18.570 178.890 ;
        RECT 22.625 178.715 22.965 179.225 ;
        RECT 14.865 177.855 16.290 178.025 ;
        RECT 14.380 177.055 14.915 177.675 ;
        RECT 15.085 176.885 15.415 177.685 ;
        RECT 15.900 177.680 16.290 177.855 ;
        RECT 20.050 177.320 20.400 178.570 ;
        RECT 16.645 176.885 21.990 177.320 ;
        RECT 22.625 177.315 22.885 178.715 ;
        RECT 23.135 178.635 23.405 179.435 ;
        RECT 23.060 178.195 23.390 178.445 ;
        RECT 23.585 178.195 23.865 179.165 ;
        RECT 24.045 178.195 24.345 179.165 ;
        RECT 24.525 178.195 24.875 179.160 ;
        RECT 25.095 178.935 25.590 179.265 ;
        RECT 23.075 178.025 23.390 178.195 ;
        RECT 25.095 178.025 25.265 178.935 ;
        RECT 23.075 177.855 25.265 178.025 ;
        RECT 22.625 177.055 22.965 177.315 ;
        RECT 23.135 176.885 23.465 177.685 ;
        RECT 23.930 177.055 24.180 177.855 ;
        RECT 24.365 176.885 24.695 177.605 ;
        RECT 24.915 177.055 25.165 177.855 ;
        RECT 25.435 177.445 25.675 178.755 ;
        RECT 26.305 178.695 26.745 179.255 ;
        RECT 26.915 178.695 27.365 179.435 ;
        RECT 27.535 178.865 27.705 179.265 ;
        RECT 27.875 179.035 28.295 179.435 ;
        RECT 28.465 178.865 28.695 179.265 ;
        RECT 27.535 178.695 28.695 178.865 ;
        RECT 28.865 178.695 29.355 179.265 ;
        RECT 26.305 177.685 26.615 178.695 ;
        RECT 26.785 178.075 26.955 178.525 ;
        RECT 27.125 178.245 27.515 178.525 ;
        RECT 27.700 178.195 27.945 178.525 ;
        RECT 26.785 177.905 27.575 178.075 ;
        RECT 25.335 176.885 25.670 177.265 ;
        RECT 26.305 177.055 26.745 177.685 ;
        RECT 26.920 176.885 27.235 177.735 ;
        RECT 27.405 177.225 27.575 177.905 ;
        RECT 27.745 177.395 27.945 178.195 ;
        RECT 28.145 177.395 28.395 178.525 ;
        RECT 28.610 178.195 29.015 178.525 ;
        RECT 29.185 178.025 29.355 178.695 ;
        RECT 29.525 178.665 31.195 179.435 ;
        RECT 31.365 178.710 31.655 179.435 ;
        RECT 32.745 178.695 33.210 179.240 ;
        RECT 29.525 178.145 30.275 178.665 ;
        RECT 28.585 177.855 29.355 178.025 ;
        RECT 30.445 177.975 31.195 178.495 ;
        RECT 28.585 177.225 28.835 177.855 ;
        RECT 27.405 177.055 28.835 177.225 ;
        RECT 29.015 176.885 29.345 177.685 ;
        RECT 29.525 176.885 31.195 177.975 ;
        RECT 31.365 176.885 31.655 178.050 ;
        RECT 32.745 177.735 32.915 178.695 ;
        RECT 33.715 178.615 33.885 179.435 ;
        RECT 34.055 178.785 34.385 179.265 ;
        RECT 34.555 179.045 34.905 179.435 ;
        RECT 35.075 178.865 35.305 179.265 ;
        RECT 34.795 178.785 35.305 178.865 ;
        RECT 34.055 178.695 35.305 178.785 ;
        RECT 35.475 178.695 35.795 179.175 ;
        RECT 34.055 178.615 34.965 178.695 ;
        RECT 33.085 178.075 33.330 178.525 ;
        RECT 33.590 178.245 34.285 178.445 ;
        RECT 34.455 178.275 35.055 178.445 ;
        RECT 34.455 178.075 34.625 178.275 ;
        RECT 35.285 178.105 35.455 178.525 ;
        RECT 33.085 177.905 34.625 178.075 ;
        RECT 34.795 177.935 35.455 178.105 ;
        RECT 34.795 177.735 34.965 177.935 ;
        RECT 35.625 177.765 35.795 178.695 ;
        RECT 35.965 178.635 36.660 179.265 ;
        RECT 36.865 178.635 37.175 179.435 ;
        RECT 37.510 178.925 37.750 179.435 ;
        RECT 37.930 178.925 38.210 179.255 ;
        RECT 38.440 178.925 38.655 179.435 ;
        RECT 36.485 178.585 36.660 178.635 ;
        RECT 35.985 178.195 36.320 178.445 ;
        RECT 36.490 178.035 36.660 178.585 ;
        RECT 36.830 178.195 37.165 178.465 ;
        RECT 37.405 178.195 37.760 178.755 ;
        RECT 32.745 177.565 34.965 177.735 ;
        RECT 35.135 177.565 35.795 177.765 ;
        RECT 32.745 176.885 33.045 177.395 ;
        RECT 33.215 177.055 33.545 177.565 ;
        RECT 35.135 177.395 35.305 177.565 ;
        RECT 33.715 176.885 34.345 177.395 ;
        RECT 34.925 177.225 35.305 177.395 ;
        RECT 35.475 176.885 35.775 177.395 ;
        RECT 35.965 176.885 36.225 178.025 ;
        RECT 36.395 177.055 36.725 178.035 ;
        RECT 37.930 178.025 38.100 178.925 ;
        RECT 38.270 178.195 38.535 178.755 ;
        RECT 38.825 178.695 39.440 179.265 ;
        RECT 39.730 178.865 39.905 179.265 ;
        RECT 40.075 179.055 40.405 179.435 ;
        RECT 40.650 178.935 40.880 179.265 ;
        RECT 39.730 178.695 40.360 178.865 ;
        RECT 38.785 178.025 38.955 178.525 ;
        RECT 36.895 176.885 37.175 178.025 ;
        RECT 37.530 177.855 38.955 178.025 ;
        RECT 37.530 177.680 37.920 177.855 ;
        RECT 38.405 176.885 38.735 177.685 ;
        RECT 39.125 177.675 39.440 178.695 ;
        RECT 40.190 178.525 40.360 178.695 ;
        RECT 39.645 177.845 40.010 178.525 ;
        RECT 40.190 178.195 40.540 178.525 ;
        RECT 40.190 177.675 40.360 178.195 ;
        RECT 38.905 177.055 39.440 177.675 ;
        RECT 39.730 177.505 40.360 177.675 ;
        RECT 40.710 177.645 40.880 178.935 ;
        RECT 41.080 177.825 41.360 179.100 ;
        RECT 41.585 179.095 41.855 179.100 ;
        RECT 41.545 178.925 41.855 179.095 ;
        RECT 42.315 179.055 42.645 179.435 ;
        RECT 42.815 179.180 43.150 179.225 ;
        RECT 41.585 177.825 41.855 178.925 ;
        RECT 42.045 177.825 42.385 178.855 ;
        RECT 42.815 178.715 43.155 179.180 ;
        RECT 43.330 178.905 43.620 179.255 ;
        RECT 43.815 179.075 44.145 179.435 ;
        RECT 44.315 178.905 44.545 179.210 ;
        RECT 43.330 178.735 44.545 178.905 ;
        RECT 44.735 179.095 44.905 179.130 ;
        RECT 44.735 178.925 44.935 179.095 ;
        RECT 42.555 178.195 42.815 178.525 ;
        RECT 42.555 177.645 42.725 178.195 ;
        RECT 42.985 178.025 43.155 178.715 ;
        RECT 44.735 178.565 44.905 178.925 ;
        RECT 45.305 178.840 45.625 179.265 ;
        RECT 45.795 179.010 46.125 179.435 ;
        RECT 46.295 179.015 47.385 179.265 ;
        RECT 47.575 179.015 48.665 179.265 ;
        RECT 46.295 178.840 46.465 179.015 ;
        RECT 45.305 178.670 46.465 178.840 ;
        RECT 46.635 178.675 48.325 178.845 ;
        RECT 48.495 178.840 48.665 179.015 ;
        RECT 48.835 179.010 49.165 179.435 ;
        RECT 49.335 178.840 49.585 179.265 ;
        RECT 43.390 178.415 43.650 178.525 ;
        RECT 43.385 178.245 43.650 178.415 ;
        RECT 43.390 178.195 43.650 178.245 ;
        RECT 43.830 178.195 44.215 178.525 ;
        RECT 44.385 178.395 44.905 178.565 ;
        RECT 45.180 178.415 46.290 178.445 ;
        RECT 39.730 177.055 39.905 177.505 ;
        RECT 40.710 177.475 42.725 177.645 ;
        RECT 40.075 176.885 40.405 177.325 ;
        RECT 40.710 177.055 40.880 177.475 ;
        RECT 41.115 176.885 41.785 177.295 ;
        RECT 42.000 177.055 42.170 177.475 ;
        RECT 42.370 176.885 42.700 177.295 ;
        RECT 42.895 177.055 43.155 178.025 ;
        RECT 43.330 176.885 43.650 178.025 ;
        RECT 43.830 177.145 44.025 178.195 ;
        RECT 44.385 178.015 44.555 178.395 ;
        RECT 45.180 178.245 46.315 178.415 ;
        RECT 46.580 178.245 47.235 178.445 ;
        RECT 44.205 177.735 44.555 178.015 ;
        RECT 44.745 177.865 44.990 178.225 ;
        RECT 47.520 178.035 47.810 178.675 ;
        RECT 48.495 178.670 49.585 178.840 ;
        RECT 49.765 178.850 50.075 179.265 ;
        RECT 50.270 179.055 50.600 179.435 ;
        RECT 50.770 179.095 52.175 179.265 ;
        RECT 50.770 178.865 50.940 179.095 ;
        RECT 47.980 178.245 48.610 178.445 ;
        RECT 48.900 178.415 49.530 178.445 ;
        RECT 48.900 178.245 49.535 178.415 ;
        RECT 45.375 177.865 47.305 178.035 ;
        RECT 44.205 177.055 44.535 177.735 ;
        RECT 44.735 176.885 44.990 177.685 ;
        RECT 45.375 177.055 45.705 177.865 ;
        RECT 45.875 176.885 46.045 177.695 ;
        RECT 46.215 177.055 46.545 177.865 ;
        RECT 46.715 176.885 46.885 177.695 ;
        RECT 47.055 177.225 47.305 177.865 ;
        RECT 47.520 177.865 49.585 178.035 ;
        RECT 47.520 177.395 47.905 177.865 ;
        RECT 48.075 177.225 48.245 177.695 ;
        RECT 48.415 177.395 48.745 177.865 ;
        RECT 48.915 177.225 49.165 177.695 ;
        RECT 47.055 177.055 49.165 177.225 ;
        RECT 49.335 177.055 49.585 177.865 ;
        RECT 49.765 177.735 49.935 178.850 ;
        RECT 50.245 178.695 50.940 178.865 ;
        RECT 52.005 178.865 52.175 179.095 ;
        RECT 52.445 179.035 52.775 179.435 ;
        RECT 53.015 178.865 53.185 179.265 ;
        RECT 50.245 178.525 50.415 178.695 ;
        RECT 50.105 178.195 50.415 178.525 ;
        RECT 50.585 178.195 50.920 178.525 ;
        RECT 51.190 178.195 51.385 178.770 ;
        RECT 51.645 178.525 51.835 178.755 ;
        RECT 52.005 178.695 53.185 178.865 ;
        RECT 53.905 178.615 54.165 179.435 ;
        RECT 54.335 178.615 54.665 179.035 ;
        RECT 54.845 178.865 55.105 179.265 ;
        RECT 55.275 179.035 55.605 179.435 ;
        RECT 55.775 178.865 55.945 179.215 ;
        RECT 56.115 179.035 56.490 179.435 ;
        RECT 54.845 178.695 56.510 178.865 ;
        RECT 56.680 178.760 56.955 179.105 ;
        RECT 54.415 178.525 54.665 178.615 ;
        RECT 56.340 178.525 56.510 178.695 ;
        RECT 51.645 178.195 51.990 178.525 ;
        RECT 52.300 178.195 52.775 178.525 ;
        RECT 53.030 178.195 53.215 178.525 ;
        RECT 53.910 178.195 54.245 178.445 ;
        RECT 54.415 178.195 55.130 178.525 ;
        RECT 55.345 178.195 56.170 178.525 ;
        RECT 56.340 178.195 56.615 178.525 ;
        RECT 50.245 178.025 50.415 178.195 ;
        RECT 50.245 177.855 53.185 178.025 ;
        RECT 49.765 177.095 50.105 177.735 ;
        RECT 50.695 177.515 52.255 177.685 ;
        RECT 50.275 176.885 50.520 177.345 ;
        RECT 50.695 177.055 50.945 177.515 ;
        RECT 51.135 176.885 51.805 177.265 ;
        RECT 52.005 177.055 52.255 177.515 ;
        RECT 53.015 177.055 53.185 177.855 ;
        RECT 53.905 176.885 54.165 178.025 ;
        RECT 54.415 177.635 54.585 178.195 ;
        RECT 54.845 177.735 55.175 178.025 ;
        RECT 55.345 177.905 55.590 178.195 ;
        RECT 56.340 178.025 56.510 178.195 ;
        RECT 56.785 178.025 56.955 178.760 ;
        RECT 57.125 178.710 57.415 179.435 ;
        RECT 57.585 178.785 57.845 179.265 ;
        RECT 58.015 178.975 58.345 179.435 ;
        RECT 58.535 178.795 58.735 179.215 ;
        RECT 55.850 177.855 56.510 178.025 ;
        RECT 55.850 177.735 56.020 177.855 ;
        RECT 54.845 177.565 56.020 177.735 ;
        RECT 54.405 177.065 56.020 177.395 ;
        RECT 56.190 176.885 56.470 177.685 ;
        RECT 56.680 177.055 56.955 178.025 ;
        RECT 57.125 176.885 57.415 178.050 ;
        RECT 57.585 177.755 57.755 178.785 ;
        RECT 57.925 178.095 58.155 178.525 ;
        RECT 58.325 178.275 58.735 178.795 ;
        RECT 58.905 178.950 59.695 179.215 ;
        RECT 58.905 178.095 59.160 178.950 ;
        RECT 59.875 178.615 60.205 179.035 ;
        RECT 60.375 178.615 60.635 179.435 ;
        RECT 60.805 179.055 61.695 179.225 ;
        RECT 59.875 178.525 60.125 178.615 ;
        RECT 59.330 178.275 60.125 178.525 ;
        RECT 60.805 178.500 61.355 178.885 ;
        RECT 57.925 177.925 59.715 178.095 ;
        RECT 57.585 177.055 57.860 177.755 ;
        RECT 58.030 177.630 58.745 177.925 ;
        RECT 58.965 177.565 59.295 177.755 ;
        RECT 58.070 176.885 58.285 177.430 ;
        RECT 58.455 177.055 58.930 177.395 ;
        RECT 59.100 177.390 59.295 177.565 ;
        RECT 59.465 177.560 59.715 177.925 ;
        RECT 59.100 176.885 59.715 177.390 ;
        RECT 59.955 177.055 60.125 178.275 ;
        RECT 60.295 177.565 60.635 178.445 ;
        RECT 61.525 178.330 61.695 179.055 ;
        RECT 60.805 178.260 61.695 178.330 ;
        RECT 61.865 178.730 62.085 179.215 ;
        RECT 62.255 178.895 62.505 179.435 ;
        RECT 62.675 178.785 62.935 179.265 ;
        RECT 61.865 178.305 62.195 178.730 ;
        RECT 60.805 178.235 61.700 178.260 ;
        RECT 60.805 178.220 61.710 178.235 ;
        RECT 60.805 178.205 61.715 178.220 ;
        RECT 60.805 178.200 61.725 178.205 ;
        RECT 60.805 178.190 61.730 178.200 ;
        RECT 60.805 178.180 61.735 178.190 ;
        RECT 60.805 178.175 61.745 178.180 ;
        RECT 60.805 178.165 61.755 178.175 ;
        RECT 60.805 178.160 61.765 178.165 ;
        RECT 60.805 177.710 61.065 178.160 ;
        RECT 61.430 178.155 61.765 178.160 ;
        RECT 61.430 178.150 61.780 178.155 ;
        RECT 61.430 178.140 61.795 178.150 ;
        RECT 61.430 178.135 61.820 178.140 ;
        RECT 62.365 178.135 62.595 178.530 ;
        RECT 61.430 178.130 62.595 178.135 ;
        RECT 61.460 178.095 62.595 178.130 ;
        RECT 61.495 178.070 62.595 178.095 ;
        RECT 61.525 178.040 62.595 178.070 ;
        RECT 61.545 178.010 62.595 178.040 ;
        RECT 61.565 177.980 62.595 178.010 ;
        RECT 61.635 177.970 62.595 177.980 ;
        RECT 61.660 177.960 62.595 177.970 ;
        RECT 61.680 177.945 62.595 177.960 ;
        RECT 61.700 177.930 62.595 177.945 ;
        RECT 61.705 177.920 62.490 177.930 ;
        RECT 61.720 177.885 62.490 177.920 ;
        RECT 61.235 177.565 61.565 177.810 ;
        RECT 61.735 177.635 62.490 177.885 ;
        RECT 62.765 177.755 62.935 178.785 ;
        RECT 63.195 178.885 63.365 179.175 ;
        RECT 63.535 179.055 63.865 179.435 ;
        RECT 63.195 178.715 63.860 178.885 ;
        RECT 63.110 177.895 63.460 178.545 ;
        RECT 61.235 177.540 61.420 177.565 ;
        RECT 60.805 177.440 61.420 177.540 ;
        RECT 60.375 176.885 60.635 177.395 ;
        RECT 60.805 176.885 61.410 177.440 ;
        RECT 61.585 177.055 62.065 177.395 ;
        RECT 62.235 176.885 62.490 177.430 ;
        RECT 62.660 177.055 62.935 177.755 ;
        RECT 63.630 177.725 63.860 178.715 ;
        RECT 63.195 177.555 63.860 177.725 ;
        RECT 63.195 177.055 63.365 177.555 ;
        RECT 63.535 176.885 63.865 177.385 ;
        RECT 64.035 177.055 64.220 179.175 ;
        RECT 64.475 178.975 64.725 179.435 ;
        RECT 64.895 178.985 65.230 179.155 ;
        RECT 65.425 178.985 66.100 179.155 ;
        RECT 64.895 178.845 65.065 178.985 ;
        RECT 64.390 177.855 64.670 178.805 ;
        RECT 64.840 178.715 65.065 178.845 ;
        RECT 64.840 177.610 65.010 178.715 ;
        RECT 65.235 178.565 65.760 178.785 ;
        RECT 65.180 177.800 65.420 178.395 ;
        RECT 65.590 177.865 65.760 178.565 ;
        RECT 65.930 178.205 66.100 178.985 ;
        RECT 66.420 178.935 66.790 179.435 ;
        RECT 66.970 178.985 67.375 179.155 ;
        RECT 67.545 178.985 68.330 179.155 ;
        RECT 66.970 178.755 67.140 178.985 ;
        RECT 66.310 178.455 67.140 178.755 ;
        RECT 67.525 178.485 67.990 178.815 ;
        RECT 66.310 178.425 66.510 178.455 ;
        RECT 66.630 178.205 66.800 178.275 ;
        RECT 65.930 178.035 66.800 178.205 ;
        RECT 66.290 177.945 66.800 178.035 ;
        RECT 64.840 177.480 65.145 177.610 ;
        RECT 65.590 177.500 66.120 177.865 ;
        RECT 64.460 176.885 64.725 177.345 ;
        RECT 64.895 177.055 65.145 177.480 ;
        RECT 66.290 177.330 66.460 177.945 ;
        RECT 65.355 177.160 66.460 177.330 ;
        RECT 66.630 176.885 66.800 177.685 ;
        RECT 66.970 177.385 67.140 178.455 ;
        RECT 67.310 177.555 67.500 178.275 ;
        RECT 67.670 177.525 67.990 178.485 ;
        RECT 68.160 178.525 68.330 178.985 ;
        RECT 68.605 178.905 68.815 179.435 ;
        RECT 69.075 178.695 69.405 179.220 ;
        RECT 69.575 178.825 69.745 179.435 ;
        RECT 69.915 178.780 70.245 179.215 ;
        RECT 70.465 178.890 75.810 179.435 ;
        RECT 75.985 178.890 81.330 179.435 ;
        RECT 69.915 178.695 70.295 178.780 ;
        RECT 69.205 178.525 69.405 178.695 ;
        RECT 70.070 178.655 70.295 178.695 ;
        RECT 68.160 178.195 69.035 178.525 ;
        RECT 69.205 178.195 69.955 178.525 ;
        RECT 66.970 177.055 67.220 177.385 ;
        RECT 68.160 177.355 68.330 178.195 ;
        RECT 69.205 177.990 69.395 178.195 ;
        RECT 70.125 178.075 70.295 178.655 ;
        RECT 70.080 178.025 70.295 178.075 ;
        RECT 72.050 178.060 72.390 178.890 ;
        RECT 68.500 177.615 69.395 177.990 ;
        RECT 69.905 177.945 70.295 178.025 ;
        RECT 67.445 177.185 68.330 177.355 ;
        RECT 68.510 176.885 68.825 177.385 ;
        RECT 69.055 177.055 69.395 177.615 ;
        RECT 69.565 176.885 69.735 177.895 ;
        RECT 69.905 177.100 70.235 177.945 ;
        RECT 73.870 177.320 74.220 178.570 ;
        RECT 77.570 178.060 77.910 178.890 ;
        RECT 81.505 178.685 82.715 179.435 ;
        RECT 82.885 178.685 84.095 179.435 ;
        RECT 79.390 177.320 79.740 178.570 ;
        RECT 81.505 178.145 82.025 178.685 ;
        RECT 82.195 177.975 82.715 178.515 ;
        RECT 70.465 176.885 75.810 177.320 ;
        RECT 75.985 176.885 81.330 177.320 ;
        RECT 81.505 176.885 82.715 177.975 ;
        RECT 82.885 177.975 83.405 178.515 ;
        RECT 83.575 178.145 84.095 178.685 ;
        RECT 82.885 176.885 84.095 177.975 ;
        RECT 5.520 176.715 84.180 176.885 ;
        RECT 5.605 175.625 6.815 176.715 ;
        RECT 6.985 175.625 10.495 176.715 ;
        RECT 11.185 175.655 11.515 176.500 ;
        RECT 11.685 175.705 11.855 176.715 ;
        RECT 12.025 175.985 12.365 176.545 ;
        RECT 12.595 176.215 12.910 176.715 ;
        RECT 13.090 176.245 13.975 176.415 ;
        RECT 5.605 174.915 6.125 175.455 ;
        RECT 6.295 175.085 6.815 175.625 ;
        RECT 6.985 174.935 8.635 175.455 ;
        RECT 8.805 175.105 10.495 175.625 ;
        RECT 11.125 175.575 11.515 175.655 ;
        RECT 12.025 175.610 12.920 175.985 ;
        RECT 11.125 175.525 11.340 175.575 ;
        RECT 11.125 174.945 11.295 175.525 ;
        RECT 12.025 175.405 12.215 175.610 ;
        RECT 13.090 175.405 13.260 176.245 ;
        RECT 14.200 176.215 14.450 176.545 ;
        RECT 11.465 175.075 12.215 175.405 ;
        RECT 12.385 175.075 13.260 175.405 ;
        RECT 5.605 174.165 6.815 174.915 ;
        RECT 6.985 174.165 10.495 174.935 ;
        RECT 11.125 174.905 11.350 174.945 ;
        RECT 12.015 174.905 12.215 175.075 ;
        RECT 11.125 174.820 11.505 174.905 ;
        RECT 11.175 174.385 11.505 174.820 ;
        RECT 11.675 174.165 11.845 174.775 ;
        RECT 12.015 174.380 12.345 174.905 ;
        RECT 12.605 174.165 12.815 174.695 ;
        RECT 13.090 174.615 13.260 175.075 ;
        RECT 13.430 175.115 13.750 176.075 ;
        RECT 13.920 175.325 14.110 176.045 ;
        RECT 14.280 175.145 14.450 176.215 ;
        RECT 14.620 175.915 14.790 176.715 ;
        RECT 14.960 176.270 16.065 176.440 ;
        RECT 14.960 175.655 15.130 176.270 ;
        RECT 16.275 176.120 16.525 176.545 ;
        RECT 16.695 176.255 16.960 176.715 ;
        RECT 15.300 175.735 15.830 176.100 ;
        RECT 16.275 175.990 16.580 176.120 ;
        RECT 14.620 175.565 15.130 175.655 ;
        RECT 14.620 175.395 15.490 175.565 ;
        RECT 14.620 175.325 14.790 175.395 ;
        RECT 14.910 175.145 15.110 175.175 ;
        RECT 13.430 174.785 13.895 175.115 ;
        RECT 14.280 174.845 15.110 175.145 ;
        RECT 14.280 174.615 14.450 174.845 ;
        RECT 13.090 174.445 13.875 174.615 ;
        RECT 14.045 174.445 14.450 174.615 ;
        RECT 14.630 174.165 15.000 174.665 ;
        RECT 15.320 174.615 15.490 175.395 ;
        RECT 15.660 175.035 15.830 175.735 ;
        RECT 16.000 175.205 16.240 175.800 ;
        RECT 15.660 174.815 16.185 175.035 ;
        RECT 16.410 174.885 16.580 175.990 ;
        RECT 16.355 174.755 16.580 174.885 ;
        RECT 16.750 174.795 17.030 175.745 ;
        RECT 16.355 174.615 16.525 174.755 ;
        RECT 15.320 174.445 15.995 174.615 ;
        RECT 16.190 174.445 16.525 174.615 ;
        RECT 16.695 174.165 16.945 174.625 ;
        RECT 17.200 174.425 17.385 176.545 ;
        RECT 17.555 176.215 17.885 176.715 ;
        RECT 18.055 176.045 18.225 176.545 ;
        RECT 17.560 175.875 18.225 176.045 ;
        RECT 17.560 174.885 17.790 175.875 ;
        RECT 17.960 175.055 18.310 175.705 ;
        RECT 18.485 175.550 18.775 176.715 ;
        RECT 18.945 176.205 19.205 176.715 ;
        RECT 18.945 175.155 19.285 176.035 ;
        RECT 19.455 175.325 19.625 176.545 ;
        RECT 19.865 176.210 20.480 176.715 ;
        RECT 19.865 175.675 20.115 176.040 ;
        RECT 20.285 176.035 20.480 176.210 ;
        RECT 20.650 176.205 21.125 176.545 ;
        RECT 21.295 176.170 21.510 176.715 ;
        RECT 20.285 175.845 20.615 176.035 ;
        RECT 20.835 175.675 21.550 175.970 ;
        RECT 21.720 175.845 21.995 176.545 ;
        RECT 22.255 176.045 22.425 176.545 ;
        RECT 22.595 176.215 22.925 176.715 ;
        RECT 22.255 175.875 22.920 176.045 ;
        RECT 19.865 175.505 21.655 175.675 ;
        RECT 19.455 175.075 20.250 175.325 ;
        RECT 19.455 174.985 19.705 175.075 ;
        RECT 17.560 174.715 18.225 174.885 ;
        RECT 17.555 174.165 17.885 174.545 ;
        RECT 18.055 174.425 18.225 174.715 ;
        RECT 18.485 174.165 18.775 174.890 ;
        RECT 18.945 174.165 19.205 174.985 ;
        RECT 19.375 174.565 19.705 174.985 ;
        RECT 20.420 174.650 20.675 175.505 ;
        RECT 19.885 174.385 20.675 174.650 ;
        RECT 20.845 174.805 21.255 175.325 ;
        RECT 21.425 175.075 21.655 175.505 ;
        RECT 21.825 174.815 21.995 175.845 ;
        RECT 22.170 175.055 22.520 175.705 ;
        RECT 22.690 174.885 22.920 175.875 ;
        RECT 20.845 174.385 21.045 174.805 ;
        RECT 21.235 174.165 21.565 174.625 ;
        RECT 21.735 174.335 21.995 174.815 ;
        RECT 22.255 174.715 22.920 174.885 ;
        RECT 22.255 174.425 22.425 174.715 ;
        RECT 22.595 174.165 22.925 174.545 ;
        RECT 23.095 174.425 23.280 176.545 ;
        RECT 23.520 176.255 23.785 176.715 ;
        RECT 23.955 176.120 24.205 176.545 ;
        RECT 24.415 176.270 25.520 176.440 ;
        RECT 23.900 175.990 24.205 176.120 ;
        RECT 23.450 174.795 23.730 175.745 ;
        RECT 23.900 174.885 24.070 175.990 ;
        RECT 24.240 175.205 24.480 175.800 ;
        RECT 24.650 175.735 25.180 176.100 ;
        RECT 24.650 175.035 24.820 175.735 ;
        RECT 25.350 175.655 25.520 176.270 ;
        RECT 25.690 175.915 25.860 176.715 ;
        RECT 26.030 176.215 26.280 176.545 ;
        RECT 26.505 176.245 27.390 176.415 ;
        RECT 25.350 175.565 25.860 175.655 ;
        RECT 23.900 174.755 24.125 174.885 ;
        RECT 24.295 174.815 24.820 175.035 ;
        RECT 24.990 175.395 25.860 175.565 ;
        RECT 23.535 174.165 23.785 174.625 ;
        RECT 23.955 174.615 24.125 174.755 ;
        RECT 24.990 174.615 25.160 175.395 ;
        RECT 25.690 175.325 25.860 175.395 ;
        RECT 25.370 175.145 25.570 175.175 ;
        RECT 26.030 175.145 26.200 176.215 ;
        RECT 26.370 175.325 26.560 176.045 ;
        RECT 25.370 174.845 26.200 175.145 ;
        RECT 26.730 175.115 27.050 176.075 ;
        RECT 23.955 174.445 24.290 174.615 ;
        RECT 24.485 174.445 25.160 174.615 ;
        RECT 25.480 174.165 25.850 174.665 ;
        RECT 26.030 174.615 26.200 174.845 ;
        RECT 26.585 174.785 27.050 175.115 ;
        RECT 27.220 175.405 27.390 176.245 ;
        RECT 27.570 176.215 27.885 176.715 ;
        RECT 28.115 175.985 28.455 176.545 ;
        RECT 27.560 175.610 28.455 175.985 ;
        RECT 28.625 175.705 28.795 176.715 ;
        RECT 28.265 175.405 28.455 175.610 ;
        RECT 28.965 175.655 29.295 176.500 ;
        RECT 30.005 175.660 30.310 176.445 ;
        RECT 30.490 176.245 31.175 176.715 ;
        RECT 30.485 175.725 31.180 176.035 ;
        RECT 28.965 175.575 29.355 175.655 ;
        RECT 29.140 175.525 29.355 175.575 ;
        RECT 27.220 175.075 28.095 175.405 ;
        RECT 28.265 175.075 29.015 175.405 ;
        RECT 27.220 174.615 27.390 175.075 ;
        RECT 28.265 174.905 28.465 175.075 ;
        RECT 29.185 174.945 29.355 175.525 ;
        RECT 29.130 174.905 29.355 174.945 ;
        RECT 26.030 174.445 26.435 174.615 ;
        RECT 26.605 174.445 27.390 174.615 ;
        RECT 27.665 174.165 27.875 174.695 ;
        RECT 28.135 174.380 28.465 174.905 ;
        RECT 28.975 174.820 29.355 174.905 ;
        RECT 30.005 174.855 30.180 175.660 ;
        RECT 31.355 175.555 31.640 176.500 ;
        RECT 31.815 176.265 32.145 176.715 ;
        RECT 32.315 176.095 32.485 176.525 ;
        RECT 32.745 176.280 38.090 176.715 ;
        RECT 30.780 175.405 31.640 175.555 ;
        RECT 30.355 175.385 31.640 175.405 ;
        RECT 31.810 175.865 32.485 176.095 ;
        RECT 30.355 175.025 31.340 175.385 ;
        RECT 31.810 175.215 32.045 175.865 ;
        RECT 28.635 174.165 28.805 174.775 ;
        RECT 28.975 174.385 29.305 174.820 ;
        RECT 30.005 174.335 30.245 174.855 ;
        RECT 31.170 174.690 31.340 175.025 ;
        RECT 31.510 174.885 32.045 175.215 ;
        RECT 31.825 174.735 32.045 174.885 ;
        RECT 32.215 174.845 32.515 175.695 ;
        RECT 30.415 174.165 30.810 174.660 ;
        RECT 31.170 174.495 31.545 174.690 ;
        RECT 31.375 174.350 31.545 174.495 ;
        RECT 31.825 174.360 32.065 174.735 ;
        RECT 34.330 174.710 34.670 175.540 ;
        RECT 36.150 175.030 36.500 176.280 ;
        RECT 38.450 175.745 38.840 175.920 ;
        RECT 39.325 175.915 39.655 176.715 ;
        RECT 39.825 175.925 40.360 176.545 ;
        RECT 41.030 176.205 42.685 176.495 ;
        RECT 38.450 175.575 39.875 175.745 ;
        RECT 38.325 174.845 38.680 175.405 ;
        RECT 32.235 174.165 32.570 174.670 ;
        RECT 32.745 174.165 38.090 174.710 ;
        RECT 38.850 174.675 39.020 175.575 ;
        RECT 39.190 174.845 39.455 175.405 ;
        RECT 39.705 175.075 39.875 175.575 ;
        RECT 40.045 174.905 40.360 175.925 ;
        RECT 41.030 175.865 42.620 176.035 ;
        RECT 42.855 175.915 43.135 176.715 ;
        RECT 41.030 175.575 41.350 175.865 ;
        RECT 42.450 175.745 42.620 175.865 ;
        RECT 41.545 175.525 42.260 175.695 ;
        RECT 42.450 175.575 43.175 175.745 ;
        RECT 43.345 175.575 43.615 176.545 ;
        RECT 38.430 174.165 38.670 174.675 ;
        RECT 38.850 174.345 39.130 174.675 ;
        RECT 39.360 174.165 39.575 174.675 ;
        RECT 39.745 174.335 40.360 174.905 ;
        RECT 41.030 174.835 41.380 175.405 ;
        RECT 41.550 175.075 42.260 175.525 ;
        RECT 43.005 175.405 43.175 175.575 ;
        RECT 42.430 175.075 42.835 175.405 ;
        RECT 43.005 175.075 43.275 175.405 ;
        RECT 43.005 174.905 43.175 175.075 ;
        RECT 41.565 174.735 43.175 174.905 ;
        RECT 43.445 174.840 43.615 175.575 ;
        RECT 44.245 175.550 44.535 176.715 ;
        RECT 41.035 174.165 41.365 174.665 ;
        RECT 41.565 174.385 41.735 174.735 ;
        RECT 41.935 174.165 42.265 174.565 ;
        RECT 42.435 174.385 42.605 174.735 ;
        RECT 42.775 174.165 43.155 174.565 ;
        RECT 43.345 174.495 43.615 174.840 ;
        RECT 44.245 174.165 44.535 174.890 ;
        RECT 44.705 174.445 44.985 176.545 ;
        RECT 45.175 175.955 45.960 176.715 ;
        RECT 46.355 175.885 46.740 176.545 ;
        RECT 46.355 175.785 46.765 175.885 ;
        RECT 45.155 175.575 46.765 175.785 ;
        RECT 47.065 175.695 47.265 176.485 ;
        RECT 45.155 174.975 45.430 175.575 ;
        RECT 46.935 175.525 47.265 175.695 ;
        RECT 47.435 175.535 47.755 176.715 ;
        RECT 48.385 175.575 48.645 176.715 ;
        RECT 48.815 175.565 49.145 176.545 ;
        RECT 49.315 175.575 49.595 176.715 ;
        RECT 49.765 175.845 50.040 176.545 ;
        RECT 50.210 176.170 50.465 176.715 ;
        RECT 50.635 176.205 51.115 176.545 ;
        RECT 51.290 176.160 51.895 176.715 ;
        RECT 51.280 176.060 51.895 176.160 ;
        RECT 51.280 176.035 51.465 176.060 ;
        RECT 46.935 175.405 47.115 175.525 ;
        RECT 45.600 175.155 45.955 175.405 ;
        RECT 46.150 175.355 46.615 175.405 ;
        RECT 46.145 175.185 46.615 175.355 ;
        RECT 46.150 175.155 46.615 175.185 ;
        RECT 46.785 175.155 47.115 175.405 ;
        RECT 47.290 175.155 47.755 175.355 ;
        RECT 48.405 175.155 48.740 175.405 ;
        RECT 45.155 174.795 46.405 174.975 ;
        RECT 48.910 174.965 49.080 175.565 ;
        RECT 49.250 175.135 49.585 175.405 ;
        RECT 46.040 174.725 46.405 174.795 ;
        RECT 46.575 174.775 47.755 174.945 ;
        RECT 45.215 174.165 45.385 174.625 ;
        RECT 46.575 174.555 46.905 174.775 ;
        RECT 45.655 174.375 46.905 174.555 ;
        RECT 47.075 174.165 47.245 174.605 ;
        RECT 47.415 174.360 47.755 174.775 ;
        RECT 48.385 174.335 49.080 174.965 ;
        RECT 49.285 174.165 49.595 174.965 ;
        RECT 49.765 174.815 49.935 175.845 ;
        RECT 50.210 175.715 50.965 175.965 ;
        RECT 51.135 175.790 51.465 176.035 ;
        RECT 52.070 175.915 52.385 176.715 ;
        RECT 52.650 176.360 53.730 176.530 ;
        RECT 50.210 175.680 50.980 175.715 ;
        RECT 50.210 175.670 50.995 175.680 ;
        RECT 50.105 175.655 51.000 175.670 ;
        RECT 50.105 175.640 51.020 175.655 ;
        RECT 50.105 175.630 51.040 175.640 ;
        RECT 50.105 175.620 51.065 175.630 ;
        RECT 50.105 175.590 51.135 175.620 ;
        RECT 50.105 175.560 51.155 175.590 ;
        RECT 50.105 175.530 51.175 175.560 ;
        RECT 50.105 175.505 51.205 175.530 ;
        RECT 50.105 175.470 51.240 175.505 ;
        RECT 50.105 175.465 51.270 175.470 ;
        RECT 50.105 175.070 50.335 175.465 ;
        RECT 50.880 175.460 51.270 175.465 ;
        RECT 50.905 175.450 51.270 175.460 ;
        RECT 50.920 175.445 51.270 175.450 ;
        RECT 50.935 175.440 51.270 175.445 ;
        RECT 51.635 175.440 51.895 175.890 ;
        RECT 52.650 175.745 52.820 176.360 ;
        RECT 50.935 175.435 51.895 175.440 ;
        RECT 50.945 175.425 51.895 175.435 ;
        RECT 50.955 175.420 51.895 175.425 ;
        RECT 50.965 175.410 51.895 175.420 ;
        RECT 50.970 175.400 51.895 175.410 ;
        RECT 50.975 175.395 51.895 175.400 ;
        RECT 50.985 175.380 51.895 175.395 ;
        RECT 50.990 175.365 51.895 175.380 ;
        RECT 51.000 175.340 51.895 175.365 ;
        RECT 50.505 174.870 50.835 175.295 ;
        RECT 49.765 174.335 50.025 174.815 ;
        RECT 50.195 174.165 50.445 174.705 ;
        RECT 50.615 174.385 50.835 174.870 ;
        RECT 51.005 175.270 51.895 175.340 ;
        RECT 51.005 174.545 51.175 175.270 ;
        RECT 51.345 174.715 51.895 175.100 ;
        RECT 52.065 174.735 52.335 175.745 ;
        RECT 52.505 175.575 52.820 175.745 ;
        RECT 52.505 174.905 52.675 175.575 ;
        RECT 52.990 175.405 53.225 176.085 ;
        RECT 53.395 175.575 53.730 176.360 ;
        RECT 54.825 175.575 55.165 176.545 ;
        RECT 55.335 175.575 55.505 176.715 ;
        RECT 55.775 175.915 56.025 176.715 ;
        RECT 56.670 175.745 57.000 176.545 ;
        RECT 57.300 175.915 57.630 176.715 ;
        RECT 57.800 175.745 58.130 176.545 ;
        RECT 55.695 175.575 58.130 175.745 ;
        RECT 58.505 175.625 62.015 176.715 ;
        RECT 52.845 175.075 53.225 175.405 ;
        RECT 53.395 175.075 53.730 175.405 ;
        RECT 54.825 174.965 55.000 175.575 ;
        RECT 55.695 175.325 55.865 175.575 ;
        RECT 55.170 175.155 55.865 175.325 ;
        RECT 56.040 175.155 56.460 175.355 ;
        RECT 56.630 175.155 56.960 175.355 ;
        RECT 57.130 175.155 57.460 175.355 ;
        RECT 52.505 174.735 53.730 174.905 ;
        RECT 51.005 174.375 51.895 174.545 ;
        RECT 52.135 174.165 52.465 174.565 ;
        RECT 52.635 174.465 52.805 174.735 ;
        RECT 52.975 174.165 53.305 174.565 ;
        RECT 53.475 174.465 53.730 174.735 ;
        RECT 54.825 174.335 55.165 174.965 ;
        RECT 55.335 174.165 55.585 174.965 ;
        RECT 55.775 174.815 57.000 174.985 ;
        RECT 55.775 174.335 56.105 174.815 ;
        RECT 56.275 174.165 56.500 174.625 ;
        RECT 56.670 174.335 57.000 174.815 ;
        RECT 57.630 174.945 57.800 175.575 ;
        RECT 57.985 175.155 58.335 175.405 ;
        RECT 57.630 174.335 58.130 174.945 ;
        RECT 58.505 174.935 60.155 175.455 ;
        RECT 60.325 175.105 62.015 175.625 ;
        RECT 62.195 175.575 62.525 176.715 ;
        RECT 63.055 175.745 63.385 176.530 ;
        RECT 62.705 175.575 63.385 175.745 ;
        RECT 63.575 175.745 63.905 176.530 ;
        RECT 63.575 175.575 64.255 175.745 ;
        RECT 64.435 175.575 64.765 176.715 ;
        RECT 64.945 175.625 68.455 176.715 ;
        RECT 68.625 175.625 69.835 176.715 ;
        RECT 62.185 175.155 62.535 175.405 ;
        RECT 62.705 174.975 62.875 175.575 ;
        RECT 63.045 175.155 63.395 175.405 ;
        RECT 63.565 175.155 63.915 175.405 ;
        RECT 64.085 174.975 64.255 175.575 ;
        RECT 64.425 175.155 64.775 175.405 ;
        RECT 58.505 174.165 62.015 174.935 ;
        RECT 62.195 174.165 62.465 174.975 ;
        RECT 62.635 174.335 62.965 174.975 ;
        RECT 63.135 174.165 63.375 174.975 ;
        RECT 63.585 174.165 63.825 174.975 ;
        RECT 63.995 174.335 64.325 174.975 ;
        RECT 64.495 174.165 64.765 174.975 ;
        RECT 64.945 174.935 66.595 175.455 ;
        RECT 66.765 175.105 68.455 175.625 ;
        RECT 64.945 174.165 68.455 174.935 ;
        RECT 68.625 174.915 69.145 175.455 ;
        RECT 69.315 175.085 69.835 175.625 ;
        RECT 70.005 175.550 70.295 176.715 ;
        RECT 70.465 176.280 75.810 176.715 ;
        RECT 75.985 176.280 81.330 176.715 ;
        RECT 68.625 174.165 69.835 174.915 ;
        RECT 70.005 174.165 70.295 174.890 ;
        RECT 72.050 174.710 72.390 175.540 ;
        RECT 73.870 175.030 74.220 176.280 ;
        RECT 77.570 174.710 77.910 175.540 ;
        RECT 79.390 175.030 79.740 176.280 ;
        RECT 81.505 175.625 82.715 176.715 ;
        RECT 81.505 174.915 82.025 175.455 ;
        RECT 82.195 175.085 82.715 175.625 ;
        RECT 82.885 175.625 84.095 176.715 ;
        RECT 82.885 175.085 83.405 175.625 ;
        RECT 83.575 174.915 84.095 175.455 ;
        RECT 70.465 174.165 75.810 174.710 ;
        RECT 75.985 174.165 81.330 174.710 ;
        RECT 81.505 174.165 82.715 174.915 ;
        RECT 82.885 174.165 84.095 174.915 ;
        RECT 5.520 173.995 84.180 174.165 ;
        RECT 5.605 173.245 6.815 173.995 ;
        RECT 6.985 173.450 12.330 173.995 ;
        RECT 12.970 173.490 13.305 173.995 ;
        RECT 5.605 172.705 6.125 173.245 ;
        RECT 6.295 172.535 6.815 173.075 ;
        RECT 8.570 172.620 8.910 173.450 ;
        RECT 13.475 173.425 13.715 173.800 ;
        RECT 13.995 173.665 14.165 173.810 ;
        RECT 13.995 173.470 14.370 173.665 ;
        RECT 14.730 173.500 15.125 173.995 ;
        RECT 5.605 171.445 6.815 172.535 ;
        RECT 10.390 171.880 10.740 173.130 ;
        RECT 13.025 172.465 13.325 173.315 ;
        RECT 13.495 173.275 13.715 173.425 ;
        RECT 13.495 172.945 14.030 173.275 ;
        RECT 14.200 173.135 14.370 173.470 ;
        RECT 15.295 173.305 15.535 173.825 ;
        RECT 15.725 173.450 21.070 173.995 ;
        RECT 21.245 173.450 26.590 173.995 ;
        RECT 13.495 172.295 13.730 172.945 ;
        RECT 14.200 172.775 15.185 173.135 ;
        RECT 13.055 172.065 13.730 172.295 ;
        RECT 13.900 172.755 15.185 172.775 ;
        RECT 13.900 172.605 14.760 172.755 ;
        RECT 6.985 171.445 12.330 171.880 ;
        RECT 13.055 171.635 13.225 172.065 ;
        RECT 13.395 171.445 13.725 171.895 ;
        RECT 13.900 171.660 14.185 172.605 ;
        RECT 15.360 172.500 15.535 173.305 ;
        RECT 17.310 172.620 17.650 173.450 ;
        RECT 14.360 172.125 15.055 172.435 ;
        RECT 14.365 171.445 15.050 171.915 ;
        RECT 15.230 171.715 15.535 172.500 ;
        RECT 19.130 171.880 19.480 173.130 ;
        RECT 22.830 172.620 23.170 173.450 ;
        RECT 26.765 173.225 30.275 173.995 ;
        RECT 31.365 173.270 31.655 173.995 ;
        RECT 31.825 173.225 35.335 173.995 ;
        RECT 35.505 173.245 36.715 173.995 ;
        RECT 24.650 171.880 25.000 173.130 ;
        RECT 26.765 172.705 28.415 173.225 ;
        RECT 28.585 172.535 30.275 173.055 ;
        RECT 31.825 172.705 33.475 173.225 ;
        RECT 15.725 171.445 21.070 171.880 ;
        RECT 21.245 171.445 26.590 171.880 ;
        RECT 26.765 171.445 30.275 172.535 ;
        RECT 31.365 171.445 31.655 172.610 ;
        RECT 33.645 172.535 35.335 173.055 ;
        RECT 35.505 172.705 36.025 173.245 ;
        RECT 36.905 173.185 37.145 173.995 ;
        RECT 37.315 173.185 37.645 173.825 ;
        RECT 37.815 173.185 38.085 173.995 ;
        RECT 38.265 173.450 43.610 173.995 ;
        RECT 43.785 173.450 49.130 173.995 ;
        RECT 49.305 173.450 54.650 173.995 ;
        RECT 36.195 172.535 36.715 173.075 ;
        RECT 36.885 172.755 37.235 173.005 ;
        RECT 37.405 172.585 37.575 173.185 ;
        RECT 37.745 172.755 38.095 173.005 ;
        RECT 39.850 172.620 40.190 173.450 ;
        RECT 31.825 171.445 35.335 172.535 ;
        RECT 35.505 171.445 36.715 172.535 ;
        RECT 36.895 172.415 37.575 172.585 ;
        RECT 36.895 171.630 37.225 172.415 ;
        RECT 37.755 171.445 38.085 172.585 ;
        RECT 41.670 171.880 42.020 173.130 ;
        RECT 45.370 172.620 45.710 173.450 ;
        RECT 47.190 171.880 47.540 173.130 ;
        RECT 50.890 172.620 51.230 173.450 ;
        RECT 54.825 173.225 56.495 173.995 ;
        RECT 57.125 173.270 57.415 173.995 ;
        RECT 57.585 173.225 60.175 173.995 ;
        RECT 52.710 171.880 53.060 173.130 ;
        RECT 54.825 172.705 55.575 173.225 ;
        RECT 55.745 172.535 56.495 173.055 ;
        RECT 57.585 172.705 58.795 173.225 ;
        RECT 60.405 173.175 60.615 173.995 ;
        RECT 60.785 173.195 61.115 173.825 ;
        RECT 38.265 171.445 43.610 171.880 ;
        RECT 43.785 171.445 49.130 171.880 ;
        RECT 49.305 171.445 54.650 171.880 ;
        RECT 54.825 171.445 56.495 172.535 ;
        RECT 57.125 171.445 57.415 172.610 ;
        RECT 58.965 172.535 60.175 173.055 ;
        RECT 60.785 172.595 61.035 173.195 ;
        RECT 61.285 173.175 61.515 173.995 ;
        RECT 62.665 173.185 62.905 173.995 ;
        RECT 63.075 173.185 63.405 173.825 ;
        RECT 63.575 173.185 63.845 173.995 ;
        RECT 64.035 173.185 64.305 173.995 ;
        RECT 64.475 173.185 64.805 173.825 ;
        RECT 64.975 173.185 65.215 173.995 ;
        RECT 65.405 173.195 66.100 173.825 ;
        RECT 66.305 173.195 66.615 173.995 ;
        RECT 66.785 173.450 72.130 173.995 ;
        RECT 72.305 173.450 77.650 173.995 ;
        RECT 61.205 172.755 61.535 173.005 ;
        RECT 62.645 172.755 62.995 173.005 ;
        RECT 57.585 171.445 60.175 172.535 ;
        RECT 60.405 171.445 60.615 172.585 ;
        RECT 60.785 171.615 61.115 172.595 ;
        RECT 63.165 172.585 63.335 173.185 ;
        RECT 63.505 172.755 63.855 173.005 ;
        RECT 64.025 172.755 64.375 173.005 ;
        RECT 64.545 172.585 64.715 173.185 ;
        RECT 65.925 173.145 66.100 173.195 ;
        RECT 64.885 172.755 65.235 173.005 ;
        RECT 65.425 172.755 65.760 173.005 ;
        RECT 65.930 172.595 66.100 173.145 ;
        RECT 66.270 172.755 66.605 173.025 ;
        RECT 68.370 172.620 68.710 173.450 ;
        RECT 61.285 171.445 61.515 172.585 ;
        RECT 62.655 172.415 63.335 172.585 ;
        RECT 62.655 171.630 62.985 172.415 ;
        RECT 63.515 171.445 63.845 172.585 ;
        RECT 64.035 171.445 64.365 172.585 ;
        RECT 64.545 172.415 65.225 172.585 ;
        RECT 64.895 171.630 65.225 172.415 ;
        RECT 65.405 171.445 65.665 172.585 ;
        RECT 65.835 171.615 66.165 172.595 ;
        RECT 66.335 171.445 66.615 172.585 ;
        RECT 70.190 171.880 70.540 173.130 ;
        RECT 73.890 172.620 74.230 173.450 ;
        RECT 77.825 173.225 81.335 173.995 ;
        RECT 81.505 173.245 82.715 173.995 ;
        RECT 82.885 173.245 84.095 173.995 ;
        RECT 75.710 171.880 76.060 173.130 ;
        RECT 77.825 172.705 79.475 173.225 ;
        RECT 79.645 172.535 81.335 173.055 ;
        RECT 81.505 172.705 82.025 173.245 ;
        RECT 82.195 172.535 82.715 173.075 ;
        RECT 66.785 171.445 72.130 171.880 ;
        RECT 72.305 171.445 77.650 171.880 ;
        RECT 77.825 171.445 81.335 172.535 ;
        RECT 81.505 171.445 82.715 172.535 ;
        RECT 82.885 172.535 83.405 173.075 ;
        RECT 83.575 172.705 84.095 173.245 ;
        RECT 82.885 171.445 84.095 172.535 ;
        RECT 5.520 171.275 84.180 171.445 ;
        RECT 5.605 170.185 6.815 171.275 ;
        RECT 6.985 170.840 12.330 171.275 ;
        RECT 12.505 170.840 17.850 171.275 ;
        RECT 5.605 169.475 6.125 170.015 ;
        RECT 6.295 169.645 6.815 170.185 ;
        RECT 5.605 168.725 6.815 169.475 ;
        RECT 8.570 169.270 8.910 170.100 ;
        RECT 10.390 169.590 10.740 170.840 ;
        RECT 14.090 169.270 14.430 170.100 ;
        RECT 15.910 169.590 16.260 170.840 ;
        RECT 18.485 170.110 18.775 171.275 ;
        RECT 18.945 170.185 21.535 171.275 ;
        RECT 22.165 170.720 22.770 171.275 ;
        RECT 22.945 170.765 23.425 171.105 ;
        RECT 23.595 170.730 23.850 171.275 ;
        RECT 22.165 170.620 22.780 170.720 ;
        RECT 22.595 170.595 22.780 170.620 ;
        RECT 18.945 169.495 20.155 170.015 ;
        RECT 20.325 169.665 21.535 170.185 ;
        RECT 22.165 170.000 22.425 170.450 ;
        RECT 22.595 170.350 22.925 170.595 ;
        RECT 23.095 170.275 23.850 170.525 ;
        RECT 24.020 170.405 24.295 171.105 ;
        RECT 23.080 170.240 23.850 170.275 ;
        RECT 23.065 170.230 23.850 170.240 ;
        RECT 23.060 170.215 23.955 170.230 ;
        RECT 23.040 170.200 23.955 170.215 ;
        RECT 23.020 170.190 23.955 170.200 ;
        RECT 22.995 170.180 23.955 170.190 ;
        RECT 22.925 170.150 23.955 170.180 ;
        RECT 22.905 170.120 23.955 170.150 ;
        RECT 22.885 170.090 23.955 170.120 ;
        RECT 22.855 170.065 23.955 170.090 ;
        RECT 22.820 170.030 23.955 170.065 ;
        RECT 22.790 170.025 23.955 170.030 ;
        RECT 22.790 170.020 23.180 170.025 ;
        RECT 22.790 170.010 23.155 170.020 ;
        RECT 22.790 170.005 23.140 170.010 ;
        RECT 22.790 170.000 23.125 170.005 ;
        RECT 22.165 169.995 23.125 170.000 ;
        RECT 22.165 169.985 23.115 169.995 ;
        RECT 22.165 169.980 23.105 169.985 ;
        RECT 22.165 169.970 23.095 169.980 ;
        RECT 22.165 169.960 23.090 169.970 ;
        RECT 22.165 169.955 23.085 169.960 ;
        RECT 22.165 169.940 23.075 169.955 ;
        RECT 22.165 169.925 23.070 169.940 ;
        RECT 22.165 169.900 23.060 169.925 ;
        RECT 22.165 169.830 23.055 169.900 ;
        RECT 6.985 168.725 12.330 169.270 ;
        RECT 12.505 168.725 17.850 169.270 ;
        RECT 18.485 168.725 18.775 169.450 ;
        RECT 18.945 168.725 21.535 169.495 ;
        RECT 22.165 169.275 22.715 169.660 ;
        RECT 22.885 169.105 23.055 169.830 ;
        RECT 22.165 168.935 23.055 169.105 ;
        RECT 23.225 169.430 23.555 169.855 ;
        RECT 23.725 169.630 23.955 170.025 ;
        RECT 23.225 168.945 23.445 169.430 ;
        RECT 24.125 169.375 24.295 170.405 ;
        RECT 23.615 168.725 23.865 169.265 ;
        RECT 24.035 168.895 24.295 169.375 ;
        RECT 24.465 170.405 24.740 171.105 ;
        RECT 24.910 170.730 25.165 171.275 ;
        RECT 25.335 170.765 25.815 171.105 ;
        RECT 25.990 170.720 26.595 171.275 ;
        RECT 25.980 170.620 26.595 170.720 ;
        RECT 25.980 170.595 26.165 170.620 ;
        RECT 24.465 169.375 24.635 170.405 ;
        RECT 24.910 170.275 25.665 170.525 ;
        RECT 25.835 170.350 26.165 170.595 ;
        RECT 24.910 170.240 25.680 170.275 ;
        RECT 24.910 170.230 25.695 170.240 ;
        RECT 24.805 170.215 25.700 170.230 ;
        RECT 24.805 170.200 25.720 170.215 ;
        RECT 24.805 170.190 25.740 170.200 ;
        RECT 24.805 170.180 25.765 170.190 ;
        RECT 24.805 170.150 25.835 170.180 ;
        RECT 24.805 170.120 25.855 170.150 ;
        RECT 24.805 170.090 25.875 170.120 ;
        RECT 24.805 170.065 25.905 170.090 ;
        RECT 24.805 170.030 25.940 170.065 ;
        RECT 24.805 170.025 25.970 170.030 ;
        RECT 24.805 169.630 25.035 170.025 ;
        RECT 25.580 170.020 25.970 170.025 ;
        RECT 25.605 170.010 25.970 170.020 ;
        RECT 25.620 170.005 25.970 170.010 ;
        RECT 25.635 170.000 25.970 170.005 ;
        RECT 26.335 170.000 26.595 170.450 ;
        RECT 26.765 170.185 29.355 171.275 ;
        RECT 30.235 170.545 30.530 171.275 ;
        RECT 30.700 170.375 30.960 171.100 ;
        RECT 31.130 170.545 31.390 171.275 ;
        RECT 31.560 170.375 31.820 171.100 ;
        RECT 31.990 170.545 32.250 171.275 ;
        RECT 32.420 170.375 32.680 171.100 ;
        RECT 32.850 170.545 33.110 171.275 ;
        RECT 33.280 170.375 33.540 171.100 ;
        RECT 25.635 169.995 26.595 170.000 ;
        RECT 25.645 169.985 26.595 169.995 ;
        RECT 25.655 169.980 26.595 169.985 ;
        RECT 25.665 169.970 26.595 169.980 ;
        RECT 25.670 169.960 26.595 169.970 ;
        RECT 25.675 169.955 26.595 169.960 ;
        RECT 25.685 169.940 26.595 169.955 ;
        RECT 25.690 169.925 26.595 169.940 ;
        RECT 25.700 169.900 26.595 169.925 ;
        RECT 25.205 169.430 25.535 169.855 ;
        RECT 25.285 169.405 25.535 169.430 ;
        RECT 24.465 168.895 24.725 169.375 ;
        RECT 24.895 168.725 25.145 169.265 ;
        RECT 25.315 168.945 25.535 169.405 ;
        RECT 25.705 169.830 26.595 169.900 ;
        RECT 25.705 169.105 25.875 169.830 ;
        RECT 26.045 169.275 26.595 169.660 ;
        RECT 26.765 169.495 27.975 170.015 ;
        RECT 28.145 169.665 29.355 170.185 ;
        RECT 30.230 170.135 33.540 170.375 ;
        RECT 33.710 170.165 33.970 171.275 ;
        RECT 30.230 169.545 31.200 170.135 ;
        RECT 34.140 169.965 34.390 171.100 ;
        RECT 34.570 170.165 34.865 171.275 ;
        RECT 35.045 170.405 35.320 171.105 ;
        RECT 35.490 170.730 35.745 171.275 ;
        RECT 35.915 170.765 36.395 171.105 ;
        RECT 36.570 170.720 37.175 171.275 ;
        RECT 36.560 170.620 37.175 170.720 ;
        RECT 36.560 170.595 36.745 170.620 ;
        RECT 31.370 169.715 34.390 169.965 ;
        RECT 25.705 168.935 26.595 169.105 ;
        RECT 26.765 168.725 29.355 169.495 ;
        RECT 30.230 169.375 33.540 169.545 ;
        RECT 30.230 168.725 30.530 169.205 ;
        RECT 30.700 168.920 30.960 169.375 ;
        RECT 31.130 168.725 31.390 169.205 ;
        RECT 31.560 168.920 31.820 169.375 ;
        RECT 31.990 168.725 32.250 169.205 ;
        RECT 32.420 168.920 32.680 169.375 ;
        RECT 32.850 168.725 33.110 169.205 ;
        RECT 33.280 168.920 33.540 169.375 ;
        RECT 33.710 168.725 33.970 169.250 ;
        RECT 34.140 168.905 34.390 169.715 ;
        RECT 34.560 169.355 34.875 169.965 ;
        RECT 35.045 169.375 35.215 170.405 ;
        RECT 35.490 170.275 36.245 170.525 ;
        RECT 36.415 170.350 36.745 170.595 ;
        RECT 35.490 170.240 36.260 170.275 ;
        RECT 35.490 170.230 36.275 170.240 ;
        RECT 35.385 170.215 36.280 170.230 ;
        RECT 35.385 170.200 36.300 170.215 ;
        RECT 35.385 170.190 36.320 170.200 ;
        RECT 35.385 170.180 36.345 170.190 ;
        RECT 35.385 170.150 36.415 170.180 ;
        RECT 35.385 170.120 36.435 170.150 ;
        RECT 35.385 170.090 36.455 170.120 ;
        RECT 35.385 170.065 36.485 170.090 ;
        RECT 35.385 170.030 36.520 170.065 ;
        RECT 35.385 170.025 36.550 170.030 ;
        RECT 35.385 169.630 35.615 170.025 ;
        RECT 36.160 170.020 36.550 170.025 ;
        RECT 36.185 170.010 36.550 170.020 ;
        RECT 36.200 170.005 36.550 170.010 ;
        RECT 36.215 170.000 36.550 170.005 ;
        RECT 36.915 170.000 37.175 170.450 ;
        RECT 36.215 169.995 37.175 170.000 ;
        RECT 36.225 169.985 37.175 169.995 ;
        RECT 36.235 169.980 37.175 169.985 ;
        RECT 36.245 169.970 37.175 169.980 ;
        RECT 36.250 169.960 37.175 169.970 ;
        RECT 36.255 169.955 37.175 169.960 ;
        RECT 36.265 169.940 37.175 169.955 ;
        RECT 36.270 169.925 37.175 169.940 ;
        RECT 36.280 169.900 37.175 169.925 ;
        RECT 35.785 169.430 36.115 169.855 ;
        RECT 34.570 168.725 34.815 169.185 ;
        RECT 35.045 168.895 35.305 169.375 ;
        RECT 35.475 168.725 35.725 169.265 ;
        RECT 35.895 168.945 36.115 169.430 ;
        RECT 36.285 169.830 37.175 169.900 ;
        RECT 37.345 170.405 37.620 171.105 ;
        RECT 37.790 170.730 38.045 171.275 ;
        RECT 38.215 170.765 38.695 171.105 ;
        RECT 38.870 170.720 39.475 171.275 ;
        RECT 38.860 170.620 39.475 170.720 ;
        RECT 39.655 170.665 39.985 171.095 ;
        RECT 40.165 170.835 40.360 171.275 ;
        RECT 40.530 170.665 40.860 171.095 ;
        RECT 38.860 170.595 39.045 170.620 ;
        RECT 36.285 169.105 36.455 169.830 ;
        RECT 36.625 169.275 37.175 169.660 ;
        RECT 37.345 169.375 37.515 170.405 ;
        RECT 37.790 170.275 38.545 170.525 ;
        RECT 38.715 170.350 39.045 170.595 ;
        RECT 39.655 170.495 40.860 170.665 ;
        RECT 37.790 170.240 38.560 170.275 ;
        RECT 37.790 170.230 38.575 170.240 ;
        RECT 37.685 170.215 38.580 170.230 ;
        RECT 37.685 170.200 38.600 170.215 ;
        RECT 37.685 170.190 38.620 170.200 ;
        RECT 37.685 170.180 38.645 170.190 ;
        RECT 37.685 170.150 38.715 170.180 ;
        RECT 37.685 170.120 38.735 170.150 ;
        RECT 37.685 170.090 38.755 170.120 ;
        RECT 37.685 170.065 38.785 170.090 ;
        RECT 37.685 170.030 38.820 170.065 ;
        RECT 37.685 170.025 38.850 170.030 ;
        RECT 37.685 169.630 37.915 170.025 ;
        RECT 38.460 170.020 38.850 170.025 ;
        RECT 38.485 170.010 38.850 170.020 ;
        RECT 38.500 170.005 38.850 170.010 ;
        RECT 38.515 170.000 38.850 170.005 ;
        RECT 39.215 170.000 39.475 170.450 ;
        RECT 39.655 170.165 40.550 170.495 ;
        RECT 41.030 170.325 41.305 171.095 ;
        RECT 38.515 169.995 39.475 170.000 ;
        RECT 38.525 169.985 39.475 169.995 ;
        RECT 38.535 169.980 39.475 169.985 ;
        RECT 38.545 169.970 39.475 169.980 ;
        RECT 38.550 169.960 39.475 169.970 ;
        RECT 40.720 170.135 41.305 170.325 ;
        RECT 41.485 170.185 44.075 171.275 ;
        RECT 38.555 169.955 39.475 169.960 ;
        RECT 38.565 169.940 39.475 169.955 ;
        RECT 38.570 169.925 39.475 169.940 ;
        RECT 38.580 169.900 39.475 169.925 ;
        RECT 38.085 169.430 38.415 169.855 ;
        RECT 36.285 168.935 37.175 169.105 ;
        RECT 37.345 168.895 37.605 169.375 ;
        RECT 37.775 168.725 38.025 169.265 ;
        RECT 38.195 168.945 38.415 169.430 ;
        RECT 38.585 169.830 39.475 169.900 ;
        RECT 38.585 169.105 38.755 169.830 ;
        RECT 38.925 169.275 39.475 169.660 ;
        RECT 39.660 169.635 39.955 169.965 ;
        RECT 40.135 169.635 40.550 169.965 ;
        RECT 38.585 168.935 39.475 169.105 ;
        RECT 39.655 168.725 39.955 169.455 ;
        RECT 40.135 169.015 40.365 169.635 ;
        RECT 40.720 169.465 40.895 170.135 ;
        RECT 40.565 169.285 40.895 169.465 ;
        RECT 41.065 169.315 41.305 169.965 ;
        RECT 41.485 169.495 42.695 170.015 ;
        RECT 42.865 169.665 44.075 170.185 ;
        RECT 44.245 170.110 44.535 171.275 ;
        RECT 44.705 170.305 44.975 171.075 ;
        RECT 45.145 170.495 45.475 171.275 ;
        RECT 45.680 170.670 45.865 171.075 ;
        RECT 46.035 170.850 46.370 171.275 ;
        RECT 46.550 170.850 46.885 171.275 ;
        RECT 47.055 170.670 47.240 171.075 ;
        RECT 45.680 170.495 46.345 170.670 ;
        RECT 44.705 170.135 45.835 170.305 ;
        RECT 40.565 168.905 40.790 169.285 ;
        RECT 40.960 168.725 41.290 169.115 ;
        RECT 41.485 168.725 44.075 169.495 ;
        RECT 44.245 168.725 44.535 169.450 ;
        RECT 44.705 169.225 44.875 170.135 ;
        RECT 45.045 169.385 45.405 169.965 ;
        RECT 45.585 169.635 45.835 170.135 ;
        RECT 46.005 169.465 46.345 170.495 ;
        RECT 45.660 169.295 46.345 169.465 ;
        RECT 46.575 170.495 47.240 170.670 ;
        RECT 47.445 170.495 47.775 171.275 ;
        RECT 46.575 169.465 46.915 170.495 ;
        RECT 47.945 170.305 48.215 171.075 ;
        RECT 47.085 170.135 48.215 170.305 ;
        RECT 48.385 170.185 49.595 171.275 ;
        RECT 47.085 169.635 47.335 170.135 ;
        RECT 46.575 169.295 47.260 169.465 ;
        RECT 47.515 169.385 47.875 169.965 ;
        RECT 44.705 168.895 44.965 169.225 ;
        RECT 45.175 168.725 45.450 169.205 ;
        RECT 45.660 168.895 45.865 169.295 ;
        RECT 46.035 168.725 46.370 169.125 ;
        RECT 46.550 168.725 46.885 169.125 ;
        RECT 47.055 168.895 47.260 169.295 ;
        RECT 48.045 169.225 48.215 170.135 ;
        RECT 47.470 168.725 47.745 169.205 ;
        RECT 47.955 168.895 48.215 169.225 ;
        RECT 48.385 169.475 48.905 170.015 ;
        RECT 49.075 169.645 49.595 170.185 ;
        RECT 49.775 170.135 50.105 171.275 ;
        RECT 50.635 170.305 50.965 171.090 ;
        RECT 50.285 170.135 50.965 170.305 ;
        RECT 51.145 170.425 51.405 171.105 ;
        RECT 51.575 170.495 51.825 171.275 ;
        RECT 52.075 170.725 52.325 171.105 ;
        RECT 52.495 170.895 52.850 171.275 ;
        RECT 53.855 170.885 54.190 171.105 ;
        RECT 53.455 170.725 53.685 170.765 ;
        RECT 52.075 170.525 53.685 170.725 ;
        RECT 52.075 170.515 52.910 170.525 ;
        RECT 53.500 170.435 53.685 170.525 ;
        RECT 49.765 169.715 50.115 169.965 ;
        RECT 50.285 169.535 50.455 170.135 ;
        RECT 50.625 169.715 50.975 169.965 ;
        RECT 48.385 168.725 49.595 169.475 ;
        RECT 49.775 168.725 50.045 169.535 ;
        RECT 50.215 168.895 50.545 169.535 ;
        RECT 50.715 168.725 50.955 169.535 ;
        RECT 51.145 169.225 51.315 170.425 ;
        RECT 53.015 170.325 53.345 170.355 ;
        RECT 51.545 170.265 53.345 170.325 ;
        RECT 53.935 170.265 54.190 170.885 ;
        RECT 54.865 170.815 55.080 171.275 ;
        RECT 55.250 170.645 55.580 171.105 ;
        RECT 51.485 170.155 54.190 170.265 ;
        RECT 51.485 170.120 51.685 170.155 ;
        RECT 51.485 169.545 51.655 170.120 ;
        RECT 53.015 170.095 54.190 170.155 ;
        RECT 54.410 170.475 55.580 170.645 ;
        RECT 55.750 170.475 56.000 171.275 ;
        RECT 51.885 169.680 52.295 169.985 ;
        RECT 52.465 169.715 52.795 169.925 ;
        RECT 51.485 169.425 51.755 169.545 ;
        RECT 51.485 169.380 52.330 169.425 ;
        RECT 51.575 169.255 52.330 169.380 ;
        RECT 52.585 169.315 52.795 169.715 ;
        RECT 53.040 169.715 53.515 169.925 ;
        RECT 53.705 169.715 54.195 169.915 ;
        RECT 53.040 169.315 53.260 169.715 ;
        RECT 51.145 168.895 51.405 169.225 ;
        RECT 52.160 169.105 52.330 169.255 ;
        RECT 51.575 168.725 51.905 169.085 ;
        RECT 52.160 168.895 53.460 169.105 ;
        RECT 53.735 168.725 54.190 169.490 ;
        RECT 54.410 169.185 54.780 170.475 ;
        RECT 56.210 170.305 56.490 170.465 ;
        RECT 55.155 170.135 56.490 170.305 ;
        RECT 56.665 170.185 58.335 171.275 ;
        RECT 55.155 169.965 55.325 170.135 ;
        RECT 54.950 169.715 55.325 169.965 ;
        RECT 55.495 169.715 55.970 169.955 ;
        RECT 56.140 169.715 56.490 169.955 ;
        RECT 55.155 169.545 55.325 169.715 ;
        RECT 55.155 169.375 56.490 169.545 ;
        RECT 54.410 168.895 55.160 169.185 ;
        RECT 55.670 168.725 56.000 169.185 ;
        RECT 56.220 169.165 56.490 169.375 ;
        RECT 56.665 169.495 57.415 170.015 ;
        RECT 57.585 169.665 58.335 170.185 ;
        RECT 58.965 170.845 59.305 171.105 ;
        RECT 56.665 168.725 58.335 169.495 ;
        RECT 58.965 169.445 59.225 170.845 ;
        RECT 59.475 170.475 59.805 171.275 ;
        RECT 60.270 170.305 60.520 171.105 ;
        RECT 60.705 170.555 61.035 171.275 ;
        RECT 61.255 170.305 61.505 171.105 ;
        RECT 61.675 170.895 62.010 171.275 ;
        RECT 59.415 170.135 61.605 170.305 ;
        RECT 59.415 169.965 59.730 170.135 ;
        RECT 59.400 169.715 59.730 169.965 ;
        RECT 58.965 168.935 59.305 169.445 ;
        RECT 59.475 168.725 59.745 169.525 ;
        RECT 59.925 168.995 60.205 169.965 ;
        RECT 60.385 168.995 60.685 169.965 ;
        RECT 60.865 169.000 61.215 169.965 ;
        RECT 61.435 169.225 61.605 170.135 ;
        RECT 61.775 169.405 62.015 170.715 ;
        RECT 62.185 170.555 62.645 171.105 ;
        RECT 62.835 170.555 63.165 171.275 ;
        RECT 61.435 168.895 61.930 169.225 ;
        RECT 62.185 169.185 62.435 170.555 ;
        RECT 63.365 170.385 63.665 170.935 ;
        RECT 63.835 170.605 64.115 171.275 ;
        RECT 64.490 170.895 64.825 171.275 ;
        RECT 62.725 170.215 63.665 170.385 ;
        RECT 62.725 169.965 62.895 170.215 ;
        RECT 64.035 169.965 64.300 170.325 ;
        RECT 62.605 169.635 62.895 169.965 ;
        RECT 63.065 169.715 63.405 169.965 ;
        RECT 63.625 169.715 64.300 169.965 ;
        RECT 62.725 169.545 62.895 169.635 ;
        RECT 62.725 169.355 64.115 169.545 ;
        RECT 64.485 169.405 64.725 170.715 ;
        RECT 64.995 170.305 65.245 171.105 ;
        RECT 65.465 170.555 65.795 171.275 ;
        RECT 65.980 170.305 66.230 171.105 ;
        RECT 66.695 170.475 67.025 171.275 ;
        RECT 67.195 170.845 67.535 171.105 ;
        RECT 64.895 170.135 67.085 170.305 ;
        RECT 62.185 168.895 62.745 169.185 ;
        RECT 62.915 168.725 63.165 169.185 ;
        RECT 63.785 168.995 64.115 169.355 ;
        RECT 64.895 169.225 65.065 170.135 ;
        RECT 66.770 169.965 67.085 170.135 ;
        RECT 64.570 168.895 65.065 169.225 ;
        RECT 65.285 169.000 65.635 169.965 ;
        RECT 65.815 168.995 66.115 169.965 ;
        RECT 66.295 168.995 66.575 169.965 ;
        RECT 66.770 169.715 67.100 169.965 ;
        RECT 66.755 168.725 67.025 169.525 ;
        RECT 67.275 169.445 67.535 170.845 ;
        RECT 67.195 168.935 67.535 169.445 ;
        RECT 67.740 170.485 68.275 171.105 ;
        RECT 67.740 169.465 68.055 170.485 ;
        RECT 68.445 170.475 68.775 171.275 ;
        RECT 69.260 170.305 69.650 170.480 ;
        RECT 68.225 170.135 69.650 170.305 ;
        RECT 68.225 169.635 68.395 170.135 ;
        RECT 67.740 168.895 68.355 169.465 ;
        RECT 68.645 169.405 68.910 169.965 ;
        RECT 69.080 169.235 69.250 170.135 ;
        RECT 70.005 170.110 70.295 171.275 ;
        RECT 70.555 170.605 70.725 171.105 ;
        RECT 70.895 170.775 71.225 171.275 ;
        RECT 70.555 170.435 71.220 170.605 ;
        RECT 69.420 169.405 69.775 169.965 ;
        RECT 70.470 169.615 70.820 170.265 ;
        RECT 68.525 168.725 68.740 169.235 ;
        RECT 68.970 168.905 69.250 169.235 ;
        RECT 69.430 168.725 69.670 169.235 ;
        RECT 70.005 168.725 70.295 169.450 ;
        RECT 70.990 169.445 71.220 170.435 ;
        RECT 70.555 169.275 71.220 169.445 ;
        RECT 70.555 168.985 70.725 169.275 ;
        RECT 70.895 168.725 71.225 169.105 ;
        RECT 71.395 168.985 71.580 171.105 ;
        RECT 71.820 170.815 72.085 171.275 ;
        RECT 72.255 170.680 72.505 171.105 ;
        RECT 72.715 170.830 73.820 171.000 ;
        RECT 72.200 170.550 72.505 170.680 ;
        RECT 71.750 169.355 72.030 170.305 ;
        RECT 72.200 169.445 72.370 170.550 ;
        RECT 72.540 169.765 72.780 170.360 ;
        RECT 72.950 170.295 73.480 170.660 ;
        RECT 72.950 169.595 73.120 170.295 ;
        RECT 73.650 170.215 73.820 170.830 ;
        RECT 73.990 170.475 74.160 171.275 ;
        RECT 74.330 170.775 74.580 171.105 ;
        RECT 74.805 170.805 75.690 170.975 ;
        RECT 73.650 170.125 74.160 170.215 ;
        RECT 72.200 169.315 72.425 169.445 ;
        RECT 72.595 169.375 73.120 169.595 ;
        RECT 73.290 169.955 74.160 170.125 ;
        RECT 71.835 168.725 72.085 169.185 ;
        RECT 72.255 169.175 72.425 169.315 ;
        RECT 73.290 169.175 73.460 169.955 ;
        RECT 73.990 169.885 74.160 169.955 ;
        RECT 73.670 169.705 73.870 169.735 ;
        RECT 74.330 169.705 74.500 170.775 ;
        RECT 74.670 169.885 74.860 170.605 ;
        RECT 73.670 169.405 74.500 169.705 ;
        RECT 75.030 169.675 75.350 170.635 ;
        RECT 72.255 169.005 72.590 169.175 ;
        RECT 72.785 169.005 73.460 169.175 ;
        RECT 73.780 168.725 74.150 169.225 ;
        RECT 74.330 169.175 74.500 169.405 ;
        RECT 74.885 169.345 75.350 169.675 ;
        RECT 75.520 169.965 75.690 170.805 ;
        RECT 75.870 170.775 76.185 171.275 ;
        RECT 76.415 170.545 76.755 171.105 ;
        RECT 75.860 170.170 76.755 170.545 ;
        RECT 76.925 170.265 77.095 171.275 ;
        RECT 76.565 169.965 76.755 170.170 ;
        RECT 77.265 170.215 77.595 171.060 ;
        RECT 77.265 170.135 77.655 170.215 ;
        RECT 77.825 170.185 81.335 171.275 ;
        RECT 81.505 170.185 82.715 171.275 ;
        RECT 77.440 170.085 77.655 170.135 ;
        RECT 75.520 169.635 76.395 169.965 ;
        RECT 76.565 169.635 77.315 169.965 ;
        RECT 75.520 169.175 75.690 169.635 ;
        RECT 76.565 169.465 76.765 169.635 ;
        RECT 77.485 169.505 77.655 170.085 ;
        RECT 77.430 169.465 77.655 169.505 ;
        RECT 74.330 169.005 74.735 169.175 ;
        RECT 74.905 169.005 75.690 169.175 ;
        RECT 75.965 168.725 76.175 169.255 ;
        RECT 76.435 168.940 76.765 169.465 ;
        RECT 77.275 169.380 77.655 169.465 ;
        RECT 77.825 169.495 79.475 170.015 ;
        RECT 79.645 169.665 81.335 170.185 ;
        RECT 76.935 168.725 77.105 169.335 ;
        RECT 77.275 168.945 77.605 169.380 ;
        RECT 77.825 168.725 81.335 169.495 ;
        RECT 81.505 169.475 82.025 170.015 ;
        RECT 82.195 169.645 82.715 170.185 ;
        RECT 82.885 170.185 84.095 171.275 ;
        RECT 82.885 169.645 83.405 170.185 ;
        RECT 83.575 169.475 84.095 170.015 ;
        RECT 81.505 168.725 82.715 169.475 ;
        RECT 82.885 168.725 84.095 169.475 ;
        RECT 5.520 168.555 84.180 168.725 ;
        RECT 5.605 167.805 6.815 168.555 ;
        RECT 6.985 168.010 12.330 168.555 ;
        RECT 5.605 167.265 6.125 167.805 ;
        RECT 6.295 167.095 6.815 167.635 ;
        RECT 8.570 167.180 8.910 168.010 ;
        RECT 12.505 167.785 14.175 168.555 ;
        RECT 14.435 168.005 14.605 168.295 ;
        RECT 14.775 168.175 15.105 168.555 ;
        RECT 14.435 167.835 15.100 168.005 ;
        RECT 5.605 166.005 6.815 167.095 ;
        RECT 10.390 166.440 10.740 167.690 ;
        RECT 12.505 167.265 13.255 167.785 ;
        RECT 13.425 167.095 14.175 167.615 ;
        RECT 6.985 166.005 12.330 166.440 ;
        RECT 12.505 166.005 14.175 167.095 ;
        RECT 14.350 167.015 14.700 167.665 ;
        RECT 14.870 166.845 15.100 167.835 ;
        RECT 14.435 166.675 15.100 166.845 ;
        RECT 14.435 166.175 14.605 166.675 ;
        RECT 14.775 166.005 15.105 166.505 ;
        RECT 15.275 166.175 15.460 168.295 ;
        RECT 15.715 168.095 15.965 168.555 ;
        RECT 16.135 168.105 16.470 168.275 ;
        RECT 16.665 168.105 17.340 168.275 ;
        RECT 16.135 167.965 16.305 168.105 ;
        RECT 15.630 166.975 15.910 167.925 ;
        RECT 16.080 167.835 16.305 167.965 ;
        RECT 16.080 166.730 16.250 167.835 ;
        RECT 16.475 167.685 17.000 167.905 ;
        RECT 16.420 166.920 16.660 167.515 ;
        RECT 16.830 166.985 17.000 167.685 ;
        RECT 17.170 167.325 17.340 168.105 ;
        RECT 17.660 168.055 18.030 168.555 ;
        RECT 18.210 168.105 18.615 168.275 ;
        RECT 18.785 168.105 19.570 168.275 ;
        RECT 18.210 167.875 18.380 168.105 ;
        RECT 17.550 167.575 18.380 167.875 ;
        RECT 18.765 167.605 19.230 167.935 ;
        RECT 17.550 167.545 17.750 167.575 ;
        RECT 17.870 167.325 18.040 167.395 ;
        RECT 17.170 167.155 18.040 167.325 ;
        RECT 17.530 167.065 18.040 167.155 ;
        RECT 16.080 166.600 16.385 166.730 ;
        RECT 16.830 166.620 17.360 166.985 ;
        RECT 15.700 166.005 15.965 166.465 ;
        RECT 16.135 166.175 16.385 166.600 ;
        RECT 17.530 166.450 17.700 167.065 ;
        RECT 16.595 166.280 17.700 166.450 ;
        RECT 17.870 166.005 18.040 166.805 ;
        RECT 18.210 166.505 18.380 167.575 ;
        RECT 18.550 166.675 18.740 167.395 ;
        RECT 18.910 166.645 19.230 167.605 ;
        RECT 19.400 167.645 19.570 168.105 ;
        RECT 19.845 168.025 20.055 168.555 ;
        RECT 20.315 167.815 20.645 168.340 ;
        RECT 20.815 167.945 20.985 168.555 ;
        RECT 21.155 167.900 21.485 168.335 ;
        RECT 21.155 167.815 21.535 167.900 ;
        RECT 20.445 167.645 20.645 167.815 ;
        RECT 21.310 167.775 21.535 167.815 ;
        RECT 19.400 167.315 20.275 167.645 ;
        RECT 20.445 167.315 21.195 167.645 ;
        RECT 18.210 166.175 18.460 166.505 ;
        RECT 19.400 166.475 19.570 167.315 ;
        RECT 20.445 167.110 20.635 167.315 ;
        RECT 21.365 167.195 21.535 167.775 ;
        RECT 21.705 167.755 22.015 168.555 ;
        RECT 22.220 167.755 22.915 168.385 ;
        RECT 23.175 168.005 23.345 168.295 ;
        RECT 23.515 168.175 23.845 168.555 ;
        RECT 23.175 167.835 23.840 168.005 ;
        RECT 21.715 167.315 22.050 167.585 ;
        RECT 21.320 167.145 21.535 167.195 ;
        RECT 22.220 167.155 22.390 167.755 ;
        RECT 22.560 167.315 22.895 167.565 ;
        RECT 19.740 166.735 20.635 167.110 ;
        RECT 21.145 167.065 21.535 167.145 ;
        RECT 18.685 166.305 19.570 166.475 ;
        RECT 19.750 166.005 20.065 166.505 ;
        RECT 20.295 166.175 20.635 166.735 ;
        RECT 20.805 166.005 20.975 167.015 ;
        RECT 21.145 166.220 21.475 167.065 ;
        RECT 21.705 166.005 21.985 167.145 ;
        RECT 22.155 166.175 22.485 167.155 ;
        RECT 22.655 166.005 22.915 167.145 ;
        RECT 23.090 167.015 23.440 167.665 ;
        RECT 23.610 166.845 23.840 167.835 ;
        RECT 23.175 166.675 23.840 166.845 ;
        RECT 23.175 166.175 23.345 166.675 ;
        RECT 23.515 166.005 23.845 166.505 ;
        RECT 24.015 166.175 24.200 168.295 ;
        RECT 24.455 168.095 24.705 168.555 ;
        RECT 24.875 168.105 25.210 168.275 ;
        RECT 25.405 168.105 26.080 168.275 ;
        RECT 24.875 167.965 25.045 168.105 ;
        RECT 24.370 166.975 24.650 167.925 ;
        RECT 24.820 167.835 25.045 167.965 ;
        RECT 24.820 166.730 24.990 167.835 ;
        RECT 25.215 167.685 25.740 167.905 ;
        RECT 25.160 166.920 25.400 167.515 ;
        RECT 25.570 166.985 25.740 167.685 ;
        RECT 25.910 167.325 26.080 168.105 ;
        RECT 26.400 168.055 26.770 168.555 ;
        RECT 26.950 168.105 27.355 168.275 ;
        RECT 27.525 168.105 28.310 168.275 ;
        RECT 26.950 167.875 27.120 168.105 ;
        RECT 26.290 167.575 27.120 167.875 ;
        RECT 27.505 167.605 27.970 167.935 ;
        RECT 26.290 167.545 26.490 167.575 ;
        RECT 26.610 167.325 26.780 167.395 ;
        RECT 25.910 167.155 26.780 167.325 ;
        RECT 26.270 167.065 26.780 167.155 ;
        RECT 24.820 166.600 25.125 166.730 ;
        RECT 25.570 166.620 26.100 166.985 ;
        RECT 24.440 166.005 24.705 166.465 ;
        RECT 24.875 166.175 25.125 166.600 ;
        RECT 26.270 166.450 26.440 167.065 ;
        RECT 25.335 166.280 26.440 166.450 ;
        RECT 26.610 166.005 26.780 166.805 ;
        RECT 26.950 166.505 27.120 167.575 ;
        RECT 27.290 166.675 27.480 167.395 ;
        RECT 27.650 166.645 27.970 167.605 ;
        RECT 28.140 167.645 28.310 168.105 ;
        RECT 28.585 168.025 28.795 168.555 ;
        RECT 29.055 167.815 29.385 168.340 ;
        RECT 29.555 167.945 29.725 168.555 ;
        RECT 29.895 167.900 30.225 168.335 ;
        RECT 29.895 167.815 30.275 167.900 ;
        RECT 31.365 167.830 31.655 168.555 ;
        RECT 31.910 168.165 33.920 168.385 ;
        RECT 29.185 167.645 29.385 167.815 ;
        RECT 30.050 167.775 30.275 167.815 ;
        RECT 28.140 167.315 29.015 167.645 ;
        RECT 29.185 167.315 29.935 167.645 ;
        RECT 26.950 166.175 27.200 166.505 ;
        RECT 28.140 166.475 28.310 167.315 ;
        RECT 29.185 167.110 29.375 167.315 ;
        RECT 30.105 167.195 30.275 167.775 ;
        RECT 30.060 167.145 30.275 167.195 ;
        RECT 31.825 167.735 33.500 167.995 ;
        RECT 33.670 167.915 33.920 168.165 ;
        RECT 34.090 168.085 34.260 168.555 ;
        RECT 34.430 167.915 34.760 168.385 ;
        RECT 34.930 168.085 35.100 168.555 ;
        RECT 35.270 167.915 35.600 168.385 ;
        RECT 33.670 167.735 35.600 167.915 ;
        RECT 35.775 167.735 36.050 168.555 ;
        RECT 36.220 167.915 36.550 168.385 ;
        RECT 36.720 168.085 36.890 168.555 ;
        RECT 37.060 167.915 37.390 168.385 ;
        RECT 37.560 168.085 37.730 168.555 ;
        RECT 37.900 167.915 38.230 168.385 ;
        RECT 38.400 168.085 38.570 168.555 ;
        RECT 38.740 167.915 39.070 168.385 ;
        RECT 39.240 168.085 39.510 168.555 ;
        RECT 39.700 168.165 41.710 168.335 ;
        RECT 36.220 167.905 39.170 167.915 ;
        RECT 39.700 167.905 39.950 168.165 ;
        RECT 42.035 168.005 42.205 168.295 ;
        RECT 42.375 168.175 42.705 168.555 ;
        RECT 36.220 167.735 39.950 167.905 ;
        RECT 40.120 167.735 41.775 167.995 ;
        RECT 42.035 167.835 42.700 168.005 ;
        RECT 31.825 167.195 32.060 167.735 ;
        RECT 32.230 167.365 33.595 167.565 ;
        RECT 33.915 167.365 37.130 167.565 ;
        RECT 37.300 167.365 39.170 167.565 ;
        RECT 39.340 167.365 41.385 167.565 ;
        RECT 33.425 167.195 33.595 167.365 ;
        RECT 37.300 167.195 37.470 167.365 ;
        RECT 39.340 167.195 39.510 167.365 ;
        RECT 41.555 167.195 41.775 167.735 ;
        RECT 28.480 166.735 29.375 167.110 ;
        RECT 29.885 167.065 30.275 167.145 ;
        RECT 27.425 166.305 28.310 166.475 ;
        RECT 28.490 166.005 28.805 166.505 ;
        RECT 29.035 166.175 29.375 166.735 ;
        RECT 29.545 166.005 29.715 167.015 ;
        RECT 29.885 166.220 30.215 167.065 ;
        RECT 31.365 166.005 31.655 167.170 ;
        RECT 31.825 167.025 33.040 167.195 ;
        RECT 33.425 167.025 37.470 167.195 ;
        RECT 37.640 167.025 39.510 167.195 ;
        RECT 31.825 166.175 32.200 167.025 ;
        RECT 32.790 166.855 33.040 167.025 ;
        RECT 39.700 166.975 41.775 167.195 ;
        RECT 41.950 167.015 42.300 167.665 ;
        RECT 39.700 166.855 39.990 166.975 ;
        RECT 32.370 166.005 32.620 166.805 ;
        RECT 32.790 166.635 35.560 166.855 ;
        RECT 32.790 166.175 33.040 166.635 ;
        RECT 33.210 166.005 33.460 166.465 ;
        RECT 33.630 166.175 33.880 166.635 ;
        RECT 34.050 166.005 34.300 166.465 ;
        RECT 34.470 166.175 34.720 166.635 ;
        RECT 34.890 166.005 35.140 166.465 ;
        RECT 35.310 166.175 35.560 166.635 ;
        RECT 35.775 166.635 37.730 166.855 ;
        RECT 35.775 166.175 36.090 166.635 ;
        RECT 36.260 166.005 36.510 166.465 ;
        RECT 36.680 166.175 36.930 166.635 ;
        RECT 37.100 166.005 37.350 166.465 ;
        RECT 37.520 166.425 37.730 166.635 ;
        RECT 37.900 166.595 39.990 166.855 ;
        RECT 37.520 166.175 39.490 166.425 ;
        RECT 39.700 166.175 39.990 166.595 ;
        RECT 40.160 166.005 40.410 166.805 ;
        RECT 40.580 166.175 40.830 166.975 ;
        RECT 41.000 166.005 41.250 166.805 ;
        RECT 41.420 166.175 41.775 166.975 ;
        RECT 42.470 166.845 42.700 167.835 ;
        RECT 42.035 166.675 42.700 166.845 ;
        RECT 42.035 166.175 42.205 166.675 ;
        RECT 42.375 166.005 42.705 166.505 ;
        RECT 42.875 166.175 43.060 168.295 ;
        RECT 43.315 168.095 43.565 168.555 ;
        RECT 43.735 168.105 44.070 168.275 ;
        RECT 44.265 168.105 44.940 168.275 ;
        RECT 43.735 167.965 43.905 168.105 ;
        RECT 43.230 166.975 43.510 167.925 ;
        RECT 43.680 167.835 43.905 167.965 ;
        RECT 43.680 166.730 43.850 167.835 ;
        RECT 44.075 167.685 44.600 167.905 ;
        RECT 44.020 166.920 44.260 167.515 ;
        RECT 44.430 166.985 44.600 167.685 ;
        RECT 44.770 167.325 44.940 168.105 ;
        RECT 45.260 168.055 45.630 168.555 ;
        RECT 45.810 168.105 46.215 168.275 ;
        RECT 46.385 168.105 47.170 168.275 ;
        RECT 45.810 167.875 45.980 168.105 ;
        RECT 45.150 167.575 45.980 167.875 ;
        RECT 46.365 167.605 46.830 167.935 ;
        RECT 45.150 167.545 45.350 167.575 ;
        RECT 45.470 167.325 45.640 167.395 ;
        RECT 44.770 167.155 45.640 167.325 ;
        RECT 45.130 167.065 45.640 167.155 ;
        RECT 43.680 166.600 43.985 166.730 ;
        RECT 44.430 166.620 44.960 166.985 ;
        RECT 43.300 166.005 43.565 166.465 ;
        RECT 43.735 166.175 43.985 166.600 ;
        RECT 45.130 166.450 45.300 167.065 ;
        RECT 44.195 166.280 45.300 166.450 ;
        RECT 45.470 166.005 45.640 166.805 ;
        RECT 45.810 166.505 45.980 167.575 ;
        RECT 46.150 166.675 46.340 167.395 ;
        RECT 46.510 166.645 46.830 167.605 ;
        RECT 47.000 167.645 47.170 168.105 ;
        RECT 47.445 168.025 47.655 168.555 ;
        RECT 47.915 167.815 48.245 168.340 ;
        RECT 48.415 167.945 48.585 168.555 ;
        RECT 48.755 167.900 49.085 168.335 ;
        RECT 49.305 167.945 49.645 168.360 ;
        RECT 49.815 168.115 49.985 168.555 ;
        RECT 50.175 168.165 51.435 168.345 ;
        RECT 50.175 167.945 50.505 168.165 ;
        RECT 48.755 167.815 49.135 167.900 ;
        RECT 48.045 167.645 48.245 167.815 ;
        RECT 48.910 167.775 49.135 167.815 ;
        RECT 49.305 167.815 50.505 167.945 ;
        RECT 50.675 167.815 51.025 167.995 ;
        RECT 49.305 167.775 50.335 167.815 ;
        RECT 47.000 167.315 47.875 167.645 ;
        RECT 48.045 167.315 48.795 167.645 ;
        RECT 45.810 166.175 46.060 166.505 ;
        RECT 47.000 166.475 47.170 167.315 ;
        RECT 48.045 167.110 48.235 167.315 ;
        RECT 48.965 167.195 49.135 167.775 ;
        RECT 49.305 167.365 49.765 167.565 ;
        RECT 49.935 167.395 50.300 167.565 ;
        RECT 49.935 167.195 50.115 167.395 ;
        RECT 50.515 167.225 50.685 167.645 ;
        RECT 48.920 167.145 49.135 167.195 ;
        RECT 47.340 166.735 48.235 167.110 ;
        RECT 48.745 167.065 49.135 167.145 ;
        RECT 46.285 166.305 47.170 166.475 ;
        RECT 47.350 166.005 47.665 166.505 ;
        RECT 47.895 166.175 48.235 166.735 ;
        RECT 48.405 166.005 48.575 167.015 ;
        RECT 48.745 166.220 49.075 167.065 ;
        RECT 49.305 166.005 49.625 167.185 ;
        RECT 49.795 167.025 50.115 167.195 ;
        RECT 49.795 166.235 49.995 167.025 ;
        RECT 50.285 166.975 50.685 167.225 ;
        RECT 50.855 166.805 51.025 167.815 ;
        RECT 50.185 166.595 51.025 166.805 ;
        RECT 51.195 166.650 51.435 167.975 ;
        RECT 52.530 167.715 52.790 168.555 ;
        RECT 52.965 167.810 53.220 168.385 ;
        RECT 53.390 168.175 53.720 168.555 ;
        RECT 53.935 168.005 54.105 168.385 ;
        RECT 53.390 167.835 54.105 168.005 ;
        RECT 50.185 166.175 50.685 166.595 ;
        RECT 51.175 166.005 51.385 166.465 ;
        RECT 52.530 166.005 52.790 167.155 ;
        RECT 52.965 167.080 53.135 167.810 ;
        RECT 53.390 167.645 53.560 167.835 ;
        RECT 54.365 167.785 56.955 168.555 ;
        RECT 57.125 167.830 57.415 168.555 ;
        RECT 57.585 167.815 57.925 168.385 ;
        RECT 58.120 167.890 58.290 168.555 ;
        RECT 58.570 168.215 58.790 168.260 ;
        RECT 58.565 168.045 58.790 168.215 ;
        RECT 58.960 168.075 59.405 168.245 ;
        RECT 58.570 167.905 58.790 168.045 ;
        RECT 53.305 167.315 53.560 167.645 ;
        RECT 53.390 167.105 53.560 167.315 ;
        RECT 53.840 167.285 54.195 167.655 ;
        RECT 54.365 167.265 55.575 167.785 ;
        RECT 52.965 166.175 53.220 167.080 ;
        RECT 53.390 166.935 54.105 167.105 ;
        RECT 55.745 167.095 56.955 167.615 ;
        RECT 53.390 166.005 53.720 166.765 ;
        RECT 53.935 166.175 54.105 166.935 ;
        RECT 54.365 166.005 56.955 167.095 ;
        RECT 57.125 166.005 57.415 167.170 ;
        RECT 57.585 166.845 57.760 167.815 ;
        RECT 58.570 167.735 59.065 167.905 ;
        RECT 57.930 167.195 58.100 167.645 ;
        RECT 58.270 167.365 58.720 167.565 ;
        RECT 58.890 167.540 59.065 167.735 ;
        RECT 59.235 167.285 59.405 168.075 ;
        RECT 59.575 167.950 59.825 168.320 ;
        RECT 59.655 167.565 59.825 167.950 ;
        RECT 59.995 167.915 60.245 168.320 ;
        RECT 60.415 168.085 60.585 168.555 ;
        RECT 60.755 167.915 61.095 168.320 ;
        RECT 59.995 167.735 61.095 167.915 ;
        RECT 61.265 167.785 62.935 168.555 ;
        RECT 63.155 167.900 63.485 168.335 ;
        RECT 63.655 167.945 63.825 168.555 ;
        RECT 63.105 167.815 63.485 167.900 ;
        RECT 63.995 167.815 64.325 168.340 ;
        RECT 64.585 168.025 64.795 168.555 ;
        RECT 65.070 168.105 65.855 168.275 ;
        RECT 66.025 168.105 66.430 168.275 ;
        RECT 59.655 167.395 59.850 167.565 ;
        RECT 57.930 167.025 58.325 167.195 ;
        RECT 59.235 167.145 59.510 167.285 ;
        RECT 57.585 166.175 57.845 166.845 ;
        RECT 58.155 166.755 58.325 167.025 ;
        RECT 58.495 166.925 59.510 167.145 ;
        RECT 59.680 167.145 59.850 167.395 ;
        RECT 60.020 167.315 60.580 167.565 ;
        RECT 59.680 166.755 60.235 167.145 ;
        RECT 58.155 166.585 60.235 166.755 ;
        RECT 58.015 166.005 58.345 166.405 ;
        RECT 59.215 166.005 59.615 166.405 ;
        RECT 59.905 166.350 60.235 166.585 ;
        RECT 60.405 166.215 60.580 167.315 ;
        RECT 60.750 166.995 61.095 167.565 ;
        RECT 61.265 167.265 62.015 167.785 ;
        RECT 63.105 167.775 63.330 167.815 ;
        RECT 62.185 167.095 62.935 167.615 ;
        RECT 60.750 166.005 61.095 166.825 ;
        RECT 61.265 166.005 62.935 167.095 ;
        RECT 63.105 167.195 63.275 167.775 ;
        RECT 63.995 167.645 64.195 167.815 ;
        RECT 65.070 167.645 65.240 168.105 ;
        RECT 63.445 167.315 64.195 167.645 ;
        RECT 64.365 167.315 65.240 167.645 ;
        RECT 63.105 167.145 63.320 167.195 ;
        RECT 63.105 167.065 63.495 167.145 ;
        RECT 63.165 166.220 63.495 167.065 ;
        RECT 64.005 167.110 64.195 167.315 ;
        RECT 63.665 166.005 63.835 167.015 ;
        RECT 64.005 166.735 64.900 167.110 ;
        RECT 64.005 166.175 64.345 166.735 ;
        RECT 64.575 166.005 64.890 166.505 ;
        RECT 65.070 166.475 65.240 167.315 ;
        RECT 65.410 167.605 65.875 167.935 ;
        RECT 66.260 167.875 66.430 168.105 ;
        RECT 66.610 168.055 66.980 168.555 ;
        RECT 67.300 168.105 67.975 168.275 ;
        RECT 68.170 168.105 68.505 168.275 ;
        RECT 65.410 166.645 65.730 167.605 ;
        RECT 66.260 167.575 67.090 167.875 ;
        RECT 65.900 166.675 66.090 167.395 ;
        RECT 66.260 166.505 66.430 167.575 ;
        RECT 66.890 167.545 67.090 167.575 ;
        RECT 66.600 167.325 66.770 167.395 ;
        RECT 67.300 167.325 67.470 168.105 ;
        RECT 68.335 167.965 68.505 168.105 ;
        RECT 68.675 168.095 68.925 168.555 ;
        RECT 66.600 167.155 67.470 167.325 ;
        RECT 67.640 167.685 68.165 167.905 ;
        RECT 68.335 167.835 68.560 167.965 ;
        RECT 66.600 167.065 67.110 167.155 ;
        RECT 65.070 166.305 65.955 166.475 ;
        RECT 66.180 166.175 66.430 166.505 ;
        RECT 66.600 166.005 66.770 166.805 ;
        RECT 66.940 166.450 67.110 167.065 ;
        RECT 67.640 166.985 67.810 167.685 ;
        RECT 67.280 166.620 67.810 166.985 ;
        RECT 67.980 166.920 68.220 167.515 ;
        RECT 68.390 166.730 68.560 167.835 ;
        RECT 68.730 166.975 69.010 167.925 ;
        RECT 68.255 166.600 68.560 166.730 ;
        RECT 66.940 166.280 68.045 166.450 ;
        RECT 68.255 166.175 68.505 166.600 ;
        RECT 68.675 166.005 68.940 166.465 ;
        RECT 69.180 166.175 69.365 168.295 ;
        RECT 69.535 168.175 69.865 168.555 ;
        RECT 70.035 168.005 70.205 168.295 ;
        RECT 70.465 168.010 75.810 168.555 ;
        RECT 75.985 168.010 81.330 168.555 ;
        RECT 69.540 167.835 70.205 168.005 ;
        RECT 69.540 166.845 69.770 167.835 ;
        RECT 69.940 167.015 70.290 167.665 ;
        RECT 72.050 167.180 72.390 168.010 ;
        RECT 69.540 166.675 70.205 166.845 ;
        RECT 69.535 166.005 69.865 166.505 ;
        RECT 70.035 166.175 70.205 166.675 ;
        RECT 73.870 166.440 74.220 167.690 ;
        RECT 77.570 167.180 77.910 168.010 ;
        RECT 81.505 167.805 82.715 168.555 ;
        RECT 82.885 167.805 84.095 168.555 ;
        RECT 79.390 166.440 79.740 167.690 ;
        RECT 81.505 167.265 82.025 167.805 ;
        RECT 82.195 167.095 82.715 167.635 ;
        RECT 70.465 166.005 75.810 166.440 ;
        RECT 75.985 166.005 81.330 166.440 ;
        RECT 81.505 166.005 82.715 167.095 ;
        RECT 82.885 167.095 83.405 167.635 ;
        RECT 83.575 167.265 84.095 167.805 ;
        RECT 82.885 166.005 84.095 167.095 ;
        RECT 5.520 165.835 84.180 166.005 ;
        RECT 5.605 164.745 6.815 165.835 ;
        RECT 6.985 165.400 12.330 165.835 ;
        RECT 5.605 164.035 6.125 164.575 ;
        RECT 6.295 164.205 6.815 164.745 ;
        RECT 5.605 163.285 6.815 164.035 ;
        RECT 8.570 163.830 8.910 164.660 ;
        RECT 10.390 164.150 10.740 165.400 ;
        RECT 12.505 164.745 14.175 165.835 ;
        RECT 12.505 164.055 13.255 164.575 ;
        RECT 13.425 164.225 14.175 164.745 ;
        RECT 14.805 164.965 15.080 165.665 ;
        RECT 15.290 165.290 15.505 165.835 ;
        RECT 15.675 165.325 16.150 165.665 ;
        RECT 16.320 165.330 16.935 165.835 ;
        RECT 16.320 165.155 16.515 165.330 ;
        RECT 6.985 163.285 12.330 163.830 ;
        RECT 12.505 163.285 14.175 164.055 ;
        RECT 14.805 163.935 14.975 164.965 ;
        RECT 15.250 164.795 15.965 165.090 ;
        RECT 16.185 164.965 16.515 165.155 ;
        RECT 16.685 164.795 16.935 165.160 ;
        RECT 15.145 164.625 16.935 164.795 ;
        RECT 15.145 164.195 15.375 164.625 ;
        RECT 14.805 163.455 15.065 163.935 ;
        RECT 15.545 163.925 15.955 164.445 ;
        RECT 15.235 163.285 15.565 163.745 ;
        RECT 15.755 163.505 15.955 163.925 ;
        RECT 16.125 163.770 16.380 164.625 ;
        RECT 17.175 164.445 17.345 165.665 ;
        RECT 17.595 165.325 17.855 165.835 ;
        RECT 16.550 164.195 17.345 164.445 ;
        RECT 17.515 164.275 17.855 165.155 ;
        RECT 18.485 164.670 18.775 165.835 ;
        RECT 17.095 164.105 17.345 164.195 ;
        RECT 16.125 163.505 16.915 163.770 ;
        RECT 17.095 163.685 17.425 164.105 ;
        RECT 17.595 163.285 17.855 164.105 ;
        RECT 18.485 163.285 18.775 164.010 ;
        RECT 18.955 163.465 19.215 165.655 ;
        RECT 19.385 165.105 19.725 165.835 ;
        RECT 19.905 164.925 20.175 165.655 ;
        RECT 19.405 164.705 20.175 164.925 ;
        RECT 20.355 164.945 20.585 165.655 ;
        RECT 20.755 165.125 21.085 165.835 ;
        RECT 21.255 164.945 21.515 165.655 ;
        RECT 21.875 165.035 22.130 165.835 ;
        RECT 20.355 164.705 21.515 164.945 ;
        RECT 22.300 164.865 22.630 165.665 ;
        RECT 22.800 165.035 22.970 165.835 ;
        RECT 23.140 164.865 23.470 165.665 ;
        RECT 23.640 165.035 23.810 165.835 ;
        RECT 23.980 164.865 24.310 165.665 ;
        RECT 24.480 165.035 24.650 165.835 ;
        RECT 24.820 164.865 25.150 165.665 ;
        RECT 25.320 165.035 25.620 165.835 ;
        RECT 19.405 164.035 19.695 164.705 ;
        RECT 21.705 164.695 25.675 164.865 ;
        RECT 25.845 164.745 27.515 165.835 ;
        RECT 19.875 164.215 20.340 164.525 ;
        RECT 20.520 164.215 21.045 164.525 ;
        RECT 19.405 163.835 20.635 164.035 ;
        RECT 19.475 163.285 20.145 163.655 ;
        RECT 20.325 163.465 20.635 163.835 ;
        RECT 20.815 163.575 21.045 164.215 ;
        RECT 21.225 164.195 21.525 164.525 ;
        RECT 21.705 164.105 22.050 164.695 ;
        RECT 22.300 164.275 25.155 164.525 ;
        RECT 25.355 164.105 25.675 164.695 ;
        RECT 21.225 163.285 21.515 164.015 ;
        RECT 21.705 163.915 25.675 164.105 ;
        RECT 25.845 164.055 26.595 164.575 ;
        RECT 26.765 164.225 27.515 164.745 ;
        RECT 27.870 164.865 28.260 165.040 ;
        RECT 28.745 165.035 29.075 165.835 ;
        RECT 29.245 165.045 29.780 165.665 ;
        RECT 27.870 164.695 29.295 164.865 ;
        RECT 21.875 163.285 22.130 163.745 ;
        RECT 22.300 163.455 22.630 163.915 ;
        RECT 22.800 163.285 22.970 163.745 ;
        RECT 23.140 163.455 23.470 163.915 ;
        RECT 23.640 163.285 23.810 163.745 ;
        RECT 23.980 163.455 24.310 163.915 ;
        RECT 24.480 163.285 24.650 163.745 ;
        RECT 24.820 163.455 25.150 163.915 ;
        RECT 25.320 163.285 25.625 163.745 ;
        RECT 25.845 163.285 27.515 164.055 ;
        RECT 27.745 163.965 28.100 164.525 ;
        RECT 28.270 163.795 28.440 164.695 ;
        RECT 28.610 163.965 28.875 164.525 ;
        RECT 29.125 164.195 29.295 164.695 ;
        RECT 29.465 164.025 29.780 165.045 ;
        RECT 30.030 164.695 30.325 165.835 ;
        RECT 30.585 164.865 30.915 165.665 ;
        RECT 31.085 165.035 31.255 165.835 ;
        RECT 31.425 164.865 31.755 165.665 ;
        RECT 31.925 165.035 32.095 165.835 ;
        RECT 32.265 164.885 32.595 165.665 ;
        RECT 32.765 165.375 32.935 165.835 ;
        RECT 33.295 165.165 33.465 165.665 ;
        RECT 33.635 165.335 33.965 165.835 ;
        RECT 33.295 164.995 33.960 165.165 ;
        RECT 32.265 164.865 33.035 164.885 ;
        RECT 30.585 164.695 33.035 164.865 ;
        RECT 30.005 164.275 32.515 164.525 ;
        RECT 32.685 164.105 33.035 164.695 ;
        RECT 33.210 164.175 33.560 164.825 ;
        RECT 27.850 163.285 28.090 163.795 ;
        RECT 28.270 163.465 28.550 163.795 ;
        RECT 28.780 163.285 28.995 163.795 ;
        RECT 29.165 163.455 29.780 164.025 ;
        RECT 30.665 163.925 33.035 164.105 ;
        RECT 33.730 164.005 33.960 164.995 ;
        RECT 30.030 163.285 30.295 163.745 ;
        RECT 30.665 163.455 30.835 163.925 ;
        RECT 31.085 163.285 31.255 163.745 ;
        RECT 31.505 163.455 31.675 163.925 ;
        RECT 31.925 163.285 32.095 163.745 ;
        RECT 32.345 163.455 32.515 163.925 ;
        RECT 33.295 163.835 33.960 164.005 ;
        RECT 32.685 163.285 32.935 163.750 ;
        RECT 33.295 163.545 33.465 163.835 ;
        RECT 33.635 163.285 33.965 163.665 ;
        RECT 34.135 163.545 34.320 165.665 ;
        RECT 34.560 165.375 34.825 165.835 ;
        RECT 34.995 165.240 35.245 165.665 ;
        RECT 35.455 165.390 36.560 165.560 ;
        RECT 34.940 165.110 35.245 165.240 ;
        RECT 34.490 163.915 34.770 164.865 ;
        RECT 34.940 164.005 35.110 165.110 ;
        RECT 35.280 164.325 35.520 164.920 ;
        RECT 35.690 164.855 36.220 165.220 ;
        RECT 35.690 164.155 35.860 164.855 ;
        RECT 36.390 164.775 36.560 165.390 ;
        RECT 36.730 165.035 36.900 165.835 ;
        RECT 37.070 165.335 37.320 165.665 ;
        RECT 37.545 165.365 38.430 165.535 ;
        RECT 36.390 164.685 36.900 164.775 ;
        RECT 34.940 163.875 35.165 164.005 ;
        RECT 35.335 163.935 35.860 164.155 ;
        RECT 36.030 164.515 36.900 164.685 ;
        RECT 34.575 163.285 34.825 163.745 ;
        RECT 34.995 163.735 35.165 163.875 ;
        RECT 36.030 163.735 36.200 164.515 ;
        RECT 36.730 164.445 36.900 164.515 ;
        RECT 36.410 164.265 36.610 164.295 ;
        RECT 37.070 164.265 37.240 165.335 ;
        RECT 37.410 164.445 37.600 165.165 ;
        RECT 36.410 163.965 37.240 164.265 ;
        RECT 37.770 164.235 38.090 165.195 ;
        RECT 34.995 163.565 35.330 163.735 ;
        RECT 35.525 163.565 36.200 163.735 ;
        RECT 36.520 163.285 36.890 163.785 ;
        RECT 37.070 163.735 37.240 163.965 ;
        RECT 37.625 163.905 38.090 164.235 ;
        RECT 38.260 164.525 38.430 165.365 ;
        RECT 38.610 165.335 38.925 165.835 ;
        RECT 39.155 165.105 39.495 165.665 ;
        RECT 38.600 164.730 39.495 165.105 ;
        RECT 39.665 164.825 39.835 165.835 ;
        RECT 39.305 164.525 39.495 164.730 ;
        RECT 40.005 164.775 40.335 165.620 ;
        RECT 40.770 164.865 41.100 165.665 ;
        RECT 41.270 165.035 41.600 165.835 ;
        RECT 41.900 164.865 42.230 165.665 ;
        RECT 42.875 165.035 43.125 165.835 ;
        RECT 40.005 164.695 40.395 164.775 ;
        RECT 40.770 164.695 43.205 164.865 ;
        RECT 43.395 164.695 43.565 165.835 ;
        RECT 43.735 164.695 44.075 165.665 ;
        RECT 40.180 164.645 40.395 164.695 ;
        RECT 38.260 164.195 39.135 164.525 ;
        RECT 39.305 164.195 40.055 164.525 ;
        RECT 38.260 163.735 38.430 164.195 ;
        RECT 39.305 164.025 39.505 164.195 ;
        RECT 40.225 164.065 40.395 164.645 ;
        RECT 40.565 164.275 40.915 164.525 ;
        RECT 41.100 164.065 41.270 164.695 ;
        RECT 41.440 164.275 41.770 164.475 ;
        RECT 41.940 164.275 42.270 164.475 ;
        RECT 42.440 164.275 42.860 164.475 ;
        RECT 43.035 164.445 43.205 164.695 ;
        RECT 43.035 164.275 43.730 164.445 ;
        RECT 40.170 164.025 40.395 164.065 ;
        RECT 37.070 163.565 37.475 163.735 ;
        RECT 37.645 163.565 38.430 163.735 ;
        RECT 38.705 163.285 38.915 163.815 ;
        RECT 39.175 163.500 39.505 164.025 ;
        RECT 40.015 163.940 40.395 164.025 ;
        RECT 39.675 163.285 39.845 163.895 ;
        RECT 40.015 163.505 40.345 163.940 ;
        RECT 40.770 163.455 41.270 164.065 ;
        RECT 41.900 163.935 43.125 164.105 ;
        RECT 43.900 164.085 44.075 164.695 ;
        RECT 44.245 164.670 44.535 165.835 ;
        RECT 44.705 164.695 44.985 165.835 ;
        RECT 45.155 164.685 45.485 165.665 ;
        RECT 45.655 164.695 45.915 165.835 ;
        RECT 46.125 164.695 46.355 165.835 ;
        RECT 46.525 164.685 46.855 165.665 ;
        RECT 47.025 164.695 47.235 165.835 ;
        RECT 47.555 165.215 47.725 165.645 ;
        RECT 47.895 165.385 48.225 165.835 ;
        RECT 47.555 164.985 48.230 165.215 ;
        RECT 44.715 164.255 45.050 164.525 ;
        RECT 45.220 164.085 45.390 164.685 ;
        RECT 45.560 164.275 45.895 164.525 ;
        RECT 46.105 164.275 46.435 164.525 ;
        RECT 41.900 163.455 42.230 163.935 ;
        RECT 42.400 163.285 42.625 163.745 ;
        RECT 42.795 163.455 43.125 163.935 ;
        RECT 43.315 163.285 43.565 164.085 ;
        RECT 43.735 163.455 44.075 164.085 ;
        RECT 44.245 163.285 44.535 164.010 ;
        RECT 44.705 163.285 45.015 164.085 ;
        RECT 45.220 163.455 45.915 164.085 ;
        RECT 46.125 163.285 46.355 164.105 ;
        RECT 46.605 164.085 46.855 164.685 ;
        RECT 46.525 163.455 46.855 164.085 ;
        RECT 47.025 163.285 47.235 164.105 ;
        RECT 47.525 163.965 47.825 164.815 ;
        RECT 47.995 164.335 48.230 164.985 ;
        RECT 48.400 164.675 48.685 165.620 ;
        RECT 48.865 165.365 49.550 165.835 ;
        RECT 48.860 164.845 49.555 165.155 ;
        RECT 49.730 164.780 50.035 165.565 ;
        RECT 48.400 164.525 49.260 164.675 ;
        RECT 49.825 164.645 50.035 164.780 ;
        RECT 50.235 164.725 50.530 165.835 ;
        RECT 48.400 164.505 49.685 164.525 ;
        RECT 47.995 164.005 48.530 164.335 ;
        RECT 48.700 164.145 49.685 164.505 ;
        RECT 47.995 163.855 48.215 164.005 ;
        RECT 47.470 163.285 47.805 163.790 ;
        RECT 47.975 163.480 48.215 163.855 ;
        RECT 48.700 163.810 48.870 164.145 ;
        RECT 49.860 163.975 50.035 164.645 ;
        RECT 50.710 164.525 50.960 165.660 ;
        RECT 51.130 164.725 51.390 165.835 ;
        RECT 51.560 164.935 51.820 165.660 ;
        RECT 51.990 165.105 52.250 165.835 ;
        RECT 52.420 164.935 52.680 165.660 ;
        RECT 52.850 165.105 53.110 165.835 ;
        RECT 53.280 164.935 53.540 165.660 ;
        RECT 53.710 165.105 53.970 165.835 ;
        RECT 54.140 164.935 54.400 165.660 ;
        RECT 54.570 165.105 54.865 165.835 ;
        RECT 55.285 164.985 55.665 165.665 ;
        RECT 56.255 164.985 56.425 165.835 ;
        RECT 56.595 165.155 56.925 165.665 ;
        RECT 57.095 165.325 57.265 165.835 ;
        RECT 57.435 165.155 57.835 165.665 ;
        RECT 56.595 164.985 57.835 165.155 ;
        RECT 51.560 164.695 54.870 164.935 ;
        RECT 48.495 163.615 48.870 163.810 ;
        RECT 48.495 163.470 48.665 163.615 ;
        RECT 49.230 163.285 49.625 163.780 ;
        RECT 49.795 163.455 50.035 163.975 ;
        RECT 50.225 163.915 50.540 164.525 ;
        RECT 50.710 164.275 53.730 164.525 ;
        RECT 50.285 163.285 50.530 163.745 ;
        RECT 50.710 163.465 50.960 164.275 ;
        RECT 53.900 164.105 54.870 164.695 ;
        RECT 51.560 163.935 54.870 164.105 ;
        RECT 55.285 164.025 55.455 164.985 ;
        RECT 55.625 164.645 56.930 164.815 ;
        RECT 58.015 164.735 58.335 165.665 ;
        RECT 58.505 164.745 60.175 165.835 ;
        RECT 55.625 164.195 55.870 164.645 ;
        RECT 56.040 164.275 56.590 164.475 ;
        RECT 56.760 164.445 56.930 164.645 ;
        RECT 57.705 164.565 58.335 164.735 ;
        RECT 56.760 164.275 57.135 164.445 ;
        RECT 57.305 164.025 57.535 164.525 ;
        RECT 51.130 163.285 51.390 163.810 ;
        RECT 51.560 163.480 51.820 163.935 ;
        RECT 51.990 163.285 52.250 163.765 ;
        RECT 52.420 163.480 52.680 163.935 ;
        RECT 52.850 163.285 53.110 163.765 ;
        RECT 53.280 163.480 53.540 163.935 ;
        RECT 53.710 163.285 53.970 163.765 ;
        RECT 54.140 163.480 54.400 163.935 ;
        RECT 55.285 163.855 57.535 164.025 ;
        RECT 54.570 163.285 54.870 163.765 ;
        RECT 55.335 163.285 55.665 163.675 ;
        RECT 55.835 163.535 56.005 163.855 ;
        RECT 57.705 163.685 57.875 164.565 ;
        RECT 56.175 163.285 56.505 163.675 ;
        RECT 56.920 163.515 57.875 163.685 ;
        RECT 58.045 163.285 58.335 164.120 ;
        RECT 58.505 164.055 59.255 164.575 ;
        RECT 59.425 164.225 60.175 164.745 ;
        RECT 60.850 164.695 61.145 165.835 ;
        RECT 61.405 164.865 61.735 165.665 ;
        RECT 61.905 165.035 62.075 165.835 ;
        RECT 62.245 164.865 62.575 165.665 ;
        RECT 62.745 165.035 62.915 165.835 ;
        RECT 63.085 164.885 63.415 165.665 ;
        RECT 63.585 165.375 63.755 165.835 ;
        RECT 64.025 164.965 64.300 165.665 ;
        RECT 64.470 165.290 64.725 165.835 ;
        RECT 64.895 165.325 65.375 165.665 ;
        RECT 65.550 165.280 66.155 165.835 ;
        RECT 65.540 165.180 66.155 165.280 ;
        RECT 65.540 165.155 65.725 165.180 ;
        RECT 63.085 164.865 63.855 164.885 ;
        RECT 61.405 164.695 63.855 164.865 ;
        RECT 60.825 164.275 63.335 164.525 ;
        RECT 63.505 164.105 63.855 164.695 ;
        RECT 58.505 163.285 60.175 164.055 ;
        RECT 61.485 163.925 63.855 164.105 ;
        RECT 64.025 163.935 64.195 164.965 ;
        RECT 64.470 164.835 65.225 165.085 ;
        RECT 65.395 164.910 65.725 165.155 ;
        RECT 64.470 164.800 65.240 164.835 ;
        RECT 64.470 164.790 65.255 164.800 ;
        RECT 64.365 164.775 65.260 164.790 ;
        RECT 64.365 164.760 65.280 164.775 ;
        RECT 64.365 164.750 65.300 164.760 ;
        RECT 64.365 164.740 65.325 164.750 ;
        RECT 64.365 164.710 65.395 164.740 ;
        RECT 64.365 164.680 65.415 164.710 ;
        RECT 64.365 164.650 65.435 164.680 ;
        RECT 64.365 164.625 65.465 164.650 ;
        RECT 64.365 164.590 65.500 164.625 ;
        RECT 64.365 164.585 65.530 164.590 ;
        RECT 64.365 164.190 64.595 164.585 ;
        RECT 65.140 164.580 65.530 164.585 ;
        RECT 65.165 164.570 65.530 164.580 ;
        RECT 65.180 164.565 65.530 164.570 ;
        RECT 65.195 164.560 65.530 164.565 ;
        RECT 65.895 164.560 66.155 165.010 ;
        RECT 66.325 164.745 69.835 165.835 ;
        RECT 65.195 164.555 66.155 164.560 ;
        RECT 65.205 164.545 66.155 164.555 ;
        RECT 65.215 164.540 66.155 164.545 ;
        RECT 65.225 164.530 66.155 164.540 ;
        RECT 65.230 164.520 66.155 164.530 ;
        RECT 65.235 164.515 66.155 164.520 ;
        RECT 65.245 164.500 66.155 164.515 ;
        RECT 65.250 164.485 66.155 164.500 ;
        RECT 65.260 164.460 66.155 164.485 ;
        RECT 64.765 163.990 65.095 164.415 ;
        RECT 64.845 163.965 65.095 163.990 ;
        RECT 60.850 163.285 61.115 163.745 ;
        RECT 61.485 163.455 61.655 163.925 ;
        RECT 61.905 163.285 62.075 163.745 ;
        RECT 62.325 163.455 62.495 163.925 ;
        RECT 62.745 163.285 62.915 163.745 ;
        RECT 63.165 163.455 63.335 163.925 ;
        RECT 63.505 163.285 63.755 163.750 ;
        RECT 64.025 163.455 64.285 163.935 ;
        RECT 64.455 163.285 64.705 163.825 ;
        RECT 64.875 163.505 65.095 163.965 ;
        RECT 65.265 164.390 66.155 164.460 ;
        RECT 65.265 163.665 65.435 164.390 ;
        RECT 65.605 163.835 66.155 164.220 ;
        RECT 66.325 164.055 67.975 164.575 ;
        RECT 68.145 164.225 69.835 164.745 ;
        RECT 70.005 164.670 70.295 165.835 ;
        RECT 70.465 165.400 75.810 165.835 ;
        RECT 75.985 165.400 81.330 165.835 ;
        RECT 65.265 163.495 66.155 163.665 ;
        RECT 66.325 163.285 69.835 164.055 ;
        RECT 70.005 163.285 70.295 164.010 ;
        RECT 72.050 163.830 72.390 164.660 ;
        RECT 73.870 164.150 74.220 165.400 ;
        RECT 77.570 163.830 77.910 164.660 ;
        RECT 79.390 164.150 79.740 165.400 ;
        RECT 81.505 164.745 82.715 165.835 ;
        RECT 81.505 164.035 82.025 164.575 ;
        RECT 82.195 164.205 82.715 164.745 ;
        RECT 82.885 164.745 84.095 165.835 ;
        RECT 82.885 164.205 83.405 164.745 ;
        RECT 83.575 164.035 84.095 164.575 ;
        RECT 70.465 163.285 75.810 163.830 ;
        RECT 75.985 163.285 81.330 163.830 ;
        RECT 81.505 163.285 82.715 164.035 ;
        RECT 82.885 163.285 84.095 164.035 ;
        RECT 5.520 163.115 84.180 163.285 ;
        RECT 5.605 162.365 6.815 163.115 ;
        RECT 6.985 162.570 12.330 163.115 ;
        RECT 5.605 161.825 6.125 162.365 ;
        RECT 6.295 161.655 6.815 162.195 ;
        RECT 8.570 161.740 8.910 162.570 ;
        RECT 12.505 162.345 16.015 163.115 ;
        RECT 16.350 162.605 16.590 163.115 ;
        RECT 16.770 162.605 17.050 162.935 ;
        RECT 17.280 162.605 17.495 163.115 ;
        RECT 5.605 160.565 6.815 161.655 ;
        RECT 10.390 161.000 10.740 162.250 ;
        RECT 12.505 161.825 14.155 162.345 ;
        RECT 14.325 161.655 16.015 162.175 ;
        RECT 16.245 161.875 16.600 162.435 ;
        RECT 16.770 161.705 16.940 162.605 ;
        RECT 17.110 161.875 17.375 162.435 ;
        RECT 17.665 162.375 18.280 162.945 ;
        RECT 17.625 161.705 17.795 162.205 ;
        RECT 6.985 160.565 12.330 161.000 ;
        RECT 12.505 160.565 16.015 161.655 ;
        RECT 16.370 161.535 17.795 161.705 ;
        RECT 16.370 161.360 16.760 161.535 ;
        RECT 17.245 160.565 17.575 161.365 ;
        RECT 17.965 161.355 18.280 162.375 ;
        RECT 17.745 160.735 18.280 161.355 ;
        RECT 18.485 162.395 18.825 162.905 ;
        RECT 18.485 160.995 18.745 162.395 ;
        RECT 18.995 162.315 19.265 163.115 ;
        RECT 18.920 161.875 19.250 162.125 ;
        RECT 19.445 161.875 19.725 162.845 ;
        RECT 19.905 161.875 20.205 162.845 ;
        RECT 20.385 161.875 20.735 162.840 ;
        RECT 20.955 162.615 21.450 162.945 ;
        RECT 21.950 162.635 22.250 163.115 ;
        RECT 18.935 161.705 19.250 161.875 ;
        RECT 20.955 161.705 21.125 162.615 ;
        RECT 22.420 162.465 22.680 162.920 ;
        RECT 22.850 162.635 23.110 163.115 ;
        RECT 23.280 162.465 23.540 162.920 ;
        RECT 23.710 162.635 23.970 163.115 ;
        RECT 24.140 162.465 24.400 162.920 ;
        RECT 24.570 162.635 24.830 163.115 ;
        RECT 25.000 162.465 25.260 162.920 ;
        RECT 25.430 162.590 25.690 163.115 ;
        RECT 18.935 161.535 21.125 161.705 ;
        RECT 18.485 160.735 18.825 160.995 ;
        RECT 18.995 160.565 19.325 161.365 ;
        RECT 19.790 160.735 20.040 161.535 ;
        RECT 20.225 160.565 20.555 161.285 ;
        RECT 20.775 160.735 21.025 161.535 ;
        RECT 21.295 161.125 21.535 162.435 ;
        RECT 21.950 162.295 25.260 162.465 ;
        RECT 21.950 161.705 22.920 162.295 ;
        RECT 25.860 162.125 26.110 162.935 ;
        RECT 26.290 162.655 26.535 163.115 ;
        RECT 23.090 161.875 26.110 162.125 ;
        RECT 26.280 161.875 26.595 162.485 ;
        RECT 21.950 161.465 25.260 161.705 ;
        RECT 21.195 160.565 21.530 160.945 ;
        RECT 21.955 160.565 22.250 161.295 ;
        RECT 22.420 160.740 22.680 161.465 ;
        RECT 22.850 160.565 23.110 161.295 ;
        RECT 23.280 160.740 23.540 161.465 ;
        RECT 23.710 160.565 23.970 161.295 ;
        RECT 24.140 160.740 24.400 161.465 ;
        RECT 24.570 160.565 24.830 161.295 ;
        RECT 25.000 160.740 25.260 161.465 ;
        RECT 25.430 160.565 25.690 161.675 ;
        RECT 25.860 160.740 26.110 161.875 ;
        RECT 26.290 160.565 26.585 161.675 ;
        RECT 26.775 160.745 27.035 162.935 ;
        RECT 27.295 162.745 27.965 163.115 ;
        RECT 28.145 162.565 28.455 162.935 ;
        RECT 27.225 162.365 28.455 162.565 ;
        RECT 27.225 161.695 27.515 162.365 ;
        RECT 28.635 162.185 28.865 162.825 ;
        RECT 29.045 162.385 29.335 163.115 ;
        RECT 29.525 162.345 31.195 163.115 ;
        RECT 31.365 162.390 31.655 163.115 ;
        RECT 31.825 162.570 37.170 163.115 ;
        RECT 37.345 162.570 42.690 163.115 ;
        RECT 42.865 162.570 48.210 163.115 ;
        RECT 27.695 161.875 28.160 162.185 ;
        RECT 28.340 161.875 28.865 162.185 ;
        RECT 29.045 161.875 29.345 162.205 ;
        RECT 29.525 161.825 30.275 162.345 ;
        RECT 27.225 161.475 27.995 161.695 ;
        RECT 27.205 160.565 27.545 161.295 ;
        RECT 27.725 160.745 27.995 161.475 ;
        RECT 28.175 161.455 29.335 161.695 ;
        RECT 30.445 161.655 31.195 162.175 ;
        RECT 33.410 161.740 33.750 162.570 ;
        RECT 28.175 160.745 28.405 161.455 ;
        RECT 28.575 160.565 28.905 161.275 ;
        RECT 29.075 160.745 29.335 161.455 ;
        RECT 29.525 160.565 31.195 161.655 ;
        RECT 31.365 160.565 31.655 161.730 ;
        RECT 35.230 161.000 35.580 162.250 ;
        RECT 38.930 161.740 39.270 162.570 ;
        RECT 40.750 161.000 41.100 162.250 ;
        RECT 44.450 161.740 44.790 162.570 ;
        RECT 48.385 162.345 50.055 163.115 ;
        RECT 50.395 162.655 50.650 163.115 ;
        RECT 50.820 162.485 51.150 162.945 ;
        RECT 51.320 162.655 51.490 163.115 ;
        RECT 51.660 162.485 51.990 162.945 ;
        RECT 52.160 162.655 52.330 163.115 ;
        RECT 52.500 162.485 52.830 162.945 ;
        RECT 53.000 162.655 53.170 163.115 ;
        RECT 53.340 162.485 53.670 162.945 ;
        RECT 53.840 162.655 54.145 163.115 ;
        RECT 46.270 161.000 46.620 162.250 ;
        RECT 48.385 161.825 49.135 162.345 ;
        RECT 50.225 162.295 54.195 162.485 ;
        RECT 54.830 162.465 55.100 162.675 ;
        RECT 55.320 162.655 55.650 163.115 ;
        RECT 56.160 162.655 56.910 162.945 ;
        RECT 54.830 162.295 56.165 162.465 ;
        RECT 49.305 161.655 50.055 162.175 ;
        RECT 31.825 160.565 37.170 161.000 ;
        RECT 37.345 160.565 42.690 161.000 ;
        RECT 42.865 160.565 48.210 161.000 ;
        RECT 48.385 160.565 50.055 161.655 ;
        RECT 50.225 161.705 50.570 162.295 ;
        RECT 50.820 162.095 53.675 162.125 ;
        RECT 50.745 161.925 53.675 162.095 ;
        RECT 50.820 161.875 53.675 161.925 ;
        RECT 53.875 161.705 54.195 162.295 ;
        RECT 55.995 162.125 56.165 162.295 ;
        RECT 54.830 161.885 55.180 162.125 ;
        RECT 55.350 161.885 55.825 162.125 ;
        RECT 55.995 161.875 56.370 162.125 ;
        RECT 55.995 161.705 56.165 161.875 ;
        RECT 50.225 161.535 54.195 161.705 ;
        RECT 54.830 161.535 56.165 161.705 ;
        RECT 50.395 160.565 50.650 161.365 ;
        RECT 50.820 160.735 51.150 161.535 ;
        RECT 51.320 160.565 51.490 161.365 ;
        RECT 51.660 160.735 51.990 161.535 ;
        RECT 52.160 160.565 52.330 161.365 ;
        RECT 52.500 160.735 52.830 161.535 ;
        RECT 53.000 160.565 53.170 161.365 ;
        RECT 53.340 160.735 53.670 161.535 ;
        RECT 54.830 161.375 55.110 161.535 ;
        RECT 56.540 161.365 56.910 162.655 ;
        RECT 57.125 162.390 57.415 163.115 ;
        RECT 57.585 162.615 57.885 162.945 ;
        RECT 58.055 162.635 58.330 163.115 ;
        RECT 53.840 160.565 54.140 161.365 ;
        RECT 55.320 160.565 55.570 161.365 ;
        RECT 55.740 161.195 56.910 161.365 ;
        RECT 55.740 160.735 56.070 161.195 ;
        RECT 56.240 160.565 56.455 161.025 ;
        RECT 57.125 160.565 57.415 161.730 ;
        RECT 57.585 161.705 57.755 162.615 ;
        RECT 58.510 162.465 58.805 162.855 ;
        RECT 58.975 162.635 59.230 163.115 ;
        RECT 59.405 162.465 59.665 162.855 ;
        RECT 59.835 162.635 60.115 163.115 ;
        RECT 60.865 162.655 61.110 163.115 ;
        RECT 57.925 161.875 58.275 162.445 ;
        RECT 58.510 162.295 60.160 162.465 ;
        RECT 58.445 161.955 59.585 162.125 ;
        RECT 58.445 161.705 58.615 161.955 ;
        RECT 59.755 161.785 60.160 162.295 ;
        RECT 60.805 161.875 61.120 162.485 ;
        RECT 61.290 162.125 61.540 162.935 ;
        RECT 61.710 162.590 61.970 163.115 ;
        RECT 62.140 162.465 62.400 162.920 ;
        RECT 62.570 162.635 62.830 163.115 ;
        RECT 63.000 162.465 63.260 162.920 ;
        RECT 63.430 162.635 63.690 163.115 ;
        RECT 63.860 162.465 64.120 162.920 ;
        RECT 64.290 162.635 64.550 163.115 ;
        RECT 64.720 162.465 64.980 162.920 ;
        RECT 65.150 162.635 65.450 163.115 ;
        RECT 65.865 162.570 71.210 163.115 ;
        RECT 71.385 162.570 76.730 163.115 ;
        RECT 76.905 162.570 82.250 163.115 ;
        RECT 62.140 162.295 65.450 162.465 ;
        RECT 61.290 161.875 64.310 162.125 ;
        RECT 57.585 161.535 58.615 161.705 ;
        RECT 59.405 161.615 60.160 161.785 ;
        RECT 57.585 160.735 57.895 161.535 ;
        RECT 59.405 161.365 59.665 161.615 ;
        RECT 58.065 160.565 58.375 161.365 ;
        RECT 58.545 161.195 59.665 161.365 ;
        RECT 58.545 160.735 58.805 161.195 ;
        RECT 58.975 160.565 59.230 161.025 ;
        RECT 59.405 160.735 59.665 161.195 ;
        RECT 59.835 160.565 60.120 161.435 ;
        RECT 60.815 160.565 61.110 161.675 ;
        RECT 61.290 160.740 61.540 161.875 ;
        RECT 64.480 161.705 65.450 162.295 ;
        RECT 67.450 161.740 67.790 162.570 ;
        RECT 61.710 160.565 61.970 161.675 ;
        RECT 62.140 161.465 65.450 161.705 ;
        RECT 62.140 160.740 62.400 161.465 ;
        RECT 62.570 160.565 62.830 161.295 ;
        RECT 63.000 160.740 63.260 161.465 ;
        RECT 63.430 160.565 63.690 161.295 ;
        RECT 63.860 160.740 64.120 161.465 ;
        RECT 64.290 160.565 64.550 161.295 ;
        RECT 64.720 160.740 64.980 161.465 ;
        RECT 65.150 160.565 65.445 161.295 ;
        RECT 69.270 161.000 69.620 162.250 ;
        RECT 72.970 161.740 73.310 162.570 ;
        RECT 74.790 161.000 75.140 162.250 ;
        RECT 78.490 161.740 78.830 162.570 ;
        RECT 82.885 162.365 84.095 163.115 ;
        RECT 80.310 161.000 80.660 162.250 ;
        RECT 82.885 161.655 83.405 162.195 ;
        RECT 83.575 161.825 84.095 162.365 ;
        RECT 65.865 160.565 71.210 161.000 ;
        RECT 71.385 160.565 76.730 161.000 ;
        RECT 76.905 160.565 82.250 161.000 ;
        RECT 82.885 160.565 84.095 161.655 ;
        RECT 5.520 160.395 84.180 160.565 ;
        RECT 5.605 159.305 6.815 160.395 ;
        RECT 6.985 159.960 12.330 160.395 ;
        RECT 12.505 159.960 17.850 160.395 ;
        RECT 5.605 158.595 6.125 159.135 ;
        RECT 6.295 158.765 6.815 159.305 ;
        RECT 5.605 157.845 6.815 158.595 ;
        RECT 8.570 158.390 8.910 159.220 ;
        RECT 10.390 158.710 10.740 159.960 ;
        RECT 14.090 158.390 14.430 159.220 ;
        RECT 15.910 158.710 16.260 159.960 ;
        RECT 18.485 159.230 18.775 160.395 ;
        RECT 18.945 159.885 19.205 160.395 ;
        RECT 18.945 158.835 19.285 159.715 ;
        RECT 19.455 159.005 19.625 160.225 ;
        RECT 19.865 159.890 20.480 160.395 ;
        RECT 19.865 159.355 20.115 159.720 ;
        RECT 20.285 159.715 20.480 159.890 ;
        RECT 20.650 159.885 21.125 160.225 ;
        RECT 21.295 159.850 21.510 160.395 ;
        RECT 20.285 159.525 20.615 159.715 ;
        RECT 20.835 159.355 21.550 159.650 ;
        RECT 21.720 159.525 21.995 160.225 ;
        RECT 19.865 159.185 21.655 159.355 ;
        RECT 19.455 158.755 20.250 159.005 ;
        RECT 19.455 158.665 19.705 158.755 ;
        RECT 6.985 157.845 12.330 158.390 ;
        RECT 12.505 157.845 17.850 158.390 ;
        RECT 18.485 157.845 18.775 158.570 ;
        RECT 18.945 157.845 19.205 158.665 ;
        RECT 19.375 158.245 19.705 158.665 ;
        RECT 20.420 158.330 20.675 159.185 ;
        RECT 19.885 158.065 20.675 158.330 ;
        RECT 20.845 158.485 21.255 159.005 ;
        RECT 21.425 158.755 21.655 159.185 ;
        RECT 21.825 158.495 21.995 159.525 ;
        RECT 22.350 159.425 22.740 159.600 ;
        RECT 23.225 159.595 23.555 160.395 ;
        RECT 23.725 159.605 24.260 160.225 ;
        RECT 22.350 159.255 23.775 159.425 ;
        RECT 22.225 158.525 22.580 159.085 ;
        RECT 20.845 158.065 21.045 158.485 ;
        RECT 21.235 157.845 21.565 158.305 ;
        RECT 21.735 158.015 21.995 158.495 ;
        RECT 22.750 158.355 22.920 159.255 ;
        RECT 23.090 158.525 23.355 159.085 ;
        RECT 23.605 158.755 23.775 159.255 ;
        RECT 23.945 158.585 24.260 159.605 ;
        RECT 25.080 159.385 25.380 160.225 ;
        RECT 25.575 159.555 25.825 160.395 ;
        RECT 26.415 159.805 27.220 160.225 ;
        RECT 25.995 159.635 27.560 159.805 ;
        RECT 25.995 159.385 26.165 159.635 ;
        RECT 25.080 159.215 26.165 159.385 ;
        RECT 24.925 158.755 25.255 159.045 ;
        RECT 25.425 158.585 25.595 159.215 ;
        RECT 26.335 159.085 26.655 159.465 ;
        RECT 26.845 159.375 27.220 159.465 ;
        RECT 26.825 159.205 27.220 159.375 ;
        RECT 27.390 159.385 27.560 159.635 ;
        RECT 27.730 159.555 28.060 160.395 ;
        RECT 28.230 159.635 28.895 160.225 ;
        RECT 27.390 159.215 28.310 159.385 ;
        RECT 25.765 158.835 26.095 159.045 ;
        RECT 26.275 158.835 26.655 159.085 ;
        RECT 26.845 159.045 27.220 159.205 ;
        RECT 28.140 159.045 28.310 159.215 ;
        RECT 26.845 158.835 27.330 159.045 ;
        RECT 27.520 158.835 27.970 159.045 ;
        RECT 28.140 158.835 28.475 159.045 ;
        RECT 28.645 158.665 28.895 159.635 ;
        RECT 22.330 157.845 22.570 158.355 ;
        RECT 22.750 158.025 23.030 158.355 ;
        RECT 23.260 157.845 23.475 158.355 ;
        RECT 23.645 158.015 24.260 158.585 ;
        RECT 25.085 158.405 25.595 158.585 ;
        RECT 26.000 158.495 27.700 158.665 ;
        RECT 26.000 158.405 26.385 158.495 ;
        RECT 25.085 158.015 25.415 158.405 ;
        RECT 25.585 158.065 26.770 158.235 ;
        RECT 27.030 157.845 27.200 158.315 ;
        RECT 27.370 158.030 27.700 158.495 ;
        RECT 27.870 157.845 28.040 158.665 ;
        RECT 28.210 158.025 28.895 158.665 ;
        RECT 29.065 158.790 29.345 160.225 ;
        RECT 29.515 159.620 30.225 160.395 ;
        RECT 30.395 159.450 30.725 160.225 ;
        RECT 29.575 159.235 30.725 159.450 ;
        RECT 29.065 158.015 29.405 158.790 ;
        RECT 29.575 158.665 29.860 159.235 ;
        RECT 30.045 158.835 30.515 159.065 ;
        RECT 30.920 159.035 31.135 160.150 ;
        RECT 31.315 159.675 31.645 160.395 ;
        RECT 32.765 159.885 33.065 160.395 ;
        RECT 33.235 159.885 33.615 160.055 ;
        RECT 34.195 159.885 34.825 160.395 ;
        RECT 33.235 159.715 33.405 159.885 ;
        RECT 34.995 159.715 35.325 160.225 ;
        RECT 35.495 159.885 35.795 160.395 ;
        RECT 32.745 159.515 33.405 159.715 ;
        RECT 33.575 159.545 35.795 159.715 ;
        RECT 31.425 159.035 31.655 159.375 ;
        RECT 30.685 158.855 31.135 159.035 ;
        RECT 30.685 158.835 31.015 158.855 ;
        RECT 31.325 158.835 31.655 159.035 ;
        RECT 29.575 158.475 30.285 158.665 ;
        RECT 29.985 158.335 30.285 158.475 ;
        RECT 30.475 158.475 31.655 158.665 ;
        RECT 30.475 158.395 30.805 158.475 ;
        RECT 29.985 158.325 30.300 158.335 ;
        RECT 29.985 158.315 30.310 158.325 ;
        RECT 29.985 158.310 30.320 158.315 ;
        RECT 29.575 157.845 29.745 158.305 ;
        RECT 29.985 158.300 30.325 158.310 ;
        RECT 29.985 158.295 30.330 158.300 ;
        RECT 29.985 158.285 30.335 158.295 ;
        RECT 29.985 158.280 30.340 158.285 ;
        RECT 29.985 158.015 30.345 158.280 ;
        RECT 30.975 157.845 31.145 158.305 ;
        RECT 31.315 158.015 31.655 158.475 ;
        RECT 32.745 158.585 32.915 159.515 ;
        RECT 33.575 159.345 33.745 159.545 ;
        RECT 33.085 159.175 33.745 159.345 ;
        RECT 33.915 159.205 35.455 159.375 ;
        RECT 33.085 158.755 33.255 159.175 ;
        RECT 33.915 159.005 34.085 159.205 ;
        RECT 33.485 158.835 34.085 159.005 ;
        RECT 34.255 158.835 34.950 159.035 ;
        RECT 35.210 158.755 35.455 159.205 ;
        RECT 33.575 158.585 34.485 158.665 ;
        RECT 32.745 158.105 33.065 158.585 ;
        RECT 33.235 158.495 34.485 158.585 ;
        RECT 33.235 158.415 33.745 158.495 ;
        RECT 33.235 158.015 33.465 158.415 ;
        RECT 33.635 157.845 33.985 158.235 ;
        RECT 34.155 158.015 34.485 158.495 ;
        RECT 34.655 157.845 34.825 158.665 ;
        RECT 35.625 158.585 35.795 159.545 ;
        RECT 35.965 159.305 38.555 160.395 ;
        RECT 39.190 159.970 39.525 160.395 ;
        RECT 39.695 159.790 39.880 160.195 ;
        RECT 35.330 158.040 35.795 158.585 ;
        RECT 35.965 158.615 37.175 159.135 ;
        RECT 37.345 158.785 38.555 159.305 ;
        RECT 39.215 159.615 39.880 159.790 ;
        RECT 40.085 159.615 40.415 160.395 ;
        RECT 35.965 157.845 38.555 158.615 ;
        RECT 39.215 158.585 39.555 159.615 ;
        RECT 40.585 159.425 40.855 160.195 ;
        RECT 39.725 159.255 40.855 159.425 ;
        RECT 39.725 158.755 39.975 159.255 ;
        RECT 39.215 158.415 39.900 158.585 ;
        RECT 40.155 158.505 40.515 159.085 ;
        RECT 39.190 157.845 39.525 158.245 ;
        RECT 39.695 158.015 39.900 158.415 ;
        RECT 40.685 158.345 40.855 159.255 ;
        RECT 40.110 157.845 40.385 158.325 ;
        RECT 40.595 158.015 40.855 158.345 ;
        RECT 41.035 159.335 41.365 160.185 ;
        RECT 41.035 158.570 41.225 159.335 ;
        RECT 41.535 159.255 41.785 160.395 ;
        RECT 41.975 159.755 42.225 160.175 ;
        RECT 42.455 159.925 42.785 160.395 ;
        RECT 43.015 159.755 43.265 160.175 ;
        RECT 41.975 159.585 43.265 159.755 ;
        RECT 43.445 159.755 43.775 160.185 ;
        RECT 43.445 159.585 43.900 159.755 ;
        RECT 41.965 159.085 42.180 159.415 ;
        RECT 41.395 158.755 41.705 159.085 ;
        RECT 41.875 158.755 42.180 159.085 ;
        RECT 42.355 158.755 42.640 159.415 ;
        RECT 42.835 158.755 43.100 159.415 ;
        RECT 43.315 158.755 43.560 159.415 ;
        RECT 41.535 158.585 41.705 158.755 ;
        RECT 43.730 158.585 43.900 159.585 ;
        RECT 44.245 159.230 44.535 160.395 ;
        RECT 44.705 159.305 45.915 160.395 ;
        RECT 41.035 158.060 41.365 158.570 ;
        RECT 41.535 158.415 43.900 158.585 ;
        RECT 44.705 158.595 45.225 159.135 ;
        RECT 45.395 158.765 45.915 159.305 ;
        RECT 46.120 159.605 46.655 160.225 ;
        RECT 41.535 157.845 41.865 158.245 ;
        RECT 42.915 158.075 43.245 158.415 ;
        RECT 43.415 157.845 43.745 158.245 ;
        RECT 44.245 157.845 44.535 158.570 ;
        RECT 44.705 157.845 45.915 158.595 ;
        RECT 46.120 158.585 46.435 159.605 ;
        RECT 46.825 159.595 47.155 160.395 ;
        RECT 47.640 159.425 48.030 159.600 ;
        RECT 46.605 159.255 48.030 159.425 ;
        RECT 48.475 159.465 48.645 160.225 ;
        RECT 48.860 159.635 49.190 160.395 ;
        RECT 48.475 159.295 49.190 159.465 ;
        RECT 49.360 159.320 49.615 160.225 ;
        RECT 46.605 158.755 46.775 159.255 ;
        RECT 46.120 158.015 46.735 158.585 ;
        RECT 47.025 158.525 47.290 159.085 ;
        RECT 47.460 158.355 47.630 159.255 ;
        RECT 47.800 158.525 48.155 159.085 ;
        RECT 48.385 158.745 48.740 159.115 ;
        RECT 49.020 159.085 49.190 159.295 ;
        RECT 49.020 158.755 49.275 159.085 ;
        RECT 49.020 158.565 49.190 158.755 ;
        RECT 49.445 158.590 49.615 159.320 ;
        RECT 49.790 159.245 50.050 160.395 ;
        RECT 51.155 159.255 51.485 160.395 ;
        RECT 52.015 159.425 52.345 160.210 ;
        RECT 51.665 159.255 52.345 159.425 ;
        RECT 52.530 160.005 52.865 160.225 ;
        RECT 53.870 160.015 54.225 160.395 ;
        RECT 52.530 159.385 52.785 160.005 ;
        RECT 53.035 159.845 53.265 159.885 ;
        RECT 54.395 159.845 54.645 160.225 ;
        RECT 53.035 159.645 54.645 159.845 ;
        RECT 53.035 159.555 53.220 159.645 ;
        RECT 53.810 159.635 54.645 159.645 ;
        RECT 54.895 159.615 55.145 160.395 ;
        RECT 55.315 159.545 55.575 160.225 ;
        RECT 56.245 159.935 56.460 160.395 ;
        RECT 56.630 159.765 56.960 160.225 ;
        RECT 53.375 159.445 53.705 159.475 ;
        RECT 53.375 159.385 55.175 159.445 ;
        RECT 52.530 159.275 55.235 159.385 ;
        RECT 51.145 158.835 51.495 159.085 ;
        RECT 48.475 158.395 49.190 158.565 ;
        RECT 46.905 157.845 47.120 158.355 ;
        RECT 47.350 158.025 47.630 158.355 ;
        RECT 47.810 157.845 48.050 158.355 ;
        RECT 48.475 158.015 48.645 158.395 ;
        RECT 48.860 157.845 49.190 158.225 ;
        RECT 49.360 158.015 49.615 158.590 ;
        RECT 49.790 157.845 50.050 158.685 ;
        RECT 51.665 158.655 51.835 159.255 ;
        RECT 52.530 159.215 53.705 159.275 ;
        RECT 55.035 159.240 55.235 159.275 ;
        RECT 52.005 158.835 52.355 159.085 ;
        RECT 52.525 158.835 53.015 159.035 ;
        RECT 53.205 158.835 53.680 159.045 ;
        RECT 51.155 157.845 51.425 158.655 ;
        RECT 51.595 158.015 51.925 158.655 ;
        RECT 52.095 157.845 52.335 158.655 ;
        RECT 52.530 157.845 52.985 158.610 ;
        RECT 53.460 158.435 53.680 158.835 ;
        RECT 53.925 158.835 54.255 159.045 ;
        RECT 53.925 158.435 54.135 158.835 ;
        RECT 54.425 158.800 54.835 159.105 ;
        RECT 55.065 158.665 55.235 159.240 ;
        RECT 54.965 158.545 55.235 158.665 ;
        RECT 54.390 158.500 55.235 158.545 ;
        RECT 54.390 158.375 55.145 158.500 ;
        RECT 54.390 158.225 54.560 158.375 ;
        RECT 55.405 158.355 55.575 159.545 ;
        RECT 55.345 158.345 55.575 158.355 ;
        RECT 53.260 158.015 54.560 158.225 ;
        RECT 54.815 157.845 55.145 158.205 ;
        RECT 55.315 158.015 55.575 158.345 ;
        RECT 55.790 159.595 56.960 159.765 ;
        RECT 57.130 159.595 57.380 160.395 ;
        RECT 55.790 158.305 56.160 159.595 ;
        RECT 57.590 159.425 57.870 159.585 ;
        RECT 56.535 159.255 57.870 159.425 ;
        RECT 58.045 159.305 59.715 160.395 ;
        RECT 56.535 159.085 56.705 159.255 ;
        RECT 56.330 158.835 56.705 159.085 ;
        RECT 56.875 158.835 57.350 159.075 ;
        RECT 57.520 158.835 57.870 159.075 ;
        RECT 56.535 158.665 56.705 158.835 ;
        RECT 56.535 158.495 57.870 158.665 ;
        RECT 55.790 158.015 56.540 158.305 ;
        RECT 57.050 157.845 57.380 158.305 ;
        RECT 57.600 158.285 57.870 158.495 ;
        RECT 58.045 158.615 58.795 159.135 ;
        RECT 58.965 158.785 59.715 159.305 ;
        RECT 59.885 159.545 60.265 160.225 ;
        RECT 60.855 159.545 61.025 160.395 ;
        RECT 61.195 159.715 61.525 160.225 ;
        RECT 61.695 159.885 61.865 160.395 ;
        RECT 62.035 159.715 62.435 160.225 ;
        RECT 61.195 159.545 62.435 159.715 ;
        RECT 58.045 157.845 59.715 158.615 ;
        RECT 59.885 158.585 60.055 159.545 ;
        RECT 60.225 159.205 61.530 159.375 ;
        RECT 62.615 159.295 62.935 160.225 ;
        RECT 63.190 159.775 63.365 160.225 ;
        RECT 63.535 159.955 63.865 160.395 ;
        RECT 64.170 159.805 64.340 160.225 ;
        RECT 64.575 159.985 65.245 160.395 ;
        RECT 65.460 159.805 65.630 160.225 ;
        RECT 65.830 159.985 66.160 160.395 ;
        RECT 63.190 159.605 63.820 159.775 ;
        RECT 60.225 158.755 60.470 159.205 ;
        RECT 60.640 158.835 61.190 159.035 ;
        RECT 61.360 159.005 61.530 159.205 ;
        RECT 62.305 159.125 62.935 159.295 ;
        RECT 61.360 158.835 61.735 159.005 ;
        RECT 61.905 158.585 62.135 159.085 ;
        RECT 59.885 158.415 62.135 158.585 ;
        RECT 59.935 157.845 60.265 158.235 ;
        RECT 60.435 158.095 60.605 158.415 ;
        RECT 62.305 158.245 62.475 159.125 ;
        RECT 63.105 158.755 63.470 159.435 ;
        RECT 63.650 159.085 63.820 159.605 ;
        RECT 64.170 159.635 66.185 159.805 ;
        RECT 63.650 158.755 64.000 159.085 ;
        RECT 60.775 157.845 61.105 158.235 ;
        RECT 61.520 158.075 62.475 158.245 ;
        RECT 62.645 157.845 62.935 158.680 ;
        RECT 63.650 158.585 63.820 158.755 ;
        RECT 63.190 158.415 63.820 158.585 ;
        RECT 63.190 158.015 63.365 158.415 ;
        RECT 64.170 158.345 64.340 159.635 ;
        RECT 63.535 157.845 63.865 158.225 ;
        RECT 64.110 158.015 64.340 158.345 ;
        RECT 64.540 158.180 64.820 159.455 ;
        RECT 65.045 159.035 65.315 159.455 ;
        RECT 65.005 158.865 65.315 159.035 ;
        RECT 65.045 158.180 65.315 158.865 ;
        RECT 65.505 158.425 65.845 159.455 ;
        RECT 66.015 159.085 66.185 159.635 ;
        RECT 66.355 159.255 66.615 160.225 ;
        RECT 66.785 159.305 69.375 160.395 ;
        RECT 66.015 158.755 66.275 159.085 ;
        RECT 66.445 158.565 66.615 159.255 ;
        RECT 65.775 157.845 66.105 158.225 ;
        RECT 66.275 158.100 66.615 158.565 ;
        RECT 66.785 158.615 67.995 159.135 ;
        RECT 68.165 158.785 69.375 159.305 ;
        RECT 70.005 159.230 70.295 160.395 ;
        RECT 70.465 159.960 75.810 160.395 ;
        RECT 75.985 159.960 81.330 160.395 ;
        RECT 66.275 158.055 66.610 158.100 ;
        RECT 66.785 157.845 69.375 158.615 ;
        RECT 70.005 157.845 70.295 158.570 ;
        RECT 72.050 158.390 72.390 159.220 ;
        RECT 73.870 158.710 74.220 159.960 ;
        RECT 77.570 158.390 77.910 159.220 ;
        RECT 79.390 158.710 79.740 159.960 ;
        RECT 81.505 159.305 82.715 160.395 ;
        RECT 81.505 158.595 82.025 159.135 ;
        RECT 82.195 158.765 82.715 159.305 ;
        RECT 82.885 159.305 84.095 160.395 ;
        RECT 82.885 158.765 83.405 159.305 ;
        RECT 83.575 158.595 84.095 159.135 ;
        RECT 70.465 157.845 75.810 158.390 ;
        RECT 75.985 157.845 81.330 158.390 ;
        RECT 81.505 157.845 82.715 158.595 ;
        RECT 82.885 157.845 84.095 158.595 ;
        RECT 5.520 157.675 84.180 157.845 ;
        RECT 5.605 156.925 6.815 157.675 ;
        RECT 6.985 157.130 12.330 157.675 ;
        RECT 5.605 156.385 6.125 156.925 ;
        RECT 6.295 156.215 6.815 156.755 ;
        RECT 8.570 156.300 8.910 157.130 ;
        RECT 12.505 156.905 16.015 157.675 ;
        RECT 16.695 157.020 17.025 157.455 ;
        RECT 17.195 157.065 17.365 157.675 ;
        RECT 16.645 156.935 17.025 157.020 ;
        RECT 17.535 156.935 17.865 157.460 ;
        RECT 18.125 157.145 18.335 157.675 ;
        RECT 18.610 157.225 19.395 157.395 ;
        RECT 19.565 157.225 19.970 157.395 ;
        RECT 5.605 155.125 6.815 156.215 ;
        RECT 10.390 155.560 10.740 156.810 ;
        RECT 12.505 156.385 14.155 156.905 ;
        RECT 16.645 156.895 16.870 156.935 ;
        RECT 14.325 156.215 16.015 156.735 ;
        RECT 6.985 155.125 12.330 155.560 ;
        RECT 12.505 155.125 16.015 156.215 ;
        RECT 16.645 156.315 16.815 156.895 ;
        RECT 17.535 156.765 17.735 156.935 ;
        RECT 18.610 156.765 18.780 157.225 ;
        RECT 16.985 156.435 17.735 156.765 ;
        RECT 17.905 156.435 18.780 156.765 ;
        RECT 16.645 156.265 16.860 156.315 ;
        RECT 16.645 156.185 17.035 156.265 ;
        RECT 16.705 155.340 17.035 156.185 ;
        RECT 17.545 156.230 17.735 156.435 ;
        RECT 17.205 155.125 17.375 156.135 ;
        RECT 17.545 155.855 18.440 156.230 ;
        RECT 17.545 155.295 17.885 155.855 ;
        RECT 18.115 155.125 18.430 155.625 ;
        RECT 18.610 155.595 18.780 156.435 ;
        RECT 18.950 156.725 19.415 157.055 ;
        RECT 19.800 156.995 19.970 157.225 ;
        RECT 20.150 157.175 20.520 157.675 ;
        RECT 20.840 157.225 21.515 157.395 ;
        RECT 21.710 157.225 22.045 157.395 ;
        RECT 18.950 155.765 19.270 156.725 ;
        RECT 19.800 156.695 20.630 156.995 ;
        RECT 19.440 155.795 19.630 156.515 ;
        RECT 19.800 155.625 19.970 156.695 ;
        RECT 20.430 156.665 20.630 156.695 ;
        RECT 20.140 156.445 20.310 156.515 ;
        RECT 20.840 156.445 21.010 157.225 ;
        RECT 21.875 157.085 22.045 157.225 ;
        RECT 22.215 157.215 22.465 157.675 ;
        RECT 20.140 156.275 21.010 156.445 ;
        RECT 21.180 156.805 21.705 157.025 ;
        RECT 21.875 156.955 22.100 157.085 ;
        RECT 20.140 156.185 20.650 156.275 ;
        RECT 18.610 155.425 19.495 155.595 ;
        RECT 19.720 155.295 19.970 155.625 ;
        RECT 20.140 155.125 20.310 155.925 ;
        RECT 20.480 155.570 20.650 156.185 ;
        RECT 21.180 156.105 21.350 156.805 ;
        RECT 20.820 155.740 21.350 156.105 ;
        RECT 21.520 156.040 21.760 156.635 ;
        RECT 21.930 155.850 22.100 156.955 ;
        RECT 22.270 156.095 22.550 157.045 ;
        RECT 21.795 155.720 22.100 155.850 ;
        RECT 20.480 155.400 21.585 155.570 ;
        RECT 21.795 155.295 22.045 155.720 ;
        RECT 22.215 155.125 22.480 155.585 ;
        RECT 22.720 155.295 22.905 157.415 ;
        RECT 23.075 157.295 23.405 157.675 ;
        RECT 23.575 157.125 23.745 157.415 ;
        RECT 23.080 156.955 23.745 157.125 ;
        RECT 23.080 155.965 23.310 156.955 ;
        RECT 23.480 156.135 23.830 156.785 ;
        RECT 24.925 156.730 25.265 157.505 ;
        RECT 25.435 157.215 25.605 157.675 ;
        RECT 25.845 157.240 26.205 157.505 ;
        RECT 25.845 157.235 26.200 157.240 ;
        RECT 25.845 157.225 26.195 157.235 ;
        RECT 25.845 157.220 26.190 157.225 ;
        RECT 25.845 157.210 26.185 157.220 ;
        RECT 26.835 157.215 27.005 157.675 ;
        RECT 25.845 157.205 26.180 157.210 ;
        RECT 25.845 157.195 26.170 157.205 ;
        RECT 25.845 157.185 26.160 157.195 ;
        RECT 25.845 157.045 26.145 157.185 ;
        RECT 25.435 156.855 26.145 157.045 ;
        RECT 26.335 157.045 26.665 157.125 ;
        RECT 27.175 157.045 27.515 157.505 ;
        RECT 26.335 156.855 27.515 157.045 ;
        RECT 27.685 156.905 29.355 157.675 ;
        RECT 23.080 155.795 23.745 155.965 ;
        RECT 23.075 155.125 23.405 155.625 ;
        RECT 23.575 155.295 23.745 155.795 ;
        RECT 24.925 155.295 25.205 156.730 ;
        RECT 25.435 156.285 25.720 156.855 ;
        RECT 25.905 156.455 26.375 156.685 ;
        RECT 26.545 156.665 26.875 156.685 ;
        RECT 26.545 156.485 26.995 156.665 ;
        RECT 27.185 156.485 27.515 156.685 ;
        RECT 25.435 156.070 26.585 156.285 ;
        RECT 25.375 155.125 26.085 155.900 ;
        RECT 26.255 155.295 26.585 156.070 ;
        RECT 26.780 155.370 26.995 156.485 ;
        RECT 27.285 156.145 27.515 156.485 ;
        RECT 27.685 156.385 28.435 156.905 ;
        RECT 29.985 156.875 30.295 157.675 ;
        RECT 30.500 156.875 31.195 157.505 ;
        RECT 31.365 156.950 31.655 157.675 ;
        RECT 32.375 157.125 32.545 157.415 ;
        RECT 32.715 157.295 33.045 157.675 ;
        RECT 32.375 156.955 33.040 157.125 ;
        RECT 28.605 156.215 29.355 156.735 ;
        RECT 29.995 156.435 30.330 156.705 ;
        RECT 30.500 156.275 30.670 156.875 ;
        RECT 30.840 156.435 31.175 156.685 ;
        RECT 27.175 155.125 27.505 155.845 ;
        RECT 27.685 155.125 29.355 156.215 ;
        RECT 29.985 155.125 30.265 156.265 ;
        RECT 30.435 155.295 30.765 156.275 ;
        RECT 30.935 155.125 31.195 156.265 ;
        RECT 31.365 155.125 31.655 156.290 ;
        RECT 32.290 156.135 32.640 156.785 ;
        RECT 32.810 155.965 33.040 156.955 ;
        RECT 32.375 155.795 33.040 155.965 ;
        RECT 32.375 155.295 32.545 155.795 ;
        RECT 32.715 155.125 33.045 155.625 ;
        RECT 33.215 155.295 33.400 157.415 ;
        RECT 33.655 157.215 33.905 157.675 ;
        RECT 34.075 157.225 34.410 157.395 ;
        RECT 34.605 157.225 35.280 157.395 ;
        RECT 34.075 157.085 34.245 157.225 ;
        RECT 33.570 156.095 33.850 157.045 ;
        RECT 34.020 156.955 34.245 157.085 ;
        RECT 34.020 155.850 34.190 156.955 ;
        RECT 34.415 156.805 34.940 157.025 ;
        RECT 34.360 156.040 34.600 156.635 ;
        RECT 34.770 156.105 34.940 156.805 ;
        RECT 35.110 156.445 35.280 157.225 ;
        RECT 35.600 157.175 35.970 157.675 ;
        RECT 36.150 157.225 36.555 157.395 ;
        RECT 36.725 157.225 37.510 157.395 ;
        RECT 36.150 156.995 36.320 157.225 ;
        RECT 35.490 156.695 36.320 156.995 ;
        RECT 36.705 156.725 37.170 157.055 ;
        RECT 35.490 156.665 35.690 156.695 ;
        RECT 35.810 156.445 35.980 156.515 ;
        RECT 35.110 156.275 35.980 156.445 ;
        RECT 35.470 156.185 35.980 156.275 ;
        RECT 34.020 155.720 34.325 155.850 ;
        RECT 34.770 155.740 35.300 156.105 ;
        RECT 33.640 155.125 33.905 155.585 ;
        RECT 34.075 155.295 34.325 155.720 ;
        RECT 35.470 155.570 35.640 156.185 ;
        RECT 34.535 155.400 35.640 155.570 ;
        RECT 35.810 155.125 35.980 155.925 ;
        RECT 36.150 155.625 36.320 156.695 ;
        RECT 36.490 155.795 36.680 156.515 ;
        RECT 36.850 155.765 37.170 156.725 ;
        RECT 37.340 156.765 37.510 157.225 ;
        RECT 37.785 157.145 37.995 157.675 ;
        RECT 38.255 156.935 38.585 157.460 ;
        RECT 38.755 157.065 38.925 157.675 ;
        RECT 39.095 157.020 39.425 157.455 ;
        RECT 39.735 157.125 39.905 157.415 ;
        RECT 40.075 157.295 40.405 157.675 ;
        RECT 39.095 156.935 39.475 157.020 ;
        RECT 39.735 156.955 40.400 157.125 ;
        RECT 38.385 156.765 38.585 156.935 ;
        RECT 39.250 156.895 39.475 156.935 ;
        RECT 37.340 156.435 38.215 156.765 ;
        RECT 38.385 156.435 39.135 156.765 ;
        RECT 36.150 155.295 36.400 155.625 ;
        RECT 37.340 155.595 37.510 156.435 ;
        RECT 38.385 156.230 38.575 156.435 ;
        RECT 39.305 156.315 39.475 156.895 ;
        RECT 39.260 156.265 39.475 156.315 ;
        RECT 37.680 155.855 38.575 156.230 ;
        RECT 39.085 156.185 39.475 156.265 ;
        RECT 36.625 155.425 37.510 155.595 ;
        RECT 37.690 155.125 38.005 155.625 ;
        RECT 38.235 155.295 38.575 155.855 ;
        RECT 38.745 155.125 38.915 156.135 ;
        RECT 39.085 155.340 39.415 156.185 ;
        RECT 39.650 156.135 40.000 156.785 ;
        RECT 40.170 155.965 40.400 156.955 ;
        RECT 39.735 155.795 40.400 155.965 ;
        RECT 39.735 155.295 39.905 155.795 ;
        RECT 40.075 155.125 40.405 155.625 ;
        RECT 40.575 155.295 40.760 157.415 ;
        RECT 41.015 157.215 41.265 157.675 ;
        RECT 41.435 157.225 41.770 157.395 ;
        RECT 41.965 157.225 42.640 157.395 ;
        RECT 41.435 157.085 41.605 157.225 ;
        RECT 40.930 156.095 41.210 157.045 ;
        RECT 41.380 156.955 41.605 157.085 ;
        RECT 41.380 155.850 41.550 156.955 ;
        RECT 41.775 156.805 42.300 157.025 ;
        RECT 41.720 156.040 41.960 156.635 ;
        RECT 42.130 156.105 42.300 156.805 ;
        RECT 42.470 156.445 42.640 157.225 ;
        RECT 42.960 157.175 43.330 157.675 ;
        RECT 43.510 157.225 43.915 157.395 ;
        RECT 44.085 157.225 44.870 157.395 ;
        RECT 43.510 156.995 43.680 157.225 ;
        RECT 42.850 156.695 43.680 156.995 ;
        RECT 44.065 156.725 44.530 157.055 ;
        RECT 42.850 156.665 43.050 156.695 ;
        RECT 43.170 156.445 43.340 156.515 ;
        RECT 42.470 156.275 43.340 156.445 ;
        RECT 42.830 156.185 43.340 156.275 ;
        RECT 41.380 155.720 41.685 155.850 ;
        RECT 42.130 155.740 42.660 156.105 ;
        RECT 41.000 155.125 41.265 155.585 ;
        RECT 41.435 155.295 41.685 155.720 ;
        RECT 42.830 155.570 43.000 156.185 ;
        RECT 41.895 155.400 43.000 155.570 ;
        RECT 43.170 155.125 43.340 155.925 ;
        RECT 43.510 155.625 43.680 156.695 ;
        RECT 43.850 155.795 44.040 156.515 ;
        RECT 44.210 155.765 44.530 156.725 ;
        RECT 44.700 156.765 44.870 157.225 ;
        RECT 45.145 157.145 45.355 157.675 ;
        RECT 45.615 156.935 45.945 157.460 ;
        RECT 46.115 157.065 46.285 157.675 ;
        RECT 46.455 157.020 46.785 157.455 ;
        RECT 46.455 156.935 46.835 157.020 ;
        RECT 45.745 156.765 45.945 156.935 ;
        RECT 46.610 156.895 46.835 156.935 ;
        RECT 44.700 156.435 45.575 156.765 ;
        RECT 45.745 156.435 46.495 156.765 ;
        RECT 43.510 155.295 43.760 155.625 ;
        RECT 44.700 155.595 44.870 156.435 ;
        RECT 45.745 156.230 45.935 156.435 ;
        RECT 46.665 156.315 46.835 156.895 ;
        RECT 47.005 156.925 48.215 157.675 ;
        RECT 47.005 156.385 47.525 156.925 ;
        RECT 46.620 156.265 46.835 156.315 ;
        RECT 45.040 155.855 45.935 156.230 ;
        RECT 46.445 156.185 46.835 156.265 ;
        RECT 47.695 156.215 48.215 156.755 ;
        RECT 43.985 155.425 44.870 155.595 ;
        RECT 45.050 155.125 45.365 155.625 ;
        RECT 45.595 155.295 45.935 155.855 ;
        RECT 46.105 155.125 46.275 156.135 ;
        RECT 46.445 155.340 46.775 156.185 ;
        RECT 47.005 155.125 48.215 156.215 ;
        RECT 48.385 156.730 48.725 157.505 ;
        RECT 48.895 157.215 49.065 157.675 ;
        RECT 49.305 157.240 49.665 157.505 ;
        RECT 49.305 157.235 49.660 157.240 ;
        RECT 49.305 157.225 49.655 157.235 ;
        RECT 49.305 157.220 49.650 157.225 ;
        RECT 49.305 157.210 49.645 157.220 ;
        RECT 50.295 157.215 50.465 157.675 ;
        RECT 49.305 157.205 49.640 157.210 ;
        RECT 49.305 157.195 49.630 157.205 ;
        RECT 49.305 157.185 49.620 157.195 ;
        RECT 49.305 157.045 49.605 157.185 ;
        RECT 48.895 156.855 49.605 157.045 ;
        RECT 49.795 157.045 50.125 157.125 ;
        RECT 50.635 157.045 50.975 157.505 ;
        RECT 51.145 157.130 56.490 157.675 ;
        RECT 49.795 156.855 50.975 157.045 ;
        RECT 48.385 155.295 48.665 156.730 ;
        RECT 48.895 156.285 49.180 156.855 ;
        RECT 49.365 156.455 49.835 156.685 ;
        RECT 50.005 156.665 50.335 156.685 ;
        RECT 50.005 156.485 50.455 156.665 ;
        RECT 50.645 156.485 50.975 156.685 ;
        RECT 48.895 156.070 50.045 156.285 ;
        RECT 48.835 155.125 49.545 155.900 ;
        RECT 49.715 155.295 50.045 156.070 ;
        RECT 50.240 155.370 50.455 156.485 ;
        RECT 50.745 156.145 50.975 156.485 ;
        RECT 52.730 156.300 53.070 157.130 ;
        RECT 57.125 156.950 57.415 157.675 ;
        RECT 57.585 157.130 62.930 157.675 ;
        RECT 50.635 155.125 50.965 155.845 ;
        RECT 54.550 155.560 54.900 156.810 ;
        RECT 59.170 156.300 59.510 157.130 ;
        RECT 63.105 156.905 64.775 157.675 ;
        RECT 65.495 157.125 65.665 157.415 ;
        RECT 65.835 157.295 66.165 157.675 ;
        RECT 65.495 156.955 66.160 157.125 ;
        RECT 51.145 155.125 56.490 155.560 ;
        RECT 57.125 155.125 57.415 156.290 ;
        RECT 60.990 155.560 61.340 156.810 ;
        RECT 63.105 156.385 63.855 156.905 ;
        RECT 64.025 156.215 64.775 156.735 ;
        RECT 57.585 155.125 62.930 155.560 ;
        RECT 63.105 155.125 64.775 156.215 ;
        RECT 65.410 156.135 65.760 156.785 ;
        RECT 65.930 155.965 66.160 156.955 ;
        RECT 65.495 155.795 66.160 155.965 ;
        RECT 65.495 155.295 65.665 155.795 ;
        RECT 65.835 155.125 66.165 155.625 ;
        RECT 66.335 155.295 66.520 157.415 ;
        RECT 66.775 157.215 67.025 157.675 ;
        RECT 67.195 157.225 67.530 157.395 ;
        RECT 67.725 157.225 68.400 157.395 ;
        RECT 67.195 157.085 67.365 157.225 ;
        RECT 66.690 156.095 66.970 157.045 ;
        RECT 67.140 156.955 67.365 157.085 ;
        RECT 67.140 155.850 67.310 156.955 ;
        RECT 67.535 156.805 68.060 157.025 ;
        RECT 67.480 156.040 67.720 156.635 ;
        RECT 67.890 156.105 68.060 156.805 ;
        RECT 68.230 156.445 68.400 157.225 ;
        RECT 68.720 157.175 69.090 157.675 ;
        RECT 69.270 157.225 69.675 157.395 ;
        RECT 69.845 157.225 70.630 157.395 ;
        RECT 69.270 156.995 69.440 157.225 ;
        RECT 68.610 156.695 69.440 156.995 ;
        RECT 69.825 156.725 70.290 157.055 ;
        RECT 68.610 156.665 68.810 156.695 ;
        RECT 68.930 156.445 69.100 156.515 ;
        RECT 68.230 156.275 69.100 156.445 ;
        RECT 68.590 156.185 69.100 156.275 ;
        RECT 67.140 155.720 67.445 155.850 ;
        RECT 67.890 155.740 68.420 156.105 ;
        RECT 66.760 155.125 67.025 155.585 ;
        RECT 67.195 155.295 67.445 155.720 ;
        RECT 68.590 155.570 68.760 156.185 ;
        RECT 67.655 155.400 68.760 155.570 ;
        RECT 68.930 155.125 69.100 155.925 ;
        RECT 69.270 155.625 69.440 156.695 ;
        RECT 69.610 155.795 69.800 156.515 ;
        RECT 69.970 155.765 70.290 156.725 ;
        RECT 70.460 156.765 70.630 157.225 ;
        RECT 70.905 157.145 71.115 157.675 ;
        RECT 71.375 156.935 71.705 157.460 ;
        RECT 71.875 157.065 72.045 157.675 ;
        RECT 72.215 157.020 72.545 157.455 ;
        RECT 72.765 157.130 78.110 157.675 ;
        RECT 72.215 156.935 72.595 157.020 ;
        RECT 71.505 156.765 71.705 156.935 ;
        RECT 72.370 156.895 72.595 156.935 ;
        RECT 70.460 156.435 71.335 156.765 ;
        RECT 71.505 156.435 72.255 156.765 ;
        RECT 69.270 155.295 69.520 155.625 ;
        RECT 70.460 155.595 70.630 156.435 ;
        RECT 71.505 156.230 71.695 156.435 ;
        RECT 72.425 156.315 72.595 156.895 ;
        RECT 72.380 156.265 72.595 156.315 ;
        RECT 74.350 156.300 74.690 157.130 ;
        RECT 78.285 156.905 81.795 157.675 ;
        RECT 82.885 156.925 84.095 157.675 ;
        RECT 70.800 155.855 71.695 156.230 ;
        RECT 72.205 156.185 72.595 156.265 ;
        RECT 69.745 155.425 70.630 155.595 ;
        RECT 70.810 155.125 71.125 155.625 ;
        RECT 71.355 155.295 71.695 155.855 ;
        RECT 71.865 155.125 72.035 156.135 ;
        RECT 72.205 155.340 72.535 156.185 ;
        RECT 76.170 155.560 76.520 156.810 ;
        RECT 78.285 156.385 79.935 156.905 ;
        RECT 80.105 156.215 81.795 156.735 ;
        RECT 72.765 155.125 78.110 155.560 ;
        RECT 78.285 155.125 81.795 156.215 ;
        RECT 82.885 156.215 83.405 156.755 ;
        RECT 83.575 156.385 84.095 156.925 ;
        RECT 82.885 155.125 84.095 156.215 ;
        RECT 5.520 154.955 84.180 155.125 ;
        RECT 5.605 153.865 6.815 154.955 ;
        RECT 6.985 154.520 12.330 154.955 ;
        RECT 12.505 154.520 17.850 154.955 ;
        RECT 5.605 153.155 6.125 153.695 ;
        RECT 6.295 153.325 6.815 153.865 ;
        RECT 5.605 152.405 6.815 153.155 ;
        RECT 8.570 152.950 8.910 153.780 ;
        RECT 10.390 153.270 10.740 154.520 ;
        RECT 14.090 152.950 14.430 153.780 ;
        RECT 15.910 153.270 16.260 154.520 ;
        RECT 18.485 153.790 18.775 154.955 ;
        RECT 18.945 153.815 19.205 154.955 ;
        RECT 19.375 153.805 19.705 154.785 ;
        RECT 19.875 153.815 20.155 154.955 ;
        RECT 20.325 153.865 23.835 154.955 ;
        RECT 24.005 153.865 25.215 154.955 ;
        RECT 18.965 153.395 19.300 153.645 ;
        RECT 19.470 153.205 19.640 153.805 ;
        RECT 19.810 153.375 20.145 153.645 ;
        RECT 6.985 152.405 12.330 152.950 ;
        RECT 12.505 152.405 17.850 152.950 ;
        RECT 18.485 152.405 18.775 153.130 ;
        RECT 18.945 152.575 19.640 153.205 ;
        RECT 19.845 152.405 20.155 153.205 ;
        RECT 20.325 153.175 21.975 153.695 ;
        RECT 22.145 153.345 23.835 153.865 ;
        RECT 20.325 152.405 23.835 153.175 ;
        RECT 24.005 153.155 24.525 153.695 ;
        RECT 24.695 153.325 25.215 153.865 ;
        RECT 25.385 154.235 25.845 154.785 ;
        RECT 26.035 154.235 26.365 154.955 ;
        RECT 24.005 152.405 25.215 153.155 ;
        RECT 25.385 152.865 25.635 154.235 ;
        RECT 26.565 154.065 26.865 154.615 ;
        RECT 27.035 154.285 27.315 154.955 ;
        RECT 25.925 153.895 26.865 154.065 ;
        RECT 25.925 153.645 26.095 153.895 ;
        RECT 27.235 153.645 27.500 154.005 ;
        RECT 27.685 153.865 31.195 154.955 ;
        RECT 31.365 153.865 32.575 154.955 ;
        RECT 25.805 153.315 26.095 153.645 ;
        RECT 26.265 153.395 26.605 153.645 ;
        RECT 26.825 153.395 27.500 153.645 ;
        RECT 25.925 153.225 26.095 153.315 ;
        RECT 25.925 153.035 27.315 153.225 ;
        RECT 25.385 152.575 25.945 152.865 ;
        RECT 26.115 152.405 26.365 152.865 ;
        RECT 26.985 152.675 27.315 153.035 ;
        RECT 27.685 153.175 29.335 153.695 ;
        RECT 29.505 153.345 31.195 153.865 ;
        RECT 27.685 152.405 31.195 153.175 ;
        RECT 31.365 153.155 31.885 153.695 ;
        RECT 32.055 153.325 32.575 153.865 ;
        RECT 32.745 153.815 33.005 154.785 ;
        RECT 33.200 154.545 33.530 154.955 ;
        RECT 33.730 154.365 33.900 154.785 ;
        RECT 34.115 154.545 34.785 154.955 ;
        RECT 35.020 154.365 35.190 154.785 ;
        RECT 35.495 154.515 35.825 154.955 ;
        RECT 33.175 154.195 35.190 154.365 ;
        RECT 35.995 154.335 36.170 154.785 ;
        RECT 31.365 152.405 32.575 153.155 ;
        RECT 32.745 153.125 32.915 153.815 ;
        RECT 33.175 153.645 33.345 154.195 ;
        RECT 33.085 153.315 33.345 153.645 ;
        RECT 32.745 152.660 33.085 153.125 ;
        RECT 33.515 152.985 33.855 154.015 ;
        RECT 34.045 152.915 34.315 154.015 ;
        RECT 32.750 152.615 33.085 152.660 ;
        RECT 33.255 152.405 33.585 152.785 ;
        RECT 34.045 152.745 34.355 152.915 ;
        RECT 34.045 152.740 34.315 152.745 ;
        RECT 34.540 152.740 34.820 154.015 ;
        RECT 35.020 152.905 35.190 154.195 ;
        RECT 35.540 154.165 36.170 154.335 ;
        RECT 35.540 153.645 35.710 154.165 ;
        RECT 35.360 153.315 35.710 153.645 ;
        RECT 35.890 153.315 36.255 153.995 ;
        RECT 36.425 153.865 37.635 154.955 ;
        RECT 37.890 154.335 38.065 154.785 ;
        RECT 38.235 154.515 38.565 154.955 ;
        RECT 38.870 154.365 39.040 154.785 ;
        RECT 39.275 154.545 39.945 154.955 ;
        RECT 40.160 154.365 40.330 154.785 ;
        RECT 40.530 154.545 40.860 154.955 ;
        RECT 37.890 154.165 38.520 154.335 ;
        RECT 35.540 153.145 35.710 153.315 ;
        RECT 36.425 153.155 36.945 153.695 ;
        RECT 37.115 153.325 37.635 153.865 ;
        RECT 37.805 153.315 38.170 153.995 ;
        RECT 38.350 153.645 38.520 154.165 ;
        RECT 38.870 154.195 40.885 154.365 ;
        RECT 38.350 153.315 38.700 153.645 ;
        RECT 35.540 152.975 36.170 153.145 ;
        RECT 35.020 152.575 35.250 152.905 ;
        RECT 35.495 152.405 35.825 152.785 ;
        RECT 35.995 152.575 36.170 152.975 ;
        RECT 36.425 152.405 37.635 153.155 ;
        RECT 38.350 153.145 38.520 153.315 ;
        RECT 37.890 152.975 38.520 153.145 ;
        RECT 37.890 152.575 38.065 152.975 ;
        RECT 38.870 152.905 39.040 154.195 ;
        RECT 38.235 152.405 38.565 152.785 ;
        RECT 38.810 152.575 39.040 152.905 ;
        RECT 39.240 152.740 39.520 154.015 ;
        RECT 39.745 152.915 40.015 154.015 ;
        RECT 40.205 152.985 40.545 154.015 ;
        RECT 40.715 153.645 40.885 154.195 ;
        RECT 41.055 153.815 41.315 154.785 ;
        RECT 41.485 153.865 44.075 154.955 ;
        RECT 40.715 153.315 40.975 153.645 ;
        RECT 41.145 153.125 41.315 153.815 ;
        RECT 39.705 152.745 40.015 152.915 ;
        RECT 39.745 152.740 40.015 152.745 ;
        RECT 40.475 152.405 40.805 152.785 ;
        RECT 40.975 152.660 41.315 153.125 ;
        RECT 41.485 153.175 42.695 153.695 ;
        RECT 42.865 153.345 44.075 153.865 ;
        RECT 44.245 153.790 44.535 154.955 ;
        RECT 44.705 153.865 46.375 154.955 ;
        RECT 44.705 153.175 45.455 153.695 ;
        RECT 45.625 153.345 46.375 153.865 ;
        RECT 46.545 154.115 46.805 154.785 ;
        RECT 46.975 154.555 47.305 154.955 ;
        RECT 48.175 154.555 48.575 154.955 ;
        RECT 48.865 154.375 49.195 154.610 ;
        RECT 47.115 154.205 49.195 154.375 ;
        RECT 40.975 152.615 41.310 152.660 ;
        RECT 41.485 152.405 44.075 153.175 ;
        RECT 44.245 152.405 44.535 153.130 ;
        RECT 44.705 152.405 46.375 153.175 ;
        RECT 46.545 153.145 46.720 154.115 ;
        RECT 47.115 153.935 47.285 154.205 ;
        RECT 46.890 153.765 47.285 153.935 ;
        RECT 47.455 153.815 48.470 154.035 ;
        RECT 46.890 153.315 47.060 153.765 ;
        RECT 48.195 153.675 48.470 153.815 ;
        RECT 48.640 153.815 49.195 154.205 ;
        RECT 47.230 153.395 47.680 153.595 ;
        RECT 47.850 153.225 48.025 153.420 ;
        RECT 46.545 152.575 46.885 153.145 ;
        RECT 47.080 152.405 47.250 153.070 ;
        RECT 47.530 153.055 48.025 153.225 ;
        RECT 47.530 152.915 47.750 153.055 ;
        RECT 47.525 152.745 47.750 152.915 ;
        RECT 48.195 152.885 48.365 153.675 ;
        RECT 48.640 153.565 48.810 153.815 ;
        RECT 49.365 153.645 49.540 154.745 ;
        RECT 49.710 154.135 50.055 154.955 ;
        RECT 48.615 153.395 48.810 153.565 ;
        RECT 48.980 153.395 49.540 153.645 ;
        RECT 49.710 153.395 50.055 153.965 ;
        RECT 50.225 153.815 50.500 154.785 ;
        RECT 50.710 154.155 50.990 154.955 ;
        RECT 51.160 154.615 53.210 154.735 ;
        RECT 51.160 154.445 53.215 154.615 ;
        RECT 51.160 154.105 52.790 154.275 ;
        RECT 51.160 153.985 51.330 154.105 ;
        RECT 50.670 153.815 51.330 153.985 ;
        RECT 48.615 153.010 48.785 153.395 ;
        RECT 47.530 152.700 47.750 152.745 ;
        RECT 47.920 152.715 48.365 152.885 ;
        RECT 48.535 152.640 48.785 153.010 ;
        RECT 48.955 153.045 50.055 153.225 ;
        RECT 48.955 152.640 49.205 153.045 ;
        RECT 49.375 152.405 49.545 152.875 ;
        RECT 49.715 152.640 50.055 153.045 ;
        RECT 50.225 153.080 50.395 153.815 ;
        RECT 50.670 153.645 50.840 153.815 ;
        RECT 50.565 153.315 50.840 153.645 ;
        RECT 51.010 153.315 51.390 153.645 ;
        RECT 51.560 153.315 52.300 153.935 ;
        RECT 52.470 153.815 52.790 154.105 ;
        RECT 52.985 153.645 53.225 154.240 ;
        RECT 53.395 153.880 53.735 154.955 ;
        RECT 53.910 154.005 54.175 154.775 ;
        RECT 54.345 154.235 54.675 154.955 ;
        RECT 54.865 154.415 55.125 154.775 ;
        RECT 55.295 154.585 55.625 154.955 ;
        RECT 55.795 154.415 56.055 154.775 ;
        RECT 54.865 154.185 56.055 154.415 ;
        RECT 56.625 154.005 56.915 154.775 ;
        RECT 57.145 154.445 57.445 154.955 ;
        RECT 57.615 154.445 57.995 154.615 ;
        RECT 58.575 154.445 59.205 154.955 ;
        RECT 57.615 154.275 57.785 154.445 ;
        RECT 59.375 154.275 59.705 154.785 ;
        RECT 59.875 154.445 60.175 154.955 ;
        RECT 60.365 154.445 60.665 154.955 ;
        RECT 60.835 154.445 61.215 154.615 ;
        RECT 61.795 154.445 62.425 154.955 ;
        RECT 60.835 154.275 61.005 154.445 ;
        RECT 62.595 154.275 62.925 154.785 ;
        RECT 63.095 154.445 63.395 154.955 ;
        RECT 52.570 153.315 53.225 153.645 ;
        RECT 50.670 153.145 50.840 153.315 ;
        RECT 50.225 152.735 50.500 153.080 ;
        RECT 50.670 152.975 52.255 153.145 ;
        RECT 50.690 152.405 51.070 152.805 ;
        RECT 51.240 152.625 51.410 152.975 ;
        RECT 51.580 152.405 51.910 152.805 ;
        RECT 52.085 152.625 52.255 152.975 ;
        RECT 52.455 152.405 52.785 152.905 ;
        RECT 52.980 152.625 53.225 153.315 ;
        RECT 53.395 153.075 53.735 153.645 ;
        RECT 53.395 152.405 53.735 152.905 ;
        RECT 53.910 152.585 54.245 154.005 ;
        RECT 54.420 153.825 56.915 154.005 ;
        RECT 57.125 154.075 57.785 154.275 ;
        RECT 57.955 154.105 60.175 154.275 ;
        RECT 54.420 153.135 54.645 153.825 ;
        RECT 54.845 153.315 55.125 153.645 ;
        RECT 55.305 153.315 55.880 153.645 ;
        RECT 56.060 153.315 56.495 153.645 ;
        RECT 56.675 153.315 56.945 153.645 ;
        RECT 57.125 153.145 57.295 154.075 ;
        RECT 57.955 153.905 58.125 154.105 ;
        RECT 57.465 153.735 58.125 153.905 ;
        RECT 58.295 153.765 59.835 153.935 ;
        RECT 57.465 153.315 57.635 153.735 ;
        RECT 58.295 153.565 58.465 153.765 ;
        RECT 57.865 153.395 58.465 153.565 ;
        RECT 58.635 153.395 59.330 153.595 ;
        RECT 59.590 153.315 59.835 153.765 ;
        RECT 57.955 153.145 58.865 153.225 ;
        RECT 54.420 152.945 56.905 153.135 ;
        RECT 54.425 152.405 55.170 152.775 ;
        RECT 55.735 152.585 55.990 152.945 ;
        RECT 56.170 152.405 56.500 152.775 ;
        RECT 56.680 152.585 56.905 152.945 ;
        RECT 57.125 152.665 57.445 153.145 ;
        RECT 57.615 153.055 58.865 153.145 ;
        RECT 57.615 152.975 58.125 153.055 ;
        RECT 57.615 152.575 57.845 152.975 ;
        RECT 58.015 152.405 58.365 152.795 ;
        RECT 58.535 152.575 58.865 153.055 ;
        RECT 59.035 152.405 59.205 153.225 ;
        RECT 60.005 153.145 60.175 154.105 ;
        RECT 59.710 152.600 60.175 153.145 ;
        RECT 60.345 154.075 61.005 154.275 ;
        RECT 61.175 154.105 63.395 154.275 ;
        RECT 60.345 153.145 60.515 154.075 ;
        RECT 61.175 153.905 61.345 154.105 ;
        RECT 60.685 153.735 61.345 153.905 ;
        RECT 61.515 153.765 63.055 153.935 ;
        RECT 60.685 153.315 60.855 153.735 ;
        RECT 61.515 153.565 61.685 153.765 ;
        RECT 61.085 153.395 61.685 153.565 ;
        RECT 61.855 153.395 62.550 153.595 ;
        RECT 62.810 153.315 63.055 153.765 ;
        RECT 61.175 153.145 62.085 153.225 ;
        RECT 60.345 152.665 60.665 153.145 ;
        RECT 60.835 153.055 62.085 153.145 ;
        RECT 60.835 152.975 61.345 153.055 ;
        RECT 60.835 152.575 61.065 152.975 ;
        RECT 61.235 152.405 61.585 152.795 ;
        RECT 61.755 152.575 62.085 153.055 ;
        RECT 62.255 152.405 62.425 153.225 ;
        RECT 63.225 153.145 63.395 154.105 ;
        RECT 64.035 153.815 64.365 154.955 ;
        RECT 64.895 153.985 65.225 154.770 ;
        RECT 65.490 154.335 65.665 154.785 ;
        RECT 65.835 154.515 66.165 154.955 ;
        RECT 66.470 154.365 66.640 154.785 ;
        RECT 66.875 154.545 67.545 154.955 ;
        RECT 67.760 154.365 67.930 154.785 ;
        RECT 68.130 154.545 68.460 154.955 ;
        RECT 65.490 154.165 66.120 154.335 ;
        RECT 64.545 153.815 65.225 153.985 ;
        RECT 64.025 153.395 64.375 153.645 ;
        RECT 64.545 153.215 64.715 153.815 ;
        RECT 64.885 153.395 65.235 153.645 ;
        RECT 65.405 153.315 65.770 153.995 ;
        RECT 65.950 153.645 66.120 154.165 ;
        RECT 66.470 154.195 68.485 154.365 ;
        RECT 65.950 153.315 66.300 153.645 ;
        RECT 62.930 152.600 63.395 153.145 ;
        RECT 64.035 152.405 64.305 153.215 ;
        RECT 64.475 152.575 64.805 153.215 ;
        RECT 64.975 152.405 65.215 153.215 ;
        RECT 65.950 153.145 66.120 153.315 ;
        RECT 65.490 152.975 66.120 153.145 ;
        RECT 65.490 152.575 65.665 152.975 ;
        RECT 66.470 152.905 66.640 154.195 ;
        RECT 65.835 152.405 66.165 152.785 ;
        RECT 66.410 152.575 66.640 152.905 ;
        RECT 66.840 152.740 67.120 154.015 ;
        RECT 67.345 153.595 67.615 154.015 ;
        RECT 67.305 153.425 67.615 153.595 ;
        RECT 67.345 152.740 67.615 153.425 ;
        RECT 67.805 152.985 68.145 154.015 ;
        RECT 68.315 153.645 68.485 154.195 ;
        RECT 68.655 153.815 68.915 154.785 ;
        RECT 68.315 153.315 68.575 153.645 ;
        RECT 68.745 153.125 68.915 153.815 ;
        RECT 70.005 153.790 70.295 154.955 ;
        RECT 70.555 154.285 70.725 154.785 ;
        RECT 70.895 154.455 71.225 154.955 ;
        RECT 70.555 154.115 71.220 154.285 ;
        RECT 70.470 153.295 70.820 153.945 ;
        RECT 68.075 152.405 68.405 152.785 ;
        RECT 68.575 152.660 68.915 153.125 ;
        RECT 68.575 152.615 68.910 152.660 ;
        RECT 70.005 152.405 70.295 153.130 ;
        RECT 70.990 153.125 71.220 154.115 ;
        RECT 70.555 152.955 71.220 153.125 ;
        RECT 70.555 152.665 70.725 152.955 ;
        RECT 70.895 152.405 71.225 152.785 ;
        RECT 71.395 152.665 71.580 154.785 ;
        RECT 71.820 154.495 72.085 154.955 ;
        RECT 72.255 154.360 72.505 154.785 ;
        RECT 72.715 154.510 73.820 154.680 ;
        RECT 72.200 154.230 72.505 154.360 ;
        RECT 71.750 153.035 72.030 153.985 ;
        RECT 72.200 153.125 72.370 154.230 ;
        RECT 72.540 153.445 72.780 154.040 ;
        RECT 72.950 153.975 73.480 154.340 ;
        RECT 72.950 153.275 73.120 153.975 ;
        RECT 73.650 153.895 73.820 154.510 ;
        RECT 73.990 154.155 74.160 154.955 ;
        RECT 74.330 154.455 74.580 154.785 ;
        RECT 74.805 154.485 75.690 154.655 ;
        RECT 73.650 153.805 74.160 153.895 ;
        RECT 72.200 152.995 72.425 153.125 ;
        RECT 72.595 153.055 73.120 153.275 ;
        RECT 73.290 153.635 74.160 153.805 ;
        RECT 71.835 152.405 72.085 152.865 ;
        RECT 72.255 152.855 72.425 152.995 ;
        RECT 73.290 152.855 73.460 153.635 ;
        RECT 73.990 153.565 74.160 153.635 ;
        RECT 73.670 153.385 73.870 153.415 ;
        RECT 74.330 153.385 74.500 154.455 ;
        RECT 74.670 153.565 74.860 154.285 ;
        RECT 73.670 153.085 74.500 153.385 ;
        RECT 75.030 153.355 75.350 154.315 ;
        RECT 72.255 152.685 72.590 152.855 ;
        RECT 72.785 152.685 73.460 152.855 ;
        RECT 73.780 152.405 74.150 152.905 ;
        RECT 74.330 152.855 74.500 153.085 ;
        RECT 74.885 153.025 75.350 153.355 ;
        RECT 75.520 153.645 75.690 154.485 ;
        RECT 75.870 154.455 76.185 154.955 ;
        RECT 76.415 154.225 76.755 154.785 ;
        RECT 75.860 153.850 76.755 154.225 ;
        RECT 76.925 153.945 77.095 154.955 ;
        RECT 76.565 153.645 76.755 153.850 ;
        RECT 77.265 153.895 77.595 154.740 ;
        RECT 77.265 153.815 77.655 153.895 ;
        RECT 77.825 153.865 81.335 154.955 ;
        RECT 81.505 153.865 82.715 154.955 ;
        RECT 77.440 153.765 77.655 153.815 ;
        RECT 75.520 153.315 76.395 153.645 ;
        RECT 76.565 153.315 77.315 153.645 ;
        RECT 75.520 152.855 75.690 153.315 ;
        RECT 76.565 153.145 76.765 153.315 ;
        RECT 77.485 153.185 77.655 153.765 ;
        RECT 77.430 153.145 77.655 153.185 ;
        RECT 74.330 152.685 74.735 152.855 ;
        RECT 74.905 152.685 75.690 152.855 ;
        RECT 75.965 152.405 76.175 152.935 ;
        RECT 76.435 152.620 76.765 153.145 ;
        RECT 77.275 153.060 77.655 153.145 ;
        RECT 77.825 153.175 79.475 153.695 ;
        RECT 79.645 153.345 81.335 153.865 ;
        RECT 76.935 152.405 77.105 153.015 ;
        RECT 77.275 152.625 77.605 153.060 ;
        RECT 77.825 152.405 81.335 153.175 ;
        RECT 81.505 153.155 82.025 153.695 ;
        RECT 82.195 153.325 82.715 153.865 ;
        RECT 82.885 153.865 84.095 154.955 ;
        RECT 82.885 153.325 83.405 153.865 ;
        RECT 83.575 153.155 84.095 153.695 ;
        RECT 81.505 152.405 82.715 153.155 ;
        RECT 82.885 152.405 84.095 153.155 ;
        RECT 5.520 152.235 84.180 152.405 ;
        RECT 5.605 151.485 6.815 152.235 ;
        RECT 6.985 151.690 12.330 152.235 ;
        RECT 5.605 150.945 6.125 151.485 ;
        RECT 6.295 150.775 6.815 151.315 ;
        RECT 8.570 150.860 8.910 151.690 ;
        RECT 12.505 151.465 14.175 152.235 ;
        RECT 14.805 151.855 15.695 152.025 ;
        RECT 5.605 149.685 6.815 150.775 ;
        RECT 10.390 150.120 10.740 151.370 ;
        RECT 12.505 150.945 13.255 151.465 ;
        RECT 14.805 151.300 15.355 151.685 ;
        RECT 13.425 150.775 14.175 151.295 ;
        RECT 15.525 151.130 15.695 151.855 ;
        RECT 6.985 149.685 12.330 150.120 ;
        RECT 12.505 149.685 14.175 150.775 ;
        RECT 14.805 151.060 15.695 151.130 ;
        RECT 15.865 151.555 16.085 152.015 ;
        RECT 16.255 151.695 16.505 152.235 ;
        RECT 16.675 151.585 16.935 152.065 ;
        RECT 15.865 151.530 16.115 151.555 ;
        RECT 15.865 151.105 16.195 151.530 ;
        RECT 14.805 151.035 15.700 151.060 ;
        RECT 14.805 151.020 15.710 151.035 ;
        RECT 14.805 151.005 15.715 151.020 ;
        RECT 14.805 151.000 15.725 151.005 ;
        RECT 14.805 150.990 15.730 151.000 ;
        RECT 14.805 150.980 15.735 150.990 ;
        RECT 14.805 150.975 15.745 150.980 ;
        RECT 14.805 150.965 15.755 150.975 ;
        RECT 14.805 150.960 15.765 150.965 ;
        RECT 14.805 150.510 15.065 150.960 ;
        RECT 15.430 150.955 15.765 150.960 ;
        RECT 15.430 150.950 15.780 150.955 ;
        RECT 15.430 150.940 15.795 150.950 ;
        RECT 15.430 150.935 15.820 150.940 ;
        RECT 16.365 150.935 16.595 151.330 ;
        RECT 15.430 150.930 16.595 150.935 ;
        RECT 15.460 150.895 16.595 150.930 ;
        RECT 15.495 150.870 16.595 150.895 ;
        RECT 15.525 150.840 16.595 150.870 ;
        RECT 15.545 150.810 16.595 150.840 ;
        RECT 15.565 150.780 16.595 150.810 ;
        RECT 15.635 150.770 16.595 150.780 ;
        RECT 15.660 150.760 16.595 150.770 ;
        RECT 15.680 150.745 16.595 150.760 ;
        RECT 15.700 150.730 16.595 150.745 ;
        RECT 15.705 150.720 16.490 150.730 ;
        RECT 15.720 150.685 16.490 150.720 ;
        RECT 15.235 150.365 15.565 150.610 ;
        RECT 15.735 150.435 16.490 150.685 ;
        RECT 16.765 150.555 16.935 151.585 ;
        RECT 15.235 150.340 15.420 150.365 ;
        RECT 14.805 150.240 15.420 150.340 ;
        RECT 14.805 149.685 15.410 150.240 ;
        RECT 15.585 149.855 16.065 150.195 ;
        RECT 16.235 149.685 16.490 150.230 ;
        RECT 16.660 149.855 16.935 150.555 ;
        RECT 17.140 151.495 17.755 152.065 ;
        RECT 17.925 151.725 18.140 152.235 ;
        RECT 18.370 151.725 18.650 152.055 ;
        RECT 18.830 151.725 19.070 152.235 ;
        RECT 17.140 150.475 17.455 151.495 ;
        RECT 17.625 150.825 17.795 151.325 ;
        RECT 18.045 150.995 18.310 151.555 ;
        RECT 18.480 150.825 18.650 151.725 ;
        RECT 19.495 151.685 19.665 151.975 ;
        RECT 19.835 151.855 20.165 152.235 ;
        RECT 18.820 150.995 19.175 151.555 ;
        RECT 19.495 151.515 20.160 151.685 ;
        RECT 17.625 150.655 19.050 150.825 ;
        RECT 19.410 150.695 19.760 151.345 ;
        RECT 17.140 149.855 17.675 150.475 ;
        RECT 17.845 149.685 18.175 150.485 ;
        RECT 18.660 150.480 19.050 150.655 ;
        RECT 19.930 150.525 20.160 151.515 ;
        RECT 19.495 150.355 20.160 150.525 ;
        RECT 19.495 149.855 19.665 150.355 ;
        RECT 19.835 149.685 20.165 150.185 ;
        RECT 20.335 149.855 20.520 151.975 ;
        RECT 20.775 151.775 21.025 152.235 ;
        RECT 21.195 151.785 21.530 151.955 ;
        RECT 21.725 151.785 22.400 151.955 ;
        RECT 21.195 151.645 21.365 151.785 ;
        RECT 20.690 150.655 20.970 151.605 ;
        RECT 21.140 151.515 21.365 151.645 ;
        RECT 21.140 150.410 21.310 151.515 ;
        RECT 21.535 151.365 22.060 151.585 ;
        RECT 21.480 150.600 21.720 151.195 ;
        RECT 21.890 150.665 22.060 151.365 ;
        RECT 22.230 151.005 22.400 151.785 ;
        RECT 22.720 151.735 23.090 152.235 ;
        RECT 23.270 151.785 23.675 151.955 ;
        RECT 23.845 151.785 24.630 151.955 ;
        RECT 23.270 151.555 23.440 151.785 ;
        RECT 22.610 151.255 23.440 151.555 ;
        RECT 23.825 151.285 24.290 151.615 ;
        RECT 22.610 151.225 22.810 151.255 ;
        RECT 22.930 151.005 23.100 151.075 ;
        RECT 22.230 150.835 23.100 151.005 ;
        RECT 22.590 150.745 23.100 150.835 ;
        RECT 21.140 150.280 21.445 150.410 ;
        RECT 21.890 150.300 22.420 150.665 ;
        RECT 20.760 149.685 21.025 150.145 ;
        RECT 21.195 149.855 21.445 150.280 ;
        RECT 22.590 150.130 22.760 150.745 ;
        RECT 21.655 149.960 22.760 150.130 ;
        RECT 22.930 149.685 23.100 150.485 ;
        RECT 23.270 150.185 23.440 151.255 ;
        RECT 23.610 150.355 23.800 151.075 ;
        RECT 23.970 150.325 24.290 151.285 ;
        RECT 24.460 151.325 24.630 151.785 ;
        RECT 24.905 151.705 25.115 152.235 ;
        RECT 25.375 151.495 25.705 152.020 ;
        RECT 25.875 151.625 26.045 152.235 ;
        RECT 26.215 151.580 26.545 152.015 ;
        RECT 26.215 151.495 26.595 151.580 ;
        RECT 25.505 151.325 25.705 151.495 ;
        RECT 26.370 151.455 26.595 151.495 ;
        RECT 24.460 150.995 25.335 151.325 ;
        RECT 25.505 150.995 26.255 151.325 ;
        RECT 23.270 149.855 23.520 150.185 ;
        RECT 24.460 150.155 24.630 150.995 ;
        RECT 25.505 150.790 25.695 150.995 ;
        RECT 26.425 150.875 26.595 151.455 ;
        RECT 26.765 151.465 30.275 152.235 ;
        RECT 31.365 151.510 31.655 152.235 ;
        RECT 31.825 151.690 37.170 152.235 ;
        RECT 26.765 150.945 28.415 151.465 ;
        RECT 26.380 150.825 26.595 150.875 ;
        RECT 24.800 150.415 25.695 150.790 ;
        RECT 26.205 150.745 26.595 150.825 ;
        RECT 28.585 150.775 30.275 151.295 ;
        RECT 33.410 150.860 33.750 151.690 ;
        RECT 37.345 151.465 40.855 152.235 ;
        RECT 41.025 151.485 42.235 152.235 ;
        RECT 23.745 149.985 24.630 150.155 ;
        RECT 24.810 149.685 25.125 150.185 ;
        RECT 25.355 149.855 25.695 150.415 ;
        RECT 25.865 149.685 26.035 150.695 ;
        RECT 26.205 149.900 26.535 150.745 ;
        RECT 26.765 149.685 30.275 150.775 ;
        RECT 31.365 149.685 31.655 150.850 ;
        RECT 35.230 150.120 35.580 151.370 ;
        RECT 37.345 150.945 38.995 151.465 ;
        RECT 39.165 150.775 40.855 151.295 ;
        RECT 41.025 150.945 41.545 151.485 ;
        RECT 42.425 151.425 42.665 152.235 ;
        RECT 42.835 151.425 43.165 152.065 ;
        RECT 43.335 151.425 43.605 152.235 ;
        RECT 43.785 151.495 44.225 152.055 ;
        RECT 44.395 151.495 44.845 152.235 ;
        RECT 45.015 151.665 45.185 152.065 ;
        RECT 45.355 151.835 45.775 152.235 ;
        RECT 45.945 151.665 46.175 152.065 ;
        RECT 45.015 151.495 46.175 151.665 ;
        RECT 46.345 151.495 46.835 152.065 ;
        RECT 47.015 151.735 47.345 152.235 ;
        RECT 47.545 151.665 47.715 152.015 ;
        RECT 47.915 151.835 48.245 152.235 ;
        RECT 48.415 151.665 48.585 152.015 ;
        RECT 48.755 151.835 49.135 152.235 ;
        RECT 41.715 150.775 42.235 151.315 ;
        RECT 42.405 150.995 42.755 151.245 ;
        RECT 42.925 150.825 43.095 151.425 ;
        RECT 43.265 150.995 43.615 151.245 ;
        RECT 31.825 149.685 37.170 150.120 ;
        RECT 37.345 149.685 40.855 150.775 ;
        RECT 41.025 149.685 42.235 150.775 ;
        RECT 42.415 150.655 43.095 150.825 ;
        RECT 42.415 149.870 42.745 150.655 ;
        RECT 43.275 149.685 43.605 150.825 ;
        RECT 43.785 150.485 44.095 151.495 ;
        RECT 44.265 150.875 44.435 151.325 ;
        RECT 44.605 151.045 44.995 151.325 ;
        RECT 45.180 150.995 45.425 151.325 ;
        RECT 44.265 150.705 45.055 150.875 ;
        RECT 43.785 149.855 44.225 150.485 ;
        RECT 44.400 149.685 44.715 150.535 ;
        RECT 44.885 150.025 45.055 150.705 ;
        RECT 45.225 150.195 45.425 150.995 ;
        RECT 45.625 150.195 45.875 151.325 ;
        RECT 46.090 150.995 46.495 151.325 ;
        RECT 46.665 150.825 46.835 151.495 ;
        RECT 47.010 150.995 47.360 151.565 ;
        RECT 47.545 151.495 49.155 151.665 ;
        RECT 49.325 151.560 49.595 151.905 ;
        RECT 48.985 151.325 49.155 151.495 ;
        RECT 47.530 150.875 48.240 151.325 ;
        RECT 48.410 150.995 48.815 151.325 ;
        RECT 48.985 150.995 49.255 151.325 ;
        RECT 46.065 150.655 46.835 150.825 ;
        RECT 46.065 150.025 46.315 150.655 ;
        RECT 47.010 150.535 47.330 150.825 ;
        RECT 47.525 150.705 48.240 150.875 ;
        RECT 48.985 150.825 49.155 150.995 ;
        RECT 49.425 150.825 49.595 151.560 ;
        RECT 49.765 151.465 53.275 152.235 ;
        RECT 54.370 151.560 54.645 151.905 ;
        RECT 54.835 151.835 55.215 152.235 ;
        RECT 55.385 151.665 55.555 152.015 ;
        RECT 55.725 151.835 56.055 152.235 ;
        RECT 56.225 151.665 56.480 152.015 ;
        RECT 49.765 150.945 51.415 151.465 ;
        RECT 48.430 150.655 49.155 150.825 ;
        RECT 48.430 150.535 48.600 150.655 ;
        RECT 44.885 149.855 46.315 150.025 ;
        RECT 46.495 149.685 46.825 150.485 ;
        RECT 47.010 150.365 48.600 150.535 ;
        RECT 47.010 149.905 48.665 150.195 ;
        RECT 48.835 149.685 49.115 150.485 ;
        RECT 49.325 149.855 49.595 150.825 ;
        RECT 51.585 150.775 53.275 151.295 ;
        RECT 49.765 149.685 53.275 150.775 ;
        RECT 54.370 150.825 54.540 151.560 ;
        RECT 54.815 151.495 56.480 151.665 ;
        RECT 57.125 151.510 57.415 152.235 ;
        RECT 58.510 151.560 58.785 151.905 ;
        RECT 58.975 151.835 59.355 152.235 ;
        RECT 59.525 151.665 59.695 152.015 ;
        RECT 59.865 151.835 60.195 152.235 ;
        RECT 60.365 151.665 60.620 152.015 ;
        RECT 54.815 151.325 54.985 151.495 ;
        RECT 54.710 150.995 54.985 151.325 ;
        RECT 55.155 150.995 55.980 151.325 ;
        RECT 56.150 150.995 56.495 151.325 ;
        RECT 54.815 150.825 54.985 150.995 ;
        RECT 54.370 149.855 54.645 150.825 ;
        RECT 54.815 150.655 55.475 150.825 ;
        RECT 55.785 150.705 55.980 150.995 ;
        RECT 55.305 150.535 55.475 150.655 ;
        RECT 56.150 150.535 56.475 150.825 ;
        RECT 54.855 149.685 55.135 150.485 ;
        RECT 55.305 150.365 56.475 150.535 ;
        RECT 55.305 149.905 56.495 150.195 ;
        RECT 57.125 149.685 57.415 150.850 ;
        RECT 58.510 150.825 58.680 151.560 ;
        RECT 58.955 151.495 60.620 151.665 ;
        RECT 61.725 151.515 62.065 152.025 ;
        RECT 58.955 151.325 59.125 151.495 ;
        RECT 58.850 150.995 59.125 151.325 ;
        RECT 59.295 150.995 60.120 151.325 ;
        RECT 60.290 150.995 60.635 151.325 ;
        RECT 58.955 150.825 59.125 150.995 ;
        RECT 58.510 149.855 58.785 150.825 ;
        RECT 58.955 150.655 59.615 150.825 ;
        RECT 59.925 150.705 60.120 150.995 ;
        RECT 59.445 150.535 59.615 150.655 ;
        RECT 60.290 150.535 60.615 150.825 ;
        RECT 58.995 149.685 59.275 150.485 ;
        RECT 59.445 150.365 60.615 150.535 ;
        RECT 59.445 149.905 60.635 150.195 ;
        RECT 61.725 150.115 61.985 151.515 ;
        RECT 62.235 151.435 62.505 152.235 ;
        RECT 62.160 150.995 62.490 151.245 ;
        RECT 62.685 150.995 62.965 151.965 ;
        RECT 63.145 150.995 63.445 151.965 ;
        RECT 63.625 150.995 63.975 151.960 ;
        RECT 64.195 151.735 64.690 152.065 ;
        RECT 62.175 150.825 62.490 150.995 ;
        RECT 64.195 150.825 64.365 151.735 ;
        RECT 62.175 150.655 64.365 150.825 ;
        RECT 61.725 149.855 62.065 150.115 ;
        RECT 62.235 149.685 62.565 150.485 ;
        RECT 63.030 149.855 63.280 150.655 ;
        RECT 63.465 149.685 63.795 150.405 ;
        RECT 64.015 149.855 64.265 150.655 ;
        RECT 64.535 150.245 64.775 151.555 ;
        RECT 64.945 151.465 66.615 152.235 ;
        RECT 66.785 151.585 67.045 152.065 ;
        RECT 67.215 151.695 67.465 152.235 ;
        RECT 64.945 150.945 65.695 151.465 ;
        RECT 65.865 150.775 66.615 151.295 ;
        RECT 64.435 149.685 64.770 150.065 ;
        RECT 64.945 149.685 66.615 150.775 ;
        RECT 66.785 150.555 66.955 151.585 ;
        RECT 67.635 151.555 67.855 152.015 ;
        RECT 67.605 151.530 67.855 151.555 ;
        RECT 67.125 150.935 67.355 151.330 ;
        RECT 67.525 151.105 67.855 151.530 ;
        RECT 68.025 151.855 68.915 152.025 ;
        RECT 68.025 151.130 68.195 151.855 ;
        RECT 68.365 151.300 68.915 151.685 ;
        RECT 69.095 151.505 69.395 152.235 ;
        RECT 69.575 151.325 69.805 151.945 ;
        RECT 70.005 151.675 70.230 152.055 ;
        RECT 70.400 151.845 70.730 152.235 ;
        RECT 70.925 151.690 76.270 152.235 ;
        RECT 76.445 151.690 81.790 152.235 ;
        RECT 70.005 151.495 70.335 151.675 ;
        RECT 68.025 151.060 68.915 151.130 ;
        RECT 68.020 151.035 68.915 151.060 ;
        RECT 68.010 151.020 68.915 151.035 ;
        RECT 68.005 151.005 68.915 151.020 ;
        RECT 67.995 151.000 68.915 151.005 ;
        RECT 67.990 150.990 68.915 151.000 ;
        RECT 69.100 150.995 69.395 151.325 ;
        RECT 69.575 150.995 69.990 151.325 ;
        RECT 67.985 150.980 68.915 150.990 ;
        RECT 67.975 150.975 68.915 150.980 ;
        RECT 67.965 150.965 68.915 150.975 ;
        RECT 67.955 150.960 68.915 150.965 ;
        RECT 67.955 150.955 68.290 150.960 ;
        RECT 67.940 150.950 68.290 150.955 ;
        RECT 67.925 150.940 68.290 150.950 ;
        RECT 67.900 150.935 68.290 150.940 ;
        RECT 67.125 150.930 68.290 150.935 ;
        RECT 67.125 150.895 68.260 150.930 ;
        RECT 67.125 150.870 68.225 150.895 ;
        RECT 67.125 150.840 68.195 150.870 ;
        RECT 67.125 150.810 68.175 150.840 ;
        RECT 67.125 150.780 68.155 150.810 ;
        RECT 67.125 150.770 68.085 150.780 ;
        RECT 67.125 150.760 68.060 150.770 ;
        RECT 67.125 150.745 68.040 150.760 ;
        RECT 67.125 150.730 68.020 150.745 ;
        RECT 67.230 150.720 68.015 150.730 ;
        RECT 67.230 150.685 68.000 150.720 ;
        RECT 66.785 149.855 67.060 150.555 ;
        RECT 67.230 150.435 67.985 150.685 ;
        RECT 68.155 150.365 68.485 150.610 ;
        RECT 68.655 150.510 68.915 150.960 ;
        RECT 70.160 150.825 70.335 151.495 ;
        RECT 70.505 150.995 70.745 151.645 ;
        RECT 72.510 150.860 72.850 151.690 ;
        RECT 68.300 150.340 68.485 150.365 ;
        RECT 69.095 150.465 69.990 150.795 ;
        RECT 70.160 150.635 70.745 150.825 ;
        RECT 68.300 150.240 68.915 150.340 ;
        RECT 67.230 149.685 67.485 150.230 ;
        RECT 67.655 149.855 68.135 150.195 ;
        RECT 68.310 149.685 68.915 150.240 ;
        RECT 69.095 150.295 70.300 150.465 ;
        RECT 69.095 149.865 69.425 150.295 ;
        RECT 69.605 149.685 69.800 150.125 ;
        RECT 69.970 149.865 70.300 150.295 ;
        RECT 70.470 149.865 70.745 150.635 ;
        RECT 74.330 150.120 74.680 151.370 ;
        RECT 78.030 150.860 78.370 151.690 ;
        RECT 82.885 151.485 84.095 152.235 ;
        RECT 79.850 150.120 80.200 151.370 ;
        RECT 82.885 150.775 83.405 151.315 ;
        RECT 83.575 150.945 84.095 151.485 ;
        RECT 70.925 149.685 76.270 150.120 ;
        RECT 76.445 149.685 81.790 150.120 ;
        RECT 82.885 149.685 84.095 150.775 ;
        RECT 5.520 149.515 84.180 149.685 ;
        RECT 5.605 148.425 6.815 149.515 ;
        RECT 6.985 148.425 10.495 149.515 ;
        RECT 11.215 148.845 11.385 149.345 ;
        RECT 11.555 149.015 11.885 149.515 ;
        RECT 11.215 148.675 11.880 148.845 ;
        RECT 5.605 147.715 6.125 148.255 ;
        RECT 6.295 147.885 6.815 148.425 ;
        RECT 6.985 147.735 8.635 148.255 ;
        RECT 8.805 147.905 10.495 148.425 ;
        RECT 11.130 147.855 11.480 148.505 ;
        RECT 5.605 146.965 6.815 147.715 ;
        RECT 6.985 146.965 10.495 147.735 ;
        RECT 11.650 147.685 11.880 148.675 ;
        RECT 11.215 147.515 11.880 147.685 ;
        RECT 11.215 147.225 11.385 147.515 ;
        RECT 11.555 146.965 11.885 147.345 ;
        RECT 12.055 147.225 12.240 149.345 ;
        RECT 12.480 149.055 12.745 149.515 ;
        RECT 12.915 148.920 13.165 149.345 ;
        RECT 13.375 149.070 14.480 149.240 ;
        RECT 12.860 148.790 13.165 148.920 ;
        RECT 12.410 147.595 12.690 148.545 ;
        RECT 12.860 147.685 13.030 148.790 ;
        RECT 13.200 148.005 13.440 148.600 ;
        RECT 13.610 148.535 14.140 148.900 ;
        RECT 13.610 147.835 13.780 148.535 ;
        RECT 14.310 148.455 14.480 149.070 ;
        RECT 14.650 148.715 14.820 149.515 ;
        RECT 14.990 149.015 15.240 149.345 ;
        RECT 15.465 149.045 16.350 149.215 ;
        RECT 14.310 148.365 14.820 148.455 ;
        RECT 12.860 147.555 13.085 147.685 ;
        RECT 13.255 147.615 13.780 147.835 ;
        RECT 13.950 148.195 14.820 148.365 ;
        RECT 12.495 146.965 12.745 147.425 ;
        RECT 12.915 147.415 13.085 147.555 ;
        RECT 13.950 147.415 14.120 148.195 ;
        RECT 14.650 148.125 14.820 148.195 ;
        RECT 14.330 147.945 14.530 147.975 ;
        RECT 14.990 147.945 15.160 149.015 ;
        RECT 15.330 148.125 15.520 148.845 ;
        RECT 14.330 147.645 15.160 147.945 ;
        RECT 15.690 147.915 16.010 148.875 ;
        RECT 12.915 147.245 13.250 147.415 ;
        RECT 13.445 147.245 14.120 147.415 ;
        RECT 14.440 146.965 14.810 147.465 ;
        RECT 14.990 147.415 15.160 147.645 ;
        RECT 15.545 147.585 16.010 147.915 ;
        RECT 16.180 148.205 16.350 149.045 ;
        RECT 16.530 149.015 16.845 149.515 ;
        RECT 17.075 148.785 17.415 149.345 ;
        RECT 16.520 148.410 17.415 148.785 ;
        RECT 17.585 148.505 17.755 149.515 ;
        RECT 17.225 148.205 17.415 148.410 ;
        RECT 17.925 148.455 18.255 149.300 ;
        RECT 17.925 148.375 18.315 148.455 ;
        RECT 18.100 148.325 18.315 148.375 ;
        RECT 18.485 148.350 18.775 149.515 ;
        RECT 16.180 147.875 17.055 148.205 ;
        RECT 17.225 147.875 17.975 148.205 ;
        RECT 16.180 147.415 16.350 147.875 ;
        RECT 17.225 147.705 17.425 147.875 ;
        RECT 18.145 147.745 18.315 148.325 ;
        RECT 18.090 147.705 18.315 147.745 ;
        RECT 14.990 147.245 15.395 147.415 ;
        RECT 15.565 147.245 16.350 147.415 ;
        RECT 16.625 146.965 16.835 147.495 ;
        RECT 17.095 147.180 17.425 147.705 ;
        RECT 17.935 147.620 18.315 147.705 ;
        RECT 17.595 146.965 17.765 147.575 ;
        RECT 17.935 147.185 18.265 147.620 ;
        RECT 18.485 146.965 18.775 147.690 ;
        RECT 18.955 147.145 19.215 149.335 ;
        RECT 19.385 148.785 19.725 149.515 ;
        RECT 19.905 148.605 20.175 149.335 ;
        RECT 19.405 148.385 20.175 148.605 ;
        RECT 20.355 148.625 20.585 149.335 ;
        RECT 20.755 148.805 21.085 149.515 ;
        RECT 21.255 148.625 21.515 149.335 ;
        RECT 20.355 148.385 21.515 148.625 ;
        RECT 21.705 148.425 24.295 149.515 ;
        RECT 19.405 147.715 19.695 148.385 ;
        RECT 19.875 147.895 20.340 148.205 ;
        RECT 20.520 147.895 21.045 148.205 ;
        RECT 19.405 147.515 20.635 147.715 ;
        RECT 19.475 146.965 20.145 147.335 ;
        RECT 20.325 147.145 20.635 147.515 ;
        RECT 20.815 147.255 21.045 147.895 ;
        RECT 21.225 147.875 21.525 148.205 ;
        RECT 21.705 147.735 22.915 148.255 ;
        RECT 23.085 147.905 24.295 148.425 ;
        RECT 24.555 148.505 24.725 149.345 ;
        RECT 24.895 149.175 26.065 149.345 ;
        RECT 24.895 148.675 25.225 149.175 ;
        RECT 25.735 149.135 26.065 149.175 ;
        RECT 26.255 149.095 26.610 149.515 ;
        RECT 25.395 148.915 25.625 149.005 ;
        RECT 26.780 148.915 27.030 149.345 ;
        RECT 25.395 148.675 27.030 148.915 ;
        RECT 27.200 148.755 27.530 149.515 ;
        RECT 27.700 148.675 27.955 149.345 ;
        RECT 24.555 148.335 27.615 148.505 ;
        RECT 24.470 147.955 24.820 148.165 ;
        RECT 24.990 147.955 25.435 148.155 ;
        RECT 25.605 147.955 26.080 148.155 ;
        RECT 21.225 146.965 21.515 147.695 ;
        RECT 21.705 146.965 24.295 147.735 ;
        RECT 24.555 147.615 25.620 147.785 ;
        RECT 24.555 147.135 24.725 147.615 ;
        RECT 24.895 146.965 25.225 147.445 ;
        RECT 25.450 147.385 25.620 147.615 ;
        RECT 25.800 147.555 26.080 147.955 ;
        RECT 26.350 147.955 26.680 148.155 ;
        RECT 26.850 147.985 27.225 148.155 ;
        RECT 26.850 147.955 27.215 147.985 ;
        RECT 26.350 147.555 26.635 147.955 ;
        RECT 27.445 147.785 27.615 148.335 ;
        RECT 26.815 147.615 27.615 147.785 ;
        RECT 26.815 147.385 26.985 147.615 ;
        RECT 27.785 147.545 27.955 148.675 ;
        RECT 28.145 148.425 29.355 149.515 ;
        RECT 30.025 149.055 30.240 149.515 ;
        RECT 30.410 148.885 30.740 149.345 ;
        RECT 27.770 147.475 27.955 147.545 ;
        RECT 27.745 147.465 27.955 147.475 ;
        RECT 25.450 147.135 26.985 147.385 ;
        RECT 27.155 146.965 27.485 147.445 ;
        RECT 27.700 147.135 27.955 147.465 ;
        RECT 28.145 147.715 28.665 148.255 ;
        RECT 28.835 147.885 29.355 148.425 ;
        RECT 29.570 148.715 30.740 148.885 ;
        RECT 30.910 148.715 31.160 149.515 ;
        RECT 28.145 146.965 29.355 147.715 ;
        RECT 29.570 147.425 29.940 148.715 ;
        RECT 31.370 148.545 31.650 148.705 ;
        RECT 30.315 148.375 31.650 148.545 ;
        RECT 32.285 148.665 32.665 149.345 ;
        RECT 33.255 148.665 33.425 149.515 ;
        RECT 33.595 148.835 33.925 149.345 ;
        RECT 34.095 149.005 34.265 149.515 ;
        RECT 34.435 148.835 34.835 149.345 ;
        RECT 33.595 148.665 34.835 148.835 ;
        RECT 30.315 148.205 30.485 148.375 ;
        RECT 30.110 147.955 30.485 148.205 ;
        RECT 30.655 147.955 31.130 148.195 ;
        RECT 31.300 147.955 31.650 148.195 ;
        RECT 30.315 147.785 30.485 147.955 ;
        RECT 30.315 147.615 31.650 147.785 ;
        RECT 29.570 147.135 30.320 147.425 ;
        RECT 30.830 146.965 31.160 147.425 ;
        RECT 31.380 147.405 31.650 147.615 ;
        RECT 32.285 147.705 32.455 148.665 ;
        RECT 32.625 148.325 33.930 148.495 ;
        RECT 35.015 148.415 35.335 149.345 ;
        RECT 35.505 148.425 36.715 149.515 ;
        RECT 36.885 149.005 37.185 149.515 ;
        RECT 37.355 148.835 37.685 149.345 ;
        RECT 37.855 149.005 38.485 149.515 ;
        RECT 39.065 149.005 39.445 149.175 ;
        RECT 39.615 149.005 39.915 149.515 ;
        RECT 39.275 148.835 39.445 149.005 ;
        RECT 32.625 147.875 32.870 148.325 ;
        RECT 33.040 147.955 33.590 148.155 ;
        RECT 33.760 148.125 33.930 148.325 ;
        RECT 34.705 148.245 35.335 148.415 ;
        RECT 33.760 147.955 34.135 148.125 ;
        RECT 34.305 147.705 34.535 148.205 ;
        RECT 32.285 147.535 34.535 147.705 ;
        RECT 32.335 146.965 32.665 147.355 ;
        RECT 32.835 147.215 33.005 147.535 ;
        RECT 34.705 147.365 34.875 148.245 ;
        RECT 33.175 146.965 33.505 147.355 ;
        RECT 33.920 147.195 34.875 147.365 ;
        RECT 35.045 146.965 35.335 147.800 ;
        RECT 35.505 147.715 36.025 148.255 ;
        RECT 36.195 147.885 36.715 148.425 ;
        RECT 36.885 148.665 39.105 148.835 ;
        RECT 35.505 146.965 36.715 147.715 ;
        RECT 36.885 147.705 37.055 148.665 ;
        RECT 37.225 148.325 38.765 148.495 ;
        RECT 37.225 147.875 37.470 148.325 ;
        RECT 37.730 147.955 38.425 148.155 ;
        RECT 38.595 148.125 38.765 148.325 ;
        RECT 38.935 148.465 39.105 148.665 ;
        RECT 39.275 148.635 39.935 148.835 ;
        RECT 38.935 148.295 39.595 148.465 ;
        RECT 38.595 147.955 39.195 148.125 ;
        RECT 39.425 147.875 39.595 148.295 ;
        RECT 36.885 147.160 37.350 147.705 ;
        RECT 37.855 146.965 38.025 147.785 ;
        RECT 38.195 147.705 39.105 147.785 ;
        RECT 39.765 147.705 39.935 148.635 ;
        RECT 40.105 148.425 41.315 149.515 ;
        RECT 41.490 149.005 43.145 149.295 ;
        RECT 38.195 147.615 39.445 147.705 ;
        RECT 38.195 147.135 38.525 147.615 ;
        RECT 38.935 147.535 39.445 147.615 ;
        RECT 38.695 146.965 39.045 147.355 ;
        RECT 39.215 147.135 39.445 147.535 ;
        RECT 39.615 147.225 39.935 147.705 ;
        RECT 40.105 147.715 40.625 148.255 ;
        RECT 40.795 147.885 41.315 148.425 ;
        RECT 41.490 148.665 43.080 148.835 ;
        RECT 43.315 148.715 43.595 149.515 ;
        RECT 41.490 148.375 41.810 148.665 ;
        RECT 42.910 148.545 43.080 148.665 ;
        RECT 40.105 146.965 41.315 147.715 ;
        RECT 41.490 147.635 41.840 148.205 ;
        RECT 42.010 147.875 42.720 148.495 ;
        RECT 42.910 148.375 43.635 148.545 ;
        RECT 43.805 148.375 44.075 149.345 ;
        RECT 43.465 148.205 43.635 148.375 ;
        RECT 42.890 147.875 43.295 148.205 ;
        RECT 43.465 147.875 43.735 148.205 ;
        RECT 43.465 147.705 43.635 147.875 ;
        RECT 42.025 147.535 43.635 147.705 ;
        RECT 43.905 147.640 44.075 148.375 ;
        RECT 44.245 148.350 44.535 149.515 ;
        RECT 44.710 148.545 45.005 149.515 ;
        RECT 45.575 149.155 45.905 149.515 ;
        RECT 46.075 149.155 48.055 149.345 ;
        RECT 45.175 148.985 45.395 149.070 ;
        RECT 46.075 148.985 46.255 149.155 ;
        RECT 48.235 149.075 48.505 149.515 ;
        RECT 49.055 149.155 49.385 149.515 ;
        RECT 49.900 149.155 50.230 149.515 ;
        RECT 50.740 149.155 51.075 149.515 ;
        RECT 51.975 149.155 52.305 149.515 ;
        RECT 45.175 148.815 46.255 148.985 ;
        RECT 46.425 148.905 48.090 148.985 ;
        RECT 48.665 148.905 52.300 148.985 ;
        RECT 45.175 148.740 45.395 148.815 ;
        RECT 46.425 148.735 52.300 148.905 ;
        RECT 45.585 148.395 48.250 148.565 ;
        RECT 45.585 148.210 46.030 148.395 ;
        RECT 45.020 147.955 46.030 148.210 ;
        RECT 46.325 147.955 47.800 148.225 ;
        RECT 47.970 147.875 48.250 148.395 ;
        RECT 48.880 148.395 51.620 148.565 ;
        RECT 48.880 148.290 49.595 148.395 ;
        RECT 48.420 147.875 49.595 148.290 ;
        RECT 49.990 147.955 51.060 148.225 ;
        RECT 51.450 147.875 51.620 148.395 ;
        RECT 51.790 148.220 52.300 148.735 ;
        RECT 52.615 148.505 52.785 149.345 ;
        RECT 52.955 149.175 54.125 149.345 ;
        RECT 52.955 148.675 53.285 149.175 ;
        RECT 53.795 149.135 54.125 149.175 ;
        RECT 54.315 149.095 54.670 149.515 ;
        RECT 53.455 148.915 53.685 149.005 ;
        RECT 54.840 148.915 55.090 149.345 ;
        RECT 53.455 148.675 55.090 148.915 ;
        RECT 55.260 148.755 55.590 149.515 ;
        RECT 55.760 148.675 56.015 149.345 ;
        RECT 52.615 148.335 55.675 148.505 ;
        RECT 44.775 147.745 46.415 147.785 ;
        RECT 41.495 146.965 41.825 147.465 ;
        RECT 42.025 147.185 42.195 147.535 ;
        RECT 42.395 146.965 42.725 147.365 ;
        RECT 42.895 147.185 43.065 147.535 ;
        RECT 43.235 146.965 43.615 147.365 ;
        RECT 43.805 147.295 44.075 147.640 ;
        RECT 44.245 146.965 44.535 147.690 ;
        RECT 44.775 147.675 47.750 147.745 ;
        RECT 51.790 147.705 51.970 148.220 ;
        RECT 52.530 147.955 52.880 148.165 ;
        RECT 53.050 147.955 53.495 148.155 ;
        RECT 53.665 147.955 54.140 148.155 ;
        RECT 44.775 147.575 48.455 147.675 ;
        RECT 44.775 147.505 45.860 147.575 ;
        RECT 46.395 147.505 48.455 147.575 ;
        RECT 48.625 147.515 50.790 147.695 ;
        RECT 51.185 147.535 51.970 147.705 ;
        RECT 52.615 147.615 53.680 147.785 ;
        RECT 44.775 147.415 44.975 147.505 ;
        RECT 45.145 146.965 45.475 147.325 ;
        RECT 45.645 147.305 45.860 147.505 ;
        RECT 46.085 146.965 46.255 147.405 ;
        RECT 48.225 147.335 48.455 147.505 ;
        RECT 46.865 146.965 47.195 147.325 ;
        RECT 47.725 146.965 48.055 147.325 ;
        RECT 48.225 147.135 49.540 147.335 ;
        RECT 51.185 147.330 51.355 147.535 ;
        RECT 52.130 147.360 52.300 147.475 ;
        RECT 49.900 147.150 51.355 147.330 ;
        RECT 51.600 147.190 52.300 147.360 ;
        RECT 52.615 147.135 52.785 147.615 ;
        RECT 52.955 146.965 53.285 147.445 ;
        RECT 53.510 147.385 53.680 147.615 ;
        RECT 53.860 147.555 54.140 147.955 ;
        RECT 54.410 147.955 54.740 148.155 ;
        RECT 54.910 147.955 55.275 148.155 ;
        RECT 54.410 147.555 54.695 147.955 ;
        RECT 55.505 147.785 55.675 148.335 ;
        RECT 54.875 147.615 55.675 147.785 ;
        RECT 54.875 147.385 55.045 147.615 ;
        RECT 55.845 147.545 56.015 148.675 ;
        RECT 56.205 148.375 56.465 149.515 ;
        RECT 56.635 148.365 56.965 149.345 ;
        RECT 57.135 148.375 57.415 149.515 ;
        RECT 57.585 149.080 62.930 149.515 ;
        RECT 56.225 147.955 56.560 148.205 ;
        RECT 56.730 147.765 56.900 148.365 ;
        RECT 57.070 147.935 57.405 148.205 ;
        RECT 55.830 147.475 56.015 147.545 ;
        RECT 55.805 147.465 56.015 147.475 ;
        RECT 53.510 147.135 55.045 147.385 ;
        RECT 55.215 146.965 55.545 147.445 ;
        RECT 55.760 147.135 56.015 147.465 ;
        RECT 56.205 147.135 56.900 147.765 ;
        RECT 57.105 146.965 57.415 147.765 ;
        RECT 59.170 147.510 59.510 148.340 ;
        RECT 60.990 147.830 61.340 149.080 ;
        RECT 63.105 148.425 65.695 149.515 ;
        RECT 63.105 147.735 64.315 148.255 ;
        RECT 64.485 147.905 65.695 148.425 ;
        RECT 65.875 148.375 66.205 149.515 ;
        RECT 66.735 148.545 67.065 149.330 ;
        RECT 66.385 148.375 67.065 148.545 ;
        RECT 67.255 148.545 67.585 149.330 ;
        RECT 67.255 148.375 67.935 148.545 ;
        RECT 68.115 148.375 68.445 149.515 ;
        RECT 68.625 148.425 69.835 149.515 ;
        RECT 65.865 147.955 66.215 148.205 ;
        RECT 66.385 147.775 66.555 148.375 ;
        RECT 66.725 147.955 67.075 148.205 ;
        RECT 67.245 147.955 67.595 148.205 ;
        RECT 67.765 147.775 67.935 148.375 ;
        RECT 68.105 147.955 68.455 148.205 ;
        RECT 57.585 146.965 62.930 147.510 ;
        RECT 63.105 146.965 65.695 147.735 ;
        RECT 65.875 146.965 66.145 147.775 ;
        RECT 66.315 147.135 66.645 147.775 ;
        RECT 66.815 146.965 67.055 147.775 ;
        RECT 67.265 146.965 67.505 147.775 ;
        RECT 67.675 147.135 68.005 147.775 ;
        RECT 68.175 146.965 68.445 147.775 ;
        RECT 68.625 147.715 69.145 148.255 ;
        RECT 69.315 147.885 69.835 148.425 ;
        RECT 70.005 148.350 70.295 149.515 ;
        RECT 70.465 149.080 75.810 149.515 ;
        RECT 75.985 149.080 81.330 149.515 ;
        RECT 68.625 146.965 69.835 147.715 ;
        RECT 70.005 146.965 70.295 147.690 ;
        RECT 72.050 147.510 72.390 148.340 ;
        RECT 73.870 147.830 74.220 149.080 ;
        RECT 77.570 147.510 77.910 148.340 ;
        RECT 79.390 147.830 79.740 149.080 ;
        RECT 81.505 148.425 82.715 149.515 ;
        RECT 81.505 147.715 82.025 148.255 ;
        RECT 82.195 147.885 82.715 148.425 ;
        RECT 82.885 148.425 84.095 149.515 ;
        RECT 82.885 147.885 83.405 148.425 ;
        RECT 83.575 147.715 84.095 148.255 ;
        RECT 70.465 146.965 75.810 147.510 ;
        RECT 75.985 146.965 81.330 147.510 ;
        RECT 81.505 146.965 82.715 147.715 ;
        RECT 82.885 146.965 84.095 147.715 ;
        RECT 5.520 146.795 84.180 146.965 ;
        RECT 5.605 146.045 6.815 146.795 ;
        RECT 6.985 146.250 12.330 146.795 ;
        RECT 5.605 145.505 6.125 146.045 ;
        RECT 6.295 145.335 6.815 145.875 ;
        RECT 8.570 145.420 8.910 146.250 ;
        RECT 12.505 146.145 12.765 146.625 ;
        RECT 12.935 146.335 13.265 146.795 ;
        RECT 13.455 146.155 13.655 146.575 ;
        RECT 5.605 144.245 6.815 145.335 ;
        RECT 10.390 144.680 10.740 145.930 ;
        RECT 12.505 145.115 12.675 146.145 ;
        RECT 12.845 145.455 13.075 145.885 ;
        RECT 13.245 145.635 13.655 146.155 ;
        RECT 13.825 146.310 14.615 146.575 ;
        RECT 13.825 145.455 14.080 146.310 ;
        RECT 14.795 145.975 15.125 146.395 ;
        RECT 15.295 145.975 15.555 146.795 ;
        RECT 16.185 146.145 16.445 146.625 ;
        RECT 16.615 146.255 16.865 146.795 ;
        RECT 14.795 145.885 15.045 145.975 ;
        RECT 14.250 145.635 15.045 145.885 ;
        RECT 12.845 145.285 14.635 145.455 ;
        RECT 6.985 144.245 12.330 144.680 ;
        RECT 12.505 144.415 12.780 145.115 ;
        RECT 12.950 144.990 13.665 145.285 ;
        RECT 13.885 144.925 14.215 145.115 ;
        RECT 12.990 144.245 13.205 144.790 ;
        RECT 13.375 144.415 13.850 144.755 ;
        RECT 14.020 144.750 14.215 144.925 ;
        RECT 14.385 144.920 14.635 145.285 ;
        RECT 14.020 144.245 14.635 144.750 ;
        RECT 14.875 144.415 15.045 145.635 ;
        RECT 15.215 144.925 15.555 145.805 ;
        RECT 16.185 145.115 16.355 146.145 ;
        RECT 17.035 146.090 17.255 146.575 ;
        RECT 16.525 145.495 16.755 145.890 ;
        RECT 16.925 145.665 17.255 146.090 ;
        RECT 17.425 146.415 18.315 146.585 ;
        RECT 17.425 145.690 17.595 146.415 ;
        RECT 18.485 146.250 23.830 146.795 ;
        RECT 17.765 145.860 18.315 146.245 ;
        RECT 17.425 145.620 18.315 145.690 ;
        RECT 17.420 145.595 18.315 145.620 ;
        RECT 17.410 145.580 18.315 145.595 ;
        RECT 17.405 145.565 18.315 145.580 ;
        RECT 17.395 145.560 18.315 145.565 ;
        RECT 17.390 145.550 18.315 145.560 ;
        RECT 17.385 145.540 18.315 145.550 ;
        RECT 17.375 145.535 18.315 145.540 ;
        RECT 17.365 145.525 18.315 145.535 ;
        RECT 17.355 145.520 18.315 145.525 ;
        RECT 17.355 145.515 17.690 145.520 ;
        RECT 17.340 145.510 17.690 145.515 ;
        RECT 17.325 145.500 17.690 145.510 ;
        RECT 17.300 145.495 17.690 145.500 ;
        RECT 16.525 145.490 17.690 145.495 ;
        RECT 16.525 145.455 17.660 145.490 ;
        RECT 16.525 145.430 17.625 145.455 ;
        RECT 16.525 145.400 17.595 145.430 ;
        RECT 16.525 145.370 17.575 145.400 ;
        RECT 16.525 145.340 17.555 145.370 ;
        RECT 16.525 145.330 17.485 145.340 ;
        RECT 16.525 145.320 17.460 145.330 ;
        RECT 16.525 145.305 17.440 145.320 ;
        RECT 16.525 145.290 17.420 145.305 ;
        RECT 16.630 145.280 17.415 145.290 ;
        RECT 16.630 145.245 17.400 145.280 ;
        RECT 15.295 144.245 15.555 144.755 ;
        RECT 16.185 144.415 16.460 145.115 ;
        RECT 16.630 144.995 17.385 145.245 ;
        RECT 17.555 144.925 17.885 145.170 ;
        RECT 18.055 145.070 18.315 145.520 ;
        RECT 20.070 145.420 20.410 146.250 ;
        RECT 24.005 146.145 24.345 146.625 ;
        RECT 24.710 146.315 25.040 146.625 ;
        RECT 25.210 146.315 25.460 146.795 ;
        RECT 24.870 146.145 25.040 146.315 ;
        RECT 25.630 146.145 25.960 146.625 ;
        RECT 26.130 146.315 26.380 146.795 ;
        RECT 26.550 146.145 26.880 146.625 ;
        RECT 24.005 145.975 24.700 146.145 ;
        RECT 24.870 145.975 26.880 146.145 ;
        RECT 27.225 146.025 30.735 146.795 ;
        RECT 31.365 146.070 31.655 146.795 ;
        RECT 31.875 146.140 32.205 146.575 ;
        RECT 32.375 146.185 32.545 146.795 ;
        RECT 31.825 146.055 32.205 146.140 ;
        RECT 32.715 146.055 33.045 146.580 ;
        RECT 33.305 146.265 33.515 146.795 ;
        RECT 33.790 146.345 34.575 146.515 ;
        RECT 34.745 146.345 35.150 146.515 ;
        RECT 17.700 144.900 17.885 144.925 ;
        RECT 17.700 144.800 18.315 144.900 ;
        RECT 16.630 144.245 16.885 144.790 ;
        RECT 17.055 144.415 17.535 144.755 ;
        RECT 17.710 144.245 18.315 144.800 ;
        RECT 21.890 144.680 22.240 145.930 ;
        RECT 24.025 145.605 24.360 145.805 ;
        RECT 18.485 144.245 23.830 144.680 ;
        RECT 24.005 144.245 24.265 145.435 ;
        RECT 24.530 145.395 24.700 145.975 ;
        RECT 24.910 145.635 25.240 145.805 ;
        RECT 24.435 144.415 24.765 145.395 ;
        RECT 24.935 144.525 25.240 145.635 ;
        RECT 25.420 145.635 25.750 145.805 ;
        RECT 25.420 144.525 25.740 145.635 ;
        RECT 25.920 145.465 26.250 145.805 ;
        RECT 26.420 145.555 27.000 145.805 ;
        RECT 27.225 145.505 28.875 146.025 ;
        RECT 31.825 146.015 32.050 146.055 ;
        RECT 25.910 144.525 26.250 145.465 ;
        RECT 26.550 144.245 26.880 145.385 ;
        RECT 29.045 145.335 30.735 145.855 ;
        RECT 31.825 145.435 31.995 146.015 ;
        RECT 32.715 145.885 32.915 146.055 ;
        RECT 33.790 145.885 33.960 146.345 ;
        RECT 32.165 145.555 32.915 145.885 ;
        RECT 33.085 145.555 33.960 145.885 ;
        RECT 27.225 144.245 30.735 145.335 ;
        RECT 31.365 144.245 31.655 145.410 ;
        RECT 31.825 145.385 32.040 145.435 ;
        RECT 31.825 145.305 32.215 145.385 ;
        RECT 31.885 144.460 32.215 145.305 ;
        RECT 32.725 145.350 32.915 145.555 ;
        RECT 32.385 144.245 32.555 145.255 ;
        RECT 32.725 144.975 33.620 145.350 ;
        RECT 32.725 144.415 33.065 144.975 ;
        RECT 33.295 144.245 33.610 144.745 ;
        RECT 33.790 144.715 33.960 145.555 ;
        RECT 34.130 145.845 34.595 146.175 ;
        RECT 34.980 146.115 35.150 146.345 ;
        RECT 35.330 146.295 35.700 146.795 ;
        RECT 36.020 146.345 36.695 146.515 ;
        RECT 36.890 146.345 37.225 146.515 ;
        RECT 34.130 144.885 34.450 145.845 ;
        RECT 34.980 145.815 35.810 146.115 ;
        RECT 34.620 144.915 34.810 145.635 ;
        RECT 34.980 144.745 35.150 145.815 ;
        RECT 35.610 145.785 35.810 145.815 ;
        RECT 35.320 145.565 35.490 145.635 ;
        RECT 36.020 145.565 36.190 146.345 ;
        RECT 37.055 146.205 37.225 146.345 ;
        RECT 37.395 146.335 37.645 146.795 ;
        RECT 35.320 145.395 36.190 145.565 ;
        RECT 36.360 145.925 36.885 146.145 ;
        RECT 37.055 146.075 37.280 146.205 ;
        RECT 35.320 145.305 35.830 145.395 ;
        RECT 33.790 144.545 34.675 144.715 ;
        RECT 34.900 144.415 35.150 144.745 ;
        RECT 35.320 144.245 35.490 145.045 ;
        RECT 35.660 144.690 35.830 145.305 ;
        RECT 36.360 145.225 36.530 145.925 ;
        RECT 36.000 144.860 36.530 145.225 ;
        RECT 36.700 145.160 36.940 145.755 ;
        RECT 37.110 144.970 37.280 146.075 ;
        RECT 37.450 145.215 37.730 146.165 ;
        RECT 36.975 144.840 37.280 144.970 ;
        RECT 35.660 144.520 36.765 144.690 ;
        RECT 36.975 144.415 37.225 144.840 ;
        RECT 37.395 144.245 37.660 144.705 ;
        RECT 37.900 144.415 38.085 146.535 ;
        RECT 38.255 146.415 38.585 146.795 ;
        RECT 38.755 146.245 38.925 146.535 ;
        RECT 38.260 146.075 38.925 146.245 ;
        RECT 38.260 145.085 38.490 146.075 ;
        RECT 39.185 146.025 40.855 146.795 ;
        RECT 41.505 146.065 41.795 146.795 ;
        RECT 38.660 145.255 39.010 145.905 ;
        RECT 39.185 145.505 39.935 146.025 ;
        RECT 40.105 145.335 40.855 145.855 ;
        RECT 41.495 145.555 41.795 145.885 ;
        RECT 41.975 145.865 42.205 146.505 ;
        RECT 42.385 146.245 42.695 146.615 ;
        RECT 42.875 146.425 43.545 146.795 ;
        RECT 42.385 146.045 43.615 146.245 ;
        RECT 41.975 145.555 42.500 145.865 ;
        RECT 42.680 145.555 43.145 145.865 ;
        RECT 43.325 145.375 43.615 146.045 ;
        RECT 38.260 144.915 38.925 145.085 ;
        RECT 38.255 144.245 38.585 144.745 ;
        RECT 38.755 144.415 38.925 144.915 ;
        RECT 39.185 144.245 40.855 145.335 ;
        RECT 41.505 145.135 42.665 145.375 ;
        RECT 41.505 144.425 41.765 145.135 ;
        RECT 41.935 144.245 42.265 144.955 ;
        RECT 42.435 144.425 42.665 145.135 ;
        RECT 42.845 145.155 43.615 145.375 ;
        RECT 42.845 144.425 43.115 145.155 ;
        RECT 43.295 144.245 43.635 144.975 ;
        RECT 43.805 144.425 44.065 146.615 ;
        RECT 44.245 146.250 49.590 146.795 ;
        RECT 45.830 145.420 46.170 146.250 ;
        RECT 49.765 146.045 50.975 146.795 ;
        RECT 51.310 146.285 51.550 146.795 ;
        RECT 51.730 146.285 52.010 146.615 ;
        RECT 52.240 146.285 52.455 146.795 ;
        RECT 47.650 144.680 48.000 145.930 ;
        RECT 49.765 145.505 50.285 146.045 ;
        RECT 50.455 145.335 50.975 145.875 ;
        RECT 51.205 145.555 51.560 146.115 ;
        RECT 51.730 145.385 51.900 146.285 ;
        RECT 52.070 145.555 52.335 146.115 ;
        RECT 52.625 146.055 53.240 146.625 ;
        RECT 52.585 145.385 52.755 145.885 ;
        RECT 44.245 144.245 49.590 144.680 ;
        RECT 49.765 144.245 50.975 145.335 ;
        RECT 51.330 145.215 52.755 145.385 ;
        RECT 51.330 145.040 51.720 145.215 ;
        RECT 52.205 144.245 52.535 145.045 ;
        RECT 52.925 145.035 53.240 146.055 ;
        RECT 52.705 144.415 53.240 145.035 ;
        RECT 53.445 145.995 53.785 146.625 ;
        RECT 53.955 145.995 54.205 146.795 ;
        RECT 54.395 146.145 54.725 146.625 ;
        RECT 54.895 146.335 55.120 146.795 ;
        RECT 55.290 146.145 55.620 146.625 ;
        RECT 53.445 145.385 53.620 145.995 ;
        RECT 54.395 145.975 55.620 146.145 ;
        RECT 56.250 146.015 56.750 146.625 ;
        RECT 57.125 146.070 57.415 146.795 ;
        RECT 53.790 145.635 54.485 145.805 ;
        RECT 54.315 145.385 54.485 145.635 ;
        RECT 54.660 145.605 55.080 145.805 ;
        RECT 55.250 145.605 55.580 145.805 ;
        RECT 55.750 145.605 56.080 145.805 ;
        RECT 56.250 145.385 56.420 146.015 ;
        RECT 57.585 145.995 57.925 146.625 ;
        RECT 58.095 145.995 58.345 146.795 ;
        RECT 58.535 146.145 58.865 146.625 ;
        RECT 59.035 146.335 59.260 146.795 ;
        RECT 59.430 146.145 59.760 146.625 ;
        RECT 57.585 145.945 57.815 145.995 ;
        RECT 58.535 145.975 59.760 146.145 ;
        RECT 60.390 146.015 60.890 146.625 ;
        RECT 61.310 146.335 62.060 146.625 ;
        RECT 62.570 146.335 62.900 146.795 ;
        RECT 56.605 145.555 56.955 145.805 ;
        RECT 53.445 144.415 53.785 145.385 ;
        RECT 53.955 144.245 54.125 145.385 ;
        RECT 54.315 145.215 56.750 145.385 ;
        RECT 54.395 144.245 54.645 145.045 ;
        RECT 55.290 144.415 55.620 145.215 ;
        RECT 55.920 144.245 56.250 145.045 ;
        RECT 56.420 144.415 56.750 145.215 ;
        RECT 57.125 144.245 57.415 145.410 ;
        RECT 57.585 145.385 57.760 145.945 ;
        RECT 57.930 145.635 58.625 145.805 ;
        RECT 58.455 145.385 58.625 145.635 ;
        RECT 58.800 145.605 59.220 145.805 ;
        RECT 59.390 145.605 59.720 145.805 ;
        RECT 59.890 145.605 60.220 145.805 ;
        RECT 60.390 145.385 60.560 146.015 ;
        RECT 60.745 145.555 61.095 145.805 ;
        RECT 57.585 144.415 57.925 145.385 ;
        RECT 58.095 144.245 58.265 145.385 ;
        RECT 58.455 145.215 60.890 145.385 ;
        RECT 58.535 144.245 58.785 145.045 ;
        RECT 59.430 144.415 59.760 145.215 ;
        RECT 60.060 144.245 60.390 145.045 ;
        RECT 60.560 144.415 60.890 145.215 ;
        RECT 61.310 145.045 61.680 146.335 ;
        RECT 63.120 146.145 63.390 146.355 ;
        RECT 62.055 145.975 63.390 146.145 ;
        RECT 63.650 146.225 63.825 146.625 ;
        RECT 63.995 146.415 64.325 146.795 ;
        RECT 64.570 146.295 64.800 146.625 ;
        RECT 63.650 146.055 64.280 146.225 ;
        RECT 62.055 145.805 62.225 145.975 ;
        RECT 64.110 145.885 64.280 146.055 ;
        RECT 61.850 145.555 62.225 145.805 ;
        RECT 62.395 145.565 62.870 145.805 ;
        RECT 63.040 145.565 63.390 145.805 ;
        RECT 62.055 145.385 62.225 145.555 ;
        RECT 62.055 145.215 63.390 145.385 ;
        RECT 63.110 145.055 63.390 145.215 ;
        RECT 63.565 145.205 63.930 145.885 ;
        RECT 64.110 145.555 64.460 145.885 ;
        RECT 61.310 144.875 62.480 145.045 ;
        RECT 61.765 144.245 61.980 144.705 ;
        RECT 62.150 144.415 62.480 144.875 ;
        RECT 62.650 144.245 62.900 145.045 ;
        RECT 64.110 145.035 64.280 145.555 ;
        RECT 63.650 144.865 64.280 145.035 ;
        RECT 64.630 145.005 64.800 146.295 ;
        RECT 65.000 145.185 65.280 146.460 ;
        RECT 65.505 146.455 65.775 146.460 ;
        RECT 65.465 146.285 65.775 146.455 ;
        RECT 66.235 146.415 66.565 146.795 ;
        RECT 66.735 146.540 67.070 146.585 ;
        RECT 65.505 145.185 65.775 146.285 ;
        RECT 65.965 145.185 66.305 146.215 ;
        RECT 66.735 146.075 67.075 146.540 ;
        RECT 67.335 146.245 67.505 146.535 ;
        RECT 67.675 146.415 68.005 146.795 ;
        RECT 67.335 146.075 68.000 146.245 ;
        RECT 66.475 145.555 66.735 145.885 ;
        RECT 66.475 145.005 66.645 145.555 ;
        RECT 66.905 145.385 67.075 146.075 ;
        RECT 63.650 144.415 63.825 144.865 ;
        RECT 64.630 144.835 66.645 145.005 ;
        RECT 63.995 144.245 64.325 144.685 ;
        RECT 64.630 144.415 64.800 144.835 ;
        RECT 65.035 144.245 65.705 144.655 ;
        RECT 65.920 144.415 66.090 144.835 ;
        RECT 66.290 144.245 66.620 144.655 ;
        RECT 66.815 144.415 67.075 145.385 ;
        RECT 67.250 145.255 67.600 145.905 ;
        RECT 67.770 145.085 68.000 146.075 ;
        RECT 67.335 144.915 68.000 145.085 ;
        RECT 67.335 144.415 67.505 144.915 ;
        RECT 67.675 144.245 68.005 144.745 ;
        RECT 68.175 144.415 68.360 146.535 ;
        RECT 68.615 146.335 68.865 146.795 ;
        RECT 69.035 146.345 69.370 146.515 ;
        RECT 69.565 146.345 70.240 146.515 ;
        RECT 69.035 146.205 69.205 146.345 ;
        RECT 68.530 145.215 68.810 146.165 ;
        RECT 68.980 146.075 69.205 146.205 ;
        RECT 68.980 144.970 69.150 146.075 ;
        RECT 69.375 145.925 69.900 146.145 ;
        RECT 69.320 145.160 69.560 145.755 ;
        RECT 69.730 145.225 69.900 145.925 ;
        RECT 70.070 145.565 70.240 146.345 ;
        RECT 70.560 146.295 70.930 146.795 ;
        RECT 71.110 146.345 71.515 146.515 ;
        RECT 71.685 146.345 72.470 146.515 ;
        RECT 71.110 146.115 71.280 146.345 ;
        RECT 70.450 145.815 71.280 146.115 ;
        RECT 71.665 145.845 72.130 146.175 ;
        RECT 70.450 145.785 70.650 145.815 ;
        RECT 70.770 145.565 70.940 145.635 ;
        RECT 70.070 145.395 70.940 145.565 ;
        RECT 70.430 145.305 70.940 145.395 ;
        RECT 68.980 144.840 69.285 144.970 ;
        RECT 69.730 144.860 70.260 145.225 ;
        RECT 68.600 144.245 68.865 144.705 ;
        RECT 69.035 144.415 69.285 144.840 ;
        RECT 70.430 144.690 70.600 145.305 ;
        RECT 69.495 144.520 70.600 144.690 ;
        RECT 70.770 144.245 70.940 145.045 ;
        RECT 71.110 144.745 71.280 145.815 ;
        RECT 71.450 144.915 71.640 145.635 ;
        RECT 71.810 144.885 72.130 145.845 ;
        RECT 72.300 145.885 72.470 146.345 ;
        RECT 72.745 146.265 72.955 146.795 ;
        RECT 73.215 146.055 73.545 146.580 ;
        RECT 73.715 146.185 73.885 146.795 ;
        RECT 74.055 146.140 74.385 146.575 ;
        RECT 74.605 146.250 79.950 146.795 ;
        RECT 74.055 146.055 74.435 146.140 ;
        RECT 73.345 145.885 73.545 146.055 ;
        RECT 74.210 146.015 74.435 146.055 ;
        RECT 72.300 145.555 73.175 145.885 ;
        RECT 73.345 145.555 74.095 145.885 ;
        RECT 71.110 144.415 71.360 144.745 ;
        RECT 72.300 144.715 72.470 145.555 ;
        RECT 73.345 145.350 73.535 145.555 ;
        RECT 74.265 145.435 74.435 146.015 ;
        RECT 74.220 145.385 74.435 145.435 ;
        RECT 76.190 145.420 76.530 146.250 ;
        RECT 80.125 146.025 82.715 146.795 ;
        RECT 82.885 146.045 84.095 146.795 ;
        RECT 72.640 144.975 73.535 145.350 ;
        RECT 74.045 145.305 74.435 145.385 ;
        RECT 71.585 144.545 72.470 144.715 ;
        RECT 72.650 144.245 72.965 144.745 ;
        RECT 73.195 144.415 73.535 144.975 ;
        RECT 73.705 144.245 73.875 145.255 ;
        RECT 74.045 144.460 74.375 145.305 ;
        RECT 78.010 144.680 78.360 145.930 ;
        RECT 80.125 145.505 81.335 146.025 ;
        RECT 81.505 145.335 82.715 145.855 ;
        RECT 74.605 144.245 79.950 144.680 ;
        RECT 80.125 144.245 82.715 145.335 ;
        RECT 82.885 145.335 83.405 145.875 ;
        RECT 83.575 145.505 84.095 146.045 ;
        RECT 82.885 144.245 84.095 145.335 ;
        RECT 5.520 144.075 84.180 144.245 ;
        RECT 5.605 142.985 6.815 144.075 ;
        RECT 6.985 143.640 12.330 144.075 ;
        RECT 12.505 143.640 17.850 144.075 ;
        RECT 5.605 142.275 6.125 142.815 ;
        RECT 6.295 142.445 6.815 142.985 ;
        RECT 5.605 141.525 6.815 142.275 ;
        RECT 8.570 142.070 8.910 142.900 ;
        RECT 10.390 142.390 10.740 143.640 ;
        RECT 14.090 142.070 14.430 142.900 ;
        RECT 15.910 142.390 16.260 143.640 ;
        RECT 18.485 142.910 18.775 144.075 ;
        RECT 18.945 142.985 20.155 144.075 ;
        RECT 18.945 142.275 19.465 142.815 ;
        RECT 19.635 142.445 20.155 142.985 ;
        RECT 20.325 142.935 20.605 144.075 ;
        RECT 20.775 142.925 21.105 143.905 ;
        RECT 21.275 142.935 21.535 144.075 ;
        RECT 20.335 142.495 20.670 142.765 ;
        RECT 20.840 142.325 21.010 142.925 ;
        RECT 21.180 142.515 21.515 142.765 ;
        RECT 6.985 141.525 12.330 142.070 ;
        RECT 12.505 141.525 17.850 142.070 ;
        RECT 18.485 141.525 18.775 142.250 ;
        RECT 18.945 141.525 20.155 142.275 ;
        RECT 20.325 141.525 20.635 142.325 ;
        RECT 20.840 141.695 21.535 142.325 ;
        RECT 22.635 141.705 22.895 143.895 ;
        RECT 23.065 143.345 23.405 144.075 ;
        RECT 23.585 143.165 23.855 143.895 ;
        RECT 23.085 142.945 23.855 143.165 ;
        RECT 24.035 143.185 24.265 143.895 ;
        RECT 24.435 143.365 24.765 144.075 ;
        RECT 24.935 143.185 25.195 143.895 ;
        RECT 25.500 143.445 25.785 143.905 ;
        RECT 25.955 143.615 26.225 144.075 ;
        RECT 25.500 143.225 26.455 143.445 ;
        RECT 24.035 142.945 25.195 143.185 ;
        RECT 23.085 142.275 23.375 142.945 ;
        RECT 23.555 142.455 24.020 142.765 ;
        RECT 24.200 142.455 24.725 142.765 ;
        RECT 23.085 142.075 24.315 142.275 ;
        RECT 23.155 141.525 23.825 141.895 ;
        RECT 24.005 141.705 24.315 142.075 ;
        RECT 24.495 141.815 24.725 142.455 ;
        RECT 24.905 142.435 25.205 142.765 ;
        RECT 25.385 142.495 26.075 143.055 ;
        RECT 26.245 142.325 26.455 143.225 ;
        RECT 24.905 141.525 25.195 142.255 ;
        RECT 25.500 142.155 26.455 142.325 ;
        RECT 26.625 143.055 27.025 143.905 ;
        RECT 27.215 143.445 27.495 143.905 ;
        RECT 28.015 143.615 28.340 144.075 ;
        RECT 27.215 143.225 28.340 143.445 ;
        RECT 26.625 142.495 27.720 143.055 ;
        RECT 27.890 142.765 28.340 143.225 ;
        RECT 28.510 142.935 28.895 143.905 ;
        RECT 29.250 143.105 29.640 143.280 ;
        RECT 30.125 143.275 30.455 144.075 ;
        RECT 30.625 143.285 31.160 143.905 ;
        RECT 29.250 142.935 30.675 143.105 ;
        RECT 25.500 141.695 25.785 142.155 ;
        RECT 25.955 141.525 26.225 141.985 ;
        RECT 26.625 141.695 27.025 142.495 ;
        RECT 27.890 142.435 28.445 142.765 ;
        RECT 27.890 142.325 28.340 142.435 ;
        RECT 27.215 142.155 28.340 142.325 ;
        RECT 28.615 142.265 28.895 142.935 ;
        RECT 27.215 141.695 27.495 142.155 ;
        RECT 28.015 141.525 28.340 141.985 ;
        RECT 28.510 141.695 28.895 142.265 ;
        RECT 29.125 142.205 29.480 142.765 ;
        RECT 29.650 142.035 29.820 142.935 ;
        RECT 29.990 142.205 30.255 142.765 ;
        RECT 30.505 142.435 30.675 142.935 ;
        RECT 30.845 142.265 31.160 143.285 ;
        RECT 31.405 142.935 31.635 144.075 ;
        RECT 31.805 142.925 32.135 143.905 ;
        RECT 32.305 142.935 32.515 144.075 ;
        RECT 32.830 143.455 33.005 143.905 ;
        RECT 33.175 143.635 33.505 144.075 ;
        RECT 33.810 143.485 33.980 143.905 ;
        RECT 34.215 143.665 34.885 144.075 ;
        RECT 35.100 143.485 35.270 143.905 ;
        RECT 35.470 143.665 35.800 144.075 ;
        RECT 32.830 143.285 33.460 143.455 ;
        RECT 31.385 142.515 31.715 142.765 ;
        RECT 29.230 141.525 29.470 142.035 ;
        RECT 29.650 141.705 29.930 142.035 ;
        RECT 30.160 141.525 30.375 142.035 ;
        RECT 30.545 141.695 31.160 142.265 ;
        RECT 31.405 141.525 31.635 142.345 ;
        RECT 31.885 142.325 32.135 142.925 ;
        RECT 32.745 142.435 33.110 143.115 ;
        RECT 33.290 142.765 33.460 143.285 ;
        RECT 33.810 143.315 35.825 143.485 ;
        RECT 33.290 142.435 33.640 142.765 ;
        RECT 31.805 141.695 32.135 142.325 ;
        RECT 32.305 141.525 32.515 142.345 ;
        RECT 33.290 142.265 33.460 142.435 ;
        RECT 32.830 142.095 33.460 142.265 ;
        RECT 32.830 141.695 33.005 142.095 ;
        RECT 33.810 142.025 33.980 143.315 ;
        RECT 33.175 141.525 33.505 141.905 ;
        RECT 33.750 141.695 33.980 142.025 ;
        RECT 34.180 141.860 34.460 143.135 ;
        RECT 34.685 143.055 34.955 143.135 ;
        RECT 34.645 142.885 34.955 143.055 ;
        RECT 34.685 141.860 34.955 142.885 ;
        RECT 35.145 142.105 35.485 143.135 ;
        RECT 35.655 142.765 35.825 143.315 ;
        RECT 35.995 142.935 36.255 143.905 ;
        RECT 36.425 143.640 41.770 144.075 ;
        RECT 35.655 142.435 35.915 142.765 ;
        RECT 36.085 142.245 36.255 142.935 ;
        RECT 35.415 141.525 35.745 141.905 ;
        RECT 35.915 141.780 36.255 142.245 ;
        RECT 38.010 142.070 38.350 142.900 ;
        RECT 39.830 142.390 40.180 143.640 ;
        RECT 41.945 142.985 43.615 144.075 ;
        RECT 41.945 142.295 42.695 142.815 ;
        RECT 42.865 142.465 43.615 142.985 ;
        RECT 44.245 142.910 44.535 144.075 ;
        RECT 44.705 143.640 50.050 144.075 ;
        RECT 35.915 141.735 36.250 141.780 ;
        RECT 36.425 141.525 41.770 142.070 ;
        RECT 41.945 141.525 43.615 142.295 ;
        RECT 44.245 141.525 44.535 142.250 ;
        RECT 46.290 142.070 46.630 142.900 ;
        RECT 48.110 142.390 48.460 143.640 ;
        RECT 50.885 143.405 51.165 144.075 ;
        RECT 51.335 143.185 51.635 143.735 ;
        RECT 51.835 143.355 52.165 144.075 ;
        RECT 52.355 143.355 52.815 143.905 ;
        RECT 50.700 142.765 50.965 143.125 ;
        RECT 51.335 143.015 52.275 143.185 ;
        RECT 52.105 142.765 52.275 143.015 ;
        RECT 50.700 142.515 51.375 142.765 ;
        RECT 51.595 142.515 51.935 142.765 ;
        RECT 52.105 142.435 52.395 142.765 ;
        RECT 52.105 142.345 52.275 142.435 ;
        RECT 50.885 142.155 52.275 142.345 ;
        RECT 44.705 141.525 50.050 142.070 ;
        RECT 50.885 141.795 51.215 142.155 ;
        RECT 52.565 141.985 52.815 143.355 ;
        RECT 52.985 142.935 53.245 144.075 ;
        RECT 53.485 143.565 55.100 143.895 ;
        RECT 53.495 142.765 53.665 143.325 ;
        RECT 53.925 143.225 55.100 143.395 ;
        RECT 55.270 143.275 55.550 144.075 ;
        RECT 53.925 142.935 54.255 143.225 ;
        RECT 54.930 143.105 55.100 143.225 ;
        RECT 54.425 142.765 54.670 143.055 ;
        RECT 54.930 142.935 55.590 143.105 ;
        RECT 55.760 142.935 56.035 143.905 ;
        RECT 56.305 143.615 56.475 144.075 ;
        RECT 56.645 143.125 56.975 143.905 ;
        RECT 57.145 143.275 57.315 144.075 ;
        RECT 55.420 142.765 55.590 142.935 ;
        RECT 52.990 142.515 53.325 142.765 ;
        RECT 53.495 142.435 54.210 142.765 ;
        RECT 54.425 142.435 55.250 142.765 ;
        RECT 55.420 142.435 55.695 142.765 ;
        RECT 53.495 142.345 53.745 142.435 ;
        RECT 51.835 141.525 52.085 141.985 ;
        RECT 52.255 141.695 52.815 141.985 ;
        RECT 52.985 141.525 53.245 142.345 ;
        RECT 53.415 141.925 53.745 142.345 ;
        RECT 55.420 142.265 55.590 142.435 ;
        RECT 53.925 142.095 55.590 142.265 ;
        RECT 55.865 142.200 56.035 142.935 ;
        RECT 53.925 141.695 54.185 142.095 ;
        RECT 54.355 141.525 54.685 141.925 ;
        RECT 54.855 141.745 55.025 142.095 ;
        RECT 55.195 141.525 55.570 141.925 ;
        RECT 55.760 141.855 56.035 142.200 ;
        RECT 56.205 143.105 56.975 143.125 ;
        RECT 57.485 143.105 57.815 143.905 ;
        RECT 57.985 143.275 58.155 144.075 ;
        RECT 58.325 143.105 58.655 143.905 ;
        RECT 56.205 142.935 58.655 143.105 ;
        RECT 58.915 142.935 59.210 144.075 ;
        RECT 59.435 142.965 59.730 144.075 ;
        RECT 56.205 142.345 56.555 142.935 ;
        RECT 59.910 142.765 60.160 143.900 ;
        RECT 60.330 142.965 60.590 144.075 ;
        RECT 60.760 143.175 61.020 143.900 ;
        RECT 61.190 143.345 61.450 144.075 ;
        RECT 61.620 143.175 61.880 143.900 ;
        RECT 62.050 143.345 62.310 144.075 ;
        RECT 62.480 143.175 62.740 143.900 ;
        RECT 62.910 143.345 63.170 144.075 ;
        RECT 63.340 143.175 63.600 143.900 ;
        RECT 63.770 143.345 64.065 144.075 ;
        RECT 60.760 142.935 64.070 143.175 ;
        RECT 56.725 142.515 59.235 142.765 ;
        RECT 56.205 142.165 58.575 142.345 ;
        RECT 56.305 141.525 56.555 141.990 ;
        RECT 56.725 141.695 56.895 142.165 ;
        RECT 57.145 141.525 57.315 141.985 ;
        RECT 57.565 141.695 57.735 142.165 ;
        RECT 57.985 141.525 58.155 141.985 ;
        RECT 58.405 141.695 58.575 142.165 ;
        RECT 59.425 142.155 59.740 142.765 ;
        RECT 59.910 142.515 62.930 142.765 ;
        RECT 58.945 141.525 59.210 141.985 ;
        RECT 59.485 141.525 59.730 141.985 ;
        RECT 59.910 141.705 60.160 142.515 ;
        RECT 63.100 142.345 64.070 142.935 ;
        RECT 60.760 142.175 64.070 142.345 ;
        RECT 60.330 141.525 60.590 142.050 ;
        RECT 60.760 141.720 61.020 142.175 ;
        RECT 61.190 141.525 61.450 142.005 ;
        RECT 61.620 141.720 61.880 142.175 ;
        RECT 62.050 141.525 62.310 142.005 ;
        RECT 62.480 141.720 62.740 142.175 ;
        RECT 62.910 141.525 63.170 142.005 ;
        RECT 63.340 141.720 63.600 142.175 ;
        RECT 63.770 141.525 64.070 142.005 ;
        RECT 64.485 141.695 64.745 143.905 ;
        RECT 64.915 143.695 65.245 144.075 ;
        RECT 65.670 143.525 65.840 143.905 ;
        RECT 66.100 143.695 66.430 144.075 ;
        RECT 66.625 143.525 66.795 143.905 ;
        RECT 67.005 143.695 67.335 144.075 ;
        RECT 67.585 143.525 67.775 143.905 ;
        RECT 68.015 143.695 68.345 144.075 ;
        RECT 68.655 143.575 68.915 143.905 ;
        RECT 64.915 143.355 66.865 143.525 ;
        RECT 64.915 142.435 65.085 143.355 ;
        RECT 65.455 142.765 65.650 143.075 ;
        RECT 65.920 142.765 66.105 143.075 ;
        RECT 65.395 142.435 65.650 142.765 ;
        RECT 65.875 142.435 66.105 142.765 ;
        RECT 64.915 141.525 65.245 141.905 ;
        RECT 65.455 141.860 65.650 142.435 ;
        RECT 65.920 141.855 66.105 142.435 ;
        RECT 66.355 141.865 66.525 142.765 ;
        RECT 66.695 142.365 66.865 143.355 ;
        RECT 67.035 143.355 67.775 143.525 ;
        RECT 67.035 142.845 67.205 143.355 ;
        RECT 67.375 143.015 67.955 143.185 ;
        RECT 68.225 143.065 68.575 143.395 ;
        RECT 67.785 142.895 67.955 143.015 ;
        RECT 68.745 142.895 68.915 143.575 ;
        RECT 70.005 142.910 70.295 144.075 ;
        RECT 70.465 143.000 70.735 143.905 ;
        RECT 70.905 143.315 71.235 144.075 ;
        RECT 71.415 143.145 71.585 143.905 ;
        RECT 71.845 143.640 77.190 144.075 ;
        RECT 77.365 143.640 82.710 144.075 ;
        RECT 67.035 142.675 67.605 142.845 ;
        RECT 67.785 142.725 68.915 142.895 ;
        RECT 66.695 142.035 67.245 142.365 ;
        RECT 67.435 142.195 67.605 142.675 ;
        RECT 67.775 142.385 68.395 142.555 ;
        RECT 68.185 142.205 68.395 142.385 ;
        RECT 67.435 141.865 67.835 142.195 ;
        RECT 68.745 142.025 68.915 142.725 ;
        RECT 66.355 141.695 67.835 141.865 ;
        RECT 68.015 141.525 68.345 141.905 ;
        RECT 68.655 141.695 68.915 142.025 ;
        RECT 70.005 141.525 70.295 142.250 ;
        RECT 70.465 142.200 70.635 143.000 ;
        RECT 70.920 142.975 71.585 143.145 ;
        RECT 70.920 142.830 71.090 142.975 ;
        RECT 70.805 142.500 71.090 142.830 ;
        RECT 70.920 142.245 71.090 142.500 ;
        RECT 71.325 142.425 71.655 142.795 ;
        RECT 70.465 141.695 70.725 142.200 ;
        RECT 70.920 142.075 71.585 142.245 ;
        RECT 70.905 141.525 71.235 141.905 ;
        RECT 71.415 141.695 71.585 142.075 ;
        RECT 73.430 142.070 73.770 142.900 ;
        RECT 75.250 142.390 75.600 143.640 ;
        RECT 78.950 142.070 79.290 142.900 ;
        RECT 80.770 142.390 81.120 143.640 ;
        RECT 82.885 142.985 84.095 144.075 ;
        RECT 82.885 142.445 83.405 142.985 ;
        RECT 83.575 142.275 84.095 142.815 ;
        RECT 71.845 141.525 77.190 142.070 ;
        RECT 77.365 141.525 82.710 142.070 ;
        RECT 82.885 141.525 84.095 142.275 ;
        RECT 5.520 141.355 84.180 141.525 ;
        RECT 5.605 140.605 6.815 141.355 ;
        RECT 6.985 140.810 12.330 141.355 ;
        RECT 5.605 140.065 6.125 140.605 ;
        RECT 6.295 139.895 6.815 140.435 ;
        RECT 8.570 139.980 8.910 140.810 ;
        RECT 12.505 140.585 15.095 141.355 ;
        RECT 15.265 140.895 15.825 141.185 ;
        RECT 15.995 140.895 16.245 141.355 ;
        RECT 5.605 138.805 6.815 139.895 ;
        RECT 10.390 139.240 10.740 140.490 ;
        RECT 12.505 140.065 13.715 140.585 ;
        RECT 13.885 139.895 15.095 140.415 ;
        RECT 6.985 138.805 12.330 139.240 ;
        RECT 12.505 138.805 15.095 139.895 ;
        RECT 15.265 139.525 15.515 140.895 ;
        RECT 16.865 140.725 17.195 141.085 ;
        RECT 17.730 140.845 17.970 141.355 ;
        RECT 18.150 140.845 18.430 141.175 ;
        RECT 18.660 140.845 18.875 141.355 ;
        RECT 15.805 140.535 17.195 140.725 ;
        RECT 15.805 140.445 15.975 140.535 ;
        RECT 15.685 140.115 15.975 140.445 ;
        RECT 16.145 140.115 16.485 140.365 ;
        RECT 16.705 140.115 17.380 140.365 ;
        RECT 17.625 140.115 17.980 140.675 ;
        RECT 15.805 139.865 15.975 140.115 ;
        RECT 15.805 139.695 16.745 139.865 ;
        RECT 17.115 139.755 17.380 140.115 ;
        RECT 18.150 139.945 18.320 140.845 ;
        RECT 18.490 140.115 18.755 140.675 ;
        RECT 19.045 140.615 19.660 141.185 ;
        RECT 19.865 140.855 20.205 141.355 ;
        RECT 19.005 139.945 19.175 140.445 ;
        RECT 17.750 139.775 19.175 139.945 ;
        RECT 15.265 138.975 15.725 139.525 ;
        RECT 15.915 138.805 16.245 139.525 ;
        RECT 16.445 139.145 16.745 139.695 ;
        RECT 17.750 139.600 18.140 139.775 ;
        RECT 16.915 138.805 17.195 139.475 ;
        RECT 18.625 138.805 18.955 139.605 ;
        RECT 19.345 139.595 19.660 140.615 ;
        RECT 19.865 140.115 20.205 140.685 ;
        RECT 20.375 140.445 20.620 141.135 ;
        RECT 20.815 140.855 21.145 141.355 ;
        RECT 21.345 140.785 21.515 141.135 ;
        RECT 21.690 140.955 22.020 141.355 ;
        RECT 22.190 140.785 22.360 141.135 ;
        RECT 22.530 140.955 22.910 141.355 ;
        RECT 21.345 140.615 22.930 140.785 ;
        RECT 23.100 140.680 23.375 141.025 ;
        RECT 23.605 140.895 23.850 141.355 ;
        RECT 22.760 140.445 22.930 140.615 ;
        RECT 20.375 140.115 21.030 140.445 ;
        RECT 19.125 138.975 19.660 139.595 ;
        RECT 19.865 138.805 20.205 139.880 ;
        RECT 20.375 139.520 20.615 140.115 ;
        RECT 20.810 139.655 21.130 139.945 ;
        RECT 21.300 139.825 22.040 140.445 ;
        RECT 22.210 140.115 22.590 140.445 ;
        RECT 22.760 140.115 23.035 140.445 ;
        RECT 22.760 139.945 22.930 140.115 ;
        RECT 23.205 139.945 23.375 140.680 ;
        RECT 23.545 140.115 23.860 140.725 ;
        RECT 24.030 140.365 24.280 141.175 ;
        RECT 24.450 140.830 24.710 141.355 ;
        RECT 24.880 140.705 25.140 141.160 ;
        RECT 25.310 140.875 25.570 141.355 ;
        RECT 25.740 140.705 26.000 141.160 ;
        RECT 26.170 140.875 26.430 141.355 ;
        RECT 26.600 140.705 26.860 141.160 ;
        RECT 27.030 140.875 27.290 141.355 ;
        RECT 27.460 140.705 27.720 141.160 ;
        RECT 27.890 140.875 28.190 141.355 ;
        RECT 28.885 140.725 29.265 141.175 ;
        RECT 24.880 140.535 28.190 140.705 ;
        RECT 24.030 140.115 27.050 140.365 ;
        RECT 22.270 139.775 22.930 139.945 ;
        RECT 22.270 139.655 22.440 139.775 ;
        RECT 20.810 139.485 22.440 139.655 ;
        RECT 20.385 139.145 22.440 139.315 ;
        RECT 20.390 139.025 22.440 139.145 ;
        RECT 22.610 138.805 22.890 139.605 ;
        RECT 23.100 138.975 23.375 139.945 ;
        RECT 23.555 138.805 23.850 139.915 ;
        RECT 24.030 138.980 24.280 140.115 ;
        RECT 27.220 139.945 28.190 140.535 ;
        RECT 24.450 138.805 24.710 139.915 ;
        RECT 24.880 139.705 28.190 139.945 ;
        RECT 28.625 139.775 28.855 140.465 ;
        RECT 29.035 140.275 29.265 140.725 ;
        RECT 29.445 140.575 29.675 141.355 ;
        RECT 29.855 140.645 30.285 141.175 ;
        RECT 29.855 140.395 30.100 140.645 ;
        RECT 30.465 140.445 30.675 141.065 ;
        RECT 30.845 140.625 31.175 141.355 ;
        RECT 31.365 140.630 31.655 141.355 ;
        RECT 31.835 140.865 32.165 141.355 ;
        RECT 32.335 140.760 32.955 141.185 ;
        RECT 24.880 138.980 25.140 139.705 ;
        RECT 25.310 138.805 25.570 139.535 ;
        RECT 25.740 138.980 26.000 139.705 ;
        RECT 26.170 138.805 26.430 139.535 ;
        RECT 26.600 138.980 26.860 139.705 ;
        RECT 27.030 138.805 27.290 139.535 ;
        RECT 27.460 138.980 27.720 139.705 ;
        RECT 29.035 139.595 29.375 140.275 ;
        RECT 27.890 138.805 28.185 139.535 ;
        RECT 28.615 139.395 29.375 139.595 ;
        RECT 29.565 140.095 30.100 140.395 ;
        RECT 30.280 140.095 30.675 140.445 ;
        RECT 30.870 140.095 31.160 140.445 ;
        RECT 31.825 140.115 32.165 140.695 ;
        RECT 32.335 140.425 32.695 140.760 ;
        RECT 33.415 140.665 33.745 141.355 ;
        RECT 34.585 140.680 34.845 141.185 ;
        RECT 35.025 140.975 35.355 141.355 ;
        RECT 35.535 140.805 35.705 141.185 ;
        RECT 32.335 140.145 33.755 140.425 ;
        RECT 28.615 139.005 28.875 139.395 ;
        RECT 29.045 138.805 29.375 139.215 ;
        RECT 29.565 138.985 29.895 140.095 ;
        RECT 30.065 139.715 31.105 139.915 ;
        RECT 30.065 138.985 30.255 139.715 ;
        RECT 30.425 138.805 30.755 139.535 ;
        RECT 30.935 138.985 31.105 139.715 ;
        RECT 31.365 138.805 31.655 139.970 ;
        RECT 31.835 138.805 32.165 139.945 ;
        RECT 32.335 138.975 32.695 140.145 ;
        RECT 32.895 138.805 33.225 139.975 ;
        RECT 33.425 138.975 33.755 140.145 ;
        RECT 33.955 138.805 34.285 139.975 ;
        RECT 34.585 139.880 34.755 140.680 ;
        RECT 35.040 140.635 35.705 140.805 ;
        RECT 35.040 140.380 35.210 140.635 ;
        RECT 36.895 140.545 37.165 141.355 ;
        RECT 37.335 140.545 37.665 141.185 ;
        RECT 37.835 140.545 38.075 141.355 ;
        RECT 38.265 140.585 39.935 141.355 ;
        RECT 34.925 140.050 35.210 140.380 ;
        RECT 35.445 140.085 35.775 140.455 ;
        RECT 36.885 140.115 37.235 140.365 ;
        RECT 35.040 139.905 35.210 140.050 ;
        RECT 37.405 139.945 37.575 140.545 ;
        RECT 37.745 140.115 38.095 140.365 ;
        RECT 38.265 140.065 39.015 140.585 ;
        RECT 40.575 140.545 40.845 141.355 ;
        RECT 41.015 140.545 41.345 141.185 ;
        RECT 41.515 140.545 41.755 141.355 ;
        RECT 41.950 140.955 42.285 141.355 ;
        RECT 42.455 140.785 42.660 141.185 ;
        RECT 42.870 140.875 43.145 141.355 ;
        RECT 43.355 140.855 43.615 141.185 ;
        RECT 41.975 140.615 42.660 140.785 ;
        RECT 34.585 138.975 34.855 139.880 ;
        RECT 35.040 139.735 35.705 139.905 ;
        RECT 35.025 138.805 35.355 139.565 ;
        RECT 35.535 138.975 35.705 139.735 ;
        RECT 36.895 138.805 37.225 139.945 ;
        RECT 37.405 139.775 38.085 139.945 ;
        RECT 39.185 139.895 39.935 140.415 ;
        RECT 40.565 140.115 40.915 140.365 ;
        RECT 41.085 139.945 41.255 140.545 ;
        RECT 41.425 140.115 41.775 140.365 ;
        RECT 37.755 138.990 38.085 139.775 ;
        RECT 38.265 138.805 39.935 139.895 ;
        RECT 40.575 138.805 40.905 139.945 ;
        RECT 41.085 139.775 41.765 139.945 ;
        RECT 41.435 138.990 41.765 139.775 ;
        RECT 41.975 139.585 42.315 140.615 ;
        RECT 42.485 139.945 42.735 140.445 ;
        RECT 42.915 140.115 43.275 140.695 ;
        RECT 43.445 139.945 43.615 140.855 ;
        RECT 43.835 140.700 44.165 141.135 ;
        RECT 44.335 140.745 44.505 141.355 ;
        RECT 42.485 139.775 43.615 139.945 ;
        RECT 43.785 140.615 44.165 140.700 ;
        RECT 44.675 140.615 45.005 141.140 ;
        RECT 45.265 140.825 45.475 141.355 ;
        RECT 45.750 140.905 46.535 141.075 ;
        RECT 46.705 140.905 47.110 141.075 ;
        RECT 43.785 140.575 44.010 140.615 ;
        RECT 43.785 139.995 43.955 140.575 ;
        RECT 44.675 140.445 44.875 140.615 ;
        RECT 45.750 140.445 45.920 140.905 ;
        RECT 44.125 140.115 44.875 140.445 ;
        RECT 45.045 140.115 45.920 140.445 ;
        RECT 43.785 139.945 44.000 139.995 ;
        RECT 43.785 139.865 44.175 139.945 ;
        RECT 41.975 139.410 42.640 139.585 ;
        RECT 41.950 138.805 42.285 139.230 ;
        RECT 42.455 139.005 42.640 139.410 ;
        RECT 42.845 138.805 43.175 139.585 ;
        RECT 43.345 139.005 43.615 139.775 ;
        RECT 43.845 139.020 44.175 139.865 ;
        RECT 44.685 139.910 44.875 140.115 ;
        RECT 44.345 138.805 44.515 139.815 ;
        RECT 44.685 139.535 45.580 139.910 ;
        RECT 44.685 138.975 45.025 139.535 ;
        RECT 45.255 138.805 45.570 139.305 ;
        RECT 45.750 139.275 45.920 140.115 ;
        RECT 46.090 140.405 46.555 140.735 ;
        RECT 46.940 140.675 47.110 140.905 ;
        RECT 47.290 140.855 47.660 141.355 ;
        RECT 47.980 140.905 48.655 141.075 ;
        RECT 48.850 140.905 49.185 141.075 ;
        RECT 46.090 139.445 46.410 140.405 ;
        RECT 46.940 140.375 47.770 140.675 ;
        RECT 46.580 139.475 46.770 140.195 ;
        RECT 46.940 139.305 47.110 140.375 ;
        RECT 47.570 140.345 47.770 140.375 ;
        RECT 47.280 140.125 47.450 140.195 ;
        RECT 47.980 140.125 48.150 140.905 ;
        RECT 49.015 140.765 49.185 140.905 ;
        RECT 49.355 140.895 49.605 141.355 ;
        RECT 47.280 139.955 48.150 140.125 ;
        RECT 48.320 140.485 48.845 140.705 ;
        RECT 49.015 140.635 49.240 140.765 ;
        RECT 47.280 139.865 47.790 139.955 ;
        RECT 45.750 139.105 46.635 139.275 ;
        RECT 46.860 138.975 47.110 139.305 ;
        RECT 47.280 138.805 47.450 139.605 ;
        RECT 47.620 139.250 47.790 139.865 ;
        RECT 48.320 139.785 48.490 140.485 ;
        RECT 47.960 139.420 48.490 139.785 ;
        RECT 48.660 139.720 48.900 140.315 ;
        RECT 49.070 139.530 49.240 140.635 ;
        RECT 49.410 139.775 49.690 140.725 ;
        RECT 48.935 139.400 49.240 139.530 ;
        RECT 47.620 139.080 48.725 139.250 ;
        RECT 48.935 138.975 49.185 139.400 ;
        RECT 49.355 138.805 49.620 139.265 ;
        RECT 49.860 138.975 50.045 141.095 ;
        RECT 50.215 140.975 50.545 141.355 ;
        RECT 50.715 140.805 50.885 141.095 ;
        RECT 50.220 140.635 50.885 140.805 ;
        RECT 50.220 139.645 50.450 140.635 ;
        RECT 50.620 139.815 50.970 140.465 ;
        RECT 50.220 139.475 50.885 139.645 ;
        RECT 50.215 138.805 50.545 139.305 ;
        RECT 50.715 138.975 50.885 139.475 ;
        RECT 52.065 138.975 52.345 141.075 ;
        RECT 52.575 140.895 52.745 141.355 ;
        RECT 53.015 140.965 54.265 141.145 ;
        RECT 53.400 140.725 53.765 140.795 ;
        RECT 52.515 140.545 53.765 140.725 ;
        RECT 53.935 140.745 54.265 140.965 ;
        RECT 54.435 140.915 54.605 141.355 ;
        RECT 54.775 140.745 55.115 141.160 ;
        RECT 53.935 140.575 55.115 140.745 ;
        RECT 55.285 140.585 56.955 141.355 ;
        RECT 57.125 140.630 57.415 141.355 ;
        RECT 52.515 139.945 52.790 140.545 ;
        RECT 52.960 140.115 53.315 140.365 ;
        RECT 53.510 140.335 53.975 140.365 ;
        RECT 53.505 140.165 53.975 140.335 ;
        RECT 53.510 140.115 53.975 140.165 ;
        RECT 54.145 140.115 54.475 140.365 ;
        RECT 54.650 140.165 55.115 140.365 ;
        RECT 54.295 139.995 54.475 140.115 ;
        RECT 55.285 140.065 56.035 140.585 ;
        RECT 52.515 139.735 54.125 139.945 ;
        RECT 54.295 139.825 54.625 139.995 ;
        RECT 53.715 139.635 54.125 139.735 ;
        RECT 52.535 138.805 53.320 139.565 ;
        RECT 53.715 138.975 54.100 139.635 ;
        RECT 54.425 139.035 54.625 139.825 ;
        RECT 54.795 138.805 55.115 139.985 ;
        RECT 56.205 139.895 56.955 140.415 ;
        RECT 57.585 140.410 57.925 141.185 ;
        RECT 58.095 140.895 58.265 141.355 ;
        RECT 58.505 140.920 58.865 141.185 ;
        RECT 58.505 140.915 58.860 140.920 ;
        RECT 58.505 140.905 58.855 140.915 ;
        RECT 58.505 140.900 58.850 140.905 ;
        RECT 58.505 140.890 58.845 140.900 ;
        RECT 59.495 140.895 59.665 141.355 ;
        RECT 58.505 140.885 58.840 140.890 ;
        RECT 58.505 140.875 58.830 140.885 ;
        RECT 58.505 140.865 58.820 140.875 ;
        RECT 58.505 140.725 58.805 140.865 ;
        RECT 58.095 140.535 58.805 140.725 ;
        RECT 58.995 140.725 59.325 140.805 ;
        RECT 59.835 140.725 60.175 141.185 ;
        RECT 58.995 140.535 60.175 140.725 ;
        RECT 60.345 140.585 62.015 141.355 ;
        RECT 62.275 140.805 62.445 141.095 ;
        RECT 62.615 140.975 62.945 141.355 ;
        RECT 62.275 140.635 62.940 140.805 ;
        RECT 55.285 138.805 56.955 139.895 ;
        RECT 57.125 138.805 57.415 139.970 ;
        RECT 57.585 138.975 57.865 140.410 ;
        RECT 58.095 139.965 58.380 140.535 ;
        RECT 58.565 140.135 59.035 140.365 ;
        RECT 59.205 140.345 59.535 140.365 ;
        RECT 59.205 140.165 59.655 140.345 ;
        RECT 59.845 140.165 60.175 140.365 ;
        RECT 58.095 139.750 59.245 139.965 ;
        RECT 58.035 138.805 58.745 139.580 ;
        RECT 58.915 138.975 59.245 139.750 ;
        RECT 59.440 139.050 59.655 140.165 ;
        RECT 59.945 139.825 60.175 140.165 ;
        RECT 60.345 140.065 61.095 140.585 ;
        RECT 61.265 139.895 62.015 140.415 ;
        RECT 59.835 138.805 60.165 139.525 ;
        RECT 60.345 138.805 62.015 139.895 ;
        RECT 62.190 139.815 62.540 140.465 ;
        RECT 62.710 139.645 62.940 140.635 ;
        RECT 62.275 139.475 62.940 139.645 ;
        RECT 62.275 138.975 62.445 139.475 ;
        RECT 62.615 138.805 62.945 139.305 ;
        RECT 63.115 138.975 63.300 141.095 ;
        RECT 63.555 140.895 63.805 141.355 ;
        RECT 63.975 140.905 64.310 141.075 ;
        RECT 64.505 140.905 65.180 141.075 ;
        RECT 63.975 140.765 64.145 140.905 ;
        RECT 63.470 139.775 63.750 140.725 ;
        RECT 63.920 140.635 64.145 140.765 ;
        RECT 63.920 139.530 64.090 140.635 ;
        RECT 64.315 140.485 64.840 140.705 ;
        RECT 64.260 139.720 64.500 140.315 ;
        RECT 64.670 139.785 64.840 140.485 ;
        RECT 65.010 140.125 65.180 140.905 ;
        RECT 65.500 140.855 65.870 141.355 ;
        RECT 66.050 140.905 66.455 141.075 ;
        RECT 66.625 140.905 67.410 141.075 ;
        RECT 66.050 140.675 66.220 140.905 ;
        RECT 65.390 140.375 66.220 140.675 ;
        RECT 66.605 140.405 67.070 140.735 ;
        RECT 65.390 140.345 65.590 140.375 ;
        RECT 65.710 140.125 65.880 140.195 ;
        RECT 65.010 139.955 65.880 140.125 ;
        RECT 65.370 139.865 65.880 139.955 ;
        RECT 63.920 139.400 64.225 139.530 ;
        RECT 64.670 139.420 65.200 139.785 ;
        RECT 63.540 138.805 63.805 139.265 ;
        RECT 63.975 138.975 64.225 139.400 ;
        RECT 65.370 139.250 65.540 139.865 ;
        RECT 64.435 139.080 65.540 139.250 ;
        RECT 65.710 138.805 65.880 139.605 ;
        RECT 66.050 139.305 66.220 140.375 ;
        RECT 66.390 139.475 66.580 140.195 ;
        RECT 66.750 139.445 67.070 140.405 ;
        RECT 67.240 140.445 67.410 140.905 ;
        RECT 67.685 140.825 67.895 141.355 ;
        RECT 68.155 140.615 68.485 141.140 ;
        RECT 68.655 140.745 68.825 141.355 ;
        RECT 68.995 140.700 69.325 141.135 ;
        RECT 69.545 140.810 74.890 141.355 ;
        RECT 75.065 140.810 80.410 141.355 ;
        RECT 68.995 140.615 69.375 140.700 ;
        RECT 68.285 140.445 68.485 140.615 ;
        RECT 69.150 140.575 69.375 140.615 ;
        RECT 67.240 140.115 68.115 140.445 ;
        RECT 68.285 140.115 69.035 140.445 ;
        RECT 66.050 138.975 66.300 139.305 ;
        RECT 67.240 139.275 67.410 140.115 ;
        RECT 68.285 139.910 68.475 140.115 ;
        RECT 69.205 139.995 69.375 140.575 ;
        RECT 69.160 139.945 69.375 139.995 ;
        RECT 71.130 139.980 71.470 140.810 ;
        RECT 67.580 139.535 68.475 139.910 ;
        RECT 68.985 139.865 69.375 139.945 ;
        RECT 66.525 139.105 67.410 139.275 ;
        RECT 67.590 138.805 67.905 139.305 ;
        RECT 68.135 138.975 68.475 139.535 ;
        RECT 68.645 138.805 68.815 139.815 ;
        RECT 68.985 139.020 69.315 139.865 ;
        RECT 72.950 139.240 73.300 140.490 ;
        RECT 76.650 139.980 76.990 140.810 ;
        RECT 80.585 140.585 82.255 141.355 ;
        RECT 82.885 140.605 84.095 141.355 ;
        RECT 78.470 139.240 78.820 140.490 ;
        RECT 80.585 140.065 81.335 140.585 ;
        RECT 81.505 139.895 82.255 140.415 ;
        RECT 69.545 138.805 74.890 139.240 ;
        RECT 75.065 138.805 80.410 139.240 ;
        RECT 80.585 138.805 82.255 139.895 ;
        RECT 82.885 139.895 83.405 140.435 ;
        RECT 83.575 140.065 84.095 140.605 ;
        RECT 82.885 138.805 84.095 139.895 ;
        RECT 5.520 138.635 84.180 138.805 ;
        RECT 5.605 137.545 6.815 138.635 ;
        RECT 6.985 137.545 10.495 138.635 ;
        RECT 11.215 137.965 11.385 138.465 ;
        RECT 11.555 138.135 11.885 138.635 ;
        RECT 11.215 137.795 11.880 137.965 ;
        RECT 5.605 136.835 6.125 137.375 ;
        RECT 6.295 137.005 6.815 137.545 ;
        RECT 6.985 136.855 8.635 137.375 ;
        RECT 8.805 137.025 10.495 137.545 ;
        RECT 11.130 136.975 11.480 137.625 ;
        RECT 5.605 136.085 6.815 136.835 ;
        RECT 6.985 136.085 10.495 136.855 ;
        RECT 11.650 136.805 11.880 137.795 ;
        RECT 11.215 136.635 11.880 136.805 ;
        RECT 11.215 136.345 11.385 136.635 ;
        RECT 11.555 136.085 11.885 136.465 ;
        RECT 12.055 136.345 12.240 138.465 ;
        RECT 12.480 138.175 12.745 138.635 ;
        RECT 12.915 138.040 13.165 138.465 ;
        RECT 13.375 138.190 14.480 138.360 ;
        RECT 12.860 137.910 13.165 138.040 ;
        RECT 12.410 136.715 12.690 137.665 ;
        RECT 12.860 136.805 13.030 137.910 ;
        RECT 13.200 137.125 13.440 137.720 ;
        RECT 13.610 137.655 14.140 138.020 ;
        RECT 13.610 136.955 13.780 137.655 ;
        RECT 14.310 137.575 14.480 138.190 ;
        RECT 14.650 137.835 14.820 138.635 ;
        RECT 14.990 138.135 15.240 138.465 ;
        RECT 15.465 138.165 16.350 138.335 ;
        RECT 14.310 137.485 14.820 137.575 ;
        RECT 12.860 136.675 13.085 136.805 ;
        RECT 13.255 136.735 13.780 136.955 ;
        RECT 13.950 137.315 14.820 137.485 ;
        RECT 12.495 136.085 12.745 136.545 ;
        RECT 12.915 136.535 13.085 136.675 ;
        RECT 13.950 136.535 14.120 137.315 ;
        RECT 14.650 137.245 14.820 137.315 ;
        RECT 14.330 137.065 14.530 137.095 ;
        RECT 14.990 137.065 15.160 138.135 ;
        RECT 15.330 137.245 15.520 137.965 ;
        RECT 14.330 136.765 15.160 137.065 ;
        RECT 15.690 137.035 16.010 137.995 ;
        RECT 12.915 136.365 13.250 136.535 ;
        RECT 13.445 136.365 14.120 136.535 ;
        RECT 14.440 136.085 14.810 136.585 ;
        RECT 14.990 136.535 15.160 136.765 ;
        RECT 15.545 136.705 16.010 137.035 ;
        RECT 16.180 137.325 16.350 138.165 ;
        RECT 16.530 138.135 16.845 138.635 ;
        RECT 17.075 137.905 17.415 138.465 ;
        RECT 16.520 137.530 17.415 137.905 ;
        RECT 17.585 137.625 17.755 138.635 ;
        RECT 17.225 137.325 17.415 137.530 ;
        RECT 17.925 137.575 18.255 138.420 ;
        RECT 17.925 137.495 18.315 137.575 ;
        RECT 18.100 137.445 18.315 137.495 ;
        RECT 18.485 137.470 18.775 138.635 ;
        RECT 19.405 137.665 19.675 138.435 ;
        RECT 19.845 137.855 20.175 138.635 ;
        RECT 20.380 138.030 20.565 138.435 ;
        RECT 20.735 138.210 21.070 138.635 ;
        RECT 20.380 137.855 21.045 138.030 ;
        RECT 19.405 137.495 20.535 137.665 ;
        RECT 16.180 136.995 17.055 137.325 ;
        RECT 17.225 136.995 17.975 137.325 ;
        RECT 16.180 136.535 16.350 136.995 ;
        RECT 17.225 136.825 17.425 136.995 ;
        RECT 18.145 136.865 18.315 137.445 ;
        RECT 18.090 136.825 18.315 136.865 ;
        RECT 14.990 136.365 15.395 136.535 ;
        RECT 15.565 136.365 16.350 136.535 ;
        RECT 16.625 136.085 16.835 136.615 ;
        RECT 17.095 136.300 17.425 136.825 ;
        RECT 17.935 136.740 18.315 136.825 ;
        RECT 17.595 136.085 17.765 136.695 ;
        RECT 17.935 136.305 18.265 136.740 ;
        RECT 18.485 136.085 18.775 136.810 ;
        RECT 19.405 136.585 19.575 137.495 ;
        RECT 19.745 136.745 20.105 137.325 ;
        RECT 20.285 136.995 20.535 137.495 ;
        RECT 20.705 136.825 21.045 137.855 ;
        RECT 21.305 137.575 21.635 138.420 ;
        RECT 21.805 137.625 21.975 138.635 ;
        RECT 22.145 137.905 22.485 138.465 ;
        RECT 22.715 138.135 23.030 138.635 ;
        RECT 23.210 138.165 24.095 138.335 ;
        RECT 20.360 136.655 21.045 136.825 ;
        RECT 21.245 137.495 21.635 137.575 ;
        RECT 22.145 137.530 23.040 137.905 ;
        RECT 21.245 137.445 21.460 137.495 ;
        RECT 21.245 136.865 21.415 137.445 ;
        RECT 22.145 137.325 22.335 137.530 ;
        RECT 23.210 137.325 23.380 138.165 ;
        RECT 24.320 138.135 24.570 138.465 ;
        RECT 21.585 136.995 22.335 137.325 ;
        RECT 22.505 136.995 23.380 137.325 ;
        RECT 21.245 136.825 21.470 136.865 ;
        RECT 22.135 136.825 22.335 136.995 ;
        RECT 21.245 136.740 21.625 136.825 ;
        RECT 19.405 136.255 19.665 136.585 ;
        RECT 19.875 136.085 20.150 136.565 ;
        RECT 20.360 136.255 20.565 136.655 ;
        RECT 20.735 136.085 21.070 136.485 ;
        RECT 21.295 136.305 21.625 136.740 ;
        RECT 21.795 136.085 21.965 136.695 ;
        RECT 22.135 136.300 22.465 136.825 ;
        RECT 22.725 136.085 22.935 136.615 ;
        RECT 23.210 136.535 23.380 136.995 ;
        RECT 23.550 137.035 23.870 137.995 ;
        RECT 24.040 137.245 24.230 137.965 ;
        RECT 24.400 137.065 24.570 138.135 ;
        RECT 24.740 137.835 24.910 138.635 ;
        RECT 25.080 138.190 26.185 138.360 ;
        RECT 25.080 137.575 25.250 138.190 ;
        RECT 26.395 138.040 26.645 138.465 ;
        RECT 26.815 138.175 27.080 138.635 ;
        RECT 25.420 137.655 25.950 138.020 ;
        RECT 26.395 137.910 26.700 138.040 ;
        RECT 24.740 137.485 25.250 137.575 ;
        RECT 24.740 137.315 25.610 137.485 ;
        RECT 24.740 137.245 24.910 137.315 ;
        RECT 25.030 137.065 25.230 137.095 ;
        RECT 23.550 136.705 24.015 137.035 ;
        RECT 24.400 136.765 25.230 137.065 ;
        RECT 24.400 136.535 24.570 136.765 ;
        RECT 23.210 136.365 23.995 136.535 ;
        RECT 24.165 136.365 24.570 136.535 ;
        RECT 24.750 136.085 25.120 136.585 ;
        RECT 25.440 136.535 25.610 137.315 ;
        RECT 25.780 136.955 25.950 137.655 ;
        RECT 26.120 137.125 26.360 137.720 ;
        RECT 25.780 136.735 26.305 136.955 ;
        RECT 26.530 136.805 26.700 137.910 ;
        RECT 26.475 136.675 26.700 136.805 ;
        RECT 26.870 136.715 27.150 137.665 ;
        RECT 26.475 136.535 26.645 136.675 ;
        RECT 25.440 136.365 26.115 136.535 ;
        RECT 26.310 136.365 26.645 136.535 ;
        RECT 26.815 136.085 27.065 136.545 ;
        RECT 27.320 136.345 27.505 138.465 ;
        RECT 27.675 138.135 28.005 138.635 ;
        RECT 28.175 137.965 28.345 138.465 ;
        RECT 27.680 137.795 28.345 137.965 ;
        RECT 27.680 136.805 27.910 137.795 ;
        RECT 28.080 136.975 28.430 137.625 ;
        RECT 28.605 137.495 28.990 138.465 ;
        RECT 29.160 138.175 29.485 138.635 ;
        RECT 30.005 138.005 30.285 138.465 ;
        RECT 29.160 137.785 30.285 138.005 ;
        RECT 28.605 136.825 28.885 137.495 ;
        RECT 29.160 137.325 29.610 137.785 ;
        RECT 30.475 137.615 30.875 138.465 ;
        RECT 31.275 138.175 31.545 138.635 ;
        RECT 31.715 138.005 32.000 138.465 ;
        RECT 29.055 136.995 29.610 137.325 ;
        RECT 29.780 137.055 30.875 137.615 ;
        RECT 29.160 136.885 29.610 136.995 ;
        RECT 27.680 136.635 28.345 136.805 ;
        RECT 27.675 136.085 28.005 136.465 ;
        RECT 28.175 136.345 28.345 136.635 ;
        RECT 28.605 136.255 28.990 136.825 ;
        RECT 29.160 136.715 30.285 136.885 ;
        RECT 29.160 136.085 29.485 136.545 ;
        RECT 30.005 136.255 30.285 136.715 ;
        RECT 30.475 136.255 30.875 137.055 ;
        RECT 31.045 137.785 32.000 138.005 ;
        RECT 31.045 136.885 31.255 137.785 ;
        RECT 31.425 137.055 32.115 137.615 ;
        RECT 32.285 137.545 33.955 138.635 ;
        RECT 34.215 137.965 34.385 138.465 ;
        RECT 34.555 138.135 34.885 138.635 ;
        RECT 34.215 137.795 34.880 137.965 ;
        RECT 31.045 136.715 32.000 136.885 ;
        RECT 31.275 136.085 31.545 136.545 ;
        RECT 31.715 136.255 32.000 136.715 ;
        RECT 32.285 136.855 33.035 137.375 ;
        RECT 33.205 137.025 33.955 137.545 ;
        RECT 34.130 136.975 34.480 137.625 ;
        RECT 32.285 136.085 33.955 136.855 ;
        RECT 34.650 136.805 34.880 137.795 ;
        RECT 34.215 136.635 34.880 136.805 ;
        RECT 34.215 136.345 34.385 136.635 ;
        RECT 34.555 136.085 34.885 136.465 ;
        RECT 35.055 136.345 35.240 138.465 ;
        RECT 35.480 138.175 35.745 138.635 ;
        RECT 35.915 138.040 36.165 138.465 ;
        RECT 36.375 138.190 37.480 138.360 ;
        RECT 35.860 137.910 36.165 138.040 ;
        RECT 35.410 136.715 35.690 137.665 ;
        RECT 35.860 136.805 36.030 137.910 ;
        RECT 36.200 137.125 36.440 137.720 ;
        RECT 36.610 137.655 37.140 138.020 ;
        RECT 36.610 136.955 36.780 137.655 ;
        RECT 37.310 137.575 37.480 138.190 ;
        RECT 37.650 137.835 37.820 138.635 ;
        RECT 37.990 138.135 38.240 138.465 ;
        RECT 38.465 138.165 39.350 138.335 ;
        RECT 37.310 137.485 37.820 137.575 ;
        RECT 35.860 136.675 36.085 136.805 ;
        RECT 36.255 136.735 36.780 136.955 ;
        RECT 36.950 137.315 37.820 137.485 ;
        RECT 35.495 136.085 35.745 136.545 ;
        RECT 35.915 136.535 36.085 136.675 ;
        RECT 36.950 136.535 37.120 137.315 ;
        RECT 37.650 137.245 37.820 137.315 ;
        RECT 37.330 137.065 37.530 137.095 ;
        RECT 37.990 137.065 38.160 138.135 ;
        RECT 38.330 137.245 38.520 137.965 ;
        RECT 37.330 136.765 38.160 137.065 ;
        RECT 38.690 137.035 39.010 137.995 ;
        RECT 35.915 136.365 36.250 136.535 ;
        RECT 36.445 136.365 37.120 136.535 ;
        RECT 37.440 136.085 37.810 136.585 ;
        RECT 37.990 136.535 38.160 136.765 ;
        RECT 38.545 136.705 39.010 137.035 ;
        RECT 39.180 137.325 39.350 138.165 ;
        RECT 39.530 138.135 39.845 138.635 ;
        RECT 40.075 137.905 40.415 138.465 ;
        RECT 39.520 137.530 40.415 137.905 ;
        RECT 40.585 137.625 40.755 138.635 ;
        RECT 40.225 137.325 40.415 137.530 ;
        RECT 40.925 137.575 41.255 138.420 ;
        RECT 41.945 138.080 42.550 138.635 ;
        RECT 42.725 138.125 43.205 138.465 ;
        RECT 43.375 138.090 43.630 138.635 ;
        RECT 41.945 137.980 42.560 138.080 ;
        RECT 42.375 137.955 42.560 137.980 ;
        RECT 40.925 137.495 41.315 137.575 ;
        RECT 41.100 137.445 41.315 137.495 ;
        RECT 39.180 136.995 40.055 137.325 ;
        RECT 40.225 136.995 40.975 137.325 ;
        RECT 39.180 136.535 39.350 136.995 ;
        RECT 40.225 136.825 40.425 136.995 ;
        RECT 41.145 136.865 41.315 137.445 ;
        RECT 41.945 137.360 42.205 137.810 ;
        RECT 42.375 137.710 42.705 137.955 ;
        RECT 42.875 137.635 43.630 137.885 ;
        RECT 43.800 137.765 44.075 138.465 ;
        RECT 42.860 137.600 43.630 137.635 ;
        RECT 42.845 137.590 43.630 137.600 ;
        RECT 42.840 137.575 43.735 137.590 ;
        RECT 42.820 137.560 43.735 137.575 ;
        RECT 42.800 137.550 43.735 137.560 ;
        RECT 42.775 137.540 43.735 137.550 ;
        RECT 42.705 137.510 43.735 137.540 ;
        RECT 42.685 137.480 43.735 137.510 ;
        RECT 42.665 137.450 43.735 137.480 ;
        RECT 42.635 137.425 43.735 137.450 ;
        RECT 42.600 137.390 43.735 137.425 ;
        RECT 42.570 137.385 43.735 137.390 ;
        RECT 42.570 137.380 42.960 137.385 ;
        RECT 42.570 137.370 42.935 137.380 ;
        RECT 42.570 137.365 42.920 137.370 ;
        RECT 42.570 137.360 42.905 137.365 ;
        RECT 41.945 137.355 42.905 137.360 ;
        RECT 41.945 137.345 42.895 137.355 ;
        RECT 41.945 137.340 42.885 137.345 ;
        RECT 41.945 137.330 42.875 137.340 ;
        RECT 41.945 137.320 42.870 137.330 ;
        RECT 41.945 137.315 42.865 137.320 ;
        RECT 41.945 137.300 42.855 137.315 ;
        RECT 41.945 137.285 42.850 137.300 ;
        RECT 41.945 137.260 42.840 137.285 ;
        RECT 41.945 137.190 42.835 137.260 ;
        RECT 41.090 136.825 41.315 136.865 ;
        RECT 37.990 136.365 38.395 136.535 ;
        RECT 38.565 136.365 39.350 136.535 ;
        RECT 39.625 136.085 39.835 136.615 ;
        RECT 40.095 136.300 40.425 136.825 ;
        RECT 40.935 136.740 41.315 136.825 ;
        RECT 40.595 136.085 40.765 136.695 ;
        RECT 40.935 136.305 41.265 136.740 ;
        RECT 41.945 136.635 42.495 137.020 ;
        RECT 42.665 136.465 42.835 137.190 ;
        RECT 41.945 136.295 42.835 136.465 ;
        RECT 43.005 136.790 43.335 137.215 ;
        RECT 43.505 136.990 43.735 137.385 ;
        RECT 43.005 136.765 43.255 136.790 ;
        RECT 43.005 136.305 43.225 136.765 ;
        RECT 43.905 136.735 44.075 137.765 ;
        RECT 44.245 137.470 44.535 138.635 ;
        RECT 44.790 138.015 44.965 138.465 ;
        RECT 45.135 138.195 45.465 138.635 ;
        RECT 45.770 138.045 45.940 138.465 ;
        RECT 46.175 138.225 46.845 138.635 ;
        RECT 47.060 138.045 47.230 138.465 ;
        RECT 47.430 138.225 47.760 138.635 ;
        RECT 44.790 137.845 45.420 138.015 ;
        RECT 44.705 136.995 45.070 137.675 ;
        RECT 45.250 137.325 45.420 137.845 ;
        RECT 45.770 137.875 47.785 138.045 ;
        RECT 45.250 136.995 45.600 137.325 ;
        RECT 45.250 136.825 45.420 136.995 ;
        RECT 43.395 136.085 43.645 136.625 ;
        RECT 43.815 136.255 44.075 136.735 ;
        RECT 44.245 136.085 44.535 136.810 ;
        RECT 44.790 136.655 45.420 136.825 ;
        RECT 44.790 136.255 44.965 136.655 ;
        RECT 45.770 136.585 45.940 137.875 ;
        RECT 45.135 136.085 45.465 136.465 ;
        RECT 45.710 136.255 45.940 136.585 ;
        RECT 46.140 136.420 46.420 137.695 ;
        RECT 46.645 136.595 46.915 137.695 ;
        RECT 47.105 136.665 47.445 137.695 ;
        RECT 47.615 137.325 47.785 137.875 ;
        RECT 47.955 137.495 48.215 138.465 ;
        RECT 48.395 137.685 48.670 138.455 ;
        RECT 48.840 138.025 49.170 138.455 ;
        RECT 49.340 138.195 49.535 138.635 ;
        RECT 49.715 138.025 50.045 138.455 ;
        RECT 48.840 137.855 50.045 138.025 ;
        RECT 50.475 137.905 50.770 138.635 ;
        RECT 48.395 137.495 48.980 137.685 ;
        RECT 49.150 137.525 50.045 137.855 ;
        RECT 50.940 137.735 51.200 138.460 ;
        RECT 51.370 137.905 51.630 138.635 ;
        RECT 51.800 137.735 52.060 138.460 ;
        RECT 52.230 137.905 52.490 138.635 ;
        RECT 52.660 137.735 52.920 138.460 ;
        RECT 53.090 137.905 53.350 138.635 ;
        RECT 53.520 137.735 53.780 138.460 ;
        RECT 47.615 136.995 47.875 137.325 ;
        RECT 48.045 136.805 48.215 137.495 ;
        RECT 46.605 136.425 46.915 136.595 ;
        RECT 46.645 136.420 46.915 136.425 ;
        RECT 47.375 136.085 47.705 136.465 ;
        RECT 47.875 136.340 48.215 136.805 ;
        RECT 48.395 136.675 48.635 137.325 ;
        RECT 48.805 136.825 48.980 137.495 ;
        RECT 50.470 137.495 53.780 137.735 ;
        RECT 53.950 137.525 54.210 138.635 ;
        RECT 49.150 136.995 49.565 137.325 ;
        RECT 49.745 136.995 50.040 137.325 ;
        RECT 48.805 136.645 49.135 136.825 ;
        RECT 47.875 136.295 48.210 136.340 ;
        RECT 48.410 136.085 48.740 136.475 ;
        RECT 48.910 136.265 49.135 136.645 ;
        RECT 49.335 136.375 49.565 136.995 ;
        RECT 50.470 136.905 51.440 137.495 ;
        RECT 54.380 137.325 54.630 138.460 ;
        RECT 54.810 137.525 55.105 138.635 ;
        RECT 55.285 137.545 56.495 138.635 ;
        RECT 51.610 137.075 54.630 137.325 ;
        RECT 49.745 136.085 50.045 136.815 ;
        RECT 50.470 136.735 53.780 136.905 ;
        RECT 50.470 136.085 50.770 136.565 ;
        RECT 50.940 136.280 51.200 136.735 ;
        RECT 51.370 136.085 51.630 136.565 ;
        RECT 51.800 136.280 52.060 136.735 ;
        RECT 52.230 136.085 52.490 136.565 ;
        RECT 52.660 136.280 52.920 136.735 ;
        RECT 53.090 136.085 53.350 136.565 ;
        RECT 53.520 136.280 53.780 136.735 ;
        RECT 53.950 136.085 54.210 136.610 ;
        RECT 54.380 136.265 54.630 137.075 ;
        RECT 54.800 136.715 55.115 137.325 ;
        RECT 55.285 136.835 55.805 137.375 ;
        RECT 55.975 137.005 56.495 137.545 ;
        RECT 56.665 138.205 57.005 138.465 ;
        RECT 54.810 136.085 55.055 136.545 ;
        RECT 55.285 136.085 56.495 136.835 ;
        RECT 56.665 136.805 56.925 138.205 ;
        RECT 57.175 137.835 57.505 138.635 ;
        RECT 57.970 137.665 58.220 138.465 ;
        RECT 58.405 137.915 58.735 138.635 ;
        RECT 58.955 137.665 59.205 138.465 ;
        RECT 59.375 138.255 59.710 138.635 ;
        RECT 59.885 138.200 65.230 138.635 ;
        RECT 57.115 137.495 59.305 137.665 ;
        RECT 57.115 137.325 57.430 137.495 ;
        RECT 57.100 137.075 57.430 137.325 ;
        RECT 56.665 136.295 57.005 136.805 ;
        RECT 57.175 136.085 57.445 136.885 ;
        RECT 57.625 136.355 57.905 137.325 ;
        RECT 58.085 136.355 58.385 137.325 ;
        RECT 58.565 136.360 58.915 137.325 ;
        RECT 59.135 136.585 59.305 137.495 ;
        RECT 59.475 136.765 59.715 138.075 ;
        RECT 61.470 136.630 61.810 137.460 ;
        RECT 63.290 136.950 63.640 138.200 ;
        RECT 65.405 137.545 68.915 138.635 ;
        RECT 65.405 136.855 67.055 137.375 ;
        RECT 67.225 137.025 68.915 137.545 ;
        RECT 70.005 137.470 70.295 138.635 ;
        RECT 70.465 138.200 75.810 138.635 ;
        RECT 75.985 138.200 81.330 138.635 ;
        RECT 59.135 136.255 59.630 136.585 ;
        RECT 59.885 136.085 65.230 136.630 ;
        RECT 65.405 136.085 68.915 136.855 ;
        RECT 70.005 136.085 70.295 136.810 ;
        RECT 72.050 136.630 72.390 137.460 ;
        RECT 73.870 136.950 74.220 138.200 ;
        RECT 77.570 136.630 77.910 137.460 ;
        RECT 79.390 136.950 79.740 138.200 ;
        RECT 81.505 137.545 82.715 138.635 ;
        RECT 81.505 136.835 82.025 137.375 ;
        RECT 82.195 137.005 82.715 137.545 ;
        RECT 82.885 137.545 84.095 138.635 ;
        RECT 82.885 137.005 83.405 137.545 ;
        RECT 83.575 136.835 84.095 137.375 ;
        RECT 70.465 136.085 75.810 136.630 ;
        RECT 75.985 136.085 81.330 136.630 ;
        RECT 81.505 136.085 82.715 136.835 ;
        RECT 82.885 136.085 84.095 136.835 ;
        RECT 5.520 135.915 84.180 136.085 ;
        RECT 5.605 135.165 6.815 135.915 ;
        RECT 5.605 134.625 6.125 135.165 ;
        RECT 6.990 135.075 7.250 135.915 ;
        RECT 7.425 135.170 7.680 135.745 ;
        RECT 7.850 135.535 8.180 135.915 ;
        RECT 8.395 135.365 8.565 135.745 ;
        RECT 7.850 135.195 8.565 135.365 ;
        RECT 6.295 134.455 6.815 134.995 ;
        RECT 5.605 133.365 6.815 134.455 ;
        RECT 6.990 133.365 7.250 134.515 ;
        RECT 7.425 134.440 7.595 135.170 ;
        RECT 7.850 135.005 8.020 135.195 ;
        RECT 8.825 135.145 12.335 135.915 ;
        RECT 13.425 135.265 13.685 135.745 ;
        RECT 13.855 135.455 14.185 135.915 ;
        RECT 14.375 135.275 14.575 135.695 ;
        RECT 7.765 134.675 8.020 135.005 ;
        RECT 7.850 134.465 8.020 134.675 ;
        RECT 8.300 134.645 8.655 135.015 ;
        RECT 8.825 134.625 10.475 135.145 ;
        RECT 7.425 133.535 7.680 134.440 ;
        RECT 7.850 134.295 8.565 134.465 ;
        RECT 10.645 134.455 12.335 134.975 ;
        RECT 7.850 133.365 8.180 134.125 ;
        RECT 8.395 133.535 8.565 134.295 ;
        RECT 8.825 133.365 12.335 134.455 ;
        RECT 13.425 134.235 13.595 135.265 ;
        RECT 13.765 134.575 13.995 135.005 ;
        RECT 14.165 134.755 14.575 135.275 ;
        RECT 14.745 135.430 15.535 135.695 ;
        RECT 14.745 134.575 15.000 135.430 ;
        RECT 15.715 135.095 16.045 135.515 ;
        RECT 16.215 135.095 16.475 135.915 ;
        RECT 16.645 135.165 17.855 135.915 ;
        RECT 18.190 135.405 18.430 135.915 ;
        RECT 18.610 135.405 18.890 135.735 ;
        RECT 19.120 135.405 19.335 135.915 ;
        RECT 15.715 135.005 15.965 135.095 ;
        RECT 15.170 134.755 15.965 135.005 ;
        RECT 13.765 134.405 15.555 134.575 ;
        RECT 13.425 133.535 13.700 134.235 ;
        RECT 13.870 134.110 14.585 134.405 ;
        RECT 14.805 134.045 15.135 134.235 ;
        RECT 13.910 133.365 14.125 133.910 ;
        RECT 14.295 133.535 14.770 133.875 ;
        RECT 14.940 133.870 15.135 134.045 ;
        RECT 15.305 134.040 15.555 134.405 ;
        RECT 14.940 133.365 15.555 133.870 ;
        RECT 15.795 133.535 15.965 134.755 ;
        RECT 16.135 134.045 16.475 134.925 ;
        RECT 16.645 134.625 17.165 135.165 ;
        RECT 17.335 134.455 17.855 134.995 ;
        RECT 18.085 134.675 18.440 135.235 ;
        RECT 18.610 134.505 18.780 135.405 ;
        RECT 18.950 134.675 19.215 135.235 ;
        RECT 19.505 135.175 20.120 135.745 ;
        RECT 20.325 135.535 21.215 135.705 ;
        RECT 19.465 134.505 19.635 135.005 ;
        RECT 16.215 133.365 16.475 133.875 ;
        RECT 16.645 133.365 17.855 134.455 ;
        RECT 18.210 134.335 19.635 134.505 ;
        RECT 18.210 134.160 18.600 134.335 ;
        RECT 19.085 133.365 19.415 134.165 ;
        RECT 19.805 134.155 20.120 135.175 ;
        RECT 20.325 134.980 20.875 135.365 ;
        RECT 21.045 134.810 21.215 135.535 ;
        RECT 20.325 134.740 21.215 134.810 ;
        RECT 21.385 135.210 21.605 135.695 ;
        RECT 21.775 135.375 22.025 135.915 ;
        RECT 22.195 135.265 22.455 135.745 ;
        RECT 21.385 134.785 21.715 135.210 ;
        RECT 20.325 134.715 21.220 134.740 ;
        RECT 20.325 134.700 21.230 134.715 ;
        RECT 20.325 134.685 21.235 134.700 ;
        RECT 20.325 134.680 21.245 134.685 ;
        RECT 20.325 134.670 21.250 134.680 ;
        RECT 20.325 134.660 21.255 134.670 ;
        RECT 20.325 134.655 21.265 134.660 ;
        RECT 20.325 134.645 21.275 134.655 ;
        RECT 20.325 134.640 21.285 134.645 ;
        RECT 20.325 134.190 20.585 134.640 ;
        RECT 20.950 134.635 21.285 134.640 ;
        RECT 20.950 134.630 21.300 134.635 ;
        RECT 20.950 134.620 21.315 134.630 ;
        RECT 20.950 134.615 21.340 134.620 ;
        RECT 21.885 134.615 22.115 135.010 ;
        RECT 20.950 134.610 22.115 134.615 ;
        RECT 20.980 134.575 22.115 134.610 ;
        RECT 21.015 134.550 22.115 134.575 ;
        RECT 21.045 134.520 22.115 134.550 ;
        RECT 21.065 134.490 22.115 134.520 ;
        RECT 21.085 134.460 22.115 134.490 ;
        RECT 21.155 134.450 22.115 134.460 ;
        RECT 21.180 134.440 22.115 134.450 ;
        RECT 21.200 134.425 22.115 134.440 ;
        RECT 21.220 134.410 22.115 134.425 ;
        RECT 21.225 134.400 22.010 134.410 ;
        RECT 21.240 134.365 22.010 134.400 ;
        RECT 19.585 133.535 20.120 134.155 ;
        RECT 20.755 134.045 21.085 134.290 ;
        RECT 21.255 134.115 22.010 134.365 ;
        RECT 22.285 134.235 22.455 135.265 ;
        RECT 22.715 135.365 22.885 135.655 ;
        RECT 23.055 135.535 23.385 135.915 ;
        RECT 22.715 135.195 23.380 135.365 ;
        RECT 22.630 134.375 22.980 135.025 ;
        RECT 20.755 134.020 20.940 134.045 ;
        RECT 20.325 133.920 20.940 134.020 ;
        RECT 20.325 133.365 20.930 133.920 ;
        RECT 21.105 133.535 21.585 133.875 ;
        RECT 21.755 133.365 22.010 133.910 ;
        RECT 22.180 133.535 22.455 134.235 ;
        RECT 23.150 134.205 23.380 135.195 ;
        RECT 22.715 134.035 23.380 134.205 ;
        RECT 22.715 133.535 22.885 134.035 ;
        RECT 23.055 133.365 23.385 133.865 ;
        RECT 23.555 133.535 23.740 135.655 ;
        RECT 23.995 135.455 24.245 135.915 ;
        RECT 24.415 135.465 24.750 135.635 ;
        RECT 24.945 135.465 25.620 135.635 ;
        RECT 24.415 135.325 24.585 135.465 ;
        RECT 23.910 134.335 24.190 135.285 ;
        RECT 24.360 135.195 24.585 135.325 ;
        RECT 24.360 134.090 24.530 135.195 ;
        RECT 24.755 135.045 25.280 135.265 ;
        RECT 24.700 134.280 24.940 134.875 ;
        RECT 25.110 134.345 25.280 135.045 ;
        RECT 25.450 134.685 25.620 135.465 ;
        RECT 25.940 135.415 26.310 135.915 ;
        RECT 26.490 135.465 26.895 135.635 ;
        RECT 27.065 135.465 27.850 135.635 ;
        RECT 26.490 135.235 26.660 135.465 ;
        RECT 25.830 134.935 26.660 135.235 ;
        RECT 27.045 134.965 27.510 135.295 ;
        RECT 25.830 134.905 26.030 134.935 ;
        RECT 26.150 134.685 26.320 134.755 ;
        RECT 25.450 134.515 26.320 134.685 ;
        RECT 25.810 134.425 26.320 134.515 ;
        RECT 24.360 133.960 24.665 134.090 ;
        RECT 25.110 133.980 25.640 134.345 ;
        RECT 23.980 133.365 24.245 133.825 ;
        RECT 24.415 133.535 24.665 133.960 ;
        RECT 25.810 133.810 25.980 134.425 ;
        RECT 24.875 133.640 25.980 133.810 ;
        RECT 26.150 133.365 26.320 134.165 ;
        RECT 26.490 133.865 26.660 134.935 ;
        RECT 26.830 134.035 27.020 134.755 ;
        RECT 27.190 134.005 27.510 134.965 ;
        RECT 27.680 135.005 27.850 135.465 ;
        RECT 28.125 135.385 28.335 135.915 ;
        RECT 28.595 135.175 28.925 135.700 ;
        RECT 29.095 135.305 29.265 135.915 ;
        RECT 29.435 135.260 29.765 135.695 ;
        RECT 29.435 135.175 29.815 135.260 ;
        RECT 28.725 135.005 28.925 135.175 ;
        RECT 29.590 135.135 29.815 135.175 ;
        RECT 27.680 134.675 28.555 135.005 ;
        RECT 28.725 134.675 29.475 135.005 ;
        RECT 26.490 133.535 26.740 133.865 ;
        RECT 27.680 133.835 27.850 134.675 ;
        RECT 28.725 134.470 28.915 134.675 ;
        RECT 29.645 134.555 29.815 135.135 ;
        RECT 29.985 135.165 31.195 135.915 ;
        RECT 31.365 135.190 31.655 135.915 ;
        RECT 32.805 135.455 33.050 135.915 ;
        RECT 29.985 134.625 30.505 135.165 ;
        RECT 29.600 134.505 29.815 134.555 ;
        RECT 28.020 134.095 28.915 134.470 ;
        RECT 29.425 134.425 29.815 134.505 ;
        RECT 30.675 134.455 31.195 134.995 ;
        RECT 32.745 134.675 33.060 135.285 ;
        RECT 33.230 134.925 33.480 135.735 ;
        RECT 33.650 135.390 33.910 135.915 ;
        RECT 34.080 135.265 34.340 135.720 ;
        RECT 34.510 135.435 34.770 135.915 ;
        RECT 34.940 135.265 35.200 135.720 ;
        RECT 35.370 135.435 35.630 135.915 ;
        RECT 35.800 135.265 36.060 135.720 ;
        RECT 36.230 135.435 36.490 135.915 ;
        RECT 36.660 135.265 36.920 135.720 ;
        RECT 37.090 135.435 37.390 135.915 ;
        RECT 37.810 135.660 38.145 135.705 ;
        RECT 34.080 135.095 37.390 135.265 ;
        RECT 33.230 134.675 36.250 134.925 ;
        RECT 26.965 133.665 27.850 133.835 ;
        RECT 28.030 133.365 28.345 133.865 ;
        RECT 28.575 133.535 28.915 134.095 ;
        RECT 29.085 133.365 29.255 134.375 ;
        RECT 29.425 133.580 29.755 134.425 ;
        RECT 29.985 133.365 31.195 134.455 ;
        RECT 31.365 133.365 31.655 134.530 ;
        RECT 32.755 133.365 33.050 134.475 ;
        RECT 33.230 133.540 33.480 134.675 ;
        RECT 36.420 134.505 37.390 135.095 ;
        RECT 33.650 133.365 33.910 134.475 ;
        RECT 34.080 134.265 37.390 134.505 ;
        RECT 37.805 135.195 38.145 135.660 ;
        RECT 38.315 135.535 38.645 135.915 ;
        RECT 39.105 135.575 39.375 135.580 ;
        RECT 39.105 135.405 39.415 135.575 ;
        RECT 37.805 134.505 37.975 135.195 ;
        RECT 38.145 134.675 38.405 135.005 ;
        RECT 34.080 133.540 34.340 134.265 ;
        RECT 34.510 133.365 34.770 134.095 ;
        RECT 34.940 133.540 35.200 134.265 ;
        RECT 35.370 133.365 35.630 134.095 ;
        RECT 35.800 133.540 36.060 134.265 ;
        RECT 36.230 133.365 36.490 134.095 ;
        RECT 36.660 133.540 36.920 134.265 ;
        RECT 37.090 133.365 37.385 134.095 ;
        RECT 37.805 133.535 38.065 134.505 ;
        RECT 38.235 134.125 38.405 134.675 ;
        RECT 38.575 134.305 38.915 135.335 ;
        RECT 39.105 134.305 39.375 135.405 ;
        RECT 39.600 134.305 39.880 135.580 ;
        RECT 40.080 135.415 40.310 135.745 ;
        RECT 40.555 135.535 40.885 135.915 ;
        RECT 40.080 134.125 40.250 135.415 ;
        RECT 41.055 135.345 41.230 135.745 ;
        RECT 40.600 135.175 41.230 135.345 ;
        RECT 41.485 135.195 41.825 135.705 ;
        RECT 40.600 135.005 40.770 135.175 ;
        RECT 40.420 134.675 40.770 135.005 ;
        RECT 38.235 133.955 40.250 134.125 ;
        RECT 40.600 134.155 40.770 134.675 ;
        RECT 40.950 134.325 41.315 135.005 ;
        RECT 40.600 133.985 41.230 134.155 ;
        RECT 38.260 133.365 38.590 133.775 ;
        RECT 38.790 133.535 38.960 133.955 ;
        RECT 39.175 133.365 39.845 133.775 ;
        RECT 40.080 133.535 40.250 133.955 ;
        RECT 40.555 133.365 40.885 133.805 ;
        RECT 41.055 133.535 41.230 133.985 ;
        RECT 41.485 133.795 41.745 135.195 ;
        RECT 41.995 135.115 42.265 135.915 ;
        RECT 41.920 134.675 42.250 134.925 ;
        RECT 42.445 134.675 42.725 135.645 ;
        RECT 42.905 134.675 43.205 135.645 ;
        RECT 43.385 134.675 43.735 135.640 ;
        RECT 43.955 135.415 44.450 135.745 ;
        RECT 41.935 134.505 42.250 134.675 ;
        RECT 43.955 134.505 44.125 135.415 ;
        RECT 41.935 134.335 44.125 134.505 ;
        RECT 41.485 133.535 41.825 133.795 ;
        RECT 41.995 133.365 42.325 134.165 ;
        RECT 42.790 133.535 43.040 134.335 ;
        RECT 43.225 133.365 43.555 134.085 ;
        RECT 43.775 133.535 44.025 134.335 ;
        RECT 44.295 133.925 44.535 135.235 ;
        RECT 44.715 135.105 44.985 135.915 ;
        RECT 45.155 135.105 45.485 135.745 ;
        RECT 45.655 135.105 45.895 135.915 ;
        RECT 46.085 135.145 49.595 135.915 ;
        RECT 50.270 135.455 50.535 135.915 ;
        RECT 50.905 135.275 51.075 135.745 ;
        RECT 51.325 135.455 51.495 135.915 ;
        RECT 51.745 135.275 51.915 135.745 ;
        RECT 52.165 135.455 52.335 135.915 ;
        RECT 52.585 135.275 52.755 135.745 ;
        RECT 52.925 135.450 53.175 135.915 ;
        RECT 44.705 134.675 45.055 134.925 ;
        RECT 45.225 134.505 45.395 135.105 ;
        RECT 45.565 134.675 45.915 134.925 ;
        RECT 46.085 134.625 47.735 135.145 ;
        RECT 50.905 135.095 53.275 135.275 ;
        RECT 44.195 133.365 44.530 133.745 ;
        RECT 44.715 133.365 45.045 134.505 ;
        RECT 45.225 134.335 45.905 134.505 ;
        RECT 47.905 134.455 49.595 134.975 ;
        RECT 50.245 134.675 52.755 134.925 ;
        RECT 52.925 134.505 53.275 135.095 ;
        RECT 53.445 135.145 56.955 135.915 ;
        RECT 57.125 135.190 57.415 135.915 ;
        RECT 57.585 135.145 59.255 135.915 ;
        RECT 53.445 134.625 55.095 135.145 ;
        RECT 45.575 133.550 45.905 134.335 ;
        RECT 46.085 133.365 49.595 134.455 ;
        RECT 50.270 133.365 50.565 134.505 ;
        RECT 50.825 134.335 53.275 134.505 ;
        RECT 55.265 134.455 56.955 134.975 ;
        RECT 57.585 134.625 58.335 135.145 ;
        RECT 59.435 135.105 59.705 135.915 ;
        RECT 59.875 135.105 60.205 135.745 ;
        RECT 60.375 135.105 60.615 135.915 ;
        RECT 60.805 135.165 62.015 135.915 ;
        RECT 62.270 135.345 62.445 135.745 ;
        RECT 62.615 135.535 62.945 135.915 ;
        RECT 63.190 135.415 63.420 135.745 ;
        RECT 62.270 135.175 62.900 135.345 ;
        RECT 50.825 133.535 51.155 134.335 ;
        RECT 51.325 133.365 51.495 134.165 ;
        RECT 51.665 133.535 51.995 134.335 ;
        RECT 52.505 134.315 53.275 134.335 ;
        RECT 52.165 133.365 52.335 134.165 ;
        RECT 52.505 133.535 52.835 134.315 ;
        RECT 53.005 133.365 53.175 133.825 ;
        RECT 53.445 133.365 56.955 134.455 ;
        RECT 57.125 133.365 57.415 134.530 ;
        RECT 58.505 134.455 59.255 134.975 ;
        RECT 59.425 134.675 59.775 134.925 ;
        RECT 59.945 134.505 60.115 135.105 ;
        RECT 60.285 134.675 60.635 134.925 ;
        RECT 60.805 134.625 61.325 135.165 ;
        RECT 62.730 135.005 62.900 135.175 ;
        RECT 57.585 133.365 59.255 134.455 ;
        RECT 59.435 133.365 59.765 134.505 ;
        RECT 59.945 134.335 60.625 134.505 ;
        RECT 61.495 134.455 62.015 134.995 ;
        RECT 60.295 133.550 60.625 134.335 ;
        RECT 60.805 133.365 62.015 134.455 ;
        RECT 62.185 134.325 62.550 135.005 ;
        RECT 62.730 134.675 63.080 135.005 ;
        RECT 62.730 134.155 62.900 134.675 ;
        RECT 62.270 133.985 62.900 134.155 ;
        RECT 63.250 134.125 63.420 135.415 ;
        RECT 63.620 134.305 63.900 135.580 ;
        RECT 64.125 135.575 64.395 135.580 ;
        RECT 64.085 135.405 64.395 135.575 ;
        RECT 64.855 135.535 65.185 135.915 ;
        RECT 65.355 135.660 65.690 135.705 ;
        RECT 64.125 134.305 64.395 135.405 ;
        RECT 64.585 134.305 64.925 135.335 ;
        RECT 65.355 135.195 65.695 135.660 ;
        RECT 65.915 135.260 66.245 135.695 ;
        RECT 66.415 135.305 66.585 135.915 ;
        RECT 65.095 134.675 65.355 135.005 ;
        RECT 65.095 134.125 65.265 134.675 ;
        RECT 65.525 134.505 65.695 135.195 ;
        RECT 62.270 133.535 62.445 133.985 ;
        RECT 63.250 133.955 65.265 134.125 ;
        RECT 62.615 133.365 62.945 133.805 ;
        RECT 63.250 133.535 63.420 133.955 ;
        RECT 63.655 133.365 64.325 133.775 ;
        RECT 64.540 133.535 64.710 133.955 ;
        RECT 64.910 133.365 65.240 133.775 ;
        RECT 65.435 133.535 65.695 134.505 ;
        RECT 65.865 135.175 66.245 135.260 ;
        RECT 66.755 135.175 67.085 135.700 ;
        RECT 67.345 135.385 67.555 135.915 ;
        RECT 67.830 135.465 68.615 135.635 ;
        RECT 68.785 135.465 69.190 135.635 ;
        RECT 65.865 135.135 66.090 135.175 ;
        RECT 65.865 134.555 66.035 135.135 ;
        RECT 66.755 135.005 66.955 135.175 ;
        RECT 67.830 135.005 68.000 135.465 ;
        RECT 66.205 134.675 66.955 135.005 ;
        RECT 67.125 134.675 68.000 135.005 ;
        RECT 65.865 134.505 66.080 134.555 ;
        RECT 65.865 134.425 66.255 134.505 ;
        RECT 65.925 133.580 66.255 134.425 ;
        RECT 66.765 134.470 66.955 134.675 ;
        RECT 66.425 133.365 66.595 134.375 ;
        RECT 66.765 134.095 67.660 134.470 ;
        RECT 66.765 133.535 67.105 134.095 ;
        RECT 67.335 133.365 67.650 133.865 ;
        RECT 67.830 133.835 68.000 134.675 ;
        RECT 68.170 134.965 68.635 135.295 ;
        RECT 69.020 135.235 69.190 135.465 ;
        RECT 69.370 135.415 69.740 135.915 ;
        RECT 70.060 135.465 70.735 135.635 ;
        RECT 70.930 135.465 71.265 135.635 ;
        RECT 68.170 134.005 68.490 134.965 ;
        RECT 69.020 134.935 69.850 135.235 ;
        RECT 68.660 134.035 68.850 134.755 ;
        RECT 69.020 133.865 69.190 134.935 ;
        RECT 69.650 134.905 69.850 134.935 ;
        RECT 69.360 134.685 69.530 134.755 ;
        RECT 70.060 134.685 70.230 135.465 ;
        RECT 71.095 135.325 71.265 135.465 ;
        RECT 71.435 135.455 71.685 135.915 ;
        RECT 69.360 134.515 70.230 134.685 ;
        RECT 70.400 135.045 70.925 135.265 ;
        RECT 71.095 135.195 71.320 135.325 ;
        RECT 69.360 134.425 69.870 134.515 ;
        RECT 67.830 133.665 68.715 133.835 ;
        RECT 68.940 133.535 69.190 133.865 ;
        RECT 69.360 133.365 69.530 134.165 ;
        RECT 69.700 133.810 69.870 134.425 ;
        RECT 70.400 134.345 70.570 135.045 ;
        RECT 70.040 133.980 70.570 134.345 ;
        RECT 70.740 134.280 70.980 134.875 ;
        RECT 71.150 134.090 71.320 135.195 ;
        RECT 71.490 134.335 71.770 135.285 ;
        RECT 71.015 133.960 71.320 134.090 ;
        RECT 69.700 133.640 70.805 133.810 ;
        RECT 71.015 133.535 71.265 133.960 ;
        RECT 71.435 133.365 71.700 133.825 ;
        RECT 71.940 133.535 72.125 135.655 ;
        RECT 72.295 135.535 72.625 135.915 ;
        RECT 72.795 135.365 72.965 135.655 ;
        RECT 73.225 135.370 78.570 135.915 ;
        RECT 72.300 135.195 72.965 135.365 ;
        RECT 72.300 134.205 72.530 135.195 ;
        RECT 72.700 134.375 73.050 135.025 ;
        RECT 74.810 134.540 75.150 135.370 ;
        RECT 78.745 135.145 82.255 135.915 ;
        RECT 82.885 135.165 84.095 135.915 ;
        RECT 72.300 134.035 72.965 134.205 ;
        RECT 72.295 133.365 72.625 133.865 ;
        RECT 72.795 133.535 72.965 134.035 ;
        RECT 76.630 133.800 76.980 135.050 ;
        RECT 78.745 134.625 80.395 135.145 ;
        RECT 80.565 134.455 82.255 134.975 ;
        RECT 73.225 133.365 78.570 133.800 ;
        RECT 78.745 133.365 82.255 134.455 ;
        RECT 82.885 134.455 83.405 134.995 ;
        RECT 83.575 134.625 84.095 135.165 ;
        RECT 82.885 133.365 84.095 134.455 ;
        RECT 5.520 133.195 84.180 133.365 ;
        RECT 5.605 132.105 6.815 133.195 ;
        RECT 6.985 132.760 12.330 133.195 ;
        RECT 12.505 132.760 17.850 133.195 ;
        RECT 5.605 131.395 6.125 131.935 ;
        RECT 6.295 131.565 6.815 132.105 ;
        RECT 5.605 130.645 6.815 131.395 ;
        RECT 8.570 131.190 8.910 132.020 ;
        RECT 10.390 131.510 10.740 132.760 ;
        RECT 14.090 131.190 14.430 132.020 ;
        RECT 15.910 131.510 16.260 132.760 ;
        RECT 18.485 132.030 18.775 133.195 ;
        RECT 18.945 132.105 22.455 133.195 ;
        RECT 18.945 131.415 20.595 131.935 ;
        RECT 20.765 131.585 22.455 132.105 ;
        RECT 23.555 132.055 23.885 133.195 ;
        RECT 6.985 130.645 12.330 131.190 ;
        RECT 12.505 130.645 17.850 131.190 ;
        RECT 18.485 130.645 18.775 131.370 ;
        RECT 18.945 130.645 22.455 131.415 ;
        RECT 23.545 131.305 23.885 131.885 ;
        RECT 24.055 131.855 24.415 133.025 ;
        RECT 24.615 132.025 24.945 133.195 ;
        RECT 25.145 131.855 25.475 133.025 ;
        RECT 25.675 132.025 26.005 133.195 ;
        RECT 26.315 132.245 26.590 133.015 ;
        RECT 26.760 132.585 27.090 133.015 ;
        RECT 27.260 132.755 27.455 133.195 ;
        RECT 27.635 132.585 27.965 133.015 ;
        RECT 26.760 132.415 27.965 132.585 ;
        RECT 26.315 132.055 26.900 132.245 ;
        RECT 27.070 132.085 27.965 132.415 ;
        RECT 28.145 132.105 29.815 133.195 ;
        RECT 30.535 132.525 30.705 133.025 ;
        RECT 30.875 132.695 31.205 133.195 ;
        RECT 30.535 132.355 31.200 132.525 ;
        RECT 24.055 131.575 25.475 131.855 ;
        RECT 24.055 131.240 24.415 131.575 ;
        RECT 23.555 130.645 23.885 131.135 ;
        RECT 24.055 130.815 24.675 131.240 ;
        RECT 25.135 130.645 25.465 131.335 ;
        RECT 26.315 131.235 26.555 131.885 ;
        RECT 26.725 131.385 26.900 132.055 ;
        RECT 27.070 131.555 27.485 131.885 ;
        RECT 27.665 131.555 27.960 131.885 ;
        RECT 26.725 131.205 27.055 131.385 ;
        RECT 26.330 130.645 26.660 131.035 ;
        RECT 26.830 130.825 27.055 131.205 ;
        RECT 27.255 130.935 27.485 131.555 ;
        RECT 28.145 131.415 28.895 131.935 ;
        RECT 29.065 131.585 29.815 132.105 ;
        RECT 30.450 131.535 30.800 132.185 ;
        RECT 27.665 130.645 27.965 131.375 ;
        RECT 28.145 130.645 29.815 131.415 ;
        RECT 30.970 131.365 31.200 132.355 ;
        RECT 30.535 131.195 31.200 131.365 ;
        RECT 30.535 130.905 30.705 131.195 ;
        RECT 30.875 130.645 31.205 131.025 ;
        RECT 31.375 130.905 31.560 133.025 ;
        RECT 31.800 132.735 32.065 133.195 ;
        RECT 32.235 132.600 32.485 133.025 ;
        RECT 32.695 132.750 33.800 132.920 ;
        RECT 32.180 132.470 32.485 132.600 ;
        RECT 31.730 131.275 32.010 132.225 ;
        RECT 32.180 131.365 32.350 132.470 ;
        RECT 32.520 131.685 32.760 132.280 ;
        RECT 32.930 132.215 33.460 132.580 ;
        RECT 32.930 131.515 33.100 132.215 ;
        RECT 33.630 132.135 33.800 132.750 ;
        RECT 33.970 132.395 34.140 133.195 ;
        RECT 34.310 132.695 34.560 133.025 ;
        RECT 34.785 132.725 35.670 132.895 ;
        RECT 33.630 132.045 34.140 132.135 ;
        RECT 32.180 131.235 32.405 131.365 ;
        RECT 32.575 131.295 33.100 131.515 ;
        RECT 33.270 131.875 34.140 132.045 ;
        RECT 31.815 130.645 32.065 131.105 ;
        RECT 32.235 131.095 32.405 131.235 ;
        RECT 33.270 131.095 33.440 131.875 ;
        RECT 33.970 131.805 34.140 131.875 ;
        RECT 33.650 131.625 33.850 131.655 ;
        RECT 34.310 131.625 34.480 132.695 ;
        RECT 34.650 131.805 34.840 132.525 ;
        RECT 33.650 131.325 34.480 131.625 ;
        RECT 35.010 131.595 35.330 132.555 ;
        RECT 32.235 130.925 32.570 131.095 ;
        RECT 32.765 130.925 33.440 131.095 ;
        RECT 33.760 130.645 34.130 131.145 ;
        RECT 34.310 131.095 34.480 131.325 ;
        RECT 34.865 131.265 35.330 131.595 ;
        RECT 35.500 131.885 35.670 132.725 ;
        RECT 35.850 132.695 36.165 133.195 ;
        RECT 36.395 132.465 36.735 133.025 ;
        RECT 35.840 132.090 36.735 132.465 ;
        RECT 36.905 132.185 37.075 133.195 ;
        RECT 36.545 131.885 36.735 132.090 ;
        RECT 37.245 132.135 37.575 132.980 ;
        RECT 37.805 132.760 43.150 133.195 ;
        RECT 37.245 132.055 37.635 132.135 ;
        RECT 37.420 132.005 37.635 132.055 ;
        RECT 35.500 131.555 36.375 131.885 ;
        RECT 36.545 131.555 37.295 131.885 ;
        RECT 35.500 131.095 35.670 131.555 ;
        RECT 36.545 131.385 36.745 131.555 ;
        RECT 37.465 131.425 37.635 132.005 ;
        RECT 37.410 131.385 37.635 131.425 ;
        RECT 34.310 130.925 34.715 131.095 ;
        RECT 34.885 130.925 35.670 131.095 ;
        RECT 35.945 130.645 36.155 131.175 ;
        RECT 36.415 130.860 36.745 131.385 ;
        RECT 37.255 131.300 37.635 131.385 ;
        RECT 36.915 130.645 37.085 131.255 ;
        RECT 37.255 130.865 37.585 131.300 ;
        RECT 39.390 131.190 39.730 132.020 ;
        RECT 41.210 131.510 41.560 132.760 ;
        RECT 44.245 132.030 44.535 133.195 ;
        RECT 44.710 132.770 45.045 133.195 ;
        RECT 45.215 132.590 45.400 132.995 ;
        RECT 44.735 132.415 45.400 132.590 ;
        RECT 45.605 132.415 45.935 133.195 ;
        RECT 44.735 131.385 45.075 132.415 ;
        RECT 46.105 132.225 46.375 132.995 ;
        RECT 45.245 132.055 46.375 132.225 ;
        RECT 46.545 132.105 50.055 133.195 ;
        RECT 50.310 132.575 50.485 133.025 ;
        RECT 50.655 132.755 50.985 133.195 ;
        RECT 51.290 132.605 51.460 133.025 ;
        RECT 51.695 132.785 52.365 133.195 ;
        RECT 52.580 132.605 52.750 133.025 ;
        RECT 52.950 132.785 53.280 133.195 ;
        RECT 50.310 132.405 50.940 132.575 ;
        RECT 45.245 131.555 45.495 132.055 ;
        RECT 37.805 130.645 43.150 131.190 ;
        RECT 44.245 130.645 44.535 131.370 ;
        RECT 44.735 131.215 45.420 131.385 ;
        RECT 45.675 131.305 46.035 131.885 ;
        RECT 44.710 130.645 45.045 131.045 ;
        RECT 45.215 130.815 45.420 131.215 ;
        RECT 46.205 131.145 46.375 132.055 ;
        RECT 45.630 130.645 45.905 131.125 ;
        RECT 46.115 130.815 46.375 131.145 ;
        RECT 46.545 131.415 48.195 131.935 ;
        RECT 48.365 131.585 50.055 132.105 ;
        RECT 50.225 131.555 50.590 132.235 ;
        RECT 50.770 131.885 50.940 132.405 ;
        RECT 51.290 132.435 53.305 132.605 ;
        RECT 50.770 131.555 51.120 131.885 ;
        RECT 46.545 130.645 50.055 131.415 ;
        RECT 50.770 131.385 50.940 131.555 ;
        RECT 50.310 131.215 50.940 131.385 ;
        RECT 50.310 130.815 50.485 131.215 ;
        RECT 51.290 131.145 51.460 132.435 ;
        RECT 50.655 130.645 50.985 131.025 ;
        RECT 51.230 130.815 51.460 131.145 ;
        RECT 51.660 130.980 51.940 132.255 ;
        RECT 52.165 132.175 52.435 132.255 ;
        RECT 52.125 132.005 52.435 132.175 ;
        RECT 52.165 130.980 52.435 132.005 ;
        RECT 52.625 131.225 52.965 132.255 ;
        RECT 53.135 131.885 53.305 132.435 ;
        RECT 53.475 132.055 53.735 133.025 ;
        RECT 53.915 132.055 54.245 133.195 ;
        RECT 54.775 132.225 55.105 133.010 ;
        RECT 54.425 132.055 55.105 132.225 ;
        RECT 55.755 132.055 56.085 133.195 ;
        RECT 56.615 132.225 56.945 133.010 ;
        RECT 56.265 132.055 56.945 132.225 ;
        RECT 58.045 132.325 58.320 133.025 ;
        RECT 58.490 132.650 58.745 133.195 ;
        RECT 58.915 132.685 59.395 133.025 ;
        RECT 59.570 132.640 60.175 133.195 ;
        RECT 59.560 132.540 60.175 132.640 ;
        RECT 59.560 132.515 59.745 132.540 ;
        RECT 53.135 131.555 53.395 131.885 ;
        RECT 53.565 131.365 53.735 132.055 ;
        RECT 53.905 131.635 54.255 131.885 ;
        RECT 54.425 131.455 54.595 132.055 ;
        RECT 54.765 131.635 55.115 131.885 ;
        RECT 55.745 131.635 56.095 131.885 ;
        RECT 56.265 131.455 56.435 132.055 ;
        RECT 56.605 131.635 56.955 131.885 ;
        RECT 52.895 130.645 53.225 131.025 ;
        RECT 53.395 130.900 53.735 131.365 ;
        RECT 53.395 130.855 53.730 130.900 ;
        RECT 53.915 130.645 54.185 131.455 ;
        RECT 54.355 130.815 54.685 131.455 ;
        RECT 54.855 130.645 55.095 131.455 ;
        RECT 55.755 130.645 56.025 131.455 ;
        RECT 56.195 130.815 56.525 131.455 ;
        RECT 56.695 130.645 56.935 131.455 ;
        RECT 58.045 131.295 58.215 132.325 ;
        RECT 58.490 132.195 59.245 132.445 ;
        RECT 59.415 132.270 59.745 132.515 ;
        RECT 58.490 132.160 59.260 132.195 ;
        RECT 58.490 132.150 59.275 132.160 ;
        RECT 58.385 132.135 59.280 132.150 ;
        RECT 58.385 132.120 59.300 132.135 ;
        RECT 58.385 132.110 59.320 132.120 ;
        RECT 58.385 132.100 59.345 132.110 ;
        RECT 58.385 132.070 59.415 132.100 ;
        RECT 58.385 132.040 59.435 132.070 ;
        RECT 58.385 132.010 59.455 132.040 ;
        RECT 58.385 131.985 59.485 132.010 ;
        RECT 58.385 131.950 59.520 131.985 ;
        RECT 58.385 131.945 59.550 131.950 ;
        RECT 58.385 131.550 58.615 131.945 ;
        RECT 59.160 131.940 59.550 131.945 ;
        RECT 59.185 131.930 59.550 131.940 ;
        RECT 59.200 131.925 59.550 131.930 ;
        RECT 59.215 131.920 59.550 131.925 ;
        RECT 59.915 131.920 60.175 132.370 ;
        RECT 60.355 132.245 60.630 133.015 ;
        RECT 60.800 132.585 61.130 133.015 ;
        RECT 61.300 132.755 61.495 133.195 ;
        RECT 61.675 132.585 62.005 133.015 ;
        RECT 60.800 132.415 62.005 132.585 ;
        RECT 60.355 132.055 60.940 132.245 ;
        RECT 61.110 132.085 62.005 132.415 ;
        RECT 63.105 132.345 63.485 133.025 ;
        RECT 64.075 132.345 64.245 133.195 ;
        RECT 64.415 132.515 64.745 133.025 ;
        RECT 64.915 132.685 65.085 133.195 ;
        RECT 65.255 132.515 65.655 133.025 ;
        RECT 64.415 132.345 65.655 132.515 ;
        RECT 59.215 131.915 60.175 131.920 ;
        RECT 59.225 131.905 60.175 131.915 ;
        RECT 59.235 131.900 60.175 131.905 ;
        RECT 59.245 131.890 60.175 131.900 ;
        RECT 59.250 131.880 60.175 131.890 ;
        RECT 59.255 131.875 60.175 131.880 ;
        RECT 59.265 131.860 60.175 131.875 ;
        RECT 59.270 131.845 60.175 131.860 ;
        RECT 59.280 131.820 60.175 131.845 ;
        RECT 58.785 131.350 59.115 131.775 ;
        RECT 58.045 130.815 58.305 131.295 ;
        RECT 58.475 130.645 58.725 131.185 ;
        RECT 58.895 130.865 59.115 131.350 ;
        RECT 59.285 131.750 60.175 131.820 ;
        RECT 59.285 131.025 59.455 131.750 ;
        RECT 59.625 131.195 60.175 131.580 ;
        RECT 60.355 131.235 60.595 131.885 ;
        RECT 60.765 131.385 60.940 132.055 ;
        RECT 61.110 131.555 61.525 131.885 ;
        RECT 61.705 131.555 62.000 131.885 ;
        RECT 60.765 131.205 61.095 131.385 ;
        RECT 59.285 130.855 60.175 131.025 ;
        RECT 60.370 130.645 60.700 131.035 ;
        RECT 60.870 130.825 61.095 131.205 ;
        RECT 61.295 130.935 61.525 131.555 ;
        RECT 63.105 131.385 63.275 132.345 ;
        RECT 63.445 132.005 64.750 132.175 ;
        RECT 65.835 132.095 66.155 133.025 ;
        RECT 66.325 132.105 69.835 133.195 ;
        RECT 63.445 131.555 63.690 132.005 ;
        RECT 63.860 131.635 64.410 131.835 ;
        RECT 64.580 131.805 64.750 132.005 ;
        RECT 65.525 131.925 66.155 132.095 ;
        RECT 64.580 131.635 64.955 131.805 ;
        RECT 65.125 131.385 65.355 131.885 ;
        RECT 61.705 130.645 62.005 131.375 ;
        RECT 63.105 131.215 65.355 131.385 ;
        RECT 63.155 130.645 63.485 131.035 ;
        RECT 63.655 130.895 63.825 131.215 ;
        RECT 65.525 131.045 65.695 131.925 ;
        RECT 63.995 130.645 64.325 131.035 ;
        RECT 64.740 130.875 65.695 131.045 ;
        RECT 65.865 130.645 66.155 131.480 ;
        RECT 66.325 131.415 67.975 131.935 ;
        RECT 68.145 131.585 69.835 132.105 ;
        RECT 70.005 132.030 70.295 133.195 ;
        RECT 70.465 132.760 75.810 133.195 ;
        RECT 75.985 132.760 81.330 133.195 ;
        RECT 66.325 130.645 69.835 131.415 ;
        RECT 70.005 130.645 70.295 131.370 ;
        RECT 72.050 131.190 72.390 132.020 ;
        RECT 73.870 131.510 74.220 132.760 ;
        RECT 77.570 131.190 77.910 132.020 ;
        RECT 79.390 131.510 79.740 132.760 ;
        RECT 81.505 132.105 82.715 133.195 ;
        RECT 81.505 131.395 82.025 131.935 ;
        RECT 82.195 131.565 82.715 132.105 ;
        RECT 82.885 132.105 84.095 133.195 ;
        RECT 82.885 131.565 83.405 132.105 ;
        RECT 83.575 131.395 84.095 131.935 ;
        RECT 70.465 130.645 75.810 131.190 ;
        RECT 75.985 130.645 81.330 131.190 ;
        RECT 81.505 130.645 82.715 131.395 ;
        RECT 82.885 130.645 84.095 131.395 ;
        RECT 5.520 130.475 84.180 130.645 ;
        RECT 5.605 129.725 6.815 130.475 ;
        RECT 6.985 129.930 12.330 130.475 ;
        RECT 12.505 129.930 17.850 130.475 ;
        RECT 5.605 129.185 6.125 129.725 ;
        RECT 6.295 129.015 6.815 129.555 ;
        RECT 8.570 129.100 8.910 129.930 ;
        RECT 5.605 127.925 6.815 129.015 ;
        RECT 10.390 128.360 10.740 129.610 ;
        RECT 14.090 129.100 14.430 129.930 ;
        RECT 18.025 129.725 19.235 130.475 ;
        RECT 19.405 129.825 19.665 130.305 ;
        RECT 19.835 130.015 20.165 130.475 ;
        RECT 20.355 129.835 20.555 130.255 ;
        RECT 15.910 128.360 16.260 129.610 ;
        RECT 18.025 129.185 18.545 129.725 ;
        RECT 18.715 129.015 19.235 129.555 ;
        RECT 6.985 127.925 12.330 128.360 ;
        RECT 12.505 127.925 17.850 128.360 ;
        RECT 18.025 127.925 19.235 129.015 ;
        RECT 19.405 128.795 19.575 129.825 ;
        RECT 19.745 129.135 19.975 129.565 ;
        RECT 20.145 129.315 20.555 129.835 ;
        RECT 20.725 129.990 21.515 130.255 ;
        RECT 20.725 129.135 20.980 129.990 ;
        RECT 21.695 129.655 22.025 130.075 ;
        RECT 22.195 129.655 22.455 130.475 ;
        RECT 23.200 129.845 23.485 130.305 ;
        RECT 23.655 130.015 23.925 130.475 ;
        RECT 23.200 129.675 24.155 129.845 ;
        RECT 21.695 129.565 21.945 129.655 ;
        RECT 21.150 129.315 21.945 129.565 ;
        RECT 19.745 128.965 21.535 129.135 ;
        RECT 19.405 128.095 19.680 128.795 ;
        RECT 19.850 128.670 20.565 128.965 ;
        RECT 20.785 128.605 21.115 128.795 ;
        RECT 19.890 127.925 20.105 128.470 ;
        RECT 20.275 128.095 20.750 128.435 ;
        RECT 20.920 128.430 21.115 128.605 ;
        RECT 21.285 128.600 21.535 128.965 ;
        RECT 20.920 127.925 21.535 128.430 ;
        RECT 21.775 128.095 21.945 129.315 ;
        RECT 22.115 128.605 22.455 129.485 ;
        RECT 23.085 128.945 23.775 129.505 ;
        RECT 23.945 128.775 24.155 129.675 ;
        RECT 23.200 128.555 24.155 128.775 ;
        RECT 24.325 129.505 24.725 130.305 ;
        RECT 24.915 129.845 25.195 130.305 ;
        RECT 25.715 130.015 26.040 130.475 ;
        RECT 24.915 129.675 26.040 129.845 ;
        RECT 26.210 129.735 26.595 130.305 ;
        RECT 25.590 129.565 26.040 129.675 ;
        RECT 24.325 128.945 25.420 129.505 ;
        RECT 25.590 129.235 26.145 129.565 ;
        RECT 22.195 127.925 22.455 128.435 ;
        RECT 23.200 128.095 23.485 128.555 ;
        RECT 23.655 127.925 23.925 128.385 ;
        RECT 24.325 128.095 24.725 128.945 ;
        RECT 25.590 128.775 26.040 129.235 ;
        RECT 26.315 129.065 26.595 129.735 ;
        RECT 27.800 129.845 28.085 130.305 ;
        RECT 28.255 130.015 28.525 130.475 ;
        RECT 27.800 129.675 28.755 129.845 ;
        RECT 24.915 128.555 26.040 128.775 ;
        RECT 24.915 128.095 25.195 128.555 ;
        RECT 25.715 127.925 26.040 128.385 ;
        RECT 26.210 128.095 26.595 129.065 ;
        RECT 27.685 128.945 28.375 129.505 ;
        RECT 28.545 128.775 28.755 129.675 ;
        RECT 27.800 128.555 28.755 128.775 ;
        RECT 28.925 129.505 29.325 130.305 ;
        RECT 29.515 129.845 29.795 130.305 ;
        RECT 30.315 130.015 30.640 130.475 ;
        RECT 29.515 129.675 30.640 129.845 ;
        RECT 30.810 129.735 31.195 130.305 ;
        RECT 31.365 129.750 31.655 130.475 ;
        RECT 31.850 130.085 32.180 130.475 ;
        RECT 32.350 129.915 32.575 130.295 ;
        RECT 30.190 129.565 30.640 129.675 ;
        RECT 28.925 128.945 30.020 129.505 ;
        RECT 30.190 129.235 30.745 129.565 ;
        RECT 27.800 128.095 28.085 128.555 ;
        RECT 28.255 127.925 28.525 128.385 ;
        RECT 28.925 128.095 29.325 128.945 ;
        RECT 30.190 128.775 30.640 129.235 ;
        RECT 30.915 129.065 31.195 129.735 ;
        RECT 31.835 129.235 32.075 129.885 ;
        RECT 32.245 129.735 32.575 129.915 ;
        RECT 29.515 128.555 30.640 128.775 ;
        RECT 29.515 128.095 29.795 128.555 ;
        RECT 30.315 127.925 30.640 128.385 ;
        RECT 30.810 128.095 31.195 129.065 ;
        RECT 31.365 127.925 31.655 129.090 ;
        RECT 32.245 129.065 32.420 129.735 ;
        RECT 32.775 129.565 33.005 130.185 ;
        RECT 33.185 129.745 33.485 130.475 ;
        RECT 33.665 129.725 34.875 130.475 ;
        RECT 35.045 129.735 35.430 130.305 ;
        RECT 35.600 130.015 35.925 130.475 ;
        RECT 36.445 129.845 36.725 130.305 ;
        RECT 32.590 129.235 33.005 129.565 ;
        RECT 33.185 129.235 33.480 129.565 ;
        RECT 33.665 129.185 34.185 129.725 ;
        RECT 31.835 128.875 32.420 129.065 ;
        RECT 31.835 128.105 32.110 128.875 ;
        RECT 32.590 128.705 33.485 129.035 ;
        RECT 34.355 129.015 34.875 129.555 ;
        RECT 32.280 128.535 33.485 128.705 ;
        RECT 32.280 128.105 32.610 128.535 ;
        RECT 32.780 127.925 32.975 128.365 ;
        RECT 33.155 128.105 33.485 128.535 ;
        RECT 33.665 127.925 34.875 129.015 ;
        RECT 35.045 129.065 35.325 129.735 ;
        RECT 35.600 129.675 36.725 129.845 ;
        RECT 35.600 129.565 36.050 129.675 ;
        RECT 35.495 129.235 36.050 129.565 ;
        RECT 36.915 129.505 37.315 130.305 ;
        RECT 37.715 130.015 37.985 130.475 ;
        RECT 38.155 129.845 38.440 130.305 ;
        RECT 35.045 128.095 35.430 129.065 ;
        RECT 35.600 128.775 36.050 129.235 ;
        RECT 36.220 128.945 37.315 129.505 ;
        RECT 35.600 128.555 36.725 128.775 ;
        RECT 35.600 127.925 35.925 128.385 ;
        RECT 36.445 128.095 36.725 128.555 ;
        RECT 36.915 128.095 37.315 128.945 ;
        RECT 37.485 129.675 38.440 129.845 ;
        RECT 38.725 129.675 39.420 130.305 ;
        RECT 39.625 129.675 39.935 130.475 ;
        RECT 41.075 130.085 41.405 130.475 ;
        RECT 41.575 129.905 41.745 130.225 ;
        RECT 41.915 130.085 42.245 130.475 ;
        RECT 42.660 130.075 43.615 130.245 ;
        RECT 41.025 129.735 43.275 129.905 ;
        RECT 37.485 128.775 37.695 129.675 ;
        RECT 37.865 128.945 38.555 129.505 ;
        RECT 38.745 129.235 39.080 129.485 ;
        RECT 39.250 129.075 39.420 129.675 ;
        RECT 39.590 129.235 39.925 129.505 ;
        RECT 37.485 128.555 38.440 128.775 ;
        RECT 37.715 127.925 37.985 128.385 ;
        RECT 38.155 128.095 38.440 128.555 ;
        RECT 38.725 127.925 38.985 129.065 ;
        RECT 39.155 128.095 39.485 129.075 ;
        RECT 39.655 127.925 39.935 129.065 ;
        RECT 41.025 128.775 41.195 129.735 ;
        RECT 41.365 129.115 41.610 129.565 ;
        RECT 41.780 129.285 42.330 129.485 ;
        RECT 42.500 129.315 42.875 129.485 ;
        RECT 42.500 129.115 42.670 129.315 ;
        RECT 43.045 129.235 43.275 129.735 ;
        RECT 41.365 128.945 42.670 129.115 ;
        RECT 43.445 129.195 43.615 130.075 ;
        RECT 43.785 129.640 44.075 130.475 ;
        RECT 44.330 129.905 44.505 130.305 ;
        RECT 44.675 130.095 45.005 130.475 ;
        RECT 45.250 129.975 45.480 130.305 ;
        RECT 44.330 129.735 44.960 129.905 ;
        RECT 44.790 129.565 44.960 129.735 ;
        RECT 43.445 129.025 44.075 129.195 ;
        RECT 41.025 128.095 41.405 128.775 ;
        RECT 41.995 127.925 42.165 128.775 ;
        RECT 42.335 128.605 43.575 128.775 ;
        RECT 42.335 128.095 42.665 128.605 ;
        RECT 42.835 127.925 43.005 128.435 ;
        RECT 43.175 128.095 43.575 128.605 ;
        RECT 43.755 128.095 44.075 129.025 ;
        RECT 44.245 128.885 44.610 129.565 ;
        RECT 44.790 129.235 45.140 129.565 ;
        RECT 44.790 128.715 44.960 129.235 ;
        RECT 44.330 128.545 44.960 128.715 ;
        RECT 45.310 128.685 45.480 129.975 ;
        RECT 45.680 128.865 45.960 130.140 ;
        RECT 46.185 130.135 46.455 130.140 ;
        RECT 46.145 129.965 46.455 130.135 ;
        RECT 46.915 130.095 47.245 130.475 ;
        RECT 47.415 130.220 47.750 130.265 ;
        RECT 46.185 128.865 46.455 129.965 ;
        RECT 46.645 128.865 46.985 129.895 ;
        RECT 47.415 129.755 47.755 130.220 ;
        RECT 47.155 129.235 47.415 129.565 ;
        RECT 47.155 128.685 47.325 129.235 ;
        RECT 47.585 129.065 47.755 129.755 ;
        RECT 47.925 129.705 49.595 130.475 ;
        RECT 49.855 129.925 50.025 130.215 ;
        RECT 50.195 130.095 50.525 130.475 ;
        RECT 49.855 129.755 50.520 129.925 ;
        RECT 47.925 129.185 48.675 129.705 ;
        RECT 44.330 128.095 44.505 128.545 ;
        RECT 45.310 128.515 47.325 128.685 ;
        RECT 44.675 127.925 45.005 128.365 ;
        RECT 45.310 128.095 45.480 128.515 ;
        RECT 45.715 127.925 46.385 128.335 ;
        RECT 46.600 128.095 46.770 128.515 ;
        RECT 46.970 127.925 47.300 128.335 ;
        RECT 47.495 128.095 47.755 129.065 ;
        RECT 48.845 129.015 49.595 129.535 ;
        RECT 47.925 127.925 49.595 129.015 ;
        RECT 49.770 128.935 50.120 129.585 ;
        RECT 50.290 128.765 50.520 129.755 ;
        RECT 49.855 128.595 50.520 128.765 ;
        RECT 49.855 128.095 50.025 128.595 ;
        RECT 50.195 127.925 50.525 128.425 ;
        RECT 50.695 128.095 50.880 130.215 ;
        RECT 51.135 130.015 51.385 130.475 ;
        RECT 51.555 130.025 51.890 130.195 ;
        RECT 52.085 130.025 52.760 130.195 ;
        RECT 51.555 129.885 51.725 130.025 ;
        RECT 51.050 128.895 51.330 129.845 ;
        RECT 51.500 129.755 51.725 129.885 ;
        RECT 51.500 128.650 51.670 129.755 ;
        RECT 51.895 129.605 52.420 129.825 ;
        RECT 51.840 128.840 52.080 129.435 ;
        RECT 52.250 128.905 52.420 129.605 ;
        RECT 52.590 129.245 52.760 130.025 ;
        RECT 53.080 129.975 53.450 130.475 ;
        RECT 53.630 130.025 54.035 130.195 ;
        RECT 54.205 130.025 54.990 130.195 ;
        RECT 53.630 129.795 53.800 130.025 ;
        RECT 52.970 129.495 53.800 129.795 ;
        RECT 54.185 129.525 54.650 129.855 ;
        RECT 52.970 129.465 53.170 129.495 ;
        RECT 53.290 129.245 53.460 129.315 ;
        RECT 52.590 129.075 53.460 129.245 ;
        RECT 52.950 128.985 53.460 129.075 ;
        RECT 51.500 128.520 51.805 128.650 ;
        RECT 52.250 128.540 52.780 128.905 ;
        RECT 51.120 127.925 51.385 128.385 ;
        RECT 51.555 128.095 51.805 128.520 ;
        RECT 52.950 128.370 53.120 128.985 ;
        RECT 52.015 128.200 53.120 128.370 ;
        RECT 53.290 127.925 53.460 128.725 ;
        RECT 53.630 128.425 53.800 129.495 ;
        RECT 53.970 128.595 54.160 129.315 ;
        RECT 54.330 128.565 54.650 129.525 ;
        RECT 54.820 129.565 54.990 130.025 ;
        RECT 55.265 129.945 55.475 130.475 ;
        RECT 55.735 129.735 56.065 130.260 ;
        RECT 56.235 129.865 56.405 130.475 ;
        RECT 56.575 129.820 56.905 130.255 ;
        RECT 56.575 129.735 56.955 129.820 ;
        RECT 57.125 129.750 57.415 130.475 ;
        RECT 58.595 129.925 58.765 130.215 ;
        RECT 58.935 130.095 59.265 130.475 ;
        RECT 58.595 129.755 59.260 129.925 ;
        RECT 55.865 129.565 56.065 129.735 ;
        RECT 56.730 129.695 56.955 129.735 ;
        RECT 54.820 129.235 55.695 129.565 ;
        RECT 55.865 129.235 56.615 129.565 ;
        RECT 53.630 128.095 53.880 128.425 ;
        RECT 54.820 128.395 54.990 129.235 ;
        RECT 55.865 129.030 56.055 129.235 ;
        RECT 56.785 129.115 56.955 129.695 ;
        RECT 56.740 129.065 56.955 129.115 ;
        RECT 55.160 128.655 56.055 129.030 ;
        RECT 56.565 128.985 56.955 129.065 ;
        RECT 54.105 128.225 54.990 128.395 ;
        RECT 55.170 127.925 55.485 128.425 ;
        RECT 55.715 128.095 56.055 128.655 ;
        RECT 56.225 127.925 56.395 128.935 ;
        RECT 56.565 128.140 56.895 128.985 ;
        RECT 57.125 127.925 57.415 129.090 ;
        RECT 58.510 128.935 58.860 129.585 ;
        RECT 59.030 128.765 59.260 129.755 ;
        RECT 58.595 128.595 59.260 128.765 ;
        RECT 58.595 128.095 58.765 128.595 ;
        RECT 58.935 127.925 59.265 128.425 ;
        RECT 59.435 128.095 59.620 130.215 ;
        RECT 59.875 130.015 60.125 130.475 ;
        RECT 60.295 130.025 60.630 130.195 ;
        RECT 60.825 130.025 61.500 130.195 ;
        RECT 60.295 129.885 60.465 130.025 ;
        RECT 59.790 128.895 60.070 129.845 ;
        RECT 60.240 129.755 60.465 129.885 ;
        RECT 60.240 128.650 60.410 129.755 ;
        RECT 60.635 129.605 61.160 129.825 ;
        RECT 60.580 128.840 60.820 129.435 ;
        RECT 60.990 128.905 61.160 129.605 ;
        RECT 61.330 129.245 61.500 130.025 ;
        RECT 61.820 129.975 62.190 130.475 ;
        RECT 62.370 130.025 62.775 130.195 ;
        RECT 62.945 130.025 63.730 130.195 ;
        RECT 62.370 129.795 62.540 130.025 ;
        RECT 61.710 129.495 62.540 129.795 ;
        RECT 62.925 129.525 63.390 129.855 ;
        RECT 61.710 129.465 61.910 129.495 ;
        RECT 62.030 129.245 62.200 129.315 ;
        RECT 61.330 129.075 62.200 129.245 ;
        RECT 61.690 128.985 62.200 129.075 ;
        RECT 60.240 128.520 60.545 128.650 ;
        RECT 60.990 128.540 61.520 128.905 ;
        RECT 59.860 127.925 60.125 128.385 ;
        RECT 60.295 128.095 60.545 128.520 ;
        RECT 61.690 128.370 61.860 128.985 ;
        RECT 60.755 128.200 61.860 128.370 ;
        RECT 62.030 127.925 62.200 128.725 ;
        RECT 62.370 128.425 62.540 129.495 ;
        RECT 62.710 128.595 62.900 129.315 ;
        RECT 63.070 128.565 63.390 129.525 ;
        RECT 63.560 129.565 63.730 130.025 ;
        RECT 64.005 129.945 64.215 130.475 ;
        RECT 64.475 129.735 64.805 130.260 ;
        RECT 64.975 129.865 65.145 130.475 ;
        RECT 65.315 129.820 65.645 130.255 ;
        RECT 65.865 129.930 71.210 130.475 ;
        RECT 71.385 129.930 76.730 130.475 ;
        RECT 76.905 129.930 82.250 130.475 ;
        RECT 65.315 129.735 65.695 129.820 ;
        RECT 64.605 129.565 64.805 129.735 ;
        RECT 65.470 129.695 65.695 129.735 ;
        RECT 63.560 129.235 64.435 129.565 ;
        RECT 64.605 129.235 65.355 129.565 ;
        RECT 62.370 128.095 62.620 128.425 ;
        RECT 63.560 128.395 63.730 129.235 ;
        RECT 64.605 129.030 64.795 129.235 ;
        RECT 65.525 129.115 65.695 129.695 ;
        RECT 65.480 129.065 65.695 129.115 ;
        RECT 67.450 129.100 67.790 129.930 ;
        RECT 63.900 128.655 64.795 129.030 ;
        RECT 65.305 128.985 65.695 129.065 ;
        RECT 62.845 128.225 63.730 128.395 ;
        RECT 63.910 127.925 64.225 128.425 ;
        RECT 64.455 128.095 64.795 128.655 ;
        RECT 64.965 127.925 65.135 128.935 ;
        RECT 65.305 128.140 65.635 128.985 ;
        RECT 69.270 128.360 69.620 129.610 ;
        RECT 72.970 129.100 73.310 129.930 ;
        RECT 74.790 128.360 75.140 129.610 ;
        RECT 78.490 129.100 78.830 129.930 ;
        RECT 82.885 129.725 84.095 130.475 ;
        RECT 80.310 128.360 80.660 129.610 ;
        RECT 82.885 129.015 83.405 129.555 ;
        RECT 83.575 129.185 84.095 129.725 ;
        RECT 65.865 127.925 71.210 128.360 ;
        RECT 71.385 127.925 76.730 128.360 ;
        RECT 76.905 127.925 82.250 128.360 ;
        RECT 82.885 127.925 84.095 129.015 ;
        RECT 5.520 127.755 84.180 127.925 ;
        RECT 5.605 126.665 6.815 127.755 ;
        RECT 6.985 127.320 12.330 127.755 ;
        RECT 12.505 127.320 17.850 127.755 ;
        RECT 5.605 125.955 6.125 126.495 ;
        RECT 6.295 126.125 6.815 126.665 ;
        RECT 5.605 125.205 6.815 125.955 ;
        RECT 8.570 125.750 8.910 126.580 ;
        RECT 10.390 126.070 10.740 127.320 ;
        RECT 14.090 125.750 14.430 126.580 ;
        RECT 15.910 126.070 16.260 127.320 ;
        RECT 18.485 126.590 18.775 127.755 ;
        RECT 19.005 126.695 19.335 127.540 ;
        RECT 19.505 126.745 19.675 127.755 ;
        RECT 19.845 127.025 20.185 127.585 ;
        RECT 20.415 127.255 20.730 127.755 ;
        RECT 20.910 127.285 21.795 127.455 ;
        RECT 18.945 126.615 19.335 126.695 ;
        RECT 19.845 126.650 20.740 127.025 ;
        RECT 18.945 126.565 19.160 126.615 ;
        RECT 18.945 125.985 19.115 126.565 ;
        RECT 19.845 126.445 20.035 126.650 ;
        RECT 20.910 126.445 21.080 127.285 ;
        RECT 22.020 127.255 22.270 127.585 ;
        RECT 19.285 126.115 20.035 126.445 ;
        RECT 20.205 126.115 21.080 126.445 ;
        RECT 18.945 125.945 19.170 125.985 ;
        RECT 19.835 125.945 20.035 126.115 ;
        RECT 6.985 125.205 12.330 125.750 ;
        RECT 12.505 125.205 17.850 125.750 ;
        RECT 18.485 125.205 18.775 125.930 ;
        RECT 18.945 125.860 19.325 125.945 ;
        RECT 18.995 125.425 19.325 125.860 ;
        RECT 19.495 125.205 19.665 125.815 ;
        RECT 19.835 125.420 20.165 125.945 ;
        RECT 20.425 125.205 20.635 125.735 ;
        RECT 20.910 125.655 21.080 126.115 ;
        RECT 21.250 126.155 21.570 127.115 ;
        RECT 21.740 126.365 21.930 127.085 ;
        RECT 22.100 126.185 22.270 127.255 ;
        RECT 22.440 126.955 22.610 127.755 ;
        RECT 22.780 127.310 23.885 127.480 ;
        RECT 22.780 126.695 22.950 127.310 ;
        RECT 24.095 127.160 24.345 127.585 ;
        RECT 24.515 127.295 24.780 127.755 ;
        RECT 23.120 126.775 23.650 127.140 ;
        RECT 24.095 127.030 24.400 127.160 ;
        RECT 22.440 126.605 22.950 126.695 ;
        RECT 22.440 126.435 23.310 126.605 ;
        RECT 22.440 126.365 22.610 126.435 ;
        RECT 22.730 126.185 22.930 126.215 ;
        RECT 21.250 125.825 21.715 126.155 ;
        RECT 22.100 125.885 22.930 126.185 ;
        RECT 22.100 125.655 22.270 125.885 ;
        RECT 20.910 125.485 21.695 125.655 ;
        RECT 21.865 125.485 22.270 125.655 ;
        RECT 22.450 125.205 22.820 125.705 ;
        RECT 23.140 125.655 23.310 126.435 ;
        RECT 23.480 126.075 23.650 126.775 ;
        RECT 23.820 126.245 24.060 126.840 ;
        RECT 23.480 125.855 24.005 126.075 ;
        RECT 24.230 125.925 24.400 127.030 ;
        RECT 24.175 125.795 24.400 125.925 ;
        RECT 24.570 125.835 24.850 126.785 ;
        RECT 24.175 125.655 24.345 125.795 ;
        RECT 23.140 125.485 23.815 125.655 ;
        RECT 24.010 125.485 24.345 125.655 ;
        RECT 24.515 125.205 24.765 125.665 ;
        RECT 25.020 125.465 25.205 127.585 ;
        RECT 25.375 127.255 25.705 127.755 ;
        RECT 25.875 127.085 26.045 127.585 ;
        RECT 25.380 126.915 26.045 127.085 ;
        RECT 26.340 126.965 26.875 127.585 ;
        RECT 25.380 125.925 25.610 126.915 ;
        RECT 25.780 126.095 26.130 126.745 ;
        RECT 26.340 125.945 26.655 126.965 ;
        RECT 27.045 126.955 27.375 127.755 ;
        RECT 28.695 127.085 28.865 127.585 ;
        RECT 29.035 127.255 29.365 127.755 ;
        RECT 27.860 126.785 28.250 126.960 ;
        RECT 28.695 126.915 29.360 127.085 ;
        RECT 26.825 126.615 28.250 126.785 ;
        RECT 26.825 126.115 26.995 126.615 ;
        RECT 25.380 125.755 26.045 125.925 ;
        RECT 25.375 125.205 25.705 125.585 ;
        RECT 25.875 125.465 26.045 125.755 ;
        RECT 26.340 125.375 26.955 125.945 ;
        RECT 27.245 125.885 27.510 126.445 ;
        RECT 27.680 125.715 27.850 126.615 ;
        RECT 28.020 125.885 28.375 126.445 ;
        RECT 28.610 126.095 28.960 126.745 ;
        RECT 29.130 125.925 29.360 126.915 ;
        RECT 28.695 125.755 29.360 125.925 ;
        RECT 27.125 125.205 27.340 125.715 ;
        RECT 27.570 125.385 27.850 125.715 ;
        RECT 28.030 125.205 28.270 125.715 ;
        RECT 28.695 125.465 28.865 125.755 ;
        RECT 29.035 125.205 29.365 125.585 ;
        RECT 29.535 125.465 29.720 127.585 ;
        RECT 29.960 127.295 30.225 127.755 ;
        RECT 30.395 127.160 30.645 127.585 ;
        RECT 30.855 127.310 31.960 127.480 ;
        RECT 30.340 127.030 30.645 127.160 ;
        RECT 29.890 125.835 30.170 126.785 ;
        RECT 30.340 125.925 30.510 127.030 ;
        RECT 30.680 126.245 30.920 126.840 ;
        RECT 31.090 126.775 31.620 127.140 ;
        RECT 31.090 126.075 31.260 126.775 ;
        RECT 31.790 126.695 31.960 127.310 ;
        RECT 32.130 126.955 32.300 127.755 ;
        RECT 32.470 127.255 32.720 127.585 ;
        RECT 32.945 127.285 33.830 127.455 ;
        RECT 31.790 126.605 32.300 126.695 ;
        RECT 30.340 125.795 30.565 125.925 ;
        RECT 30.735 125.855 31.260 126.075 ;
        RECT 31.430 126.435 32.300 126.605 ;
        RECT 29.975 125.205 30.225 125.665 ;
        RECT 30.395 125.655 30.565 125.795 ;
        RECT 31.430 125.655 31.600 126.435 ;
        RECT 32.130 126.365 32.300 126.435 ;
        RECT 31.810 126.185 32.010 126.215 ;
        RECT 32.470 126.185 32.640 127.255 ;
        RECT 32.810 126.365 33.000 127.085 ;
        RECT 31.810 125.885 32.640 126.185 ;
        RECT 33.170 126.155 33.490 127.115 ;
        RECT 30.395 125.485 30.730 125.655 ;
        RECT 30.925 125.485 31.600 125.655 ;
        RECT 31.920 125.205 32.290 125.705 ;
        RECT 32.470 125.655 32.640 125.885 ;
        RECT 33.025 125.825 33.490 126.155 ;
        RECT 33.660 126.445 33.830 127.285 ;
        RECT 34.010 127.255 34.325 127.755 ;
        RECT 34.555 127.025 34.895 127.585 ;
        RECT 34.000 126.650 34.895 127.025 ;
        RECT 35.065 126.745 35.235 127.755 ;
        RECT 34.705 126.445 34.895 126.650 ;
        RECT 35.405 126.695 35.735 127.540 ;
        RECT 36.045 127.125 36.225 127.585 ;
        RECT 36.395 127.295 36.645 127.755 ;
        RECT 36.815 127.375 37.145 127.545 ;
        RECT 37.315 127.490 37.570 127.585 ;
        RECT 36.815 127.125 36.985 127.375 ;
        RECT 37.315 127.320 38.455 127.490 ;
        RECT 38.715 127.355 39.045 127.755 ;
        RECT 37.315 127.185 37.570 127.320 ;
        RECT 36.045 126.955 36.985 127.125 ;
        RECT 37.160 127.015 37.570 127.185 ;
        RECT 38.285 127.095 38.455 127.320 ;
        RECT 35.405 126.615 35.795 126.695 ;
        RECT 35.580 126.565 35.795 126.615 ;
        RECT 33.660 126.115 34.535 126.445 ;
        RECT 34.705 126.115 35.455 126.445 ;
        RECT 33.660 125.655 33.830 126.115 ;
        RECT 34.705 125.945 34.905 126.115 ;
        RECT 35.625 125.985 35.795 126.565 ;
        RECT 35.570 125.945 35.795 125.985 ;
        RECT 32.470 125.485 32.875 125.655 ;
        RECT 33.045 125.485 33.830 125.655 ;
        RECT 34.105 125.205 34.315 125.735 ;
        RECT 34.575 125.420 34.905 125.945 ;
        RECT 35.415 125.860 35.795 125.945 ;
        RECT 36.020 125.885 36.280 126.775 ;
        RECT 36.480 126.475 36.960 126.775 ;
        RECT 36.480 125.885 36.740 126.475 ;
        RECT 37.160 125.990 37.330 127.015 ;
        RECT 37.850 126.835 38.020 127.025 ;
        RECT 38.285 126.925 39.045 127.095 ;
        RECT 35.075 125.205 35.245 125.815 ;
        RECT 35.415 125.425 35.745 125.860 ;
        RECT 36.980 125.820 37.330 125.990 ;
        RECT 37.500 126.665 38.020 126.835 ;
        RECT 37.500 125.945 37.670 126.665 ;
        RECT 37.860 126.115 38.150 126.495 ;
        RECT 38.320 126.115 38.650 126.735 ;
        RECT 38.875 126.445 39.045 126.925 ;
        RECT 39.215 126.645 39.475 127.585 ;
        RECT 38.875 126.115 39.130 126.445 ;
        RECT 36.005 125.205 36.405 125.715 ;
        RECT 36.980 125.375 37.150 125.820 ;
        RECT 37.500 125.775 38.380 125.945 ;
        RECT 39.300 125.930 39.475 126.645 ;
        RECT 37.320 125.205 38.040 125.605 ;
        RECT 38.210 125.375 38.380 125.775 ;
        RECT 38.615 125.205 39.045 125.650 ;
        RECT 39.215 125.375 39.475 125.930 ;
        RECT 39.645 126.615 40.030 127.585 ;
        RECT 40.200 127.295 40.525 127.755 ;
        RECT 41.045 127.125 41.325 127.585 ;
        RECT 40.200 126.905 41.325 127.125 ;
        RECT 39.645 125.945 39.925 126.615 ;
        RECT 40.200 126.445 40.650 126.905 ;
        RECT 41.515 126.735 41.915 127.585 ;
        RECT 42.315 127.295 42.585 127.755 ;
        RECT 42.755 127.125 43.040 127.585 ;
        RECT 40.095 126.115 40.650 126.445 ;
        RECT 40.820 126.175 41.915 126.735 ;
        RECT 40.200 126.005 40.650 126.115 ;
        RECT 39.645 125.375 40.030 125.945 ;
        RECT 40.200 125.835 41.325 126.005 ;
        RECT 40.200 125.205 40.525 125.665 ;
        RECT 41.045 125.375 41.325 125.835 ;
        RECT 41.515 125.375 41.915 126.175 ;
        RECT 42.085 126.905 43.040 127.125 ;
        RECT 42.085 126.005 42.295 126.905 ;
        RECT 42.465 126.175 43.155 126.735 ;
        RECT 44.245 126.590 44.535 127.755 ;
        RECT 44.705 126.615 44.965 127.755 ;
        RECT 45.135 126.605 45.465 127.585 ;
        RECT 45.635 126.615 45.915 127.755 ;
        RECT 46.175 127.085 46.345 127.585 ;
        RECT 46.515 127.255 46.845 127.755 ;
        RECT 46.175 126.915 46.840 127.085 ;
        RECT 44.725 126.195 45.060 126.445 ;
        RECT 45.230 126.005 45.400 126.605 ;
        RECT 45.570 126.175 45.905 126.445 ;
        RECT 46.090 126.095 46.440 126.745 ;
        RECT 42.085 125.835 43.040 126.005 ;
        RECT 42.315 125.205 42.585 125.665 ;
        RECT 42.755 125.375 43.040 125.835 ;
        RECT 44.245 125.205 44.535 125.930 ;
        RECT 44.705 125.375 45.400 126.005 ;
        RECT 45.605 125.205 45.915 126.005 ;
        RECT 46.610 125.925 46.840 126.915 ;
        RECT 46.175 125.755 46.840 125.925 ;
        RECT 46.175 125.465 46.345 125.755 ;
        RECT 46.515 125.205 46.845 125.585 ;
        RECT 47.015 125.465 47.200 127.585 ;
        RECT 47.440 127.295 47.705 127.755 ;
        RECT 47.875 127.160 48.125 127.585 ;
        RECT 48.335 127.310 49.440 127.480 ;
        RECT 47.820 127.030 48.125 127.160 ;
        RECT 47.370 125.835 47.650 126.785 ;
        RECT 47.820 125.925 47.990 127.030 ;
        RECT 48.160 126.245 48.400 126.840 ;
        RECT 48.570 126.775 49.100 127.140 ;
        RECT 48.570 126.075 48.740 126.775 ;
        RECT 49.270 126.695 49.440 127.310 ;
        RECT 49.610 126.955 49.780 127.755 ;
        RECT 49.950 127.255 50.200 127.585 ;
        RECT 50.425 127.285 51.310 127.455 ;
        RECT 49.270 126.605 49.780 126.695 ;
        RECT 47.820 125.795 48.045 125.925 ;
        RECT 48.215 125.855 48.740 126.075 ;
        RECT 48.910 126.435 49.780 126.605 ;
        RECT 47.455 125.205 47.705 125.665 ;
        RECT 47.875 125.655 48.045 125.795 ;
        RECT 48.910 125.655 49.080 126.435 ;
        RECT 49.610 126.365 49.780 126.435 ;
        RECT 49.290 126.185 49.490 126.215 ;
        RECT 49.950 126.185 50.120 127.255 ;
        RECT 50.290 126.365 50.480 127.085 ;
        RECT 49.290 125.885 50.120 126.185 ;
        RECT 50.650 126.155 50.970 127.115 ;
        RECT 47.875 125.485 48.210 125.655 ;
        RECT 48.405 125.485 49.080 125.655 ;
        RECT 49.400 125.205 49.770 125.705 ;
        RECT 49.950 125.655 50.120 125.885 ;
        RECT 50.505 125.825 50.970 126.155 ;
        RECT 51.140 126.445 51.310 127.285 ;
        RECT 51.490 127.255 51.805 127.755 ;
        RECT 52.035 127.025 52.375 127.585 ;
        RECT 51.480 126.650 52.375 127.025 ;
        RECT 52.545 126.745 52.715 127.755 ;
        RECT 52.185 126.445 52.375 126.650 ;
        RECT 52.885 126.695 53.215 127.540 ;
        RECT 52.885 126.615 53.275 126.695 ;
        RECT 53.445 126.665 56.955 127.755 ;
        RECT 57.670 127.135 57.845 127.585 ;
        RECT 58.015 127.315 58.345 127.755 ;
        RECT 58.650 127.165 58.820 127.585 ;
        RECT 59.055 127.345 59.725 127.755 ;
        RECT 59.940 127.165 60.110 127.585 ;
        RECT 60.310 127.345 60.640 127.755 ;
        RECT 57.670 126.965 58.300 127.135 ;
        RECT 53.060 126.565 53.275 126.615 ;
        RECT 51.140 126.115 52.015 126.445 ;
        RECT 52.185 126.115 52.935 126.445 ;
        RECT 51.140 125.655 51.310 126.115 ;
        RECT 52.185 125.945 52.385 126.115 ;
        RECT 53.105 125.985 53.275 126.565 ;
        RECT 53.050 125.945 53.275 125.985 ;
        RECT 49.950 125.485 50.355 125.655 ;
        RECT 50.525 125.485 51.310 125.655 ;
        RECT 51.585 125.205 51.795 125.735 ;
        RECT 52.055 125.420 52.385 125.945 ;
        RECT 52.895 125.860 53.275 125.945 ;
        RECT 53.445 125.975 55.095 126.495 ;
        RECT 55.265 126.145 56.955 126.665 ;
        RECT 57.585 126.115 57.950 126.795 ;
        RECT 58.130 126.445 58.300 126.965 ;
        RECT 58.650 126.995 60.665 127.165 ;
        RECT 58.130 126.115 58.480 126.445 ;
        RECT 52.555 125.205 52.725 125.815 ;
        RECT 52.895 125.425 53.225 125.860 ;
        RECT 53.445 125.205 56.955 125.975 ;
        RECT 58.130 125.945 58.300 126.115 ;
        RECT 57.670 125.775 58.300 125.945 ;
        RECT 57.670 125.375 57.845 125.775 ;
        RECT 58.650 125.705 58.820 126.995 ;
        RECT 58.015 125.205 58.345 125.585 ;
        RECT 58.590 125.375 58.820 125.705 ;
        RECT 59.020 125.540 59.300 126.815 ;
        RECT 59.525 125.715 59.795 126.815 ;
        RECT 59.985 125.785 60.325 126.815 ;
        RECT 60.495 126.445 60.665 126.995 ;
        RECT 60.835 126.615 61.095 127.585 ;
        RECT 61.265 127.320 66.610 127.755 ;
        RECT 60.495 126.115 60.755 126.445 ;
        RECT 60.925 125.925 61.095 126.615 ;
        RECT 59.485 125.545 59.795 125.715 ;
        RECT 59.525 125.540 59.795 125.545 ;
        RECT 60.255 125.205 60.585 125.585 ;
        RECT 60.755 125.460 61.095 125.925 ;
        RECT 62.850 125.750 63.190 126.580 ;
        RECT 64.670 126.070 65.020 127.320 ;
        RECT 66.785 126.665 69.375 127.755 ;
        RECT 66.785 125.975 67.995 126.495 ;
        RECT 68.165 126.145 69.375 126.665 ;
        RECT 70.005 126.590 70.295 127.755 ;
        RECT 70.465 127.320 75.810 127.755 ;
        RECT 75.985 127.320 81.330 127.755 ;
        RECT 60.755 125.415 61.090 125.460 ;
        RECT 61.265 125.205 66.610 125.750 ;
        RECT 66.785 125.205 69.375 125.975 ;
        RECT 70.005 125.205 70.295 125.930 ;
        RECT 72.050 125.750 72.390 126.580 ;
        RECT 73.870 126.070 74.220 127.320 ;
        RECT 77.570 125.750 77.910 126.580 ;
        RECT 79.390 126.070 79.740 127.320 ;
        RECT 81.505 126.665 82.715 127.755 ;
        RECT 81.505 125.955 82.025 126.495 ;
        RECT 82.195 126.125 82.715 126.665 ;
        RECT 82.885 126.665 84.095 127.755 ;
        RECT 82.885 126.125 83.405 126.665 ;
        RECT 83.575 125.955 84.095 126.495 ;
        RECT 70.465 125.205 75.810 125.750 ;
        RECT 75.985 125.205 81.330 125.750 ;
        RECT 81.505 125.205 82.715 125.955 ;
        RECT 82.885 125.205 84.095 125.955 ;
        RECT 5.520 125.035 84.180 125.205 ;
        RECT 5.605 124.285 6.815 125.035 ;
        RECT 6.985 124.490 12.330 125.035 ;
        RECT 12.505 124.490 17.850 125.035 ;
        RECT 5.605 123.745 6.125 124.285 ;
        RECT 6.295 123.575 6.815 124.115 ;
        RECT 8.570 123.660 8.910 124.490 ;
        RECT 5.605 122.485 6.815 123.575 ;
        RECT 10.390 122.920 10.740 124.170 ;
        RECT 14.090 123.660 14.430 124.490 ;
        RECT 18.025 124.265 20.615 125.035 ;
        RECT 20.835 124.380 21.165 124.815 ;
        RECT 21.335 124.425 21.505 125.035 ;
        RECT 20.785 124.295 21.165 124.380 ;
        RECT 21.675 124.295 22.005 124.820 ;
        RECT 22.265 124.505 22.475 125.035 ;
        RECT 22.750 124.585 23.535 124.755 ;
        RECT 23.705 124.585 24.110 124.755 ;
        RECT 15.910 122.920 16.260 124.170 ;
        RECT 18.025 123.745 19.235 124.265 ;
        RECT 20.785 124.255 21.010 124.295 ;
        RECT 19.405 123.575 20.615 124.095 ;
        RECT 6.985 122.485 12.330 122.920 ;
        RECT 12.505 122.485 17.850 122.920 ;
        RECT 18.025 122.485 20.615 123.575 ;
        RECT 20.785 123.675 20.955 124.255 ;
        RECT 21.675 124.125 21.875 124.295 ;
        RECT 22.750 124.125 22.920 124.585 ;
        RECT 21.125 123.795 21.875 124.125 ;
        RECT 22.045 123.795 22.920 124.125 ;
        RECT 20.785 123.625 21.000 123.675 ;
        RECT 20.785 123.545 21.175 123.625 ;
        RECT 20.845 122.700 21.175 123.545 ;
        RECT 21.685 123.590 21.875 123.795 ;
        RECT 21.345 122.485 21.515 123.495 ;
        RECT 21.685 123.215 22.580 123.590 ;
        RECT 21.685 122.655 22.025 123.215 ;
        RECT 22.255 122.485 22.570 122.985 ;
        RECT 22.750 122.955 22.920 123.795 ;
        RECT 23.090 124.085 23.555 124.415 ;
        RECT 23.940 124.355 24.110 124.585 ;
        RECT 24.290 124.535 24.660 125.035 ;
        RECT 24.980 124.585 25.655 124.755 ;
        RECT 25.850 124.585 26.185 124.755 ;
        RECT 23.090 123.125 23.410 124.085 ;
        RECT 23.940 124.055 24.770 124.355 ;
        RECT 23.580 123.155 23.770 123.875 ;
        RECT 23.940 122.985 24.110 124.055 ;
        RECT 24.570 124.025 24.770 124.055 ;
        RECT 24.280 123.805 24.450 123.875 ;
        RECT 24.980 123.805 25.150 124.585 ;
        RECT 26.015 124.445 26.185 124.585 ;
        RECT 26.355 124.575 26.605 125.035 ;
        RECT 24.280 123.635 25.150 123.805 ;
        RECT 25.320 124.165 25.845 124.385 ;
        RECT 26.015 124.315 26.240 124.445 ;
        RECT 24.280 123.545 24.790 123.635 ;
        RECT 22.750 122.785 23.635 122.955 ;
        RECT 23.860 122.655 24.110 122.985 ;
        RECT 24.280 122.485 24.450 123.285 ;
        RECT 24.620 122.930 24.790 123.545 ;
        RECT 25.320 123.465 25.490 124.165 ;
        RECT 24.960 123.100 25.490 123.465 ;
        RECT 25.660 123.400 25.900 123.995 ;
        RECT 26.070 123.210 26.240 124.315 ;
        RECT 26.410 123.455 26.690 124.405 ;
        RECT 25.935 123.080 26.240 123.210 ;
        RECT 24.620 122.760 25.725 122.930 ;
        RECT 25.935 122.655 26.185 123.080 ;
        RECT 26.355 122.485 26.620 122.945 ;
        RECT 26.860 122.655 27.045 124.775 ;
        RECT 27.215 124.655 27.545 125.035 ;
        RECT 27.715 124.485 27.885 124.775 ;
        RECT 27.220 124.315 27.885 124.485 ;
        RECT 27.220 123.325 27.450 124.315 ;
        RECT 28.145 124.295 28.465 124.775 ;
        RECT 28.635 124.465 28.865 124.865 ;
        RECT 29.035 124.645 29.385 125.035 ;
        RECT 28.635 124.385 29.145 124.465 ;
        RECT 29.555 124.385 29.885 124.865 ;
        RECT 28.635 124.295 29.885 124.385 ;
        RECT 27.620 123.495 27.970 124.145 ;
        RECT 28.145 123.365 28.315 124.295 ;
        RECT 28.975 124.215 29.885 124.295 ;
        RECT 30.055 124.215 30.225 125.035 ;
        RECT 30.730 124.295 31.195 124.840 ;
        RECT 31.365 124.310 31.655 125.035 ;
        RECT 32.860 124.405 33.145 124.865 ;
        RECT 33.315 124.575 33.585 125.035 ;
        RECT 28.485 123.705 28.655 124.125 ;
        RECT 28.885 123.875 29.485 124.045 ;
        RECT 28.485 123.535 29.145 123.705 ;
        RECT 27.220 123.155 27.885 123.325 ;
        RECT 28.145 123.165 28.805 123.365 ;
        RECT 28.975 123.335 29.145 123.535 ;
        RECT 29.315 123.675 29.485 123.875 ;
        RECT 29.655 123.845 30.350 124.045 ;
        RECT 30.610 123.675 30.855 124.125 ;
        RECT 29.315 123.505 30.855 123.675 ;
        RECT 31.025 123.335 31.195 124.295 ;
        RECT 32.860 124.235 33.815 124.405 ;
        RECT 28.975 123.165 31.195 123.335 ;
        RECT 27.215 122.485 27.545 122.985 ;
        RECT 27.715 122.655 27.885 123.155 ;
        RECT 28.635 122.995 28.805 123.165 ;
        RECT 28.165 122.485 28.465 122.995 ;
        RECT 28.635 122.825 29.015 122.995 ;
        RECT 29.595 122.485 30.225 122.995 ;
        RECT 30.395 122.655 30.725 123.165 ;
        RECT 30.895 122.485 31.195 122.995 ;
        RECT 31.365 122.485 31.655 123.650 ;
        RECT 32.745 123.505 33.435 124.065 ;
        RECT 33.605 123.335 33.815 124.235 ;
        RECT 32.860 123.115 33.815 123.335 ;
        RECT 33.985 124.065 34.385 124.865 ;
        RECT 34.575 124.405 34.855 124.865 ;
        RECT 35.375 124.575 35.700 125.035 ;
        RECT 34.575 124.235 35.700 124.405 ;
        RECT 35.870 124.295 36.255 124.865 ;
        RECT 36.465 124.525 36.865 125.035 ;
        RECT 37.440 124.420 37.610 124.865 ;
        RECT 37.780 124.635 38.500 125.035 ;
        RECT 38.670 124.465 38.840 124.865 ;
        RECT 39.075 124.590 39.505 125.035 ;
        RECT 35.250 124.125 35.700 124.235 ;
        RECT 33.985 123.505 35.080 124.065 ;
        RECT 35.250 123.795 35.805 124.125 ;
        RECT 32.860 122.655 33.145 123.115 ;
        RECT 33.315 122.485 33.585 122.945 ;
        RECT 33.985 122.655 34.385 123.505 ;
        RECT 35.250 123.335 35.700 123.795 ;
        RECT 35.975 123.625 36.255 124.295 ;
        RECT 34.575 123.115 35.700 123.335 ;
        RECT 34.575 122.655 34.855 123.115 ;
        RECT 35.375 122.485 35.700 122.945 ;
        RECT 35.870 122.655 36.255 123.625 ;
        RECT 36.480 123.465 36.740 124.355 ;
        RECT 36.940 123.765 37.200 124.355 ;
        RECT 37.440 124.250 37.790 124.420 ;
        RECT 36.940 123.465 37.420 123.765 ;
        RECT 36.505 123.115 37.445 123.285 ;
        RECT 36.505 122.655 36.685 123.115 ;
        RECT 36.855 122.485 37.105 122.945 ;
        RECT 37.275 122.865 37.445 123.115 ;
        RECT 37.620 123.225 37.790 124.250 ;
        RECT 37.960 124.295 38.840 124.465 ;
        RECT 39.675 124.310 39.935 124.865 ;
        RECT 40.195 124.485 40.365 124.775 ;
        RECT 40.535 124.655 40.865 125.035 ;
        RECT 40.195 124.315 40.860 124.485 ;
        RECT 37.960 123.575 38.130 124.295 ;
        RECT 38.320 123.745 38.610 124.125 ;
        RECT 37.960 123.405 38.480 123.575 ;
        RECT 38.780 123.505 39.110 124.125 ;
        RECT 39.335 123.795 39.590 124.125 ;
        RECT 37.620 123.055 38.030 123.225 ;
        RECT 38.310 123.215 38.480 123.405 ;
        RECT 39.335 123.315 39.505 123.795 ;
        RECT 39.760 123.595 39.935 124.310 ;
        RECT 37.775 122.920 38.030 123.055 ;
        RECT 38.745 123.145 39.505 123.315 ;
        RECT 38.745 122.920 38.915 123.145 ;
        RECT 37.275 122.695 37.605 122.865 ;
        RECT 37.775 122.750 38.915 122.920 ;
        RECT 37.775 122.655 38.030 122.750 ;
        RECT 39.175 122.485 39.505 122.885 ;
        RECT 39.675 122.655 39.935 123.595 ;
        RECT 40.110 123.495 40.460 124.145 ;
        RECT 40.630 123.325 40.860 124.315 ;
        RECT 40.195 123.155 40.860 123.325 ;
        RECT 40.195 122.655 40.365 123.155 ;
        RECT 40.535 122.485 40.865 122.985 ;
        RECT 41.035 122.655 41.220 124.775 ;
        RECT 41.475 124.575 41.725 125.035 ;
        RECT 41.895 124.585 42.230 124.755 ;
        RECT 42.425 124.585 43.100 124.755 ;
        RECT 41.895 124.445 42.065 124.585 ;
        RECT 41.390 123.455 41.670 124.405 ;
        RECT 41.840 124.315 42.065 124.445 ;
        RECT 41.840 123.210 42.010 124.315 ;
        RECT 42.235 124.165 42.760 124.385 ;
        RECT 42.180 123.400 42.420 123.995 ;
        RECT 42.590 123.465 42.760 124.165 ;
        RECT 42.930 123.805 43.100 124.585 ;
        RECT 43.420 124.535 43.790 125.035 ;
        RECT 43.970 124.585 44.375 124.755 ;
        RECT 44.545 124.585 45.330 124.755 ;
        RECT 43.970 124.355 44.140 124.585 ;
        RECT 43.310 124.055 44.140 124.355 ;
        RECT 44.525 124.085 44.990 124.415 ;
        RECT 43.310 124.025 43.510 124.055 ;
        RECT 43.630 123.805 43.800 123.875 ;
        RECT 42.930 123.635 43.800 123.805 ;
        RECT 43.290 123.545 43.800 123.635 ;
        RECT 41.840 123.080 42.145 123.210 ;
        RECT 42.590 123.100 43.120 123.465 ;
        RECT 41.460 122.485 41.725 122.945 ;
        RECT 41.895 122.655 42.145 123.080 ;
        RECT 43.290 122.930 43.460 123.545 ;
        RECT 42.355 122.760 43.460 122.930 ;
        RECT 43.630 122.485 43.800 123.285 ;
        RECT 43.970 122.985 44.140 124.055 ;
        RECT 44.310 123.155 44.500 123.875 ;
        RECT 44.670 123.125 44.990 124.085 ;
        RECT 45.160 124.125 45.330 124.585 ;
        RECT 45.605 124.505 45.815 125.035 ;
        RECT 46.075 124.295 46.405 124.820 ;
        RECT 46.575 124.425 46.745 125.035 ;
        RECT 46.915 124.380 47.245 124.815 ;
        RECT 47.465 124.490 52.810 125.035 ;
        RECT 46.915 124.295 47.295 124.380 ;
        RECT 46.205 124.125 46.405 124.295 ;
        RECT 47.070 124.255 47.295 124.295 ;
        RECT 45.160 123.795 46.035 124.125 ;
        RECT 46.205 123.795 46.955 124.125 ;
        RECT 43.970 122.655 44.220 122.985 ;
        RECT 45.160 122.955 45.330 123.795 ;
        RECT 46.205 123.590 46.395 123.795 ;
        RECT 47.125 123.675 47.295 124.255 ;
        RECT 47.080 123.625 47.295 123.675 ;
        RECT 49.050 123.660 49.390 124.490 ;
        RECT 52.985 124.265 56.495 125.035 ;
        RECT 57.125 124.310 57.415 125.035 ;
        RECT 57.585 124.490 62.930 125.035 ;
        RECT 63.105 124.490 68.450 125.035 ;
        RECT 68.625 124.490 73.970 125.035 ;
        RECT 74.145 124.490 79.490 125.035 ;
        RECT 45.500 123.215 46.395 123.590 ;
        RECT 46.905 123.545 47.295 123.625 ;
        RECT 44.445 122.785 45.330 122.955 ;
        RECT 45.510 122.485 45.825 122.985 ;
        RECT 46.055 122.655 46.395 123.215 ;
        RECT 46.565 122.485 46.735 123.495 ;
        RECT 46.905 122.700 47.235 123.545 ;
        RECT 50.870 122.920 51.220 124.170 ;
        RECT 52.985 123.745 54.635 124.265 ;
        RECT 54.805 123.575 56.495 124.095 ;
        RECT 59.170 123.660 59.510 124.490 ;
        RECT 47.465 122.485 52.810 122.920 ;
        RECT 52.985 122.485 56.495 123.575 ;
        RECT 57.125 122.485 57.415 123.650 ;
        RECT 60.990 122.920 61.340 124.170 ;
        RECT 64.690 123.660 65.030 124.490 ;
        RECT 66.510 122.920 66.860 124.170 ;
        RECT 70.210 123.660 70.550 124.490 ;
        RECT 72.030 122.920 72.380 124.170 ;
        RECT 75.730 123.660 76.070 124.490 ;
        RECT 79.665 124.265 82.255 125.035 ;
        RECT 82.885 124.285 84.095 125.035 ;
        RECT 77.550 122.920 77.900 124.170 ;
        RECT 79.665 123.745 80.875 124.265 ;
        RECT 81.045 123.575 82.255 124.095 ;
        RECT 57.585 122.485 62.930 122.920 ;
        RECT 63.105 122.485 68.450 122.920 ;
        RECT 68.625 122.485 73.970 122.920 ;
        RECT 74.145 122.485 79.490 122.920 ;
        RECT 79.665 122.485 82.255 123.575 ;
        RECT 82.885 123.575 83.405 124.115 ;
        RECT 83.575 123.745 84.095 124.285 ;
        RECT 82.885 122.485 84.095 123.575 ;
        RECT 5.520 122.315 84.180 122.485 ;
        RECT 5.605 121.225 6.815 122.315 ;
        RECT 6.985 121.880 12.330 122.315 ;
        RECT 12.505 121.880 17.850 122.315 ;
        RECT 5.605 120.515 6.125 121.055 ;
        RECT 6.295 120.685 6.815 121.225 ;
        RECT 5.605 119.765 6.815 120.515 ;
        RECT 8.570 120.310 8.910 121.140 ;
        RECT 10.390 120.630 10.740 121.880 ;
        RECT 14.090 120.310 14.430 121.140 ;
        RECT 15.910 120.630 16.260 121.880 ;
        RECT 18.485 121.150 18.775 122.315 ;
        RECT 18.945 121.225 20.155 122.315 ;
        RECT 20.440 121.685 20.725 122.145 ;
        RECT 20.895 121.855 21.165 122.315 ;
        RECT 20.440 121.465 21.395 121.685 ;
        RECT 18.945 120.515 19.465 121.055 ;
        RECT 19.635 120.685 20.155 121.225 ;
        RECT 20.325 120.735 21.015 121.295 ;
        RECT 21.185 120.565 21.395 121.465 ;
        RECT 6.985 119.765 12.330 120.310 ;
        RECT 12.505 119.765 17.850 120.310 ;
        RECT 18.485 119.765 18.775 120.490 ;
        RECT 18.945 119.765 20.155 120.515 ;
        RECT 20.440 120.395 21.395 120.565 ;
        RECT 21.565 121.295 21.965 122.145 ;
        RECT 22.155 121.685 22.435 122.145 ;
        RECT 22.955 121.855 23.280 122.315 ;
        RECT 22.155 121.465 23.280 121.685 ;
        RECT 21.565 120.735 22.660 121.295 ;
        RECT 22.830 121.005 23.280 121.465 ;
        RECT 23.450 121.175 23.835 122.145 ;
        RECT 24.005 121.225 26.595 122.315 ;
        RECT 20.440 119.935 20.725 120.395 ;
        RECT 20.895 119.765 21.165 120.225 ;
        RECT 21.565 119.935 21.965 120.735 ;
        RECT 22.830 120.675 23.385 121.005 ;
        RECT 22.830 120.565 23.280 120.675 ;
        RECT 22.155 120.395 23.280 120.565 ;
        RECT 23.555 120.505 23.835 121.175 ;
        RECT 22.155 119.935 22.435 120.395 ;
        RECT 22.955 119.765 23.280 120.225 ;
        RECT 23.450 119.935 23.835 120.505 ;
        RECT 24.005 120.535 25.215 121.055 ;
        RECT 25.385 120.705 26.595 121.225 ;
        RECT 27.225 120.750 27.575 122.145 ;
        RECT 27.745 121.515 28.150 122.315 ;
        RECT 28.320 121.975 29.855 122.145 ;
        RECT 28.320 121.345 28.490 121.975 ;
        RECT 27.745 121.175 28.490 121.345 ;
        RECT 24.005 119.765 26.595 120.535 ;
        RECT 27.225 119.935 27.495 120.750 ;
        RECT 27.745 120.675 27.915 121.175 ;
        RECT 28.660 121.005 28.930 121.750 ;
        RECT 28.085 120.675 28.420 121.005 ;
        RECT 28.590 120.675 28.930 121.005 ;
        RECT 29.120 121.005 29.355 121.750 ;
        RECT 29.525 121.345 29.855 121.975 ;
        RECT 30.040 121.515 30.275 122.315 ;
        RECT 30.445 121.345 30.735 122.145 ;
        RECT 29.525 121.175 30.735 121.345 ;
        RECT 30.905 121.725 31.605 122.145 ;
        RECT 31.805 121.955 32.135 122.315 ;
        RECT 32.305 121.725 32.635 122.125 ;
        RECT 30.905 121.495 32.635 121.725 ;
        RECT 29.120 120.675 29.410 121.005 ;
        RECT 29.580 120.675 29.980 121.005 ;
        RECT 30.150 120.505 30.320 121.175 ;
        RECT 30.490 120.675 30.735 121.005 ;
        RECT 30.905 120.525 31.110 121.495 ;
        RECT 31.280 120.755 31.610 121.295 ;
        RECT 31.785 121.005 32.110 121.295 ;
        RECT 32.305 121.275 32.635 121.495 ;
        RECT 32.805 121.005 32.975 121.975 ;
        RECT 33.155 121.255 33.485 122.315 ;
        RECT 33.755 121.645 33.925 122.145 ;
        RECT 34.095 121.815 34.425 122.315 ;
        RECT 33.755 121.475 34.420 121.645 ;
        RECT 31.785 120.675 32.280 121.005 ;
        RECT 32.600 120.675 32.975 121.005 ;
        RECT 33.185 120.675 33.495 121.005 ;
        RECT 33.670 120.655 34.020 121.305 ;
        RECT 27.665 119.765 28.335 120.505 ;
        RECT 28.505 120.335 29.900 120.505 ;
        RECT 28.505 119.990 28.800 120.335 ;
        RECT 28.980 119.765 29.355 120.165 ;
        RECT 29.570 119.990 29.900 120.335 ;
        RECT 30.150 119.935 30.735 120.505 ;
        RECT 30.905 119.935 31.615 120.525 ;
        RECT 32.125 120.295 33.485 120.505 ;
        RECT 34.190 120.485 34.420 121.475 ;
        RECT 32.125 119.935 32.455 120.295 ;
        RECT 32.655 119.765 32.985 120.125 ;
        RECT 33.155 119.935 33.485 120.295 ;
        RECT 33.755 120.315 34.420 120.485 ;
        RECT 33.755 120.025 33.925 120.315 ;
        RECT 34.095 119.765 34.425 120.145 ;
        RECT 34.595 120.025 34.780 122.145 ;
        RECT 35.020 121.855 35.285 122.315 ;
        RECT 35.455 121.720 35.705 122.145 ;
        RECT 35.915 121.870 37.020 122.040 ;
        RECT 35.400 121.590 35.705 121.720 ;
        RECT 34.950 120.395 35.230 121.345 ;
        RECT 35.400 120.485 35.570 121.590 ;
        RECT 35.740 120.805 35.980 121.400 ;
        RECT 36.150 121.335 36.680 121.700 ;
        RECT 36.150 120.635 36.320 121.335 ;
        RECT 36.850 121.255 37.020 121.870 ;
        RECT 37.190 121.515 37.360 122.315 ;
        RECT 37.530 121.815 37.780 122.145 ;
        RECT 38.005 121.845 38.890 122.015 ;
        RECT 36.850 121.165 37.360 121.255 ;
        RECT 35.400 120.355 35.625 120.485 ;
        RECT 35.795 120.415 36.320 120.635 ;
        RECT 36.490 120.995 37.360 121.165 ;
        RECT 35.035 119.765 35.285 120.225 ;
        RECT 35.455 120.215 35.625 120.355 ;
        RECT 36.490 120.215 36.660 120.995 ;
        RECT 37.190 120.925 37.360 120.995 ;
        RECT 36.870 120.745 37.070 120.775 ;
        RECT 37.530 120.745 37.700 121.815 ;
        RECT 37.870 120.925 38.060 121.645 ;
        RECT 36.870 120.445 37.700 120.745 ;
        RECT 38.230 120.715 38.550 121.675 ;
        RECT 35.455 120.045 35.790 120.215 ;
        RECT 35.985 120.045 36.660 120.215 ;
        RECT 36.980 119.765 37.350 120.265 ;
        RECT 37.530 120.215 37.700 120.445 ;
        RECT 38.085 120.385 38.550 120.715 ;
        RECT 38.720 121.005 38.890 121.845 ;
        RECT 39.070 121.815 39.385 122.315 ;
        RECT 39.615 121.585 39.955 122.145 ;
        RECT 39.060 121.210 39.955 121.585 ;
        RECT 40.125 121.305 40.295 122.315 ;
        RECT 39.765 121.005 39.955 121.210 ;
        RECT 40.465 121.255 40.795 122.100 ;
        RECT 41.025 121.805 42.215 122.095 ;
        RECT 41.045 121.465 42.215 121.635 ;
        RECT 42.385 121.515 42.665 122.315 ;
        RECT 40.465 121.175 40.855 121.255 ;
        RECT 41.045 121.175 41.370 121.465 ;
        RECT 42.045 121.345 42.215 121.465 ;
        RECT 40.640 121.125 40.855 121.175 ;
        RECT 38.720 120.675 39.595 121.005 ;
        RECT 39.765 120.675 40.515 121.005 ;
        RECT 38.720 120.215 38.890 120.675 ;
        RECT 39.765 120.505 39.965 120.675 ;
        RECT 40.685 120.545 40.855 121.125 ;
        RECT 41.540 121.005 41.735 121.295 ;
        RECT 42.045 121.175 42.705 121.345 ;
        RECT 42.875 121.175 43.150 122.145 ;
        RECT 42.535 121.005 42.705 121.175 ;
        RECT 41.025 120.675 41.370 121.005 ;
        RECT 41.540 120.675 42.365 121.005 ;
        RECT 42.535 120.675 42.810 121.005 ;
        RECT 40.630 120.505 40.855 120.545 ;
        RECT 42.535 120.505 42.705 120.675 ;
        RECT 37.530 120.045 37.935 120.215 ;
        RECT 38.105 120.045 38.890 120.215 ;
        RECT 39.165 119.765 39.375 120.295 ;
        RECT 39.635 119.980 39.965 120.505 ;
        RECT 40.475 120.420 40.855 120.505 ;
        RECT 40.135 119.765 40.305 120.375 ;
        RECT 40.475 119.985 40.805 120.420 ;
        RECT 41.040 120.335 42.705 120.505 ;
        RECT 42.980 120.440 43.150 121.175 ;
        RECT 44.245 121.150 44.535 122.315 ;
        RECT 44.705 121.345 45.015 122.145 ;
        RECT 45.185 121.515 45.495 122.315 ;
        RECT 45.665 121.685 45.925 122.145 ;
        RECT 46.095 121.855 46.350 122.315 ;
        RECT 46.525 121.685 46.785 122.145 ;
        RECT 45.665 121.515 46.785 121.685 ;
        RECT 46.145 121.465 46.315 121.515 ;
        RECT 44.705 121.175 45.735 121.345 ;
        RECT 41.040 119.985 41.295 120.335 ;
        RECT 41.465 119.765 41.795 120.165 ;
        RECT 41.965 119.985 42.135 120.335 ;
        RECT 42.305 119.765 42.685 120.165 ;
        RECT 42.875 120.095 43.150 120.440 ;
        RECT 44.245 119.765 44.535 120.490 ;
        RECT 44.705 120.265 44.875 121.175 ;
        RECT 45.045 120.435 45.395 121.005 ;
        RECT 45.565 120.925 45.735 121.175 ;
        RECT 46.525 121.265 46.785 121.515 ;
        RECT 46.955 121.445 47.240 122.315 ;
        RECT 46.525 121.095 47.280 121.265 ;
        RECT 47.465 121.225 49.135 122.315 ;
        RECT 45.565 120.755 46.705 120.925 ;
        RECT 46.875 120.585 47.280 121.095 ;
        RECT 45.630 120.415 47.280 120.585 ;
        RECT 47.465 120.535 48.215 121.055 ;
        RECT 48.385 120.705 49.135 121.225 ;
        RECT 49.305 121.175 49.690 122.145 ;
        RECT 49.860 121.855 50.185 122.315 ;
        RECT 50.705 121.685 50.985 122.145 ;
        RECT 49.860 121.465 50.985 121.685 ;
        RECT 44.705 119.935 45.005 120.265 ;
        RECT 45.175 119.765 45.450 120.245 ;
        RECT 45.630 120.025 45.925 120.415 ;
        RECT 46.095 119.765 46.350 120.245 ;
        RECT 46.525 120.025 46.785 120.415 ;
        RECT 46.955 119.765 47.235 120.245 ;
        RECT 47.465 119.765 49.135 120.535 ;
        RECT 49.305 120.505 49.585 121.175 ;
        RECT 49.860 121.005 50.310 121.465 ;
        RECT 51.175 121.295 51.575 122.145 ;
        RECT 51.975 121.855 52.245 122.315 ;
        RECT 52.415 121.685 52.700 122.145 ;
        RECT 49.755 120.675 50.310 121.005 ;
        RECT 50.480 120.735 51.575 121.295 ;
        RECT 49.860 120.565 50.310 120.675 ;
        RECT 49.305 119.935 49.690 120.505 ;
        RECT 49.860 120.395 50.985 120.565 ;
        RECT 49.860 119.765 50.185 120.225 ;
        RECT 50.705 119.935 50.985 120.395 ;
        RECT 51.175 119.935 51.575 120.735 ;
        RECT 51.745 121.465 52.700 121.685 ;
        RECT 51.745 120.565 51.955 121.465 ;
        RECT 52.125 120.735 52.815 121.295 ;
        RECT 52.985 121.225 54.655 122.315 ;
        RECT 51.745 120.395 52.700 120.565 ;
        RECT 51.975 119.765 52.245 120.225 ;
        RECT 52.415 119.935 52.700 120.395 ;
        RECT 52.985 120.535 53.735 121.055 ;
        RECT 53.905 120.705 54.655 121.225 ;
        RECT 54.825 121.175 55.210 122.145 ;
        RECT 55.380 121.855 55.705 122.315 ;
        RECT 56.225 121.685 56.505 122.145 ;
        RECT 55.380 121.465 56.505 121.685 ;
        RECT 52.985 119.765 54.655 120.535 ;
        RECT 54.825 120.505 55.105 121.175 ;
        RECT 55.380 121.005 55.830 121.465 ;
        RECT 56.695 121.295 57.095 122.145 ;
        RECT 57.495 121.855 57.765 122.315 ;
        RECT 57.935 121.685 58.220 122.145 ;
        RECT 55.275 120.675 55.830 121.005 ;
        RECT 56.000 120.735 57.095 121.295 ;
        RECT 55.380 120.565 55.830 120.675 ;
        RECT 54.825 119.935 55.210 120.505 ;
        RECT 55.380 120.395 56.505 120.565 ;
        RECT 55.380 119.765 55.705 120.225 ;
        RECT 56.225 119.935 56.505 120.395 ;
        RECT 56.695 119.935 57.095 120.735 ;
        RECT 57.265 121.465 58.220 121.685 ;
        RECT 57.265 120.565 57.475 121.465 ;
        RECT 57.645 120.735 58.335 121.295 ;
        RECT 58.505 121.175 58.845 122.145 ;
        RECT 59.015 121.175 59.185 122.315 ;
        RECT 59.455 121.515 59.705 122.315 ;
        RECT 60.350 121.345 60.680 122.145 ;
        RECT 60.980 121.515 61.310 122.315 ;
        RECT 61.480 121.345 61.810 122.145 ;
        RECT 62.185 121.880 67.530 122.315 ;
        RECT 59.375 121.175 61.810 121.345 ;
        RECT 58.505 121.125 58.735 121.175 ;
        RECT 58.505 120.565 58.680 121.125 ;
        RECT 59.375 120.925 59.545 121.175 ;
        RECT 58.850 120.755 59.545 120.925 ;
        RECT 59.720 120.755 60.140 120.955 ;
        RECT 60.310 120.755 60.640 120.955 ;
        RECT 60.810 120.755 61.140 120.955 ;
        RECT 57.265 120.395 58.220 120.565 ;
        RECT 57.495 119.765 57.765 120.225 ;
        RECT 57.935 119.935 58.220 120.395 ;
        RECT 58.505 119.935 58.845 120.565 ;
        RECT 59.015 119.765 59.265 120.565 ;
        RECT 59.455 120.415 60.680 120.585 ;
        RECT 59.455 119.935 59.785 120.415 ;
        RECT 59.955 119.765 60.180 120.225 ;
        RECT 60.350 119.935 60.680 120.415 ;
        RECT 61.310 120.545 61.480 121.175 ;
        RECT 61.665 120.755 62.015 121.005 ;
        RECT 61.310 119.935 61.810 120.545 ;
        RECT 63.770 120.310 64.110 121.140 ;
        RECT 65.590 120.630 65.940 121.880 ;
        RECT 67.705 121.225 69.375 122.315 ;
        RECT 67.705 120.535 68.455 121.055 ;
        RECT 68.625 120.705 69.375 121.225 ;
        RECT 70.005 121.150 70.295 122.315 ;
        RECT 70.465 121.880 75.810 122.315 ;
        RECT 75.985 121.880 81.330 122.315 ;
        RECT 62.185 119.765 67.530 120.310 ;
        RECT 67.705 119.765 69.375 120.535 ;
        RECT 70.005 119.765 70.295 120.490 ;
        RECT 72.050 120.310 72.390 121.140 ;
        RECT 73.870 120.630 74.220 121.880 ;
        RECT 77.570 120.310 77.910 121.140 ;
        RECT 79.390 120.630 79.740 121.880 ;
        RECT 81.505 121.225 82.715 122.315 ;
        RECT 81.505 120.515 82.025 121.055 ;
        RECT 82.195 120.685 82.715 121.225 ;
        RECT 82.885 121.225 84.095 122.315 ;
        RECT 82.885 120.685 83.405 121.225 ;
        RECT 83.575 120.515 84.095 121.055 ;
        RECT 70.465 119.765 75.810 120.310 ;
        RECT 75.985 119.765 81.330 120.310 ;
        RECT 81.505 119.765 82.715 120.515 ;
        RECT 82.885 119.765 84.095 120.515 ;
        RECT 5.520 119.595 84.180 119.765 ;
        RECT 5.605 118.845 6.815 119.595 ;
        RECT 6.985 119.050 12.330 119.595 ;
        RECT 5.605 118.305 6.125 118.845 ;
        RECT 6.295 118.135 6.815 118.675 ;
        RECT 8.570 118.220 8.910 119.050 ;
        RECT 12.505 118.825 15.095 119.595 ;
        RECT 15.355 119.045 15.525 119.335 ;
        RECT 15.695 119.215 16.025 119.595 ;
        RECT 15.355 118.875 16.020 119.045 ;
        RECT 5.605 117.045 6.815 118.135 ;
        RECT 10.390 117.480 10.740 118.730 ;
        RECT 12.505 118.305 13.715 118.825 ;
        RECT 13.885 118.135 15.095 118.655 ;
        RECT 6.985 117.045 12.330 117.480 ;
        RECT 12.505 117.045 15.095 118.135 ;
        RECT 15.270 118.055 15.620 118.705 ;
        RECT 15.790 117.885 16.020 118.875 ;
        RECT 15.355 117.715 16.020 117.885 ;
        RECT 15.355 117.215 15.525 117.715 ;
        RECT 15.695 117.045 16.025 117.545 ;
        RECT 16.195 117.215 16.380 119.335 ;
        RECT 16.635 119.135 16.885 119.595 ;
        RECT 17.055 119.145 17.390 119.315 ;
        RECT 17.585 119.145 18.260 119.315 ;
        RECT 17.055 119.005 17.225 119.145 ;
        RECT 16.550 118.015 16.830 118.965 ;
        RECT 17.000 118.875 17.225 119.005 ;
        RECT 17.000 117.770 17.170 118.875 ;
        RECT 17.395 118.725 17.920 118.945 ;
        RECT 17.340 117.960 17.580 118.555 ;
        RECT 17.750 118.025 17.920 118.725 ;
        RECT 18.090 118.365 18.260 119.145 ;
        RECT 18.580 119.095 18.950 119.595 ;
        RECT 19.130 119.145 19.535 119.315 ;
        RECT 19.705 119.145 20.490 119.315 ;
        RECT 19.130 118.915 19.300 119.145 ;
        RECT 18.470 118.615 19.300 118.915 ;
        RECT 19.685 118.645 20.150 118.975 ;
        RECT 18.470 118.585 18.670 118.615 ;
        RECT 18.790 118.365 18.960 118.435 ;
        RECT 18.090 118.195 18.960 118.365 ;
        RECT 18.450 118.105 18.960 118.195 ;
        RECT 17.000 117.640 17.305 117.770 ;
        RECT 17.750 117.660 18.280 118.025 ;
        RECT 16.620 117.045 16.885 117.505 ;
        RECT 17.055 117.215 17.305 117.640 ;
        RECT 18.450 117.490 18.620 118.105 ;
        RECT 17.515 117.320 18.620 117.490 ;
        RECT 18.790 117.045 18.960 117.845 ;
        RECT 19.130 117.545 19.300 118.615 ;
        RECT 19.470 117.715 19.660 118.435 ;
        RECT 19.830 117.685 20.150 118.645 ;
        RECT 20.320 118.685 20.490 119.145 ;
        RECT 20.765 119.065 20.975 119.595 ;
        RECT 21.235 118.855 21.565 119.380 ;
        RECT 21.735 118.985 21.905 119.595 ;
        RECT 22.075 118.940 22.405 119.375 ;
        RECT 22.625 119.050 27.970 119.595 ;
        RECT 22.075 118.855 22.455 118.940 ;
        RECT 21.365 118.685 21.565 118.855 ;
        RECT 22.230 118.815 22.455 118.855 ;
        RECT 20.320 118.355 21.195 118.685 ;
        RECT 21.365 118.355 22.115 118.685 ;
        RECT 19.130 117.215 19.380 117.545 ;
        RECT 20.320 117.515 20.490 118.355 ;
        RECT 21.365 118.150 21.555 118.355 ;
        RECT 22.285 118.235 22.455 118.815 ;
        RECT 22.240 118.185 22.455 118.235 ;
        RECT 24.210 118.220 24.550 119.050 ;
        RECT 28.145 118.825 30.735 119.595 ;
        RECT 31.365 118.870 31.655 119.595 ;
        RECT 31.825 119.050 37.170 119.595 ;
        RECT 20.660 117.775 21.555 118.150 ;
        RECT 22.065 118.105 22.455 118.185 ;
        RECT 19.605 117.345 20.490 117.515 ;
        RECT 20.670 117.045 20.985 117.545 ;
        RECT 21.215 117.215 21.555 117.775 ;
        RECT 21.725 117.045 21.895 118.055 ;
        RECT 22.065 117.260 22.395 118.105 ;
        RECT 26.030 117.480 26.380 118.730 ;
        RECT 28.145 118.305 29.355 118.825 ;
        RECT 29.525 118.135 30.735 118.655 ;
        RECT 33.410 118.220 33.750 119.050 ;
        RECT 37.380 118.855 37.995 119.425 ;
        RECT 38.165 119.085 38.380 119.595 ;
        RECT 38.610 119.085 38.890 119.415 ;
        RECT 39.070 119.085 39.310 119.595 ;
        RECT 22.625 117.045 27.970 117.480 ;
        RECT 28.145 117.045 30.735 118.135 ;
        RECT 31.365 117.045 31.655 118.210 ;
        RECT 35.230 117.480 35.580 118.730 ;
        RECT 37.380 117.835 37.695 118.855 ;
        RECT 37.865 118.185 38.035 118.685 ;
        RECT 38.285 118.355 38.550 118.915 ;
        RECT 38.720 118.185 38.890 119.085 ;
        RECT 39.060 118.355 39.415 118.915 ;
        RECT 39.705 118.775 39.915 119.595 ;
        RECT 40.085 118.795 40.415 119.425 ;
        RECT 40.085 118.195 40.335 118.795 ;
        RECT 40.585 118.775 40.815 119.595 ;
        RECT 41.035 118.785 41.305 119.595 ;
        RECT 41.475 118.785 41.805 119.425 ;
        RECT 41.975 118.785 42.215 119.595 ;
        RECT 42.405 118.825 45.915 119.595 ;
        RECT 46.085 118.845 47.295 119.595 ;
        RECT 47.555 119.045 47.725 119.335 ;
        RECT 47.895 119.215 48.225 119.595 ;
        RECT 47.555 118.875 48.220 119.045 ;
        RECT 40.505 118.355 40.835 118.605 ;
        RECT 41.025 118.355 41.375 118.605 ;
        RECT 37.865 118.015 39.290 118.185 ;
        RECT 31.825 117.045 37.170 117.480 ;
        RECT 37.380 117.215 37.915 117.835 ;
        RECT 38.085 117.045 38.415 117.845 ;
        RECT 38.900 117.840 39.290 118.015 ;
        RECT 39.705 117.045 39.915 118.185 ;
        RECT 40.085 117.215 40.415 118.195 ;
        RECT 41.545 118.185 41.715 118.785 ;
        RECT 41.885 118.355 42.235 118.605 ;
        RECT 42.405 118.305 44.055 118.825 ;
        RECT 40.585 117.045 40.815 118.185 ;
        RECT 41.035 117.045 41.365 118.185 ;
        RECT 41.545 118.015 42.225 118.185 ;
        RECT 44.225 118.135 45.915 118.655 ;
        RECT 46.085 118.305 46.605 118.845 ;
        RECT 46.775 118.135 47.295 118.675 ;
        RECT 41.895 117.230 42.225 118.015 ;
        RECT 42.405 117.045 45.915 118.135 ;
        RECT 46.085 117.045 47.295 118.135 ;
        RECT 47.470 118.055 47.820 118.705 ;
        RECT 47.990 117.885 48.220 118.875 ;
        RECT 47.555 117.715 48.220 117.885 ;
        RECT 47.555 117.215 47.725 117.715 ;
        RECT 47.895 117.045 48.225 117.545 ;
        RECT 48.395 117.215 48.580 119.335 ;
        RECT 48.835 119.135 49.085 119.595 ;
        RECT 49.255 119.145 49.590 119.315 ;
        RECT 49.785 119.145 50.460 119.315 ;
        RECT 49.255 119.005 49.425 119.145 ;
        RECT 48.750 118.015 49.030 118.965 ;
        RECT 49.200 118.875 49.425 119.005 ;
        RECT 49.200 117.770 49.370 118.875 ;
        RECT 49.595 118.725 50.120 118.945 ;
        RECT 49.540 117.960 49.780 118.555 ;
        RECT 49.950 118.025 50.120 118.725 ;
        RECT 50.290 118.365 50.460 119.145 ;
        RECT 50.780 119.095 51.150 119.595 ;
        RECT 51.330 119.145 51.735 119.315 ;
        RECT 51.905 119.145 52.690 119.315 ;
        RECT 51.330 118.915 51.500 119.145 ;
        RECT 50.670 118.615 51.500 118.915 ;
        RECT 51.885 118.645 52.350 118.975 ;
        RECT 50.670 118.585 50.870 118.615 ;
        RECT 50.990 118.365 51.160 118.435 ;
        RECT 50.290 118.195 51.160 118.365 ;
        RECT 50.650 118.105 51.160 118.195 ;
        RECT 49.200 117.640 49.505 117.770 ;
        RECT 49.950 117.660 50.480 118.025 ;
        RECT 48.820 117.045 49.085 117.505 ;
        RECT 49.255 117.215 49.505 117.640 ;
        RECT 50.650 117.490 50.820 118.105 ;
        RECT 49.715 117.320 50.820 117.490 ;
        RECT 50.990 117.045 51.160 117.845 ;
        RECT 51.330 117.545 51.500 118.615 ;
        RECT 51.670 117.715 51.860 118.435 ;
        RECT 52.030 117.685 52.350 118.645 ;
        RECT 52.520 118.685 52.690 119.145 ;
        RECT 52.965 119.065 53.175 119.595 ;
        RECT 53.435 118.855 53.765 119.380 ;
        RECT 53.935 118.985 54.105 119.595 ;
        RECT 54.275 118.940 54.605 119.375 ;
        RECT 54.275 118.855 54.655 118.940 ;
        RECT 53.565 118.685 53.765 118.855 ;
        RECT 54.430 118.815 54.655 118.855 ;
        RECT 52.520 118.355 53.395 118.685 ;
        RECT 53.565 118.355 54.315 118.685 ;
        RECT 51.330 117.215 51.580 117.545 ;
        RECT 52.520 117.515 52.690 118.355 ;
        RECT 53.565 118.150 53.755 118.355 ;
        RECT 54.485 118.235 54.655 118.815 ;
        RECT 54.845 118.785 55.085 119.595 ;
        RECT 55.255 118.785 55.585 119.425 ;
        RECT 55.755 118.785 56.025 119.595 ;
        RECT 57.125 118.870 57.415 119.595 ;
        RECT 57.585 118.825 59.255 119.595 ;
        RECT 59.475 118.940 59.805 119.375 ;
        RECT 59.975 118.985 60.145 119.595 ;
        RECT 59.425 118.855 59.805 118.940 ;
        RECT 60.315 118.855 60.645 119.380 ;
        RECT 60.905 119.065 61.115 119.595 ;
        RECT 61.390 119.145 62.175 119.315 ;
        RECT 62.345 119.145 62.750 119.315 ;
        RECT 54.825 118.355 55.175 118.605 ;
        RECT 54.440 118.185 54.655 118.235 ;
        RECT 55.345 118.185 55.515 118.785 ;
        RECT 55.685 118.355 56.035 118.605 ;
        RECT 57.585 118.305 58.335 118.825 ;
        RECT 59.425 118.815 59.650 118.855 ;
        RECT 52.860 117.775 53.755 118.150 ;
        RECT 54.265 118.105 54.655 118.185 ;
        RECT 51.805 117.345 52.690 117.515 ;
        RECT 52.870 117.045 53.185 117.545 ;
        RECT 53.415 117.215 53.755 117.775 ;
        RECT 53.925 117.045 54.095 118.055 ;
        RECT 54.265 117.260 54.595 118.105 ;
        RECT 54.835 118.015 55.515 118.185 ;
        RECT 54.835 117.230 55.165 118.015 ;
        RECT 55.695 117.045 56.025 118.185 ;
        RECT 57.125 117.045 57.415 118.210 ;
        RECT 58.505 118.135 59.255 118.655 ;
        RECT 57.585 117.045 59.255 118.135 ;
        RECT 59.425 118.235 59.595 118.815 ;
        RECT 60.315 118.685 60.515 118.855 ;
        RECT 61.390 118.685 61.560 119.145 ;
        RECT 59.765 118.355 60.515 118.685 ;
        RECT 60.685 118.355 61.560 118.685 ;
        RECT 59.425 118.185 59.640 118.235 ;
        RECT 59.425 118.105 59.815 118.185 ;
        RECT 59.485 117.260 59.815 118.105 ;
        RECT 60.325 118.150 60.515 118.355 ;
        RECT 59.985 117.045 60.155 118.055 ;
        RECT 60.325 117.775 61.220 118.150 ;
        RECT 60.325 117.215 60.665 117.775 ;
        RECT 60.895 117.045 61.210 117.545 ;
        RECT 61.390 117.515 61.560 118.355 ;
        RECT 61.730 118.645 62.195 118.975 ;
        RECT 62.580 118.915 62.750 119.145 ;
        RECT 62.930 119.095 63.300 119.595 ;
        RECT 63.620 119.145 64.295 119.315 ;
        RECT 64.490 119.145 64.825 119.315 ;
        RECT 61.730 117.685 62.050 118.645 ;
        RECT 62.580 118.615 63.410 118.915 ;
        RECT 62.220 117.715 62.410 118.435 ;
        RECT 62.580 117.545 62.750 118.615 ;
        RECT 63.210 118.585 63.410 118.615 ;
        RECT 62.920 118.365 63.090 118.435 ;
        RECT 63.620 118.365 63.790 119.145 ;
        RECT 64.655 119.005 64.825 119.145 ;
        RECT 64.995 119.135 65.245 119.595 ;
        RECT 62.920 118.195 63.790 118.365 ;
        RECT 63.960 118.725 64.485 118.945 ;
        RECT 64.655 118.875 64.880 119.005 ;
        RECT 62.920 118.105 63.430 118.195 ;
        RECT 61.390 117.345 62.275 117.515 ;
        RECT 62.500 117.215 62.750 117.545 ;
        RECT 62.920 117.045 63.090 117.845 ;
        RECT 63.260 117.490 63.430 118.105 ;
        RECT 63.960 118.025 64.130 118.725 ;
        RECT 63.600 117.660 64.130 118.025 ;
        RECT 64.300 117.960 64.540 118.555 ;
        RECT 64.710 117.770 64.880 118.875 ;
        RECT 65.050 118.015 65.330 118.965 ;
        RECT 64.575 117.640 64.880 117.770 ;
        RECT 63.260 117.320 64.365 117.490 ;
        RECT 64.575 117.215 64.825 117.640 ;
        RECT 64.995 117.045 65.260 117.505 ;
        RECT 65.500 117.215 65.685 119.335 ;
        RECT 65.855 119.215 66.185 119.595 ;
        RECT 66.355 119.045 66.525 119.335 ;
        RECT 66.785 119.050 72.130 119.595 ;
        RECT 72.305 119.050 77.650 119.595 ;
        RECT 65.860 118.875 66.525 119.045 ;
        RECT 65.860 117.885 66.090 118.875 ;
        RECT 66.260 118.055 66.610 118.705 ;
        RECT 68.370 118.220 68.710 119.050 ;
        RECT 65.860 117.715 66.525 117.885 ;
        RECT 65.855 117.045 66.185 117.545 ;
        RECT 66.355 117.215 66.525 117.715 ;
        RECT 70.190 117.480 70.540 118.730 ;
        RECT 73.890 118.220 74.230 119.050 ;
        RECT 77.825 118.825 81.335 119.595 ;
        RECT 81.505 118.845 82.715 119.595 ;
        RECT 82.885 118.845 84.095 119.595 ;
        RECT 75.710 117.480 76.060 118.730 ;
        RECT 77.825 118.305 79.475 118.825 ;
        RECT 79.645 118.135 81.335 118.655 ;
        RECT 81.505 118.305 82.025 118.845 ;
        RECT 82.195 118.135 82.715 118.675 ;
        RECT 66.785 117.045 72.130 117.480 ;
        RECT 72.305 117.045 77.650 117.480 ;
        RECT 77.825 117.045 81.335 118.135 ;
        RECT 81.505 117.045 82.715 118.135 ;
        RECT 82.885 118.135 83.405 118.675 ;
        RECT 83.575 118.305 84.095 118.845 ;
        RECT 82.885 117.045 84.095 118.135 ;
        RECT 5.520 116.875 84.180 117.045 ;
        RECT 5.605 115.785 6.815 116.875 ;
        RECT 6.985 115.785 8.195 116.875 ;
        RECT 8.425 115.815 8.755 116.660 ;
        RECT 8.925 115.865 9.095 116.875 ;
        RECT 9.265 116.145 9.605 116.705 ;
        RECT 9.835 116.375 10.150 116.875 ;
        RECT 10.330 116.405 11.215 116.575 ;
        RECT 5.605 115.075 6.125 115.615 ;
        RECT 6.295 115.245 6.815 115.785 ;
        RECT 6.985 115.075 7.505 115.615 ;
        RECT 7.675 115.245 8.195 115.785 ;
        RECT 8.365 115.735 8.755 115.815 ;
        RECT 9.265 115.770 10.160 116.145 ;
        RECT 8.365 115.685 8.580 115.735 ;
        RECT 8.365 115.105 8.535 115.685 ;
        RECT 9.265 115.565 9.455 115.770 ;
        RECT 10.330 115.565 10.500 116.405 ;
        RECT 11.440 116.375 11.690 116.705 ;
        RECT 8.705 115.235 9.455 115.565 ;
        RECT 9.625 115.235 10.500 115.565 ;
        RECT 5.605 114.325 6.815 115.075 ;
        RECT 6.985 114.325 8.195 115.075 ;
        RECT 8.365 115.065 8.590 115.105 ;
        RECT 9.255 115.065 9.455 115.235 ;
        RECT 8.365 114.980 8.745 115.065 ;
        RECT 8.415 114.545 8.745 114.980 ;
        RECT 8.915 114.325 9.085 114.935 ;
        RECT 9.255 114.540 9.585 115.065 ;
        RECT 9.845 114.325 10.055 114.855 ;
        RECT 10.330 114.775 10.500 115.235 ;
        RECT 10.670 115.275 10.990 116.235 ;
        RECT 11.160 115.485 11.350 116.205 ;
        RECT 11.520 115.305 11.690 116.375 ;
        RECT 11.860 116.075 12.030 116.875 ;
        RECT 12.200 116.430 13.305 116.600 ;
        RECT 12.200 115.815 12.370 116.430 ;
        RECT 13.515 116.280 13.765 116.705 ;
        RECT 13.935 116.415 14.200 116.875 ;
        RECT 12.540 115.895 13.070 116.260 ;
        RECT 13.515 116.150 13.820 116.280 ;
        RECT 11.860 115.725 12.370 115.815 ;
        RECT 11.860 115.555 12.730 115.725 ;
        RECT 11.860 115.485 12.030 115.555 ;
        RECT 12.150 115.305 12.350 115.335 ;
        RECT 10.670 114.945 11.135 115.275 ;
        RECT 11.520 115.005 12.350 115.305 ;
        RECT 11.520 114.775 11.690 115.005 ;
        RECT 10.330 114.605 11.115 114.775 ;
        RECT 11.285 114.605 11.690 114.775 ;
        RECT 11.870 114.325 12.240 114.825 ;
        RECT 12.560 114.775 12.730 115.555 ;
        RECT 12.900 115.195 13.070 115.895 ;
        RECT 13.240 115.365 13.480 115.960 ;
        RECT 12.900 114.975 13.425 115.195 ;
        RECT 13.650 115.045 13.820 116.150 ;
        RECT 13.595 114.915 13.820 115.045 ;
        RECT 13.990 114.955 14.270 115.905 ;
        RECT 13.595 114.775 13.765 114.915 ;
        RECT 12.560 114.605 13.235 114.775 ;
        RECT 13.430 114.605 13.765 114.775 ;
        RECT 13.935 114.325 14.185 114.785 ;
        RECT 14.440 114.585 14.625 116.705 ;
        RECT 14.795 116.375 15.125 116.875 ;
        RECT 15.295 116.205 15.465 116.705 ;
        RECT 14.800 116.035 15.465 116.205 ;
        RECT 14.800 115.045 15.030 116.035 ;
        RECT 15.200 115.215 15.550 115.865 ;
        RECT 15.725 115.270 16.005 116.705 ;
        RECT 16.175 116.100 16.885 116.875 ;
        RECT 17.055 115.930 17.385 116.705 ;
        RECT 16.235 115.715 17.385 115.930 ;
        RECT 14.800 114.875 15.465 115.045 ;
        RECT 14.795 114.325 15.125 114.705 ;
        RECT 15.295 114.585 15.465 114.875 ;
        RECT 15.725 114.495 16.065 115.270 ;
        RECT 16.235 115.145 16.520 115.715 ;
        RECT 16.705 115.315 17.175 115.545 ;
        RECT 17.580 115.515 17.795 116.630 ;
        RECT 17.975 116.155 18.305 116.875 ;
        RECT 18.085 115.515 18.315 115.855 ;
        RECT 18.485 115.710 18.775 116.875 ;
        RECT 19.035 116.205 19.205 116.705 ;
        RECT 19.375 116.375 19.705 116.875 ;
        RECT 19.035 116.035 19.700 116.205 ;
        RECT 17.345 115.335 17.795 115.515 ;
        RECT 17.345 115.315 17.675 115.335 ;
        RECT 17.985 115.315 18.315 115.515 ;
        RECT 18.950 115.215 19.300 115.865 ;
        RECT 16.235 114.955 16.945 115.145 ;
        RECT 16.645 114.815 16.945 114.955 ;
        RECT 17.135 114.955 18.315 115.145 ;
        RECT 17.135 114.875 17.465 114.955 ;
        RECT 16.645 114.805 16.960 114.815 ;
        RECT 16.645 114.795 16.970 114.805 ;
        RECT 16.645 114.790 16.980 114.795 ;
        RECT 16.235 114.325 16.405 114.785 ;
        RECT 16.645 114.780 16.985 114.790 ;
        RECT 16.645 114.775 16.990 114.780 ;
        RECT 16.645 114.765 16.995 114.775 ;
        RECT 16.645 114.760 17.000 114.765 ;
        RECT 16.645 114.495 17.005 114.760 ;
        RECT 17.635 114.325 17.805 114.785 ;
        RECT 17.975 114.495 18.315 114.955 ;
        RECT 18.485 114.325 18.775 115.050 ;
        RECT 19.470 115.045 19.700 116.035 ;
        RECT 19.035 114.875 19.700 115.045 ;
        RECT 19.035 114.585 19.205 114.875 ;
        RECT 19.375 114.325 19.705 114.705 ;
        RECT 19.875 114.585 20.060 116.705 ;
        RECT 20.300 116.415 20.565 116.875 ;
        RECT 20.735 116.280 20.985 116.705 ;
        RECT 21.195 116.430 22.300 116.600 ;
        RECT 20.680 116.150 20.985 116.280 ;
        RECT 20.230 114.955 20.510 115.905 ;
        RECT 20.680 115.045 20.850 116.150 ;
        RECT 21.020 115.365 21.260 115.960 ;
        RECT 21.430 115.895 21.960 116.260 ;
        RECT 21.430 115.195 21.600 115.895 ;
        RECT 22.130 115.815 22.300 116.430 ;
        RECT 22.470 116.075 22.640 116.875 ;
        RECT 22.810 116.375 23.060 116.705 ;
        RECT 23.285 116.405 24.170 116.575 ;
        RECT 22.130 115.725 22.640 115.815 ;
        RECT 20.680 114.915 20.905 115.045 ;
        RECT 21.075 114.975 21.600 115.195 ;
        RECT 21.770 115.555 22.640 115.725 ;
        RECT 20.315 114.325 20.565 114.785 ;
        RECT 20.735 114.775 20.905 114.915 ;
        RECT 21.770 114.775 21.940 115.555 ;
        RECT 22.470 115.485 22.640 115.555 ;
        RECT 22.150 115.305 22.350 115.335 ;
        RECT 22.810 115.305 22.980 116.375 ;
        RECT 23.150 115.485 23.340 116.205 ;
        RECT 22.150 115.005 22.980 115.305 ;
        RECT 23.510 115.275 23.830 116.235 ;
        RECT 20.735 114.605 21.070 114.775 ;
        RECT 21.265 114.605 21.940 114.775 ;
        RECT 22.260 114.325 22.630 114.825 ;
        RECT 22.810 114.775 22.980 115.005 ;
        RECT 23.365 114.945 23.830 115.275 ;
        RECT 24.000 115.565 24.170 116.405 ;
        RECT 24.350 116.375 24.665 116.875 ;
        RECT 24.895 116.145 25.235 116.705 ;
        RECT 24.340 115.770 25.235 116.145 ;
        RECT 25.405 115.865 25.575 116.875 ;
        RECT 25.045 115.565 25.235 115.770 ;
        RECT 25.745 115.815 26.075 116.660 ;
        RECT 25.745 115.735 26.135 115.815 ;
        RECT 25.920 115.685 26.135 115.735 ;
        RECT 24.000 115.235 24.875 115.565 ;
        RECT 25.045 115.235 25.795 115.565 ;
        RECT 24.000 114.775 24.170 115.235 ;
        RECT 25.045 115.065 25.245 115.235 ;
        RECT 25.965 115.105 26.135 115.685 ;
        RECT 25.910 115.065 26.135 115.105 ;
        RECT 22.810 114.605 23.215 114.775 ;
        RECT 23.385 114.605 24.170 114.775 ;
        RECT 24.445 114.325 24.655 114.855 ;
        RECT 24.915 114.540 25.245 115.065 ;
        RECT 25.755 114.980 26.135 115.065 ;
        RECT 26.305 115.735 26.690 116.705 ;
        RECT 26.860 116.415 27.185 116.875 ;
        RECT 27.705 116.245 27.985 116.705 ;
        RECT 26.860 116.025 27.985 116.245 ;
        RECT 26.305 115.065 26.585 115.735 ;
        RECT 26.860 115.565 27.310 116.025 ;
        RECT 28.175 115.855 28.575 116.705 ;
        RECT 28.975 116.415 29.245 116.875 ;
        RECT 29.415 116.245 29.700 116.705 ;
        RECT 26.755 115.235 27.310 115.565 ;
        RECT 27.480 115.295 28.575 115.855 ;
        RECT 26.860 115.125 27.310 115.235 ;
        RECT 25.415 114.325 25.585 114.935 ;
        RECT 25.755 114.545 26.085 114.980 ;
        RECT 26.305 114.495 26.690 115.065 ;
        RECT 26.860 114.955 27.985 115.125 ;
        RECT 26.860 114.325 27.185 114.785 ;
        RECT 27.705 114.495 27.985 114.955 ;
        RECT 28.175 114.495 28.575 115.295 ;
        RECT 28.745 116.025 29.700 116.245 ;
        RECT 28.745 115.125 28.955 116.025 ;
        RECT 29.125 115.295 29.815 115.855 ;
        RECT 30.445 115.735 30.830 116.705 ;
        RECT 31.000 116.415 31.325 116.875 ;
        RECT 31.845 116.245 32.125 116.705 ;
        RECT 31.000 116.025 32.125 116.245 ;
        RECT 28.745 114.955 29.700 115.125 ;
        RECT 28.975 114.325 29.245 114.785 ;
        RECT 29.415 114.495 29.700 114.955 ;
        RECT 30.445 115.065 30.725 115.735 ;
        RECT 31.000 115.565 31.450 116.025 ;
        RECT 32.315 115.855 32.715 116.705 ;
        RECT 33.115 116.415 33.385 116.875 ;
        RECT 33.555 116.245 33.840 116.705 ;
        RECT 34.125 116.440 39.470 116.875 ;
        RECT 30.895 115.235 31.450 115.565 ;
        RECT 31.620 115.295 32.715 115.855 ;
        RECT 31.000 115.125 31.450 115.235 ;
        RECT 30.445 114.495 30.830 115.065 ;
        RECT 31.000 114.955 32.125 115.125 ;
        RECT 31.000 114.325 31.325 114.785 ;
        RECT 31.845 114.495 32.125 114.955 ;
        RECT 32.315 114.495 32.715 115.295 ;
        RECT 32.885 116.025 33.840 116.245 ;
        RECT 32.885 115.125 33.095 116.025 ;
        RECT 33.265 115.295 33.955 115.855 ;
        RECT 32.885 114.955 33.840 115.125 ;
        RECT 33.115 114.325 33.385 114.785 ;
        RECT 33.555 114.495 33.840 114.955 ;
        RECT 35.710 114.870 36.050 115.700 ;
        RECT 37.530 115.190 37.880 116.440 ;
        RECT 39.645 115.785 43.155 116.875 ;
        RECT 39.645 115.095 41.295 115.615 ;
        RECT 41.465 115.265 43.155 115.785 ;
        RECT 44.245 115.710 44.535 116.875 ;
        RECT 44.795 116.205 44.965 116.705 ;
        RECT 45.135 116.375 45.465 116.875 ;
        RECT 44.795 116.035 45.460 116.205 ;
        RECT 44.710 115.215 45.060 115.865 ;
        RECT 34.125 114.325 39.470 114.870 ;
        RECT 39.645 114.325 43.155 115.095 ;
        RECT 44.245 114.325 44.535 115.050 ;
        RECT 45.230 115.045 45.460 116.035 ;
        RECT 44.795 114.875 45.460 115.045 ;
        RECT 44.795 114.585 44.965 114.875 ;
        RECT 45.135 114.325 45.465 114.705 ;
        RECT 45.635 114.585 45.820 116.705 ;
        RECT 46.060 116.415 46.325 116.875 ;
        RECT 46.495 116.280 46.745 116.705 ;
        RECT 46.955 116.430 48.060 116.600 ;
        RECT 46.440 116.150 46.745 116.280 ;
        RECT 45.990 114.955 46.270 115.905 ;
        RECT 46.440 115.045 46.610 116.150 ;
        RECT 46.780 115.365 47.020 115.960 ;
        RECT 47.190 115.895 47.720 116.260 ;
        RECT 47.190 115.195 47.360 115.895 ;
        RECT 47.890 115.815 48.060 116.430 ;
        RECT 48.230 116.075 48.400 116.875 ;
        RECT 48.570 116.375 48.820 116.705 ;
        RECT 49.045 116.405 49.930 116.575 ;
        RECT 47.890 115.725 48.400 115.815 ;
        RECT 46.440 114.915 46.665 115.045 ;
        RECT 46.835 114.975 47.360 115.195 ;
        RECT 47.530 115.555 48.400 115.725 ;
        RECT 46.075 114.325 46.325 114.785 ;
        RECT 46.495 114.775 46.665 114.915 ;
        RECT 47.530 114.775 47.700 115.555 ;
        RECT 48.230 115.485 48.400 115.555 ;
        RECT 47.910 115.305 48.110 115.335 ;
        RECT 48.570 115.305 48.740 116.375 ;
        RECT 48.910 115.485 49.100 116.205 ;
        RECT 47.910 115.005 48.740 115.305 ;
        RECT 49.270 115.275 49.590 116.235 ;
        RECT 46.495 114.605 46.830 114.775 ;
        RECT 47.025 114.605 47.700 114.775 ;
        RECT 48.020 114.325 48.390 114.825 ;
        RECT 48.570 114.775 48.740 115.005 ;
        RECT 49.125 114.945 49.590 115.275 ;
        RECT 49.760 115.565 49.930 116.405 ;
        RECT 50.110 116.375 50.425 116.875 ;
        RECT 50.655 116.145 50.995 116.705 ;
        RECT 50.100 115.770 50.995 116.145 ;
        RECT 51.165 115.865 51.335 116.875 ;
        RECT 50.805 115.565 50.995 115.770 ;
        RECT 51.505 115.815 51.835 116.660 ;
        RECT 52.615 116.205 52.785 116.705 ;
        RECT 52.955 116.375 53.285 116.875 ;
        RECT 52.615 116.035 53.280 116.205 ;
        RECT 51.505 115.735 51.895 115.815 ;
        RECT 51.680 115.685 51.895 115.735 ;
        RECT 49.760 115.235 50.635 115.565 ;
        RECT 50.805 115.235 51.555 115.565 ;
        RECT 49.760 114.775 49.930 115.235 ;
        RECT 50.805 115.065 51.005 115.235 ;
        RECT 51.725 115.105 51.895 115.685 ;
        RECT 52.530 115.215 52.880 115.865 ;
        RECT 51.670 115.065 51.895 115.105 ;
        RECT 48.570 114.605 48.975 114.775 ;
        RECT 49.145 114.605 49.930 114.775 ;
        RECT 50.205 114.325 50.415 114.855 ;
        RECT 50.675 114.540 51.005 115.065 ;
        RECT 51.515 114.980 51.895 115.065 ;
        RECT 53.050 115.045 53.280 116.035 ;
        RECT 51.175 114.325 51.345 114.935 ;
        RECT 51.515 114.545 51.845 114.980 ;
        RECT 52.615 114.875 53.280 115.045 ;
        RECT 52.615 114.585 52.785 114.875 ;
        RECT 52.955 114.325 53.285 114.705 ;
        RECT 53.455 114.585 53.640 116.705 ;
        RECT 53.880 116.415 54.145 116.875 ;
        RECT 54.315 116.280 54.565 116.705 ;
        RECT 54.775 116.430 55.880 116.600 ;
        RECT 54.260 116.150 54.565 116.280 ;
        RECT 53.810 114.955 54.090 115.905 ;
        RECT 54.260 115.045 54.430 116.150 ;
        RECT 54.600 115.365 54.840 115.960 ;
        RECT 55.010 115.895 55.540 116.260 ;
        RECT 55.010 115.195 55.180 115.895 ;
        RECT 55.710 115.815 55.880 116.430 ;
        RECT 56.050 116.075 56.220 116.875 ;
        RECT 56.390 116.375 56.640 116.705 ;
        RECT 56.865 116.405 57.750 116.575 ;
        RECT 55.710 115.725 56.220 115.815 ;
        RECT 54.260 114.915 54.485 115.045 ;
        RECT 54.655 114.975 55.180 115.195 ;
        RECT 55.350 115.555 56.220 115.725 ;
        RECT 53.895 114.325 54.145 114.785 ;
        RECT 54.315 114.775 54.485 114.915 ;
        RECT 55.350 114.775 55.520 115.555 ;
        RECT 56.050 115.485 56.220 115.555 ;
        RECT 55.730 115.305 55.930 115.335 ;
        RECT 56.390 115.305 56.560 116.375 ;
        RECT 56.730 115.485 56.920 116.205 ;
        RECT 55.730 115.005 56.560 115.305 ;
        RECT 57.090 115.275 57.410 116.235 ;
        RECT 54.315 114.605 54.650 114.775 ;
        RECT 54.845 114.605 55.520 114.775 ;
        RECT 55.840 114.325 56.210 114.825 ;
        RECT 56.390 114.775 56.560 115.005 ;
        RECT 56.945 114.945 57.410 115.275 ;
        RECT 57.580 115.565 57.750 116.405 ;
        RECT 57.930 116.375 58.245 116.875 ;
        RECT 58.475 116.145 58.815 116.705 ;
        RECT 57.920 115.770 58.815 116.145 ;
        RECT 58.985 115.865 59.155 116.875 ;
        RECT 58.625 115.565 58.815 115.770 ;
        RECT 59.325 115.815 59.655 116.660 ;
        RECT 59.325 115.735 59.715 115.815 ;
        RECT 59.500 115.685 59.715 115.735 ;
        RECT 57.580 115.235 58.455 115.565 ;
        RECT 58.625 115.235 59.375 115.565 ;
        RECT 57.580 114.775 57.750 115.235 ;
        RECT 58.625 115.065 58.825 115.235 ;
        RECT 59.545 115.105 59.715 115.685 ;
        RECT 59.490 115.065 59.715 115.105 ;
        RECT 56.390 114.605 56.795 114.775 ;
        RECT 56.965 114.605 57.750 114.775 ;
        RECT 58.025 114.325 58.235 114.855 ;
        RECT 58.495 114.540 58.825 115.065 ;
        RECT 59.335 114.980 59.715 115.065 ;
        RECT 59.885 115.735 60.270 116.705 ;
        RECT 60.440 116.415 60.765 116.875 ;
        RECT 61.285 116.245 61.565 116.705 ;
        RECT 60.440 116.025 61.565 116.245 ;
        RECT 59.885 115.065 60.165 115.735 ;
        RECT 60.440 115.565 60.890 116.025 ;
        RECT 61.755 115.855 62.155 116.705 ;
        RECT 62.555 116.415 62.825 116.875 ;
        RECT 62.995 116.245 63.280 116.705 ;
        RECT 60.335 115.235 60.890 115.565 ;
        RECT 61.060 115.295 62.155 115.855 ;
        RECT 60.440 115.125 60.890 115.235 ;
        RECT 58.995 114.325 59.165 114.935 ;
        RECT 59.335 114.545 59.665 114.980 ;
        RECT 59.885 114.495 60.270 115.065 ;
        RECT 60.440 114.955 61.565 115.125 ;
        RECT 60.440 114.325 60.765 114.785 ;
        RECT 61.285 114.495 61.565 114.955 ;
        RECT 61.755 114.495 62.155 115.295 ;
        RECT 62.325 116.025 63.280 116.245 ;
        RECT 63.570 116.485 63.905 116.705 ;
        RECT 64.910 116.495 65.265 116.875 ;
        RECT 62.325 115.125 62.535 116.025 ;
        RECT 63.570 115.865 63.825 116.485 ;
        RECT 64.075 116.325 64.305 116.365 ;
        RECT 65.435 116.325 65.685 116.705 ;
        RECT 64.075 116.125 65.685 116.325 ;
        RECT 64.075 116.035 64.260 116.125 ;
        RECT 64.850 116.115 65.685 116.125 ;
        RECT 65.935 116.095 66.185 116.875 ;
        RECT 66.355 116.025 66.615 116.705 ;
        RECT 64.415 115.925 64.745 115.955 ;
        RECT 64.415 115.865 66.215 115.925 ;
        RECT 62.705 115.295 63.395 115.855 ;
        RECT 63.570 115.755 66.275 115.865 ;
        RECT 63.570 115.695 64.745 115.755 ;
        RECT 66.075 115.720 66.275 115.755 ;
        RECT 63.565 115.315 64.055 115.515 ;
        RECT 64.245 115.315 64.720 115.525 ;
        RECT 62.325 114.955 63.280 115.125 ;
        RECT 62.555 114.325 62.825 114.785 ;
        RECT 62.995 114.495 63.280 114.955 ;
        RECT 63.570 114.325 64.025 115.090 ;
        RECT 64.500 114.915 64.720 115.315 ;
        RECT 64.965 115.315 65.295 115.525 ;
        RECT 64.965 114.915 65.175 115.315 ;
        RECT 65.465 115.280 65.875 115.585 ;
        RECT 66.105 115.145 66.275 115.720 ;
        RECT 66.005 115.025 66.275 115.145 ;
        RECT 65.430 114.980 66.275 115.025 ;
        RECT 65.430 114.855 66.185 114.980 ;
        RECT 65.430 114.705 65.600 114.855 ;
        RECT 66.445 114.825 66.615 116.025 ;
        RECT 66.785 115.785 69.375 116.875 ;
        RECT 64.300 114.495 65.600 114.705 ;
        RECT 65.855 114.325 66.185 114.685 ;
        RECT 66.355 114.495 66.615 114.825 ;
        RECT 66.785 115.095 67.995 115.615 ;
        RECT 68.165 115.265 69.375 115.785 ;
        RECT 70.005 115.710 70.295 116.875 ;
        RECT 70.465 116.440 75.810 116.875 ;
        RECT 75.985 116.440 81.330 116.875 ;
        RECT 66.785 114.325 69.375 115.095 ;
        RECT 70.005 114.325 70.295 115.050 ;
        RECT 72.050 114.870 72.390 115.700 ;
        RECT 73.870 115.190 74.220 116.440 ;
        RECT 77.570 114.870 77.910 115.700 ;
        RECT 79.390 115.190 79.740 116.440 ;
        RECT 81.505 115.785 82.715 116.875 ;
        RECT 81.505 115.075 82.025 115.615 ;
        RECT 82.195 115.245 82.715 115.785 ;
        RECT 82.885 115.785 84.095 116.875 ;
        RECT 82.885 115.245 83.405 115.785 ;
        RECT 83.575 115.075 84.095 115.615 ;
        RECT 70.465 114.325 75.810 114.870 ;
        RECT 75.985 114.325 81.330 114.870 ;
        RECT 81.505 114.325 82.715 115.075 ;
        RECT 82.885 114.325 84.095 115.075 ;
        RECT 5.520 114.155 84.180 114.325 ;
        RECT 5.605 113.405 6.815 114.155 ;
        RECT 6.985 113.655 7.245 113.985 ;
        RECT 7.455 113.675 7.730 114.155 ;
        RECT 5.605 112.865 6.125 113.405 ;
        RECT 6.295 112.695 6.815 113.235 ;
        RECT 5.605 111.605 6.815 112.695 ;
        RECT 6.985 112.745 7.155 113.655 ;
        RECT 7.940 113.585 8.145 113.985 ;
        RECT 8.315 113.755 8.650 114.155 ;
        RECT 8.825 113.610 14.170 114.155 ;
        RECT 7.325 112.915 7.685 113.495 ;
        RECT 7.940 113.415 8.625 113.585 ;
        RECT 7.865 112.745 8.115 113.245 ;
        RECT 6.985 112.575 8.115 112.745 ;
        RECT 6.985 111.805 7.255 112.575 ;
        RECT 8.285 112.385 8.625 113.415 ;
        RECT 10.410 112.780 10.750 113.610 ;
        RECT 14.345 113.385 16.015 114.155 ;
        RECT 16.210 113.765 16.540 114.155 ;
        RECT 16.710 113.595 16.935 113.975 ;
        RECT 7.425 111.605 7.755 112.385 ;
        RECT 7.960 112.210 8.625 112.385 ;
        RECT 7.960 111.805 8.145 112.210 ;
        RECT 12.230 112.040 12.580 113.290 ;
        RECT 14.345 112.865 15.095 113.385 ;
        RECT 15.265 112.695 16.015 113.215 ;
        RECT 16.195 112.915 16.435 113.565 ;
        RECT 16.605 113.415 16.935 113.595 ;
        RECT 16.605 112.745 16.780 113.415 ;
        RECT 17.135 113.245 17.365 113.865 ;
        RECT 17.545 113.425 17.845 114.155 ;
        RECT 18.025 113.505 18.285 113.985 ;
        RECT 18.455 113.615 18.705 114.155 ;
        RECT 16.950 112.915 17.365 113.245 ;
        RECT 17.545 112.915 17.840 113.245 ;
        RECT 8.315 111.605 8.650 112.030 ;
        RECT 8.825 111.605 14.170 112.040 ;
        RECT 14.345 111.605 16.015 112.695 ;
        RECT 16.195 112.555 16.780 112.745 ;
        RECT 16.195 111.785 16.470 112.555 ;
        RECT 16.950 112.385 17.845 112.715 ;
        RECT 16.640 112.215 17.845 112.385 ;
        RECT 16.640 111.785 16.970 112.215 ;
        RECT 17.140 111.605 17.335 112.045 ;
        RECT 17.515 111.785 17.845 112.215 ;
        RECT 18.025 112.475 18.195 113.505 ;
        RECT 18.875 113.450 19.095 113.935 ;
        RECT 18.365 112.855 18.595 113.250 ;
        RECT 18.765 113.025 19.095 113.450 ;
        RECT 19.265 113.775 20.155 113.945 ;
        RECT 19.265 113.050 19.435 113.775 ;
        RECT 19.605 113.220 20.155 113.605 ;
        RECT 20.325 113.415 20.710 113.985 ;
        RECT 20.880 113.695 21.205 114.155 ;
        RECT 21.725 113.525 22.005 113.985 ;
        RECT 19.265 112.980 20.155 113.050 ;
        RECT 19.260 112.955 20.155 112.980 ;
        RECT 19.250 112.940 20.155 112.955 ;
        RECT 19.245 112.925 20.155 112.940 ;
        RECT 19.235 112.920 20.155 112.925 ;
        RECT 19.230 112.910 20.155 112.920 ;
        RECT 19.225 112.900 20.155 112.910 ;
        RECT 19.215 112.895 20.155 112.900 ;
        RECT 19.205 112.885 20.155 112.895 ;
        RECT 19.195 112.880 20.155 112.885 ;
        RECT 19.195 112.875 19.530 112.880 ;
        RECT 19.180 112.870 19.530 112.875 ;
        RECT 19.165 112.860 19.530 112.870 ;
        RECT 19.140 112.855 19.530 112.860 ;
        RECT 18.365 112.850 19.530 112.855 ;
        RECT 18.365 112.815 19.500 112.850 ;
        RECT 18.365 112.790 19.465 112.815 ;
        RECT 18.365 112.760 19.435 112.790 ;
        RECT 18.365 112.730 19.415 112.760 ;
        RECT 18.365 112.700 19.395 112.730 ;
        RECT 18.365 112.690 19.325 112.700 ;
        RECT 18.365 112.680 19.300 112.690 ;
        RECT 18.365 112.665 19.280 112.680 ;
        RECT 18.365 112.650 19.260 112.665 ;
        RECT 18.470 112.640 19.255 112.650 ;
        RECT 18.470 112.605 19.240 112.640 ;
        RECT 18.025 111.775 18.300 112.475 ;
        RECT 18.470 112.355 19.225 112.605 ;
        RECT 19.395 112.285 19.725 112.530 ;
        RECT 19.895 112.430 20.155 112.880 ;
        RECT 20.325 112.745 20.605 113.415 ;
        RECT 20.880 113.355 22.005 113.525 ;
        RECT 20.880 113.245 21.330 113.355 ;
        RECT 20.775 112.915 21.330 113.245 ;
        RECT 22.195 113.185 22.595 113.985 ;
        RECT 22.995 113.695 23.265 114.155 ;
        RECT 23.435 113.525 23.720 113.985 ;
        RECT 19.540 112.260 19.725 112.285 ;
        RECT 19.540 112.160 20.155 112.260 ;
        RECT 18.470 111.605 18.725 112.150 ;
        RECT 18.895 111.775 19.375 112.115 ;
        RECT 19.550 111.605 20.155 112.160 ;
        RECT 20.325 111.775 20.710 112.745 ;
        RECT 20.880 112.455 21.330 112.915 ;
        RECT 21.500 112.625 22.595 113.185 ;
        RECT 20.880 112.235 22.005 112.455 ;
        RECT 20.880 111.605 21.205 112.065 ;
        RECT 21.725 111.775 22.005 112.235 ;
        RECT 22.195 111.775 22.595 112.625 ;
        RECT 22.765 113.355 23.720 113.525 ;
        RECT 22.765 112.455 22.975 113.355 ;
        RECT 24.025 113.345 24.265 114.155 ;
        RECT 24.435 113.345 24.765 113.985 ;
        RECT 24.935 113.345 25.205 114.155 ;
        RECT 25.385 113.385 27.975 114.155 ;
        RECT 28.155 113.430 28.485 113.940 ;
        RECT 28.655 113.755 28.985 114.155 ;
        RECT 30.035 113.585 30.365 113.925 ;
        RECT 30.535 113.755 30.865 114.155 ;
        RECT 23.145 112.625 23.835 113.185 ;
        RECT 24.005 112.915 24.355 113.165 ;
        RECT 24.525 112.745 24.695 113.345 ;
        RECT 24.865 112.915 25.215 113.165 ;
        RECT 25.385 112.865 26.595 113.385 ;
        RECT 24.015 112.575 24.695 112.745 ;
        RECT 22.765 112.235 23.720 112.455 ;
        RECT 22.995 111.605 23.265 112.065 ;
        RECT 23.435 111.775 23.720 112.235 ;
        RECT 24.015 111.790 24.345 112.575 ;
        RECT 24.875 111.605 25.205 112.745 ;
        RECT 26.765 112.695 27.975 113.215 ;
        RECT 25.385 111.605 27.975 112.695 ;
        RECT 28.155 112.665 28.345 113.430 ;
        RECT 28.655 113.415 31.020 113.585 ;
        RECT 31.365 113.430 31.655 114.155 ;
        RECT 28.655 113.245 28.825 113.415 ;
        RECT 28.515 112.915 28.825 113.245 ;
        RECT 28.995 112.915 29.300 113.245 ;
        RECT 28.155 111.815 28.485 112.665 ;
        RECT 28.655 111.605 28.905 112.745 ;
        RECT 29.085 112.585 29.300 112.915 ;
        RECT 29.475 112.585 29.760 113.245 ;
        RECT 29.955 112.585 30.220 113.245 ;
        RECT 30.435 112.585 30.680 113.245 ;
        RECT 30.850 112.415 31.020 113.415 ;
        RECT 32.285 113.355 32.980 113.985 ;
        RECT 33.185 113.355 33.495 114.155 ;
        RECT 33.780 113.525 34.065 113.985 ;
        RECT 34.235 113.695 34.505 114.155 ;
        RECT 33.780 113.355 34.735 113.525 ;
        RECT 32.305 112.915 32.640 113.165 ;
        RECT 29.095 112.245 30.385 112.415 ;
        RECT 29.095 111.825 29.345 112.245 ;
        RECT 29.575 111.605 29.905 112.075 ;
        RECT 30.135 111.825 30.385 112.245 ;
        RECT 30.565 112.245 31.020 112.415 ;
        RECT 30.565 111.815 30.895 112.245 ;
        RECT 31.365 111.605 31.655 112.770 ;
        RECT 32.810 112.755 32.980 113.355 ;
        RECT 33.150 112.915 33.485 113.185 ;
        RECT 32.285 111.605 32.545 112.745 ;
        RECT 32.715 111.775 33.045 112.755 ;
        RECT 33.215 111.605 33.495 112.745 ;
        RECT 33.665 112.625 34.355 113.185 ;
        RECT 34.525 112.455 34.735 113.355 ;
        RECT 33.780 112.235 34.735 112.455 ;
        RECT 34.905 113.185 35.305 113.985 ;
        RECT 35.495 113.525 35.775 113.985 ;
        RECT 36.295 113.695 36.620 114.155 ;
        RECT 35.495 113.355 36.620 113.525 ;
        RECT 36.790 113.415 37.175 113.985 ;
        RECT 36.170 113.245 36.620 113.355 ;
        RECT 34.905 112.625 36.000 113.185 ;
        RECT 36.170 112.915 36.725 113.245 ;
        RECT 33.780 111.775 34.065 112.235 ;
        RECT 34.235 111.605 34.505 112.065 ;
        RECT 34.905 111.775 35.305 112.625 ;
        RECT 36.170 112.455 36.620 112.915 ;
        RECT 36.895 112.745 37.175 113.415 ;
        RECT 37.345 113.355 37.655 114.155 ;
        RECT 37.860 113.355 38.555 113.985 ;
        RECT 38.725 113.415 39.110 113.985 ;
        RECT 39.280 113.695 39.605 114.155 ;
        RECT 40.125 113.525 40.405 113.985 ;
        RECT 37.355 112.915 37.690 113.185 ;
        RECT 37.860 112.755 38.030 113.355 ;
        RECT 38.200 112.915 38.535 113.165 ;
        RECT 35.495 112.235 36.620 112.455 ;
        RECT 35.495 111.775 35.775 112.235 ;
        RECT 36.295 111.605 36.620 112.065 ;
        RECT 36.790 111.775 37.175 112.745 ;
        RECT 37.345 111.605 37.625 112.745 ;
        RECT 37.795 111.775 38.125 112.755 ;
        RECT 38.725 112.745 39.005 113.415 ;
        RECT 39.280 113.355 40.405 113.525 ;
        RECT 39.280 113.245 39.730 113.355 ;
        RECT 39.175 112.915 39.730 113.245 ;
        RECT 40.595 113.185 40.995 113.985 ;
        RECT 41.395 113.695 41.665 114.155 ;
        RECT 41.835 113.525 42.120 113.985 ;
        RECT 38.295 111.605 38.555 112.745 ;
        RECT 38.725 111.775 39.110 112.745 ;
        RECT 39.280 112.455 39.730 112.915 ;
        RECT 39.900 112.625 40.995 113.185 ;
        RECT 39.280 112.235 40.405 112.455 ;
        RECT 39.280 111.605 39.605 112.065 ;
        RECT 40.125 111.775 40.405 112.235 ;
        RECT 40.595 111.775 40.995 112.625 ;
        RECT 41.165 113.355 42.120 113.525 ;
        RECT 42.495 113.605 42.665 113.895 ;
        RECT 42.835 113.775 43.165 114.155 ;
        RECT 42.495 113.435 43.160 113.605 ;
        RECT 41.165 112.455 41.375 113.355 ;
        RECT 41.545 112.625 42.235 113.185 ;
        RECT 42.410 112.615 42.760 113.265 ;
        RECT 41.165 112.235 42.120 112.455 ;
        RECT 42.930 112.445 43.160 113.435 ;
        RECT 41.395 111.605 41.665 112.065 ;
        RECT 41.835 111.775 42.120 112.235 ;
        RECT 42.495 112.275 43.160 112.445 ;
        RECT 42.495 111.775 42.665 112.275 ;
        RECT 42.835 111.605 43.165 112.105 ;
        RECT 43.335 111.775 43.520 113.895 ;
        RECT 43.775 113.695 44.025 114.155 ;
        RECT 44.195 113.705 44.530 113.875 ;
        RECT 44.725 113.705 45.400 113.875 ;
        RECT 44.195 113.565 44.365 113.705 ;
        RECT 43.690 112.575 43.970 113.525 ;
        RECT 44.140 113.435 44.365 113.565 ;
        RECT 44.140 112.330 44.310 113.435 ;
        RECT 44.535 113.285 45.060 113.505 ;
        RECT 44.480 112.520 44.720 113.115 ;
        RECT 44.890 112.585 45.060 113.285 ;
        RECT 45.230 112.925 45.400 113.705 ;
        RECT 45.720 113.655 46.090 114.155 ;
        RECT 46.270 113.705 46.675 113.875 ;
        RECT 46.845 113.705 47.630 113.875 ;
        RECT 46.270 113.475 46.440 113.705 ;
        RECT 45.610 113.175 46.440 113.475 ;
        RECT 46.825 113.205 47.290 113.535 ;
        RECT 45.610 113.145 45.810 113.175 ;
        RECT 45.930 112.925 46.100 112.995 ;
        RECT 45.230 112.755 46.100 112.925 ;
        RECT 45.590 112.665 46.100 112.755 ;
        RECT 44.140 112.200 44.445 112.330 ;
        RECT 44.890 112.220 45.420 112.585 ;
        RECT 43.760 111.605 44.025 112.065 ;
        RECT 44.195 111.775 44.445 112.200 ;
        RECT 45.590 112.050 45.760 112.665 ;
        RECT 44.655 111.880 45.760 112.050 ;
        RECT 45.930 111.605 46.100 112.405 ;
        RECT 46.270 112.105 46.440 113.175 ;
        RECT 46.610 112.275 46.800 112.995 ;
        RECT 46.970 112.245 47.290 113.205 ;
        RECT 47.460 113.245 47.630 113.705 ;
        RECT 47.905 113.625 48.115 114.155 ;
        RECT 48.375 113.415 48.705 113.940 ;
        RECT 48.875 113.545 49.045 114.155 ;
        RECT 49.215 113.500 49.545 113.935 ;
        RECT 49.765 113.610 55.110 114.155 ;
        RECT 49.215 113.415 49.595 113.500 ;
        RECT 48.505 113.245 48.705 113.415 ;
        RECT 49.370 113.375 49.595 113.415 ;
        RECT 47.460 112.915 48.335 113.245 ;
        RECT 48.505 112.915 49.255 113.245 ;
        RECT 46.270 111.775 46.520 112.105 ;
        RECT 47.460 112.075 47.630 112.915 ;
        RECT 48.505 112.710 48.695 112.915 ;
        RECT 49.425 112.795 49.595 113.375 ;
        RECT 49.380 112.745 49.595 112.795 ;
        RECT 51.350 112.780 51.690 113.610 ;
        RECT 55.285 113.385 56.955 114.155 ;
        RECT 57.125 113.430 57.415 114.155 ;
        RECT 47.800 112.335 48.695 112.710 ;
        RECT 49.205 112.665 49.595 112.745 ;
        RECT 46.745 111.905 47.630 112.075 ;
        RECT 47.810 111.605 48.125 112.105 ;
        RECT 48.355 111.775 48.695 112.335 ;
        RECT 48.865 111.605 49.035 112.615 ;
        RECT 49.205 111.820 49.535 112.665 ;
        RECT 53.170 112.040 53.520 113.290 ;
        RECT 55.285 112.865 56.035 113.385 ;
        RECT 58.045 113.355 58.740 113.985 ;
        RECT 58.945 113.355 59.255 114.155 ;
        RECT 59.425 113.405 60.635 114.155 ;
        RECT 56.205 112.695 56.955 113.215 ;
        RECT 58.065 112.915 58.400 113.165 ;
        RECT 49.765 111.605 55.110 112.040 ;
        RECT 55.285 111.605 56.955 112.695 ;
        RECT 57.125 111.605 57.415 112.770 ;
        RECT 58.570 112.755 58.740 113.355 ;
        RECT 58.910 112.915 59.245 113.185 ;
        RECT 59.425 112.865 59.945 113.405 ;
        RECT 60.825 113.345 61.065 114.155 ;
        RECT 61.235 113.345 61.565 113.985 ;
        RECT 61.735 113.345 62.005 114.155 ;
        RECT 62.185 113.385 63.855 114.155 ;
        RECT 64.490 113.650 64.825 114.155 ;
        RECT 64.995 113.585 65.235 113.960 ;
        RECT 65.515 113.825 65.685 113.970 ;
        RECT 65.515 113.630 65.890 113.825 ;
        RECT 66.250 113.660 66.645 114.155 ;
        RECT 58.045 111.605 58.305 112.745 ;
        RECT 58.475 111.775 58.805 112.755 ;
        RECT 58.975 111.605 59.255 112.745 ;
        RECT 60.115 112.695 60.635 113.235 ;
        RECT 60.805 112.915 61.155 113.165 ;
        RECT 61.325 112.745 61.495 113.345 ;
        RECT 61.665 112.915 62.015 113.165 ;
        RECT 62.185 112.865 62.935 113.385 ;
        RECT 59.425 111.605 60.635 112.695 ;
        RECT 60.815 112.575 61.495 112.745 ;
        RECT 60.815 111.790 61.145 112.575 ;
        RECT 61.675 111.605 62.005 112.745 ;
        RECT 63.105 112.695 63.855 113.215 ;
        RECT 62.185 111.605 63.855 112.695 ;
        RECT 64.545 112.625 64.845 113.475 ;
        RECT 65.015 113.435 65.235 113.585 ;
        RECT 65.015 113.105 65.550 113.435 ;
        RECT 65.720 113.295 65.890 113.630 ;
        RECT 66.815 113.465 67.055 113.985 ;
        RECT 67.245 113.610 72.590 114.155 ;
        RECT 72.765 113.610 78.110 114.155 ;
        RECT 65.015 112.455 65.250 113.105 ;
        RECT 65.720 112.935 66.705 113.295 ;
        RECT 64.575 112.225 65.250 112.455 ;
        RECT 65.420 112.915 66.705 112.935 ;
        RECT 65.420 112.765 66.280 112.915 ;
        RECT 64.575 111.795 64.745 112.225 ;
        RECT 64.915 111.605 65.245 112.055 ;
        RECT 65.420 111.820 65.705 112.765 ;
        RECT 66.880 112.660 67.055 113.465 ;
        RECT 68.830 112.780 69.170 113.610 ;
        RECT 65.880 112.285 66.575 112.595 ;
        RECT 65.885 111.605 66.570 112.075 ;
        RECT 66.750 111.875 67.055 112.660 ;
        RECT 70.650 112.040 71.000 113.290 ;
        RECT 74.350 112.780 74.690 113.610 ;
        RECT 78.285 113.385 80.875 114.155 ;
        RECT 81.135 113.605 81.305 113.985 ;
        RECT 81.520 113.775 81.850 114.155 ;
        RECT 81.135 113.435 81.850 113.605 ;
        RECT 76.170 112.040 76.520 113.290 ;
        RECT 78.285 112.865 79.495 113.385 ;
        RECT 79.665 112.695 80.875 113.215 ;
        RECT 81.045 112.885 81.400 113.255 ;
        RECT 81.680 113.245 81.850 113.435 ;
        RECT 82.020 113.410 82.275 113.985 ;
        RECT 81.680 112.915 81.935 113.245 ;
        RECT 81.680 112.705 81.850 112.915 ;
        RECT 67.245 111.605 72.590 112.040 ;
        RECT 72.765 111.605 78.110 112.040 ;
        RECT 78.285 111.605 80.875 112.695 ;
        RECT 81.135 112.535 81.850 112.705 ;
        RECT 82.105 112.680 82.275 113.410 ;
        RECT 82.450 113.315 82.710 114.155 ;
        RECT 82.885 113.405 84.095 114.155 ;
        RECT 81.135 111.775 81.305 112.535 ;
        RECT 81.520 111.605 81.850 112.365 ;
        RECT 82.020 111.775 82.275 112.680 ;
        RECT 82.450 111.605 82.710 112.755 ;
        RECT 82.885 112.695 83.405 113.235 ;
        RECT 83.575 112.865 84.095 113.405 ;
        RECT 82.885 111.605 84.095 112.695 ;
        RECT 5.520 111.435 84.180 111.605 ;
        RECT 5.605 110.345 6.815 111.435 ;
        RECT 6.985 110.840 7.420 111.265 ;
        RECT 7.590 111.010 7.975 111.435 ;
        RECT 6.985 110.670 7.975 110.840 ;
        RECT 5.605 109.635 6.125 110.175 ;
        RECT 6.295 109.805 6.815 110.345 ;
        RECT 6.985 109.795 7.470 110.500 ;
        RECT 7.640 110.125 7.975 110.670 ;
        RECT 8.145 110.475 8.570 111.265 ;
        RECT 8.740 110.840 9.015 111.265 ;
        RECT 9.185 111.010 9.570 111.435 ;
        RECT 8.740 110.645 9.570 110.840 ;
        RECT 8.145 110.295 9.050 110.475 ;
        RECT 7.640 109.795 8.050 110.125 ;
        RECT 8.220 109.795 9.050 110.295 ;
        RECT 9.220 110.125 9.570 110.645 ;
        RECT 9.740 110.475 9.985 111.265 ;
        RECT 10.175 110.840 10.430 111.265 ;
        RECT 10.600 111.010 10.985 111.435 ;
        RECT 10.175 110.645 10.985 110.840 ;
        RECT 9.740 110.295 10.465 110.475 ;
        RECT 9.220 109.795 9.645 110.125 ;
        RECT 9.815 109.795 10.465 110.295 ;
        RECT 10.635 110.125 10.985 110.645 ;
        RECT 11.155 110.295 11.415 111.265 ;
        RECT 10.635 109.795 11.060 110.125 ;
        RECT 5.605 108.885 6.815 109.635 ;
        RECT 7.640 109.625 7.975 109.795 ;
        RECT 8.220 109.625 8.570 109.795 ;
        RECT 9.220 109.625 9.570 109.795 ;
        RECT 9.815 109.625 9.985 109.795 ;
        RECT 10.635 109.625 10.985 109.795 ;
        RECT 11.230 109.625 11.415 110.295 ;
        RECT 6.985 109.455 7.975 109.625 ;
        RECT 6.985 109.055 7.420 109.455 ;
        RECT 7.590 108.885 7.975 109.285 ;
        RECT 8.145 109.055 8.570 109.625 ;
        RECT 8.760 109.455 9.570 109.625 ;
        RECT 8.760 109.055 9.015 109.455 ;
        RECT 9.185 108.885 9.570 109.285 ;
        RECT 9.740 109.055 9.985 109.625 ;
        RECT 10.175 109.455 10.985 109.625 ;
        RECT 10.175 109.055 10.430 109.455 ;
        RECT 10.600 108.885 10.985 109.285 ;
        RECT 11.155 109.055 11.415 109.625 ;
        RECT 11.585 110.295 11.970 111.265 ;
        RECT 12.140 110.975 12.465 111.435 ;
        RECT 12.985 110.805 13.265 111.265 ;
        RECT 12.140 110.585 13.265 110.805 ;
        RECT 11.585 109.625 11.865 110.295 ;
        RECT 12.140 110.125 12.590 110.585 ;
        RECT 13.455 110.415 13.855 111.265 ;
        RECT 14.255 110.975 14.525 111.435 ;
        RECT 14.695 110.805 14.980 111.265 ;
        RECT 12.035 109.795 12.590 110.125 ;
        RECT 12.760 109.855 13.855 110.415 ;
        RECT 12.140 109.685 12.590 109.795 ;
        RECT 11.585 109.055 11.970 109.625 ;
        RECT 12.140 109.515 13.265 109.685 ;
        RECT 12.140 108.885 12.465 109.345 ;
        RECT 12.985 109.055 13.265 109.515 ;
        RECT 13.455 109.055 13.855 109.855 ;
        RECT 14.025 110.585 14.980 110.805 ;
        RECT 14.025 109.685 14.235 110.585 ;
        RECT 14.405 109.855 15.095 110.415 ;
        RECT 15.265 110.345 17.855 111.435 ;
        RECT 14.025 109.515 14.980 109.685 ;
        RECT 14.255 108.885 14.525 109.345 ;
        RECT 14.695 109.055 14.980 109.515 ;
        RECT 15.265 109.655 16.475 110.175 ;
        RECT 16.645 109.825 17.855 110.345 ;
        RECT 18.485 110.270 18.775 111.435 ;
        RECT 18.945 111.000 24.290 111.435 ;
        RECT 15.265 108.885 17.855 109.655 ;
        RECT 18.485 108.885 18.775 109.610 ;
        RECT 20.530 109.430 20.870 110.260 ;
        RECT 22.350 109.750 22.700 111.000 ;
        RECT 24.465 110.345 26.135 111.435 ;
        RECT 26.855 110.765 27.025 111.265 ;
        RECT 27.195 110.935 27.525 111.435 ;
        RECT 26.855 110.595 27.520 110.765 ;
        RECT 24.465 109.655 25.215 110.175 ;
        RECT 25.385 109.825 26.135 110.345 ;
        RECT 26.770 109.775 27.120 110.425 ;
        RECT 18.945 108.885 24.290 109.430 ;
        RECT 24.465 108.885 26.135 109.655 ;
        RECT 27.290 109.605 27.520 110.595 ;
        RECT 26.855 109.435 27.520 109.605 ;
        RECT 26.855 109.145 27.025 109.435 ;
        RECT 27.195 108.885 27.525 109.265 ;
        RECT 27.695 109.145 27.880 111.265 ;
        RECT 28.120 110.975 28.385 111.435 ;
        RECT 28.555 110.840 28.805 111.265 ;
        RECT 29.015 110.990 30.120 111.160 ;
        RECT 28.500 110.710 28.805 110.840 ;
        RECT 28.050 109.515 28.330 110.465 ;
        RECT 28.500 109.605 28.670 110.710 ;
        RECT 28.840 109.925 29.080 110.520 ;
        RECT 29.250 110.455 29.780 110.820 ;
        RECT 29.250 109.755 29.420 110.455 ;
        RECT 29.950 110.375 30.120 110.990 ;
        RECT 30.290 110.635 30.460 111.435 ;
        RECT 30.630 110.935 30.880 111.265 ;
        RECT 31.105 110.965 31.990 111.135 ;
        RECT 29.950 110.285 30.460 110.375 ;
        RECT 28.500 109.475 28.725 109.605 ;
        RECT 28.895 109.535 29.420 109.755 ;
        RECT 29.590 110.115 30.460 110.285 ;
        RECT 28.135 108.885 28.385 109.345 ;
        RECT 28.555 109.335 28.725 109.475 ;
        RECT 29.590 109.335 29.760 110.115 ;
        RECT 30.290 110.045 30.460 110.115 ;
        RECT 29.970 109.865 30.170 109.895 ;
        RECT 30.630 109.865 30.800 110.935 ;
        RECT 30.970 110.045 31.160 110.765 ;
        RECT 29.970 109.565 30.800 109.865 ;
        RECT 31.330 109.835 31.650 110.795 ;
        RECT 28.555 109.165 28.890 109.335 ;
        RECT 29.085 109.165 29.760 109.335 ;
        RECT 30.080 108.885 30.450 109.385 ;
        RECT 30.630 109.335 30.800 109.565 ;
        RECT 31.185 109.505 31.650 109.835 ;
        RECT 31.820 110.125 31.990 110.965 ;
        RECT 32.170 110.935 32.485 111.435 ;
        RECT 32.715 110.705 33.055 111.265 ;
        RECT 32.160 110.330 33.055 110.705 ;
        RECT 33.225 110.425 33.395 111.435 ;
        RECT 32.865 110.125 33.055 110.330 ;
        RECT 33.565 110.375 33.895 111.220 ;
        RECT 33.565 110.295 33.955 110.375 ;
        RECT 33.740 110.245 33.955 110.295 ;
        RECT 31.820 109.795 32.695 110.125 ;
        RECT 32.865 109.795 33.615 110.125 ;
        RECT 31.820 109.335 31.990 109.795 ;
        RECT 32.865 109.625 33.065 109.795 ;
        RECT 33.785 109.665 33.955 110.245 ;
        RECT 33.730 109.625 33.955 109.665 ;
        RECT 30.630 109.165 31.035 109.335 ;
        RECT 31.205 109.165 31.990 109.335 ;
        RECT 32.265 108.885 32.475 109.415 ;
        RECT 32.735 109.100 33.065 109.625 ;
        RECT 33.575 109.540 33.955 109.625 ;
        RECT 33.235 108.885 33.405 109.495 ;
        RECT 33.575 109.105 33.905 109.540 ;
        RECT 34.135 109.065 34.395 111.255 ;
        RECT 34.565 110.705 34.905 111.435 ;
        RECT 35.085 110.525 35.355 111.255 ;
        RECT 34.585 110.305 35.355 110.525 ;
        RECT 35.535 110.545 35.765 111.255 ;
        RECT 35.935 110.725 36.265 111.435 ;
        RECT 36.435 110.545 36.695 111.255 ;
        RECT 36.975 110.765 37.145 111.265 ;
        RECT 37.315 110.935 37.645 111.435 ;
        RECT 36.975 110.595 37.640 110.765 ;
        RECT 35.535 110.305 36.695 110.545 ;
        RECT 34.585 109.635 34.875 110.305 ;
        RECT 35.055 109.815 35.520 110.125 ;
        RECT 35.700 109.815 36.225 110.125 ;
        RECT 34.585 109.435 35.815 109.635 ;
        RECT 34.655 108.885 35.325 109.255 ;
        RECT 35.505 109.065 35.815 109.435 ;
        RECT 35.995 109.175 36.225 109.815 ;
        RECT 36.405 109.795 36.705 110.125 ;
        RECT 36.890 109.775 37.240 110.425 ;
        RECT 36.405 108.885 36.695 109.615 ;
        RECT 37.410 109.605 37.640 110.595 ;
        RECT 36.975 109.435 37.640 109.605 ;
        RECT 36.975 109.145 37.145 109.435 ;
        RECT 37.315 108.885 37.645 109.265 ;
        RECT 37.815 109.145 38.000 111.265 ;
        RECT 38.240 110.975 38.505 111.435 ;
        RECT 38.675 110.840 38.925 111.265 ;
        RECT 39.135 110.990 40.240 111.160 ;
        RECT 38.620 110.710 38.925 110.840 ;
        RECT 38.170 109.515 38.450 110.465 ;
        RECT 38.620 109.605 38.790 110.710 ;
        RECT 38.960 109.925 39.200 110.520 ;
        RECT 39.370 110.455 39.900 110.820 ;
        RECT 39.370 109.755 39.540 110.455 ;
        RECT 40.070 110.375 40.240 110.990 ;
        RECT 40.410 110.635 40.580 111.435 ;
        RECT 40.750 110.935 41.000 111.265 ;
        RECT 41.225 110.965 42.110 111.135 ;
        RECT 40.070 110.285 40.580 110.375 ;
        RECT 38.620 109.475 38.845 109.605 ;
        RECT 39.015 109.535 39.540 109.755 ;
        RECT 39.710 110.115 40.580 110.285 ;
        RECT 38.255 108.885 38.505 109.345 ;
        RECT 38.675 109.335 38.845 109.475 ;
        RECT 39.710 109.335 39.880 110.115 ;
        RECT 40.410 110.045 40.580 110.115 ;
        RECT 40.090 109.865 40.290 109.895 ;
        RECT 40.750 109.865 40.920 110.935 ;
        RECT 41.090 110.045 41.280 110.765 ;
        RECT 40.090 109.565 40.920 109.865 ;
        RECT 41.450 109.835 41.770 110.795 ;
        RECT 38.675 109.165 39.010 109.335 ;
        RECT 39.205 109.165 39.880 109.335 ;
        RECT 40.200 108.885 40.570 109.385 ;
        RECT 40.750 109.335 40.920 109.565 ;
        RECT 41.305 109.505 41.770 109.835 ;
        RECT 41.940 110.125 42.110 110.965 ;
        RECT 42.290 110.935 42.605 111.435 ;
        RECT 42.835 110.705 43.175 111.265 ;
        RECT 42.280 110.330 43.175 110.705 ;
        RECT 43.345 110.425 43.515 111.435 ;
        RECT 42.985 110.125 43.175 110.330 ;
        RECT 43.685 110.375 44.015 111.220 ;
        RECT 43.685 110.295 44.075 110.375 ;
        RECT 43.860 110.245 44.075 110.295 ;
        RECT 44.245 110.270 44.535 111.435 ;
        RECT 44.705 110.345 47.295 111.435 ;
        RECT 47.465 110.925 47.725 111.435 ;
        RECT 41.940 109.795 42.815 110.125 ;
        RECT 42.985 109.795 43.735 110.125 ;
        RECT 41.940 109.335 42.110 109.795 ;
        RECT 42.985 109.625 43.185 109.795 ;
        RECT 43.905 109.665 44.075 110.245 ;
        RECT 43.850 109.625 44.075 109.665 ;
        RECT 40.750 109.165 41.155 109.335 ;
        RECT 41.325 109.165 42.110 109.335 ;
        RECT 42.385 108.885 42.595 109.415 ;
        RECT 42.855 109.100 43.185 109.625 ;
        RECT 43.695 109.540 44.075 109.625 ;
        RECT 44.705 109.655 45.915 110.175 ;
        RECT 46.085 109.825 47.295 110.345 ;
        RECT 47.465 109.875 47.805 110.755 ;
        RECT 47.975 110.045 48.145 111.265 ;
        RECT 48.385 110.930 49.000 111.435 ;
        RECT 48.385 110.395 48.635 110.760 ;
        RECT 48.805 110.755 49.000 110.930 ;
        RECT 49.170 110.925 49.645 111.265 ;
        RECT 49.815 110.890 50.030 111.435 ;
        RECT 48.805 110.565 49.135 110.755 ;
        RECT 49.355 110.395 50.070 110.690 ;
        RECT 50.240 110.565 50.515 111.265 ;
        RECT 50.775 110.765 50.945 111.265 ;
        RECT 51.115 110.935 51.445 111.435 ;
        RECT 50.775 110.595 51.440 110.765 ;
        RECT 48.385 110.225 50.175 110.395 ;
        RECT 47.975 109.795 48.770 110.045 ;
        RECT 47.975 109.705 48.225 109.795 ;
        RECT 43.355 108.885 43.525 109.495 ;
        RECT 43.695 109.105 44.025 109.540 ;
        RECT 44.245 108.885 44.535 109.610 ;
        RECT 44.705 108.885 47.295 109.655 ;
        RECT 47.465 108.885 47.725 109.705 ;
        RECT 47.895 109.285 48.225 109.705 ;
        RECT 48.940 109.370 49.195 110.225 ;
        RECT 48.405 109.105 49.195 109.370 ;
        RECT 49.365 109.525 49.775 110.045 ;
        RECT 49.945 109.795 50.175 110.225 ;
        RECT 50.345 109.535 50.515 110.565 ;
        RECT 50.690 109.775 51.040 110.425 ;
        RECT 51.210 109.605 51.440 110.595 ;
        RECT 49.365 109.105 49.565 109.525 ;
        RECT 49.755 108.885 50.085 109.345 ;
        RECT 50.255 109.055 50.515 109.535 ;
        RECT 50.775 109.435 51.440 109.605 ;
        RECT 50.775 109.145 50.945 109.435 ;
        RECT 51.115 108.885 51.445 109.265 ;
        RECT 51.615 109.145 51.800 111.265 ;
        RECT 52.040 110.975 52.305 111.435 ;
        RECT 52.475 110.840 52.725 111.265 ;
        RECT 52.935 110.990 54.040 111.160 ;
        RECT 52.420 110.710 52.725 110.840 ;
        RECT 51.970 109.515 52.250 110.465 ;
        RECT 52.420 109.605 52.590 110.710 ;
        RECT 52.760 109.925 53.000 110.520 ;
        RECT 53.170 110.455 53.700 110.820 ;
        RECT 53.170 109.755 53.340 110.455 ;
        RECT 53.870 110.375 54.040 110.990 ;
        RECT 54.210 110.635 54.380 111.435 ;
        RECT 54.550 110.935 54.800 111.265 ;
        RECT 55.025 110.965 55.910 111.135 ;
        RECT 53.870 110.285 54.380 110.375 ;
        RECT 52.420 109.475 52.645 109.605 ;
        RECT 52.815 109.535 53.340 109.755 ;
        RECT 53.510 110.115 54.380 110.285 ;
        RECT 52.055 108.885 52.305 109.345 ;
        RECT 52.475 109.335 52.645 109.475 ;
        RECT 53.510 109.335 53.680 110.115 ;
        RECT 54.210 110.045 54.380 110.115 ;
        RECT 53.890 109.865 54.090 109.895 ;
        RECT 54.550 109.865 54.720 110.935 ;
        RECT 54.890 110.045 55.080 110.765 ;
        RECT 53.890 109.565 54.720 109.865 ;
        RECT 55.250 109.835 55.570 110.795 ;
        RECT 52.475 109.165 52.810 109.335 ;
        RECT 53.005 109.165 53.680 109.335 ;
        RECT 54.000 108.885 54.370 109.385 ;
        RECT 54.550 109.335 54.720 109.565 ;
        RECT 55.105 109.505 55.570 109.835 ;
        RECT 55.740 110.125 55.910 110.965 ;
        RECT 56.090 110.935 56.405 111.435 ;
        RECT 56.635 110.705 56.975 111.265 ;
        RECT 56.080 110.330 56.975 110.705 ;
        RECT 57.145 110.425 57.315 111.435 ;
        RECT 56.785 110.125 56.975 110.330 ;
        RECT 57.485 110.375 57.815 111.220 ;
        RECT 58.055 110.465 58.385 111.250 ;
        RECT 57.485 110.295 57.875 110.375 ;
        RECT 58.055 110.295 58.735 110.465 ;
        RECT 58.915 110.295 59.245 111.435 ;
        RECT 59.425 110.345 60.635 111.435 ;
        RECT 57.660 110.245 57.875 110.295 ;
        RECT 55.740 109.795 56.615 110.125 ;
        RECT 56.785 109.795 57.535 110.125 ;
        RECT 55.740 109.335 55.910 109.795 ;
        RECT 56.785 109.625 56.985 109.795 ;
        RECT 57.705 109.665 57.875 110.245 ;
        RECT 58.045 109.875 58.395 110.125 ;
        RECT 58.565 109.695 58.735 110.295 ;
        RECT 58.905 109.875 59.255 110.125 ;
        RECT 57.650 109.625 57.875 109.665 ;
        RECT 54.550 109.165 54.955 109.335 ;
        RECT 55.125 109.165 55.910 109.335 ;
        RECT 56.185 108.885 56.395 109.415 ;
        RECT 56.655 109.100 56.985 109.625 ;
        RECT 57.495 109.540 57.875 109.625 ;
        RECT 57.155 108.885 57.325 109.495 ;
        RECT 57.495 109.105 57.825 109.540 ;
        RECT 58.065 108.885 58.305 109.695 ;
        RECT 58.475 109.055 58.805 109.695 ;
        RECT 58.975 108.885 59.245 109.695 ;
        RECT 59.425 109.635 59.945 110.175 ;
        RECT 60.115 109.805 60.635 110.345 ;
        RECT 60.865 110.295 61.075 111.435 ;
        RECT 61.245 110.285 61.575 111.265 ;
        RECT 61.745 110.295 61.975 111.435 ;
        RECT 62.245 110.375 62.575 111.220 ;
        RECT 62.745 110.425 62.915 111.435 ;
        RECT 63.085 110.705 63.425 111.265 ;
        RECT 63.655 110.935 63.970 111.435 ;
        RECT 64.150 110.965 65.035 111.135 ;
        RECT 62.185 110.295 62.575 110.375 ;
        RECT 63.085 110.330 63.980 110.705 ;
        RECT 59.425 108.885 60.635 109.635 ;
        RECT 60.865 108.885 61.075 109.705 ;
        RECT 61.245 109.685 61.495 110.285 ;
        RECT 62.185 110.245 62.400 110.295 ;
        RECT 61.665 109.875 61.995 110.125 ;
        RECT 61.245 109.055 61.575 109.685 ;
        RECT 61.745 108.885 61.975 109.705 ;
        RECT 62.185 109.665 62.355 110.245 ;
        RECT 63.085 110.125 63.275 110.330 ;
        RECT 64.150 110.125 64.320 110.965 ;
        RECT 65.260 110.935 65.510 111.265 ;
        RECT 62.525 109.795 63.275 110.125 ;
        RECT 63.445 109.795 64.320 110.125 ;
        RECT 62.185 109.625 62.410 109.665 ;
        RECT 63.075 109.625 63.275 109.795 ;
        RECT 62.185 109.540 62.565 109.625 ;
        RECT 62.235 109.105 62.565 109.540 ;
        RECT 62.735 108.885 62.905 109.495 ;
        RECT 63.075 109.100 63.405 109.625 ;
        RECT 63.665 108.885 63.875 109.415 ;
        RECT 64.150 109.335 64.320 109.795 ;
        RECT 64.490 109.835 64.810 110.795 ;
        RECT 64.980 110.045 65.170 110.765 ;
        RECT 65.340 109.865 65.510 110.935 ;
        RECT 65.680 110.635 65.850 111.435 ;
        RECT 66.020 110.990 67.125 111.160 ;
        RECT 66.020 110.375 66.190 110.990 ;
        RECT 67.335 110.840 67.585 111.265 ;
        RECT 67.755 110.975 68.020 111.435 ;
        RECT 66.360 110.455 66.890 110.820 ;
        RECT 67.335 110.710 67.640 110.840 ;
        RECT 65.680 110.285 66.190 110.375 ;
        RECT 65.680 110.115 66.550 110.285 ;
        RECT 65.680 110.045 65.850 110.115 ;
        RECT 65.970 109.865 66.170 109.895 ;
        RECT 64.490 109.505 64.955 109.835 ;
        RECT 65.340 109.565 66.170 109.865 ;
        RECT 65.340 109.335 65.510 109.565 ;
        RECT 64.150 109.165 64.935 109.335 ;
        RECT 65.105 109.165 65.510 109.335 ;
        RECT 65.690 108.885 66.060 109.385 ;
        RECT 66.380 109.335 66.550 110.115 ;
        RECT 66.720 109.755 66.890 110.455 ;
        RECT 67.060 109.925 67.300 110.520 ;
        RECT 66.720 109.535 67.245 109.755 ;
        RECT 67.470 109.605 67.640 110.710 ;
        RECT 67.415 109.475 67.640 109.605 ;
        RECT 67.810 109.515 68.090 110.465 ;
        RECT 67.415 109.335 67.585 109.475 ;
        RECT 66.380 109.165 67.055 109.335 ;
        RECT 67.250 109.165 67.585 109.335 ;
        RECT 67.755 108.885 68.005 109.345 ;
        RECT 68.260 109.145 68.445 111.265 ;
        RECT 68.615 110.935 68.945 111.435 ;
        RECT 69.115 110.765 69.285 111.265 ;
        RECT 68.620 110.595 69.285 110.765 ;
        RECT 68.620 109.605 68.850 110.595 ;
        RECT 69.020 109.775 69.370 110.425 ;
        RECT 70.005 110.270 70.295 111.435 ;
        RECT 70.465 111.000 75.810 111.435 ;
        RECT 68.620 109.435 69.285 109.605 ;
        RECT 68.615 108.885 68.945 109.265 ;
        RECT 69.115 109.145 69.285 109.435 ;
        RECT 70.005 108.885 70.295 109.610 ;
        RECT 72.050 109.430 72.390 110.260 ;
        RECT 73.870 109.750 74.220 111.000 ;
        RECT 75.985 110.345 79.495 111.435 ;
        RECT 75.985 109.655 77.635 110.175 ;
        RECT 77.805 109.825 79.495 110.345 ;
        RECT 79.755 110.505 79.925 111.265 ;
        RECT 80.105 110.675 80.435 111.435 ;
        RECT 79.755 110.335 80.420 110.505 ;
        RECT 80.605 110.360 80.875 111.265 ;
        RECT 80.250 110.190 80.420 110.335 ;
        RECT 79.685 109.785 80.015 110.155 ;
        RECT 80.250 109.860 80.535 110.190 ;
        RECT 70.465 108.885 75.810 109.430 ;
        RECT 75.985 108.885 79.495 109.655 ;
        RECT 80.250 109.605 80.420 109.860 ;
        RECT 79.755 109.435 80.420 109.605 ;
        RECT 80.705 109.560 80.875 110.360 ;
        RECT 81.135 110.505 81.305 111.265 ;
        RECT 81.520 110.675 81.850 111.435 ;
        RECT 81.135 110.335 81.850 110.505 ;
        RECT 82.020 110.360 82.275 111.265 ;
        RECT 81.045 109.785 81.400 110.155 ;
        RECT 81.680 110.125 81.850 110.335 ;
        RECT 81.680 109.795 81.935 110.125 ;
        RECT 81.680 109.605 81.850 109.795 ;
        RECT 82.105 109.630 82.275 110.360 ;
        RECT 82.450 110.285 82.710 111.435 ;
        RECT 82.885 110.345 84.095 111.435 ;
        RECT 82.885 109.805 83.405 110.345 ;
        RECT 79.755 109.055 79.925 109.435 ;
        RECT 80.105 108.885 80.435 109.265 ;
        RECT 80.615 109.055 80.875 109.560 ;
        RECT 81.135 109.435 81.850 109.605 ;
        RECT 81.135 109.055 81.305 109.435 ;
        RECT 81.520 108.885 81.850 109.265 ;
        RECT 82.020 109.055 82.275 109.630 ;
        RECT 82.450 108.885 82.710 109.725 ;
        RECT 83.575 109.635 84.095 110.175 ;
        RECT 82.885 108.885 84.095 109.635 ;
        RECT 5.520 108.715 84.180 108.885 ;
        RECT 5.605 107.965 6.815 108.715 ;
        RECT 6.985 107.965 8.195 108.715 ;
        RECT 8.370 108.185 8.660 108.535 ;
        RECT 8.855 108.355 9.185 108.715 ;
        RECT 9.355 108.185 9.585 108.490 ;
        RECT 8.370 108.015 9.585 108.185 ;
        RECT 5.605 107.425 6.125 107.965 ;
        RECT 6.295 107.255 6.815 107.795 ;
        RECT 6.985 107.425 7.505 107.965 ;
        RECT 9.775 107.845 9.945 108.410 ;
        RECT 10.320 108.085 10.605 108.545 ;
        RECT 10.775 108.255 11.045 108.715 ;
        RECT 10.320 107.915 11.275 108.085 ;
        RECT 7.675 107.255 8.195 107.795 ;
        RECT 8.430 107.695 8.690 107.805 ;
        RECT 8.425 107.525 8.690 107.695 ;
        RECT 8.430 107.475 8.690 107.525 ;
        RECT 8.870 107.475 9.255 107.805 ;
        RECT 9.425 107.675 9.945 107.845 ;
        RECT 5.605 106.165 6.815 107.255 ;
        RECT 6.985 106.165 8.195 107.255 ;
        RECT 8.370 106.165 8.690 107.305 ;
        RECT 8.870 106.425 9.065 107.475 ;
        RECT 9.425 107.295 9.595 107.675 ;
        RECT 9.245 107.015 9.595 107.295 ;
        RECT 9.785 107.145 10.030 107.505 ;
        RECT 10.205 107.185 10.895 107.745 ;
        RECT 11.065 107.015 11.275 107.915 ;
        RECT 9.245 106.335 9.575 107.015 ;
        RECT 9.775 106.165 10.030 106.965 ;
        RECT 10.320 106.795 11.275 107.015 ;
        RECT 11.445 107.745 11.845 108.545 ;
        RECT 12.035 108.085 12.315 108.545 ;
        RECT 12.835 108.255 13.160 108.715 ;
        RECT 12.035 107.915 13.160 108.085 ;
        RECT 13.330 107.975 13.715 108.545 ;
        RECT 13.975 108.165 14.145 108.455 ;
        RECT 14.315 108.335 14.645 108.715 ;
        RECT 13.975 107.995 14.640 108.165 ;
        RECT 12.710 107.805 13.160 107.915 ;
        RECT 11.445 107.185 12.540 107.745 ;
        RECT 12.710 107.475 13.265 107.805 ;
        RECT 10.320 106.335 10.605 106.795 ;
        RECT 10.775 106.165 11.045 106.625 ;
        RECT 11.445 106.335 11.845 107.185 ;
        RECT 12.710 107.015 13.160 107.475 ;
        RECT 13.435 107.305 13.715 107.975 ;
        RECT 12.035 106.795 13.160 107.015 ;
        RECT 12.035 106.335 12.315 106.795 ;
        RECT 12.835 106.165 13.160 106.625 ;
        RECT 13.330 106.335 13.715 107.305 ;
        RECT 13.890 107.175 14.240 107.825 ;
        RECT 14.410 107.005 14.640 107.995 ;
        RECT 13.975 106.835 14.640 107.005 ;
        RECT 13.975 106.335 14.145 106.835 ;
        RECT 14.315 106.165 14.645 106.665 ;
        RECT 14.815 106.335 15.000 108.455 ;
        RECT 15.255 108.255 15.505 108.715 ;
        RECT 15.675 108.265 16.010 108.435 ;
        RECT 16.205 108.265 16.880 108.435 ;
        RECT 15.675 108.125 15.845 108.265 ;
        RECT 15.170 107.135 15.450 108.085 ;
        RECT 15.620 107.995 15.845 108.125 ;
        RECT 15.620 106.890 15.790 107.995 ;
        RECT 16.015 107.845 16.540 108.065 ;
        RECT 15.960 107.080 16.200 107.675 ;
        RECT 16.370 107.145 16.540 107.845 ;
        RECT 16.710 107.485 16.880 108.265 ;
        RECT 17.200 108.215 17.570 108.715 ;
        RECT 17.750 108.265 18.155 108.435 ;
        RECT 18.325 108.265 19.110 108.435 ;
        RECT 17.750 108.035 17.920 108.265 ;
        RECT 17.090 107.735 17.920 108.035 ;
        RECT 18.305 107.765 18.770 108.095 ;
        RECT 17.090 107.705 17.290 107.735 ;
        RECT 17.410 107.485 17.580 107.555 ;
        RECT 16.710 107.315 17.580 107.485 ;
        RECT 17.070 107.225 17.580 107.315 ;
        RECT 15.620 106.760 15.925 106.890 ;
        RECT 16.370 106.780 16.900 107.145 ;
        RECT 15.240 106.165 15.505 106.625 ;
        RECT 15.675 106.335 15.925 106.760 ;
        RECT 17.070 106.610 17.240 107.225 ;
        RECT 16.135 106.440 17.240 106.610 ;
        RECT 17.410 106.165 17.580 106.965 ;
        RECT 17.750 106.665 17.920 107.735 ;
        RECT 18.090 106.835 18.280 107.555 ;
        RECT 18.450 106.805 18.770 107.765 ;
        RECT 18.940 107.805 19.110 108.265 ;
        RECT 19.385 108.185 19.595 108.715 ;
        RECT 19.855 107.975 20.185 108.500 ;
        RECT 20.355 108.105 20.525 108.715 ;
        RECT 20.695 108.060 21.025 108.495 ;
        RECT 20.695 107.975 21.075 108.060 ;
        RECT 19.985 107.805 20.185 107.975 ;
        RECT 20.850 107.935 21.075 107.975 ;
        RECT 18.940 107.475 19.815 107.805 ;
        RECT 19.985 107.475 20.735 107.805 ;
        RECT 17.750 106.335 18.000 106.665 ;
        RECT 18.940 106.635 19.110 107.475 ;
        RECT 19.985 107.270 20.175 107.475 ;
        RECT 20.905 107.355 21.075 107.935 ;
        RECT 21.265 107.905 21.505 108.715 ;
        RECT 21.675 107.905 22.005 108.545 ;
        RECT 22.175 107.905 22.445 108.715 ;
        RECT 23.635 108.165 23.805 108.455 ;
        RECT 23.975 108.335 24.305 108.715 ;
        RECT 23.635 107.995 24.300 108.165 ;
        RECT 21.245 107.475 21.595 107.725 ;
        RECT 20.860 107.305 21.075 107.355 ;
        RECT 21.765 107.305 21.935 107.905 ;
        RECT 22.105 107.475 22.455 107.725 ;
        RECT 19.280 106.895 20.175 107.270 ;
        RECT 20.685 107.225 21.075 107.305 ;
        RECT 18.225 106.465 19.110 106.635 ;
        RECT 19.290 106.165 19.605 106.665 ;
        RECT 19.835 106.335 20.175 106.895 ;
        RECT 20.345 106.165 20.515 107.175 ;
        RECT 20.685 106.380 21.015 107.225 ;
        RECT 21.255 107.135 21.935 107.305 ;
        RECT 21.255 106.350 21.585 107.135 ;
        RECT 22.115 106.165 22.445 107.305 ;
        RECT 23.550 107.175 23.900 107.825 ;
        RECT 24.070 107.005 24.300 107.995 ;
        RECT 23.635 106.835 24.300 107.005 ;
        RECT 23.635 106.335 23.805 106.835 ;
        RECT 23.975 106.165 24.305 106.665 ;
        RECT 24.475 106.335 24.660 108.455 ;
        RECT 24.915 108.255 25.165 108.715 ;
        RECT 25.335 108.265 25.670 108.435 ;
        RECT 25.865 108.265 26.540 108.435 ;
        RECT 25.335 108.125 25.505 108.265 ;
        RECT 24.830 107.135 25.110 108.085 ;
        RECT 25.280 107.995 25.505 108.125 ;
        RECT 25.280 106.890 25.450 107.995 ;
        RECT 25.675 107.845 26.200 108.065 ;
        RECT 25.620 107.080 25.860 107.675 ;
        RECT 26.030 107.145 26.200 107.845 ;
        RECT 26.370 107.485 26.540 108.265 ;
        RECT 26.860 108.215 27.230 108.715 ;
        RECT 27.410 108.265 27.815 108.435 ;
        RECT 27.985 108.265 28.770 108.435 ;
        RECT 27.410 108.035 27.580 108.265 ;
        RECT 26.750 107.735 27.580 108.035 ;
        RECT 27.965 107.765 28.430 108.095 ;
        RECT 26.750 107.705 26.950 107.735 ;
        RECT 27.070 107.485 27.240 107.555 ;
        RECT 26.370 107.315 27.240 107.485 ;
        RECT 26.730 107.225 27.240 107.315 ;
        RECT 25.280 106.760 25.585 106.890 ;
        RECT 26.030 106.780 26.560 107.145 ;
        RECT 24.900 106.165 25.165 106.625 ;
        RECT 25.335 106.335 25.585 106.760 ;
        RECT 26.730 106.610 26.900 107.225 ;
        RECT 25.795 106.440 26.900 106.610 ;
        RECT 27.070 106.165 27.240 106.965 ;
        RECT 27.410 106.665 27.580 107.735 ;
        RECT 27.750 106.835 27.940 107.555 ;
        RECT 28.110 106.805 28.430 107.765 ;
        RECT 28.600 107.805 28.770 108.265 ;
        RECT 29.045 108.185 29.255 108.715 ;
        RECT 29.515 107.975 29.845 108.500 ;
        RECT 30.015 108.105 30.185 108.715 ;
        RECT 30.355 108.060 30.685 108.495 ;
        RECT 30.355 107.975 30.735 108.060 ;
        RECT 31.365 107.990 31.655 108.715 ;
        RECT 31.840 108.145 32.095 108.495 ;
        RECT 32.265 108.315 32.595 108.715 ;
        RECT 32.765 108.145 32.935 108.495 ;
        RECT 33.105 108.315 33.485 108.715 ;
        RECT 31.840 107.975 33.505 108.145 ;
        RECT 33.675 108.040 33.950 108.385 ;
        RECT 34.750 108.205 34.990 108.715 ;
        RECT 35.170 108.205 35.450 108.535 ;
        RECT 35.680 108.205 35.895 108.715 ;
        RECT 29.645 107.805 29.845 107.975 ;
        RECT 30.510 107.935 30.735 107.975 ;
        RECT 28.600 107.475 29.475 107.805 ;
        RECT 29.645 107.475 30.395 107.805 ;
        RECT 27.410 106.335 27.660 106.665 ;
        RECT 28.600 106.635 28.770 107.475 ;
        RECT 29.645 107.270 29.835 107.475 ;
        RECT 30.565 107.355 30.735 107.935 ;
        RECT 33.335 107.805 33.505 107.975 ;
        RECT 31.825 107.475 32.170 107.805 ;
        RECT 32.340 107.475 33.165 107.805 ;
        RECT 33.335 107.475 33.610 107.805 ;
        RECT 30.520 107.305 30.735 107.355 ;
        RECT 28.940 106.895 29.835 107.270 ;
        RECT 30.345 107.225 30.735 107.305 ;
        RECT 27.885 106.465 28.770 106.635 ;
        RECT 28.950 106.165 29.265 106.665 ;
        RECT 29.495 106.335 29.835 106.895 ;
        RECT 30.005 106.165 30.175 107.175 ;
        RECT 30.345 106.380 30.675 107.225 ;
        RECT 31.365 106.165 31.655 107.330 ;
        RECT 31.845 107.015 32.170 107.305 ;
        RECT 32.340 107.185 32.535 107.475 ;
        RECT 33.335 107.305 33.505 107.475 ;
        RECT 33.780 107.305 33.950 108.040 ;
        RECT 34.645 107.475 35.000 108.035 ;
        RECT 35.170 107.305 35.340 108.205 ;
        RECT 35.510 107.475 35.775 108.035 ;
        RECT 36.065 107.975 36.680 108.545 ;
        RECT 36.890 108.185 37.180 108.535 ;
        RECT 37.375 108.355 37.705 108.715 ;
        RECT 37.875 108.185 38.105 108.490 ;
        RECT 36.890 108.015 38.105 108.185 ;
        RECT 38.295 108.375 38.465 108.410 ;
        RECT 38.295 108.205 38.495 108.375 ;
        RECT 36.025 107.305 36.195 107.805 ;
        RECT 32.845 107.135 33.505 107.305 ;
        RECT 32.845 107.015 33.015 107.135 ;
        RECT 31.845 106.845 33.015 107.015 ;
        RECT 31.825 106.385 33.015 106.675 ;
        RECT 33.185 106.165 33.465 106.965 ;
        RECT 33.675 106.335 33.950 107.305 ;
        RECT 34.770 107.135 36.195 107.305 ;
        RECT 34.770 106.960 35.160 107.135 ;
        RECT 35.645 106.165 35.975 106.965 ;
        RECT 36.365 106.955 36.680 107.975 ;
        RECT 38.295 107.845 38.465 108.205 ;
        RECT 38.765 107.895 38.995 108.715 ;
        RECT 39.165 107.915 39.495 108.545 ;
        RECT 36.950 107.695 37.210 107.805 ;
        RECT 36.945 107.525 37.210 107.695 ;
        RECT 36.950 107.475 37.210 107.525 ;
        RECT 37.390 107.475 37.775 107.805 ;
        RECT 37.945 107.675 38.465 107.845 ;
        RECT 36.145 106.335 36.680 106.955 ;
        RECT 36.890 106.165 37.210 107.305 ;
        RECT 37.390 106.425 37.585 107.475 ;
        RECT 37.945 107.295 38.115 107.675 ;
        RECT 37.765 107.015 38.115 107.295 ;
        RECT 38.305 107.145 38.550 107.505 ;
        RECT 38.745 107.475 39.075 107.725 ;
        RECT 39.245 107.315 39.495 107.915 ;
        RECT 39.665 107.895 39.875 108.715 ;
        RECT 40.105 108.170 45.450 108.715 ;
        RECT 41.690 107.340 42.030 108.170 ;
        RECT 45.625 107.945 47.295 108.715 ;
        RECT 47.930 108.145 48.250 108.545 ;
        RECT 37.765 106.335 38.095 107.015 ;
        RECT 38.295 106.165 38.550 106.965 ;
        RECT 38.765 106.165 38.995 107.305 ;
        RECT 39.165 106.335 39.495 107.315 ;
        RECT 39.665 106.165 39.875 107.305 ;
        RECT 43.510 106.600 43.860 107.850 ;
        RECT 45.625 107.425 46.375 107.945 ;
        RECT 46.545 107.255 47.295 107.775 ;
        RECT 40.105 106.165 45.450 106.600 ;
        RECT 45.625 106.165 47.295 107.255 ;
        RECT 47.930 107.355 48.100 108.145 ;
        RECT 48.420 107.895 48.730 108.715 ;
        RECT 48.900 108.085 49.230 108.545 ;
        RECT 49.400 108.255 49.650 108.715 ;
        RECT 49.840 108.335 51.890 108.545 ;
        RECT 49.840 108.085 50.590 108.165 ;
        RECT 48.900 107.895 50.590 108.085 ;
        RECT 50.760 107.895 50.930 108.335 ;
        RECT 51.100 107.895 51.890 108.165 ;
        RECT 48.270 107.525 48.620 107.725 ;
        RECT 48.900 107.525 49.580 107.725 ;
        RECT 49.790 107.525 50.980 107.725 ;
        RECT 51.160 107.355 51.490 107.725 ;
        RECT 47.930 107.185 51.490 107.355 ;
        RECT 47.930 106.735 48.100 107.185 ;
        RECT 51.690 107.015 51.890 107.895 ;
        RECT 52.065 107.945 53.735 108.715 ;
        RECT 54.365 108.085 54.705 108.545 ;
        RECT 54.875 108.255 55.045 108.715 ;
        RECT 55.675 108.280 56.035 108.545 ;
        RECT 55.680 108.275 56.035 108.280 ;
        RECT 55.685 108.265 56.035 108.275 ;
        RECT 55.690 108.260 56.035 108.265 ;
        RECT 55.695 108.250 56.035 108.260 ;
        RECT 56.275 108.255 56.445 108.715 ;
        RECT 55.700 108.245 56.035 108.250 ;
        RECT 55.710 108.235 56.035 108.245 ;
        RECT 55.720 108.225 56.035 108.235 ;
        RECT 55.215 108.085 55.545 108.165 ;
        RECT 52.065 107.425 52.815 107.945 ;
        RECT 54.365 107.895 55.545 108.085 ;
        RECT 55.735 108.085 56.035 108.225 ;
        RECT 55.735 107.895 56.445 108.085 ;
        RECT 52.985 107.255 53.735 107.775 ;
        RECT 47.930 106.335 48.250 106.735 ;
        RECT 48.420 106.165 48.730 106.965 ;
        RECT 48.900 106.845 51.890 107.015 ;
        RECT 48.900 106.795 50.070 106.845 ;
        RECT 48.900 106.335 49.230 106.795 ;
        RECT 49.400 106.165 49.570 106.625 ;
        RECT 49.740 106.335 50.070 106.795 ;
        RECT 51.100 106.795 51.890 106.845 ;
        RECT 50.240 106.165 50.490 106.625 ;
        RECT 50.680 106.165 50.930 106.625 ;
        RECT 51.100 106.335 51.350 106.795 ;
        RECT 51.600 106.165 51.890 106.625 ;
        RECT 52.065 106.165 53.735 107.255 ;
        RECT 54.365 107.525 54.695 107.725 ;
        RECT 55.005 107.705 55.335 107.725 ;
        RECT 54.885 107.525 55.335 107.705 ;
        RECT 54.365 107.185 54.595 107.525 ;
        RECT 54.375 106.165 54.705 106.885 ;
        RECT 54.885 106.410 55.100 107.525 ;
        RECT 55.505 107.495 55.975 107.725 ;
        RECT 56.160 107.325 56.445 107.895 ;
        RECT 56.615 107.770 56.955 108.545 ;
        RECT 57.125 107.990 57.415 108.715 ;
        RECT 57.670 108.145 57.845 108.545 ;
        RECT 58.015 108.335 58.345 108.715 ;
        RECT 58.590 108.215 58.820 108.545 ;
        RECT 57.670 107.975 58.300 108.145 ;
        RECT 58.130 107.805 58.300 107.975 ;
        RECT 55.295 107.110 56.445 107.325 ;
        RECT 55.295 106.335 55.625 107.110 ;
        RECT 55.795 106.165 56.505 106.940 ;
        RECT 56.675 106.335 56.955 107.770 ;
        RECT 57.125 106.165 57.415 107.330 ;
        RECT 57.585 107.125 57.950 107.805 ;
        RECT 58.130 107.475 58.480 107.805 ;
        RECT 58.130 106.955 58.300 107.475 ;
        RECT 57.670 106.785 58.300 106.955 ;
        RECT 58.650 106.925 58.820 108.215 ;
        RECT 59.020 107.105 59.300 108.380 ;
        RECT 59.525 108.375 59.795 108.380 ;
        RECT 59.485 108.205 59.795 108.375 ;
        RECT 60.255 108.335 60.585 108.715 ;
        RECT 60.755 108.460 61.090 108.505 ;
        RECT 59.525 107.105 59.795 108.205 ;
        RECT 59.985 107.105 60.325 108.135 ;
        RECT 60.755 107.995 61.095 108.460 ;
        RECT 60.495 107.475 60.755 107.805 ;
        RECT 60.495 106.925 60.665 107.475 ;
        RECT 60.925 107.305 61.095 107.995 ;
        RECT 57.670 106.335 57.845 106.785 ;
        RECT 58.650 106.755 60.665 106.925 ;
        RECT 58.015 106.165 58.345 106.605 ;
        RECT 58.650 106.335 58.820 106.755 ;
        RECT 59.055 106.165 59.725 106.575 ;
        RECT 59.940 106.335 60.110 106.755 ;
        RECT 60.310 106.165 60.640 106.575 ;
        RECT 60.835 106.335 61.095 107.305 ;
        RECT 62.185 107.975 62.570 108.545 ;
        RECT 62.740 108.255 63.065 108.715 ;
        RECT 63.585 108.085 63.865 108.545 ;
        RECT 62.185 107.305 62.465 107.975 ;
        RECT 62.740 107.915 63.865 108.085 ;
        RECT 62.740 107.805 63.190 107.915 ;
        RECT 62.635 107.475 63.190 107.805 ;
        RECT 64.055 107.745 64.455 108.545 ;
        RECT 64.855 108.255 65.125 108.715 ;
        RECT 65.295 108.085 65.580 108.545 ;
        RECT 65.865 108.325 67.125 108.505 ;
        RECT 62.185 106.335 62.570 107.305 ;
        RECT 62.740 107.015 63.190 107.475 ;
        RECT 63.360 107.185 64.455 107.745 ;
        RECT 62.740 106.795 63.865 107.015 ;
        RECT 62.740 106.165 63.065 106.625 ;
        RECT 63.585 106.335 63.865 106.795 ;
        RECT 64.055 106.335 64.455 107.185 ;
        RECT 64.625 107.915 65.580 108.085 ;
        RECT 64.625 107.015 64.835 107.915 ;
        RECT 65.005 107.185 65.695 107.745 ;
        RECT 64.625 106.795 65.580 107.015 ;
        RECT 65.865 106.810 66.105 108.135 ;
        RECT 66.275 107.975 66.625 108.155 ;
        RECT 66.795 108.105 67.125 108.325 ;
        RECT 67.315 108.275 67.485 108.715 ;
        RECT 67.655 108.105 67.995 108.520 ;
        RECT 66.795 107.975 67.995 108.105 ;
        RECT 66.275 106.965 66.445 107.975 ;
        RECT 66.965 107.935 67.995 107.975 ;
        RECT 68.165 107.945 71.675 108.715 ;
        RECT 71.935 108.165 72.105 108.455 ;
        RECT 72.275 108.335 72.605 108.715 ;
        RECT 71.935 107.995 72.600 108.165 ;
        RECT 66.615 107.385 66.785 107.805 ;
        RECT 67.000 107.555 67.365 107.725 ;
        RECT 66.615 107.135 67.015 107.385 ;
        RECT 67.185 107.355 67.365 107.555 ;
        RECT 67.535 107.525 67.995 107.725 ;
        RECT 68.165 107.425 69.815 107.945 ;
        RECT 67.185 107.185 67.505 107.355 ;
        RECT 64.855 106.165 65.125 106.625 ;
        RECT 65.295 106.335 65.580 106.795 ;
        RECT 66.275 106.755 67.115 106.965 ;
        RECT 65.915 106.165 66.125 106.625 ;
        RECT 66.615 106.335 67.115 106.755 ;
        RECT 67.305 106.395 67.505 107.185 ;
        RECT 67.675 106.165 67.995 107.345 ;
        RECT 69.985 107.255 71.675 107.775 ;
        RECT 68.165 106.165 71.675 107.255 ;
        RECT 71.850 107.175 72.200 107.825 ;
        RECT 72.370 107.005 72.600 107.995 ;
        RECT 71.935 106.835 72.600 107.005 ;
        RECT 71.935 106.335 72.105 106.835 ;
        RECT 72.275 106.165 72.605 106.665 ;
        RECT 72.775 106.335 72.960 108.455 ;
        RECT 73.215 108.255 73.465 108.715 ;
        RECT 73.635 108.265 73.970 108.435 ;
        RECT 74.165 108.265 74.840 108.435 ;
        RECT 73.635 108.125 73.805 108.265 ;
        RECT 73.130 107.135 73.410 108.085 ;
        RECT 73.580 107.995 73.805 108.125 ;
        RECT 73.580 106.890 73.750 107.995 ;
        RECT 73.975 107.845 74.500 108.065 ;
        RECT 73.920 107.080 74.160 107.675 ;
        RECT 74.330 107.145 74.500 107.845 ;
        RECT 74.670 107.485 74.840 108.265 ;
        RECT 75.160 108.215 75.530 108.715 ;
        RECT 75.710 108.265 76.115 108.435 ;
        RECT 76.285 108.265 77.070 108.435 ;
        RECT 75.710 108.035 75.880 108.265 ;
        RECT 75.050 107.735 75.880 108.035 ;
        RECT 76.265 107.765 76.730 108.095 ;
        RECT 75.050 107.705 75.250 107.735 ;
        RECT 75.370 107.485 75.540 107.555 ;
        RECT 74.670 107.315 75.540 107.485 ;
        RECT 75.030 107.225 75.540 107.315 ;
        RECT 73.580 106.760 73.885 106.890 ;
        RECT 74.330 106.780 74.860 107.145 ;
        RECT 73.200 106.165 73.465 106.625 ;
        RECT 73.635 106.335 73.885 106.760 ;
        RECT 75.030 106.610 75.200 107.225 ;
        RECT 74.095 106.440 75.200 106.610 ;
        RECT 75.370 106.165 75.540 106.965 ;
        RECT 75.710 106.665 75.880 107.735 ;
        RECT 76.050 106.835 76.240 107.555 ;
        RECT 76.410 106.805 76.730 107.765 ;
        RECT 76.900 107.805 77.070 108.265 ;
        RECT 77.345 108.185 77.555 108.715 ;
        RECT 77.815 107.975 78.145 108.500 ;
        RECT 78.315 108.105 78.485 108.715 ;
        RECT 78.655 108.060 78.985 108.495 ;
        RECT 78.655 107.975 79.035 108.060 ;
        RECT 77.945 107.805 78.145 107.975 ;
        RECT 78.810 107.935 79.035 107.975 ;
        RECT 76.900 107.475 77.775 107.805 ;
        RECT 77.945 107.475 78.695 107.805 ;
        RECT 75.710 106.335 75.960 106.665 ;
        RECT 76.900 106.635 77.070 107.475 ;
        RECT 77.945 107.270 78.135 107.475 ;
        RECT 78.865 107.355 79.035 107.935 ;
        RECT 78.820 107.305 79.035 107.355 ;
        RECT 77.240 106.895 78.135 107.270 ;
        RECT 78.645 107.225 79.035 107.305 ;
        RECT 79.205 107.975 79.590 108.545 ;
        RECT 79.760 108.255 80.085 108.715 ;
        RECT 80.605 108.085 80.885 108.545 ;
        RECT 79.205 107.305 79.485 107.975 ;
        RECT 79.760 107.915 80.885 108.085 ;
        RECT 79.760 107.805 80.210 107.915 ;
        RECT 79.655 107.475 80.210 107.805 ;
        RECT 81.075 107.745 81.475 108.545 ;
        RECT 81.875 108.255 82.145 108.715 ;
        RECT 82.315 108.085 82.600 108.545 ;
        RECT 76.185 106.465 77.070 106.635 ;
        RECT 77.250 106.165 77.565 106.665 ;
        RECT 77.795 106.335 78.135 106.895 ;
        RECT 78.305 106.165 78.475 107.175 ;
        RECT 78.645 106.380 78.975 107.225 ;
        RECT 79.205 106.335 79.590 107.305 ;
        RECT 79.760 107.015 80.210 107.475 ;
        RECT 80.380 107.185 81.475 107.745 ;
        RECT 79.760 106.795 80.885 107.015 ;
        RECT 79.760 106.165 80.085 106.625 ;
        RECT 80.605 106.335 80.885 106.795 ;
        RECT 81.075 106.335 81.475 107.185 ;
        RECT 81.645 107.915 82.600 108.085 ;
        RECT 82.885 107.965 84.095 108.715 ;
        RECT 81.645 107.015 81.855 107.915 ;
        RECT 82.025 107.185 82.715 107.745 ;
        RECT 82.885 107.255 83.405 107.795 ;
        RECT 83.575 107.425 84.095 107.965 ;
        RECT 81.645 106.795 82.600 107.015 ;
        RECT 81.875 106.165 82.145 106.625 ;
        RECT 82.315 106.335 82.600 106.795 ;
        RECT 82.885 106.165 84.095 107.255 ;
        RECT 5.520 105.995 84.180 106.165 ;
        RECT 5.605 104.905 6.815 105.995 ;
        RECT 7.075 105.325 7.245 105.825 ;
        RECT 7.415 105.495 7.745 105.995 ;
        RECT 7.075 105.155 7.740 105.325 ;
        RECT 5.605 104.195 6.125 104.735 ;
        RECT 6.295 104.365 6.815 104.905 ;
        RECT 6.990 104.335 7.340 104.985 ;
        RECT 5.605 103.445 6.815 104.195 ;
        RECT 7.510 104.165 7.740 105.155 ;
        RECT 7.075 103.995 7.740 104.165 ;
        RECT 7.075 103.705 7.245 103.995 ;
        RECT 7.415 103.445 7.745 103.825 ;
        RECT 7.915 103.705 8.100 105.825 ;
        RECT 8.340 105.535 8.605 105.995 ;
        RECT 8.775 105.400 9.025 105.825 ;
        RECT 9.235 105.550 10.340 105.720 ;
        RECT 8.720 105.270 9.025 105.400 ;
        RECT 8.270 104.075 8.550 105.025 ;
        RECT 8.720 104.165 8.890 105.270 ;
        RECT 9.060 104.485 9.300 105.080 ;
        RECT 9.470 105.015 10.000 105.380 ;
        RECT 9.470 104.315 9.640 105.015 ;
        RECT 10.170 104.935 10.340 105.550 ;
        RECT 10.510 105.195 10.680 105.995 ;
        RECT 10.850 105.495 11.100 105.825 ;
        RECT 11.325 105.525 12.210 105.695 ;
        RECT 10.170 104.845 10.680 104.935 ;
        RECT 8.720 104.035 8.945 104.165 ;
        RECT 9.115 104.095 9.640 104.315 ;
        RECT 9.810 104.675 10.680 104.845 ;
        RECT 8.355 103.445 8.605 103.905 ;
        RECT 8.775 103.895 8.945 104.035 ;
        RECT 9.810 103.895 9.980 104.675 ;
        RECT 10.510 104.605 10.680 104.675 ;
        RECT 10.190 104.425 10.390 104.455 ;
        RECT 10.850 104.425 11.020 105.495 ;
        RECT 11.190 104.605 11.380 105.325 ;
        RECT 10.190 104.125 11.020 104.425 ;
        RECT 11.550 104.395 11.870 105.355 ;
        RECT 8.775 103.725 9.110 103.895 ;
        RECT 9.305 103.725 9.980 103.895 ;
        RECT 10.300 103.445 10.670 103.945 ;
        RECT 10.850 103.895 11.020 104.125 ;
        RECT 11.405 104.065 11.870 104.395 ;
        RECT 12.040 104.685 12.210 105.525 ;
        RECT 12.390 105.495 12.705 105.995 ;
        RECT 12.935 105.265 13.275 105.825 ;
        RECT 12.380 104.890 13.275 105.265 ;
        RECT 13.445 104.985 13.615 105.995 ;
        RECT 13.085 104.685 13.275 104.890 ;
        RECT 13.785 104.935 14.115 105.780 ;
        RECT 13.785 104.855 14.175 104.935 ;
        RECT 14.350 104.855 14.670 105.995 ;
        RECT 13.960 104.805 14.175 104.855 ;
        RECT 12.040 104.355 12.915 104.685 ;
        RECT 13.085 104.355 13.835 104.685 ;
        RECT 12.040 103.895 12.210 104.355 ;
        RECT 13.085 104.185 13.285 104.355 ;
        RECT 14.005 104.225 14.175 104.805 ;
        RECT 14.850 104.685 15.045 105.735 ;
        RECT 15.225 105.145 15.555 105.825 ;
        RECT 15.755 105.195 16.010 105.995 ;
        RECT 16.220 105.205 16.755 105.825 ;
        RECT 15.225 104.865 15.575 105.145 ;
        RECT 14.410 104.635 14.670 104.685 ;
        RECT 14.405 104.465 14.670 104.635 ;
        RECT 14.410 104.355 14.670 104.465 ;
        RECT 14.850 104.355 15.235 104.685 ;
        RECT 15.405 104.485 15.575 104.865 ;
        RECT 15.765 104.655 16.010 105.015 ;
        RECT 15.405 104.315 15.925 104.485 ;
        RECT 13.950 104.185 14.175 104.225 ;
        RECT 10.850 103.725 11.255 103.895 ;
        RECT 11.425 103.725 12.210 103.895 ;
        RECT 12.485 103.445 12.695 103.975 ;
        RECT 12.955 103.660 13.285 104.185 ;
        RECT 13.795 104.100 14.175 104.185 ;
        RECT 13.455 103.445 13.625 104.055 ;
        RECT 13.795 103.665 14.125 104.100 ;
        RECT 14.350 103.975 15.565 104.145 ;
        RECT 14.350 103.625 14.640 103.975 ;
        RECT 14.835 103.445 15.165 103.805 ;
        RECT 15.335 103.670 15.565 103.975 ;
        RECT 15.755 103.750 15.925 104.315 ;
        RECT 16.220 104.185 16.535 105.205 ;
        RECT 16.925 105.195 17.255 105.995 ;
        RECT 17.740 105.025 18.130 105.200 ;
        RECT 16.705 104.855 18.130 105.025 ;
        RECT 16.705 104.355 16.875 104.855 ;
        RECT 16.220 103.615 16.835 104.185 ;
        RECT 17.125 104.125 17.390 104.685 ;
        RECT 17.560 103.955 17.730 104.855 ;
        RECT 18.485 104.830 18.775 105.995 ;
        RECT 19.865 105.485 21.065 105.725 ;
        RECT 21.245 105.570 21.575 105.995 ;
        RECT 22.090 105.570 22.450 105.995 ;
        RECT 22.655 105.400 22.915 105.580 ;
        RECT 21.280 105.315 22.915 105.400 ;
        RECT 19.865 104.855 20.170 105.285 ;
        RECT 20.340 105.230 22.915 105.315 ;
        RECT 20.340 105.145 21.450 105.230 ;
        RECT 22.235 105.170 22.915 105.230 ;
        RECT 17.900 104.125 18.255 104.685 ;
        RECT 19.865 104.185 20.035 104.855 ;
        RECT 20.340 104.685 20.510 105.145 ;
        RECT 20.210 104.355 20.510 104.685 ;
        RECT 20.770 104.435 21.305 104.975 ;
        RECT 21.670 104.855 22.065 105.060 ;
        RECT 21.555 104.295 21.725 104.685 ;
        RECT 21.405 104.265 21.725 104.295 ;
        RECT 20.840 104.185 21.725 104.265 ;
        RECT 17.005 103.445 17.220 103.955 ;
        RECT 17.450 103.625 17.730 103.955 ;
        RECT 17.910 103.445 18.150 103.955 ;
        RECT 18.485 103.445 18.775 104.170 ;
        RECT 19.865 104.125 21.725 104.185 ;
        RECT 19.865 104.095 21.575 104.125 ;
        RECT 19.865 104.015 21.010 104.095 ;
        RECT 19.865 103.965 20.170 104.015 ;
        RECT 19.915 103.665 20.170 103.965 ;
        RECT 20.340 103.445 20.670 103.845 ;
        RECT 20.840 103.665 21.010 104.015 ;
        RECT 21.895 103.955 22.065 104.855 ;
        RECT 22.235 104.265 22.405 105.170 ;
        RECT 22.575 104.435 22.915 105.000 ;
        RECT 23.090 104.855 23.365 105.825 ;
        RECT 23.575 105.195 23.855 105.995 ;
        RECT 24.025 105.485 25.215 105.775 ;
        RECT 24.025 105.145 25.195 105.315 ;
        RECT 24.025 105.025 24.195 105.145 ;
        RECT 23.535 104.855 24.195 105.025 ;
        RECT 22.235 104.095 22.915 104.265 ;
        RECT 21.310 103.445 21.480 103.925 ;
        RECT 21.715 103.625 22.065 103.955 ;
        RECT 22.235 103.445 22.405 103.925 ;
        RECT 22.655 103.650 22.915 104.095 ;
        RECT 23.090 104.120 23.260 104.855 ;
        RECT 23.535 104.685 23.705 104.855 ;
        RECT 24.505 104.685 24.700 104.975 ;
        RECT 24.870 104.855 25.195 105.145 ;
        RECT 25.385 104.905 27.055 105.995 ;
        RECT 23.430 104.355 23.705 104.685 ;
        RECT 23.875 104.355 24.700 104.685 ;
        RECT 24.870 104.355 25.215 104.685 ;
        RECT 23.535 104.185 23.705 104.355 ;
        RECT 25.385 104.215 26.135 104.735 ;
        RECT 26.305 104.385 27.055 104.905 ;
        RECT 27.685 104.855 27.965 105.995 ;
        RECT 28.135 104.845 28.465 105.825 ;
        RECT 28.635 104.855 28.895 105.995 ;
        RECT 29.065 104.855 29.340 105.825 ;
        RECT 29.550 105.195 29.830 105.995 ;
        RECT 30.000 105.485 31.615 105.815 ;
        RECT 30.000 105.145 31.175 105.315 ;
        RECT 30.000 105.025 30.170 105.145 ;
        RECT 29.510 104.855 30.170 105.025 ;
        RECT 27.695 104.415 28.030 104.685 ;
        RECT 28.200 104.245 28.370 104.845 ;
        RECT 28.540 104.435 28.875 104.685 ;
        RECT 23.090 103.775 23.365 104.120 ;
        RECT 23.535 104.015 25.200 104.185 ;
        RECT 23.555 103.445 23.935 103.845 ;
        RECT 24.105 103.665 24.275 104.015 ;
        RECT 24.445 103.445 24.775 103.845 ;
        RECT 24.945 103.665 25.200 104.015 ;
        RECT 25.385 103.445 27.055 104.215 ;
        RECT 27.685 103.445 27.995 104.245 ;
        RECT 28.200 103.615 28.895 104.245 ;
        RECT 29.065 104.120 29.235 104.855 ;
        RECT 29.510 104.685 29.680 104.855 ;
        RECT 30.430 104.685 30.675 104.975 ;
        RECT 30.845 104.855 31.175 105.145 ;
        RECT 31.435 104.685 31.605 105.245 ;
        RECT 31.855 104.855 32.115 105.995 ;
        RECT 32.285 104.855 32.670 105.825 ;
        RECT 32.840 105.535 33.165 105.995 ;
        RECT 33.685 105.365 33.965 105.825 ;
        RECT 32.840 105.145 33.965 105.365 ;
        RECT 29.405 104.355 29.680 104.685 ;
        RECT 29.850 104.355 30.675 104.685 ;
        RECT 30.890 104.355 31.605 104.685 ;
        RECT 31.775 104.435 32.110 104.685 ;
        RECT 29.510 104.185 29.680 104.355 ;
        RECT 31.355 104.265 31.605 104.355 ;
        RECT 29.065 103.775 29.340 104.120 ;
        RECT 29.510 104.015 31.175 104.185 ;
        RECT 29.530 103.445 29.905 103.845 ;
        RECT 30.075 103.665 30.245 104.015 ;
        RECT 30.415 103.445 30.745 103.845 ;
        RECT 30.915 103.615 31.175 104.015 ;
        RECT 31.355 103.845 31.685 104.265 ;
        RECT 31.855 103.445 32.115 104.265 ;
        RECT 32.285 104.185 32.565 104.855 ;
        RECT 32.840 104.685 33.290 105.145 ;
        RECT 34.155 104.975 34.555 105.825 ;
        RECT 34.955 105.535 35.225 105.995 ;
        RECT 35.395 105.365 35.680 105.825 ;
        RECT 32.735 104.355 33.290 104.685 ;
        RECT 33.460 104.415 34.555 104.975 ;
        RECT 32.840 104.245 33.290 104.355 ;
        RECT 32.285 103.615 32.670 104.185 ;
        RECT 32.840 104.075 33.965 104.245 ;
        RECT 32.840 103.445 33.165 103.905 ;
        RECT 33.685 103.615 33.965 104.075 ;
        RECT 34.155 103.615 34.555 104.415 ;
        RECT 34.725 105.145 35.680 105.365 ;
        RECT 36.165 105.325 36.445 105.995 ;
        RECT 34.725 104.245 34.935 105.145 ;
        RECT 36.615 105.105 36.915 105.655 ;
        RECT 37.115 105.275 37.445 105.995 ;
        RECT 37.635 105.275 38.095 105.825 ;
        RECT 35.105 104.415 35.795 104.975 ;
        RECT 35.980 104.685 36.245 105.045 ;
        RECT 36.615 104.935 37.555 105.105 ;
        RECT 37.385 104.685 37.555 104.935 ;
        RECT 35.980 104.435 36.655 104.685 ;
        RECT 36.875 104.435 37.215 104.685 ;
        RECT 37.385 104.355 37.675 104.685 ;
        RECT 37.385 104.265 37.555 104.355 ;
        RECT 34.725 104.075 35.680 104.245 ;
        RECT 34.955 103.445 35.225 103.905 ;
        RECT 35.395 103.615 35.680 104.075 ;
        RECT 36.165 104.075 37.555 104.265 ;
        RECT 36.165 103.715 36.495 104.075 ;
        RECT 37.845 103.905 38.095 105.275 ;
        RECT 38.265 104.905 41.775 105.995 ;
        RECT 41.945 105.440 42.550 105.995 ;
        RECT 42.725 105.485 43.205 105.825 ;
        RECT 43.375 105.450 43.630 105.995 ;
        RECT 41.945 105.340 42.560 105.440 ;
        RECT 42.375 105.315 42.560 105.340 ;
        RECT 37.115 103.445 37.365 103.905 ;
        RECT 37.535 103.615 38.095 103.905 ;
        RECT 38.265 104.215 39.915 104.735 ;
        RECT 40.085 104.385 41.775 104.905 ;
        RECT 41.945 104.720 42.205 105.170 ;
        RECT 42.375 105.070 42.705 105.315 ;
        RECT 42.875 104.995 43.630 105.245 ;
        RECT 43.800 105.125 44.075 105.825 ;
        RECT 42.860 104.960 43.630 104.995 ;
        RECT 42.845 104.950 43.630 104.960 ;
        RECT 42.840 104.935 43.735 104.950 ;
        RECT 42.820 104.920 43.735 104.935 ;
        RECT 42.800 104.910 43.735 104.920 ;
        RECT 42.775 104.900 43.735 104.910 ;
        RECT 42.705 104.870 43.735 104.900 ;
        RECT 42.685 104.840 43.735 104.870 ;
        RECT 42.665 104.810 43.735 104.840 ;
        RECT 42.635 104.785 43.735 104.810 ;
        RECT 42.600 104.750 43.735 104.785 ;
        RECT 42.570 104.745 43.735 104.750 ;
        RECT 42.570 104.740 42.960 104.745 ;
        RECT 42.570 104.730 42.935 104.740 ;
        RECT 42.570 104.725 42.920 104.730 ;
        RECT 42.570 104.720 42.905 104.725 ;
        RECT 41.945 104.715 42.905 104.720 ;
        RECT 41.945 104.705 42.895 104.715 ;
        RECT 41.945 104.700 42.885 104.705 ;
        RECT 41.945 104.690 42.875 104.700 ;
        RECT 41.945 104.680 42.870 104.690 ;
        RECT 41.945 104.675 42.865 104.680 ;
        RECT 41.945 104.660 42.855 104.675 ;
        RECT 41.945 104.645 42.850 104.660 ;
        RECT 41.945 104.620 42.840 104.645 ;
        RECT 41.945 104.550 42.835 104.620 ;
        RECT 38.265 103.445 41.775 104.215 ;
        RECT 41.945 103.995 42.495 104.380 ;
        RECT 42.665 103.825 42.835 104.550 ;
        RECT 41.945 103.655 42.835 103.825 ;
        RECT 43.005 104.150 43.335 104.575 ;
        RECT 43.505 104.350 43.735 104.745 ;
        RECT 43.005 103.665 43.225 104.150 ;
        RECT 43.905 104.095 44.075 105.125 ;
        RECT 44.245 104.830 44.535 105.995 ;
        RECT 44.715 105.185 45.010 105.995 ;
        RECT 45.190 104.685 45.435 105.825 ;
        RECT 45.610 105.185 45.870 105.995 ;
        RECT 46.470 105.990 52.745 105.995 ;
        RECT 46.050 104.685 46.300 105.820 ;
        RECT 46.470 105.195 46.730 105.990 ;
        RECT 46.900 105.095 47.160 105.820 ;
        RECT 47.330 105.265 47.590 105.990 ;
        RECT 47.760 105.095 48.020 105.820 ;
        RECT 48.190 105.265 48.450 105.990 ;
        RECT 48.620 105.095 48.880 105.820 ;
        RECT 49.050 105.265 49.310 105.990 ;
        RECT 49.480 105.095 49.740 105.820 ;
        RECT 49.910 105.265 50.155 105.990 ;
        RECT 50.325 105.095 50.585 105.820 ;
        RECT 50.770 105.265 51.015 105.990 ;
        RECT 51.185 105.095 51.445 105.820 ;
        RECT 51.630 105.265 51.875 105.990 ;
        RECT 52.045 105.095 52.305 105.820 ;
        RECT 52.490 105.265 52.745 105.990 ;
        RECT 46.900 105.080 52.305 105.095 ;
        RECT 52.915 105.080 53.205 105.820 ;
        RECT 53.375 105.250 53.645 105.995 ;
        RECT 46.900 104.855 53.645 105.080 ;
        RECT 53.905 104.905 57.415 105.995 ;
        RECT 43.395 103.445 43.645 103.985 ;
        RECT 43.815 103.615 44.075 104.095 ;
        RECT 44.245 103.445 44.535 104.170 ;
        RECT 44.705 104.125 45.020 104.685 ;
        RECT 45.190 104.435 52.310 104.685 ;
        RECT 44.705 103.445 45.010 103.955 ;
        RECT 45.190 103.625 45.440 104.435 ;
        RECT 45.610 103.445 45.870 103.970 ;
        RECT 46.050 103.625 46.300 104.435 ;
        RECT 52.480 104.265 53.645 104.855 ;
        RECT 46.900 104.095 53.645 104.265 ;
        RECT 53.905 104.215 55.555 104.735 ;
        RECT 55.725 104.385 57.415 104.905 ;
        RECT 58.545 104.855 58.775 105.995 ;
        RECT 58.945 104.845 59.275 105.825 ;
        RECT 59.445 104.855 59.655 105.995 ;
        RECT 59.885 104.905 61.095 105.995 ;
        RECT 58.525 104.435 58.855 104.685 ;
        RECT 46.470 103.445 46.730 104.005 ;
        RECT 46.900 103.640 47.160 104.095 ;
        RECT 47.330 103.445 47.590 103.925 ;
        RECT 47.760 103.640 48.020 104.095 ;
        RECT 48.190 103.445 48.450 103.925 ;
        RECT 48.620 103.640 48.880 104.095 ;
        RECT 49.050 103.445 49.295 103.925 ;
        RECT 49.465 103.640 49.740 104.095 ;
        RECT 49.910 103.445 50.155 103.925 ;
        RECT 50.325 103.640 50.585 104.095 ;
        RECT 50.765 103.445 51.015 103.925 ;
        RECT 51.185 103.640 51.445 104.095 ;
        RECT 51.625 103.445 51.875 103.925 ;
        RECT 52.045 103.640 52.305 104.095 ;
        RECT 52.485 103.445 52.745 103.925 ;
        RECT 52.915 103.640 53.175 104.095 ;
        RECT 53.345 103.445 53.645 103.925 ;
        RECT 53.905 103.445 57.415 104.215 ;
        RECT 58.545 103.445 58.775 104.265 ;
        RECT 59.025 104.245 59.275 104.845 ;
        RECT 58.945 103.615 59.275 104.245 ;
        RECT 59.445 103.445 59.655 104.265 ;
        RECT 59.885 104.195 60.405 104.735 ;
        RECT 60.575 104.365 61.095 104.905 ;
        RECT 61.265 105.125 61.540 105.825 ;
        RECT 61.750 105.450 61.965 105.995 ;
        RECT 62.135 105.485 62.610 105.825 ;
        RECT 62.780 105.490 63.395 105.995 ;
        RECT 62.780 105.315 62.975 105.490 ;
        RECT 59.885 103.445 61.095 104.195 ;
        RECT 61.265 104.095 61.435 105.125 ;
        RECT 61.710 104.955 62.425 105.250 ;
        RECT 62.645 105.125 62.975 105.315 ;
        RECT 63.145 104.955 63.395 105.320 ;
        RECT 61.605 104.785 63.395 104.955 ;
        RECT 61.605 104.355 61.835 104.785 ;
        RECT 61.265 103.615 61.525 104.095 ;
        RECT 62.005 104.085 62.415 104.605 ;
        RECT 61.695 103.445 62.025 103.905 ;
        RECT 62.215 103.665 62.415 104.085 ;
        RECT 62.585 103.930 62.840 104.785 ;
        RECT 63.635 104.605 63.805 105.825 ;
        RECT 64.055 105.485 64.315 105.995 ;
        RECT 64.485 105.485 65.675 105.775 ;
        RECT 63.010 104.355 63.805 104.605 ;
        RECT 63.975 104.435 64.315 105.315 ;
        RECT 64.505 105.145 65.675 105.315 ;
        RECT 65.845 105.195 66.125 105.995 ;
        RECT 64.505 104.855 64.830 105.145 ;
        RECT 65.505 105.025 65.675 105.145 ;
        RECT 65.000 104.685 65.195 104.975 ;
        RECT 65.505 104.855 66.165 105.025 ;
        RECT 66.335 104.855 66.610 105.825 ;
        RECT 66.785 104.855 67.045 105.995 ;
        RECT 67.215 105.025 67.545 105.825 ;
        RECT 67.715 105.195 67.885 105.995 ;
        RECT 68.055 105.025 68.385 105.825 ;
        RECT 68.555 105.195 68.810 105.995 ;
        RECT 67.215 104.855 68.915 105.025 ;
        RECT 65.995 104.685 66.165 104.855 ;
        RECT 64.485 104.355 64.830 104.685 ;
        RECT 65.000 104.355 65.825 104.685 ;
        RECT 65.995 104.355 66.270 104.685 ;
        RECT 63.555 104.265 63.805 104.355 ;
        RECT 62.585 103.665 63.375 103.930 ;
        RECT 63.555 103.845 63.885 104.265 ;
        RECT 64.055 103.445 64.315 104.265 ;
        RECT 65.995 104.185 66.165 104.355 ;
        RECT 64.500 104.015 66.165 104.185 ;
        RECT 66.440 104.120 66.610 104.855 ;
        RECT 66.785 104.435 67.545 104.685 ;
        RECT 67.715 104.435 68.465 104.685 ;
        RECT 68.635 104.265 68.915 104.855 ;
        RECT 70.005 104.830 70.295 105.995 ;
        RECT 70.960 105.195 71.210 105.995 ;
        RECT 71.380 105.365 71.710 105.825 ;
        RECT 71.880 105.535 72.095 105.995 ;
        RECT 71.380 105.195 72.550 105.365 ;
        RECT 70.470 105.025 70.750 105.185 ;
        RECT 70.470 104.855 71.805 105.025 ;
        RECT 71.635 104.685 71.805 104.855 ;
        RECT 70.470 104.435 70.820 104.675 ;
        RECT 70.990 104.435 71.465 104.675 ;
        RECT 71.635 104.435 72.010 104.685 ;
        RECT 71.635 104.265 71.805 104.435 ;
        RECT 64.500 103.665 64.755 104.015 ;
        RECT 64.925 103.445 65.255 103.845 ;
        RECT 65.425 103.665 65.595 104.015 ;
        RECT 65.765 103.445 66.145 103.845 ;
        RECT 66.335 103.775 66.610 104.120 ;
        RECT 66.785 104.075 67.885 104.245 ;
        RECT 66.785 103.615 67.125 104.075 ;
        RECT 67.295 103.445 67.465 103.905 ;
        RECT 67.635 103.825 67.885 104.075 ;
        RECT 68.055 104.015 68.915 104.265 ;
        RECT 68.475 103.825 68.805 103.845 ;
        RECT 67.635 103.615 68.805 103.825 ;
        RECT 70.005 103.445 70.295 104.170 ;
        RECT 70.470 104.095 71.805 104.265 ;
        RECT 70.470 103.885 70.740 104.095 ;
        RECT 72.180 103.905 72.550 105.195 ;
        RECT 72.765 104.905 73.975 105.995 ;
        RECT 70.960 103.445 71.290 103.905 ;
        RECT 71.800 103.615 72.550 103.905 ;
        RECT 72.765 104.195 73.285 104.735 ;
        RECT 73.455 104.365 73.975 104.905 ;
        RECT 74.150 104.855 74.485 105.825 ;
        RECT 74.655 104.855 74.825 105.995 ;
        RECT 74.995 105.655 77.025 105.825 ;
        RECT 72.765 103.445 73.975 104.195 ;
        RECT 74.150 104.185 74.320 104.855 ;
        RECT 74.995 104.685 75.165 105.655 ;
        RECT 74.490 104.355 74.745 104.685 ;
        RECT 74.970 104.355 75.165 104.685 ;
        RECT 75.335 105.315 76.460 105.485 ;
        RECT 74.575 104.185 74.745 104.355 ;
        RECT 75.335 104.185 75.505 105.315 ;
        RECT 74.150 103.615 74.405 104.185 ;
        RECT 74.575 104.015 75.505 104.185 ;
        RECT 75.675 104.975 76.685 105.145 ;
        RECT 75.675 104.175 75.845 104.975 ;
        RECT 76.050 104.635 76.325 104.775 ;
        RECT 76.045 104.465 76.325 104.635 ;
        RECT 75.330 103.980 75.505 104.015 ;
        RECT 74.575 103.445 74.905 103.845 ;
        RECT 75.330 103.615 75.860 103.980 ;
        RECT 76.050 103.615 76.325 104.465 ;
        RECT 76.495 103.615 76.685 104.975 ;
        RECT 76.855 104.990 77.025 105.655 ;
        RECT 77.195 105.235 77.365 105.995 ;
        RECT 77.600 105.235 78.115 105.645 ;
        RECT 76.855 104.800 77.605 104.990 ;
        RECT 77.775 104.425 78.115 105.235 ;
        RECT 78.285 104.905 79.495 105.995 ;
        RECT 76.885 104.255 78.115 104.425 ;
        RECT 76.865 103.445 77.375 103.980 ;
        RECT 77.595 103.650 77.840 104.255 ;
        RECT 78.285 104.195 78.805 104.735 ;
        RECT 78.975 104.365 79.495 104.905 ;
        RECT 79.755 105.065 79.925 105.825 ;
        RECT 80.105 105.235 80.435 105.995 ;
        RECT 79.755 104.895 80.420 105.065 ;
        RECT 80.605 104.920 80.875 105.825 ;
        RECT 80.250 104.750 80.420 104.895 ;
        RECT 79.685 104.345 80.015 104.715 ;
        RECT 80.250 104.420 80.535 104.750 ;
        RECT 78.285 103.445 79.495 104.195 ;
        RECT 80.250 104.165 80.420 104.420 ;
        RECT 79.755 103.995 80.420 104.165 ;
        RECT 80.705 104.120 80.875 104.920 ;
        RECT 81.045 104.905 82.715 105.995 ;
        RECT 79.755 103.615 79.925 103.995 ;
        RECT 80.105 103.445 80.435 103.825 ;
        RECT 80.615 103.615 80.875 104.120 ;
        RECT 81.045 104.215 81.795 104.735 ;
        RECT 81.965 104.385 82.715 104.905 ;
        RECT 82.885 104.905 84.095 105.995 ;
        RECT 82.885 104.365 83.405 104.905 ;
        RECT 81.045 103.445 82.715 104.215 ;
        RECT 83.575 104.195 84.095 104.735 ;
        RECT 82.885 103.445 84.095 104.195 ;
        RECT 5.520 103.275 84.180 103.445 ;
        RECT 5.605 102.525 6.815 103.275 ;
        RECT 7.450 102.800 7.785 103.060 ;
        RECT 7.955 102.875 8.285 103.275 ;
        RECT 8.455 102.875 10.070 103.045 ;
        RECT 5.605 101.985 6.125 102.525 ;
        RECT 6.295 101.815 6.815 102.355 ;
        RECT 5.605 100.725 6.815 101.815 ;
        RECT 7.450 101.445 7.705 102.800 ;
        RECT 8.455 102.705 8.625 102.875 ;
        RECT 8.065 102.535 8.625 102.705 ;
        RECT 8.890 102.595 9.160 102.695 ;
        RECT 9.350 102.595 9.640 102.695 ;
        RECT 8.065 102.365 8.235 102.535 ;
        RECT 8.885 102.425 9.160 102.595 ;
        RECT 9.345 102.425 9.640 102.595 ;
        RECT 7.930 102.035 8.235 102.365 ;
        RECT 8.430 102.255 8.680 102.365 ;
        RECT 8.425 102.085 8.680 102.255 ;
        RECT 8.430 102.035 8.680 102.085 ;
        RECT 8.890 102.035 9.160 102.425 ;
        RECT 9.350 102.035 9.640 102.425 ;
        RECT 9.810 102.035 10.230 102.700 ;
        RECT 10.615 102.555 10.945 103.275 ;
        RECT 11.130 102.435 11.390 103.275 ;
        RECT 11.565 102.530 11.820 103.105 ;
        RECT 11.990 102.895 12.320 103.275 ;
        RECT 12.535 102.725 12.705 103.105 ;
        RECT 11.990 102.555 12.705 102.725 ;
        RECT 10.540 102.255 10.890 102.365 ;
        RECT 10.540 102.085 10.895 102.255 ;
        RECT 10.540 102.035 10.890 102.085 ;
        RECT 8.065 101.865 8.235 102.035 ;
        RECT 8.065 101.695 10.435 101.865 ;
        RECT 10.685 101.745 10.890 102.035 ;
        RECT 7.450 100.935 7.785 101.445 ;
        RECT 8.035 100.725 8.365 101.525 ;
        RECT 8.610 101.315 10.035 101.485 ;
        RECT 8.610 100.895 8.895 101.315 ;
        RECT 9.150 100.725 9.480 101.145 ;
        RECT 9.705 101.065 10.035 101.315 ;
        RECT 10.265 101.235 10.435 101.695 ;
        RECT 10.695 101.065 10.865 101.565 ;
        RECT 9.705 100.895 10.865 101.065 ;
        RECT 11.130 100.725 11.390 101.875 ;
        RECT 11.565 101.800 11.735 102.530 ;
        RECT 11.990 102.365 12.160 102.555 ;
        RECT 13.885 102.475 14.195 103.275 ;
        RECT 14.400 102.475 15.095 103.105 ;
        RECT 15.355 102.725 15.525 103.105 ;
        RECT 15.705 102.895 16.035 103.275 ;
        RECT 15.355 102.555 16.020 102.725 ;
        RECT 16.215 102.600 16.475 103.105 ;
        RECT 17.195 102.935 17.365 102.970 ;
        RECT 17.165 102.765 17.365 102.935 ;
        RECT 11.905 102.035 12.160 102.365 ;
        RECT 11.990 101.825 12.160 102.035 ;
        RECT 12.440 102.005 12.795 102.375 ;
        RECT 13.895 102.035 14.230 102.305 ;
        RECT 14.400 101.915 14.570 102.475 ;
        RECT 14.740 102.035 15.075 102.285 ;
        RECT 15.285 102.005 15.625 102.375 ;
        RECT 15.850 102.300 16.020 102.555 ;
        RECT 15.850 101.970 16.125 102.300 ;
        RECT 14.400 101.875 14.575 101.915 ;
        RECT 11.565 100.895 11.820 101.800 ;
        RECT 11.990 101.655 12.705 101.825 ;
        RECT 11.990 100.725 12.320 101.485 ;
        RECT 12.535 100.895 12.705 101.655 ;
        RECT 13.885 100.725 14.165 101.865 ;
        RECT 14.335 100.895 14.665 101.875 ;
        RECT 14.835 100.725 15.095 101.865 ;
        RECT 15.850 101.825 16.020 101.970 ;
        RECT 15.345 101.655 16.020 101.825 ;
        RECT 16.295 101.800 16.475 102.600 ;
        RECT 17.195 102.405 17.365 102.765 ;
        RECT 17.555 102.745 17.785 103.050 ;
        RECT 17.955 102.915 18.285 103.275 ;
        RECT 18.480 102.745 18.770 103.095 ;
        RECT 17.555 102.575 18.770 102.745 ;
        RECT 18.945 102.525 20.155 103.275 ;
        RECT 20.325 102.535 20.710 103.105 ;
        RECT 20.880 102.815 21.205 103.275 ;
        RECT 21.725 102.645 22.005 103.105 ;
        RECT 17.195 102.235 17.715 102.405 ;
        RECT 15.345 100.895 15.525 101.655 ;
        RECT 15.705 100.725 16.035 101.485 ;
        RECT 16.205 100.895 16.475 101.800 ;
        RECT 17.110 101.705 17.355 102.065 ;
        RECT 17.545 101.855 17.715 102.235 ;
        RECT 17.885 102.035 18.270 102.365 ;
        RECT 18.450 102.255 18.710 102.365 ;
        RECT 18.450 102.085 18.715 102.255 ;
        RECT 18.450 102.035 18.710 102.085 ;
        RECT 17.545 101.575 17.895 101.855 ;
        RECT 17.110 100.725 17.365 101.525 ;
        RECT 17.565 100.895 17.895 101.575 ;
        RECT 18.075 100.985 18.270 102.035 ;
        RECT 18.945 101.985 19.465 102.525 ;
        RECT 18.450 100.725 18.770 101.865 ;
        RECT 19.635 101.815 20.155 102.355 ;
        RECT 18.945 100.725 20.155 101.815 ;
        RECT 20.325 101.865 20.605 102.535 ;
        RECT 20.880 102.475 22.005 102.645 ;
        RECT 20.880 102.365 21.330 102.475 ;
        RECT 20.775 102.035 21.330 102.365 ;
        RECT 22.195 102.305 22.595 103.105 ;
        RECT 22.995 102.815 23.265 103.275 ;
        RECT 23.435 102.645 23.720 103.105 ;
        RECT 20.325 100.895 20.710 101.865 ;
        RECT 20.880 101.575 21.330 102.035 ;
        RECT 21.500 101.745 22.595 102.305 ;
        RECT 20.880 101.355 22.005 101.575 ;
        RECT 20.880 100.725 21.205 101.185 ;
        RECT 21.725 100.895 22.005 101.355 ;
        RECT 22.195 100.895 22.595 101.745 ;
        RECT 22.765 102.475 23.720 102.645 ;
        RECT 24.095 102.725 24.265 103.015 ;
        RECT 24.435 102.895 24.765 103.275 ;
        RECT 24.095 102.555 24.760 102.725 ;
        RECT 22.765 101.575 22.975 102.475 ;
        RECT 23.145 101.745 23.835 102.305 ;
        RECT 24.010 101.735 24.360 102.385 ;
        RECT 22.765 101.355 23.720 101.575 ;
        RECT 24.530 101.565 24.760 102.555 ;
        RECT 22.995 100.725 23.265 101.185 ;
        RECT 23.435 100.895 23.720 101.355 ;
        RECT 24.095 101.395 24.760 101.565 ;
        RECT 24.095 100.895 24.265 101.395 ;
        RECT 24.435 100.725 24.765 101.225 ;
        RECT 24.935 100.895 25.120 103.015 ;
        RECT 25.375 102.815 25.625 103.275 ;
        RECT 25.795 102.825 26.130 102.995 ;
        RECT 26.325 102.825 27.000 102.995 ;
        RECT 25.795 102.685 25.965 102.825 ;
        RECT 25.290 101.695 25.570 102.645 ;
        RECT 25.740 102.555 25.965 102.685 ;
        RECT 25.740 101.450 25.910 102.555 ;
        RECT 26.135 102.405 26.660 102.625 ;
        RECT 26.080 101.640 26.320 102.235 ;
        RECT 26.490 101.705 26.660 102.405 ;
        RECT 26.830 102.045 27.000 102.825 ;
        RECT 27.320 102.775 27.690 103.275 ;
        RECT 27.870 102.825 28.275 102.995 ;
        RECT 28.445 102.825 29.230 102.995 ;
        RECT 27.870 102.595 28.040 102.825 ;
        RECT 27.210 102.295 28.040 102.595 ;
        RECT 28.425 102.325 28.890 102.655 ;
        RECT 27.210 102.265 27.410 102.295 ;
        RECT 27.530 102.045 27.700 102.115 ;
        RECT 26.830 101.875 27.700 102.045 ;
        RECT 27.190 101.785 27.700 101.875 ;
        RECT 25.740 101.320 26.045 101.450 ;
        RECT 26.490 101.340 27.020 101.705 ;
        RECT 25.360 100.725 25.625 101.185 ;
        RECT 25.795 100.895 26.045 101.320 ;
        RECT 27.190 101.170 27.360 101.785 ;
        RECT 26.255 101.000 27.360 101.170 ;
        RECT 27.530 100.725 27.700 101.525 ;
        RECT 27.870 101.225 28.040 102.295 ;
        RECT 28.210 101.395 28.400 102.115 ;
        RECT 28.570 101.365 28.890 102.325 ;
        RECT 29.060 102.365 29.230 102.825 ;
        RECT 29.505 102.745 29.715 103.275 ;
        RECT 29.975 102.535 30.305 103.060 ;
        RECT 30.475 102.665 30.645 103.275 ;
        RECT 30.815 102.620 31.145 103.055 ;
        RECT 30.815 102.535 31.195 102.620 ;
        RECT 31.365 102.550 31.655 103.275 ;
        RECT 31.845 102.545 32.135 103.275 ;
        RECT 30.105 102.365 30.305 102.535 ;
        RECT 30.970 102.495 31.195 102.535 ;
        RECT 29.060 102.035 29.935 102.365 ;
        RECT 30.105 102.035 30.855 102.365 ;
        RECT 27.870 100.895 28.120 101.225 ;
        RECT 29.060 101.195 29.230 102.035 ;
        RECT 30.105 101.830 30.295 102.035 ;
        RECT 31.025 101.915 31.195 102.495 ;
        RECT 31.835 102.035 32.135 102.365 ;
        RECT 32.315 102.345 32.545 102.985 ;
        RECT 32.725 102.725 33.035 103.095 ;
        RECT 33.215 102.905 33.885 103.275 ;
        RECT 32.725 102.525 33.955 102.725 ;
        RECT 32.315 102.035 32.840 102.345 ;
        RECT 33.020 102.035 33.485 102.345 ;
        RECT 30.980 101.865 31.195 101.915 ;
        RECT 29.400 101.455 30.295 101.830 ;
        RECT 30.805 101.785 31.195 101.865 ;
        RECT 28.345 101.025 29.230 101.195 ;
        RECT 29.410 100.725 29.725 101.225 ;
        RECT 29.955 100.895 30.295 101.455 ;
        RECT 30.465 100.725 30.635 101.735 ;
        RECT 30.805 100.940 31.135 101.785 ;
        RECT 31.365 100.725 31.655 101.890 ;
        RECT 33.665 101.855 33.955 102.525 ;
        RECT 31.845 101.615 33.005 101.855 ;
        RECT 31.845 100.905 32.105 101.615 ;
        RECT 32.275 100.725 32.605 101.435 ;
        RECT 32.775 100.905 33.005 101.615 ;
        RECT 33.185 101.635 33.955 101.855 ;
        RECT 33.185 100.905 33.455 101.635 ;
        RECT 33.635 100.725 33.975 101.455 ;
        RECT 34.145 100.905 34.405 103.095 ;
        RECT 34.595 102.465 34.865 103.275 ;
        RECT 35.035 102.465 35.365 103.105 ;
        RECT 35.535 102.465 35.775 103.275 ;
        RECT 36.055 102.725 36.225 103.015 ;
        RECT 36.395 102.895 36.725 103.275 ;
        RECT 36.055 102.555 36.720 102.725 ;
        RECT 34.585 102.035 34.935 102.285 ;
        RECT 35.105 101.865 35.275 102.465 ;
        RECT 35.445 102.035 35.795 102.285 ;
        RECT 34.595 100.725 34.925 101.865 ;
        RECT 35.105 101.695 35.785 101.865 ;
        RECT 35.970 101.735 36.320 102.385 ;
        RECT 35.455 100.910 35.785 101.695 ;
        RECT 36.490 101.565 36.720 102.555 ;
        RECT 36.055 101.395 36.720 101.565 ;
        RECT 36.055 100.895 36.225 101.395 ;
        RECT 36.395 100.725 36.725 101.225 ;
        RECT 36.895 100.895 37.080 103.015 ;
        RECT 37.335 102.815 37.585 103.275 ;
        RECT 37.755 102.825 38.090 102.995 ;
        RECT 38.285 102.825 38.960 102.995 ;
        RECT 37.755 102.685 37.925 102.825 ;
        RECT 37.250 101.695 37.530 102.645 ;
        RECT 37.700 102.555 37.925 102.685 ;
        RECT 37.700 101.450 37.870 102.555 ;
        RECT 38.095 102.405 38.620 102.625 ;
        RECT 38.040 101.640 38.280 102.235 ;
        RECT 38.450 101.705 38.620 102.405 ;
        RECT 38.790 102.045 38.960 102.825 ;
        RECT 39.280 102.775 39.650 103.275 ;
        RECT 39.830 102.825 40.235 102.995 ;
        RECT 40.405 102.825 41.190 102.995 ;
        RECT 39.830 102.595 40.000 102.825 ;
        RECT 39.170 102.295 40.000 102.595 ;
        RECT 40.385 102.325 40.850 102.655 ;
        RECT 39.170 102.265 39.370 102.295 ;
        RECT 39.490 102.045 39.660 102.115 ;
        RECT 38.790 101.875 39.660 102.045 ;
        RECT 39.150 101.785 39.660 101.875 ;
        RECT 37.700 101.320 38.005 101.450 ;
        RECT 38.450 101.340 38.980 101.705 ;
        RECT 37.320 100.725 37.585 101.185 ;
        RECT 37.755 100.895 38.005 101.320 ;
        RECT 39.150 101.170 39.320 101.785 ;
        RECT 38.215 101.000 39.320 101.170 ;
        RECT 39.490 100.725 39.660 101.525 ;
        RECT 39.830 101.225 40.000 102.295 ;
        RECT 40.170 101.395 40.360 102.115 ;
        RECT 40.530 101.365 40.850 102.325 ;
        RECT 41.020 102.365 41.190 102.825 ;
        RECT 41.465 102.745 41.675 103.275 ;
        RECT 41.935 102.535 42.265 103.060 ;
        RECT 42.435 102.665 42.605 103.275 ;
        RECT 42.775 102.620 43.105 103.055 ;
        RECT 42.775 102.535 43.155 102.620 ;
        RECT 42.065 102.365 42.265 102.535 ;
        RECT 42.930 102.495 43.155 102.535 ;
        RECT 41.020 102.035 41.895 102.365 ;
        RECT 42.065 102.035 42.815 102.365 ;
        RECT 39.830 100.895 40.080 101.225 ;
        RECT 41.020 101.195 41.190 102.035 ;
        RECT 42.065 101.830 42.255 102.035 ;
        RECT 42.985 101.915 43.155 102.495 ;
        RECT 42.940 101.865 43.155 101.915 ;
        RECT 41.360 101.455 42.255 101.830 ;
        RECT 42.765 101.785 43.155 101.865 ;
        RECT 44.245 102.535 44.630 103.105 ;
        RECT 44.800 102.815 45.125 103.275 ;
        RECT 45.645 102.645 45.925 103.105 ;
        RECT 44.245 101.865 44.525 102.535 ;
        RECT 44.800 102.475 45.925 102.645 ;
        RECT 44.800 102.365 45.250 102.475 ;
        RECT 44.695 102.035 45.250 102.365 ;
        RECT 46.115 102.305 46.515 103.105 ;
        RECT 46.915 102.815 47.185 103.275 ;
        RECT 47.355 102.645 47.640 103.105 ;
        RECT 48.385 102.895 49.275 103.065 ;
        RECT 40.305 101.025 41.190 101.195 ;
        RECT 41.370 100.725 41.685 101.225 ;
        RECT 41.915 100.895 42.255 101.455 ;
        RECT 42.425 100.725 42.595 101.735 ;
        RECT 42.765 100.940 43.095 101.785 ;
        RECT 44.245 100.895 44.630 101.865 ;
        RECT 44.800 101.575 45.250 102.035 ;
        RECT 45.420 101.745 46.515 102.305 ;
        RECT 44.800 101.355 45.925 101.575 ;
        RECT 44.800 100.725 45.125 101.185 ;
        RECT 45.645 100.895 45.925 101.355 ;
        RECT 46.115 100.895 46.515 101.745 ;
        RECT 46.685 102.475 47.640 102.645 ;
        RECT 46.685 101.575 46.895 102.475 ;
        RECT 48.385 102.340 48.935 102.725 ;
        RECT 47.065 101.745 47.755 102.305 ;
        RECT 49.105 102.170 49.275 102.895 ;
        RECT 48.385 102.100 49.275 102.170 ;
        RECT 49.445 102.570 49.665 103.055 ;
        RECT 49.835 102.735 50.085 103.275 ;
        RECT 50.255 102.625 50.515 103.105 ;
        RECT 49.445 102.145 49.775 102.570 ;
        RECT 48.385 102.075 49.280 102.100 ;
        RECT 48.385 102.060 49.290 102.075 ;
        RECT 48.385 102.045 49.295 102.060 ;
        RECT 48.385 102.040 49.305 102.045 ;
        RECT 48.385 102.030 49.310 102.040 ;
        RECT 48.385 102.020 49.315 102.030 ;
        RECT 48.385 102.015 49.325 102.020 ;
        RECT 48.385 102.005 49.335 102.015 ;
        RECT 48.385 102.000 49.345 102.005 ;
        RECT 46.685 101.355 47.640 101.575 ;
        RECT 48.385 101.550 48.645 102.000 ;
        RECT 49.010 101.995 49.345 102.000 ;
        RECT 49.010 101.990 49.360 101.995 ;
        RECT 49.010 101.980 49.375 101.990 ;
        RECT 49.010 101.975 49.400 101.980 ;
        RECT 49.945 101.975 50.175 102.370 ;
        RECT 49.010 101.970 50.175 101.975 ;
        RECT 49.040 101.935 50.175 101.970 ;
        RECT 49.075 101.910 50.175 101.935 ;
        RECT 49.105 101.880 50.175 101.910 ;
        RECT 49.125 101.850 50.175 101.880 ;
        RECT 49.145 101.820 50.175 101.850 ;
        RECT 49.215 101.810 50.175 101.820 ;
        RECT 49.240 101.800 50.175 101.810 ;
        RECT 49.260 101.785 50.175 101.800 ;
        RECT 49.280 101.770 50.175 101.785 ;
        RECT 49.285 101.760 50.070 101.770 ;
        RECT 49.300 101.725 50.070 101.760 ;
        RECT 48.815 101.405 49.145 101.650 ;
        RECT 49.315 101.475 50.070 101.725 ;
        RECT 50.345 101.595 50.515 102.625 ;
        RECT 50.800 102.645 51.085 103.105 ;
        RECT 51.255 102.815 51.525 103.275 ;
        RECT 50.800 102.475 51.755 102.645 ;
        RECT 50.685 101.745 51.375 102.305 ;
        RECT 48.815 101.380 49.000 101.405 ;
        RECT 46.915 100.725 47.185 101.185 ;
        RECT 47.355 100.895 47.640 101.355 ;
        RECT 48.385 101.280 49.000 101.380 ;
        RECT 48.385 100.725 48.990 101.280 ;
        RECT 49.165 100.895 49.645 101.235 ;
        RECT 49.815 100.725 50.070 101.270 ;
        RECT 50.240 100.895 50.515 101.595 ;
        RECT 51.545 101.575 51.755 102.475 ;
        RECT 50.800 101.355 51.755 101.575 ;
        RECT 51.925 102.305 52.325 103.105 ;
        RECT 52.515 102.645 52.795 103.105 ;
        RECT 53.315 102.815 53.640 103.275 ;
        RECT 52.515 102.475 53.640 102.645 ;
        RECT 53.810 102.535 54.195 103.105 ;
        RECT 53.190 102.365 53.640 102.475 ;
        RECT 51.925 101.745 53.020 102.305 ;
        RECT 53.190 102.035 53.745 102.365 ;
        RECT 50.800 100.895 51.085 101.355 ;
        RECT 51.255 100.725 51.525 101.185 ;
        RECT 51.925 100.895 52.325 101.745 ;
        RECT 53.190 101.575 53.640 102.035 ;
        RECT 53.915 101.865 54.195 102.535 ;
        RECT 54.365 102.505 56.955 103.275 ;
        RECT 57.125 102.550 57.415 103.275 ;
        RECT 57.590 102.745 57.880 103.095 ;
        RECT 58.075 102.915 58.405 103.275 ;
        RECT 58.575 102.745 58.805 103.050 ;
        RECT 57.590 102.575 58.805 102.745 ;
        RECT 54.365 101.985 55.575 102.505 ;
        RECT 58.995 102.405 59.165 102.970 ;
        RECT 59.425 102.730 64.770 103.275 ;
        RECT 65.425 102.765 65.665 103.275 ;
        RECT 65.835 102.765 66.125 103.105 ;
        RECT 66.355 102.765 66.670 103.275 ;
        RECT 52.515 101.355 53.640 101.575 ;
        RECT 52.515 100.895 52.795 101.355 ;
        RECT 53.315 100.725 53.640 101.185 ;
        RECT 53.810 100.895 54.195 101.865 ;
        RECT 55.745 101.815 56.955 102.335 ;
        RECT 57.650 102.255 57.910 102.365 ;
        RECT 57.645 102.085 57.910 102.255 ;
        RECT 57.650 102.035 57.910 102.085 ;
        RECT 58.090 102.035 58.475 102.365 ;
        RECT 58.645 102.235 59.165 102.405 ;
        RECT 54.365 100.725 56.955 101.815 ;
        RECT 57.125 100.725 57.415 101.890 ;
        RECT 57.590 100.725 57.910 101.865 ;
        RECT 58.090 100.985 58.285 102.035 ;
        RECT 58.645 101.855 58.815 102.235 ;
        RECT 58.465 101.575 58.815 101.855 ;
        RECT 59.005 101.705 59.250 102.065 ;
        RECT 61.010 101.900 61.350 102.730 ;
        RECT 58.465 100.895 58.795 101.575 ;
        RECT 58.995 100.725 59.250 101.525 ;
        RECT 62.830 101.160 63.180 102.410 ;
        RECT 65.470 102.255 65.665 102.595 ;
        RECT 65.465 102.085 65.665 102.255 ;
        RECT 65.470 102.035 65.665 102.085 ;
        RECT 65.835 101.865 66.015 102.765 ;
        RECT 66.840 102.705 67.010 102.975 ;
        RECT 67.180 102.875 67.510 103.275 ;
        RECT 66.185 102.035 66.595 102.595 ;
        RECT 66.840 102.535 67.535 102.705 ;
        RECT 66.765 101.865 66.935 102.365 ;
        RECT 65.475 101.695 66.935 101.865 ;
        RECT 65.475 101.520 65.835 101.695 ;
        RECT 67.105 101.525 67.535 102.535 ;
        RECT 67.910 102.495 68.410 103.105 ;
        RECT 67.705 102.035 68.055 102.285 ;
        RECT 68.240 101.865 68.410 102.495 ;
        RECT 69.040 102.625 69.370 103.105 ;
        RECT 69.540 102.815 69.765 103.275 ;
        RECT 69.935 102.625 70.265 103.105 ;
        RECT 69.040 102.455 70.265 102.625 ;
        RECT 70.455 102.475 70.705 103.275 ;
        RECT 70.875 102.475 71.215 103.105 ;
        RECT 68.580 102.085 68.910 102.285 ;
        RECT 69.080 102.085 69.410 102.285 ;
        RECT 69.580 102.085 70.000 102.285 ;
        RECT 70.175 102.115 70.870 102.285 ;
        RECT 70.175 101.865 70.345 102.115 ;
        RECT 71.040 101.865 71.215 102.475 ;
        RECT 71.390 102.435 71.650 103.275 ;
        RECT 71.825 102.530 72.080 103.105 ;
        RECT 72.250 102.895 72.580 103.275 ;
        RECT 72.795 102.725 72.965 103.105 ;
        RECT 72.250 102.555 72.965 102.725 ;
        RECT 59.425 100.725 64.770 101.160 ;
        RECT 66.420 100.725 66.590 101.525 ;
        RECT 66.760 101.355 67.535 101.525 ;
        RECT 67.910 101.695 70.345 101.865 ;
        RECT 66.760 100.895 67.090 101.355 ;
        RECT 67.260 100.725 67.430 101.185 ;
        RECT 67.910 100.895 68.240 101.695 ;
        RECT 68.410 100.725 68.740 101.525 ;
        RECT 69.040 100.895 69.370 101.695 ;
        RECT 70.015 100.725 70.265 101.525 ;
        RECT 70.535 100.725 70.705 101.865 ;
        RECT 70.875 100.895 71.215 101.865 ;
        RECT 71.390 100.725 71.650 101.875 ;
        RECT 71.825 101.800 71.995 102.530 ;
        RECT 72.250 102.365 72.420 102.555 ;
        RECT 73.225 102.505 76.735 103.275 ;
        RECT 76.905 102.525 78.115 103.275 ;
        RECT 78.285 102.535 78.670 103.105 ;
        RECT 78.840 102.815 79.165 103.275 ;
        RECT 79.685 102.645 79.965 103.105 ;
        RECT 72.165 102.035 72.420 102.365 ;
        RECT 72.250 101.825 72.420 102.035 ;
        RECT 72.700 102.005 73.055 102.375 ;
        RECT 73.225 101.985 74.875 102.505 ;
        RECT 71.825 100.895 72.080 101.800 ;
        RECT 72.250 101.655 72.965 101.825 ;
        RECT 75.045 101.815 76.735 102.335 ;
        RECT 76.905 101.985 77.425 102.525 ;
        RECT 77.595 101.815 78.115 102.355 ;
        RECT 72.250 100.725 72.580 101.485 ;
        RECT 72.795 100.895 72.965 101.655 ;
        RECT 73.225 100.725 76.735 101.815 ;
        RECT 76.905 100.725 78.115 101.815 ;
        RECT 78.285 101.865 78.565 102.535 ;
        RECT 78.840 102.475 79.965 102.645 ;
        RECT 78.840 102.365 79.290 102.475 ;
        RECT 78.735 102.035 79.290 102.365 ;
        RECT 80.155 102.305 80.555 103.105 ;
        RECT 80.955 102.815 81.225 103.275 ;
        RECT 81.395 102.645 81.680 103.105 ;
        RECT 78.285 100.895 78.670 101.865 ;
        RECT 78.840 101.575 79.290 102.035 ;
        RECT 79.460 101.745 80.555 102.305 ;
        RECT 78.840 101.355 79.965 101.575 ;
        RECT 78.840 100.725 79.165 101.185 ;
        RECT 79.685 100.895 79.965 101.355 ;
        RECT 80.155 100.895 80.555 101.745 ;
        RECT 80.725 102.475 81.680 102.645 ;
        RECT 82.885 102.525 84.095 103.275 ;
        RECT 80.725 101.575 80.935 102.475 ;
        RECT 81.105 101.745 81.795 102.305 ;
        RECT 82.885 101.815 83.405 102.355 ;
        RECT 83.575 101.985 84.095 102.525 ;
        RECT 80.725 101.355 81.680 101.575 ;
        RECT 80.955 100.725 81.225 101.185 ;
        RECT 81.395 100.895 81.680 101.355 ;
        RECT 82.885 100.725 84.095 101.815 ;
        RECT 5.520 100.555 84.180 100.725 ;
        RECT 5.605 99.465 6.815 100.555 ;
        RECT 5.605 98.755 6.125 99.295 ;
        RECT 6.295 98.925 6.815 99.465 ;
        RECT 6.985 99.585 7.255 100.355 ;
        RECT 7.425 99.775 7.755 100.555 ;
        RECT 7.960 99.950 8.145 100.355 ;
        RECT 8.315 100.130 8.650 100.555 ;
        RECT 7.960 99.775 8.625 99.950 ;
        RECT 6.985 99.415 8.115 99.585 ;
        RECT 5.605 98.005 6.815 98.755 ;
        RECT 6.985 98.505 7.155 99.415 ;
        RECT 7.325 98.665 7.685 99.245 ;
        RECT 7.865 98.915 8.115 99.415 ;
        RECT 8.285 98.745 8.625 99.775 ;
        RECT 9.745 99.415 10.025 100.555 ;
        RECT 10.195 99.405 10.525 100.385 ;
        RECT 10.695 99.415 10.955 100.555 ;
        RECT 11.240 99.925 11.525 100.385 ;
        RECT 11.695 100.095 11.965 100.555 ;
        RECT 11.240 99.705 12.195 99.925 ;
        RECT 9.755 98.975 10.090 99.245 ;
        RECT 10.260 98.805 10.430 99.405 ;
        RECT 10.600 98.995 10.935 99.245 ;
        RECT 11.125 98.975 11.815 99.535 ;
        RECT 11.985 98.805 12.195 99.705 ;
        RECT 7.940 98.575 8.625 98.745 ;
        RECT 6.985 98.175 7.245 98.505 ;
        RECT 7.455 98.005 7.730 98.485 ;
        RECT 7.940 98.175 8.145 98.575 ;
        RECT 8.315 98.005 8.650 98.405 ;
        RECT 9.745 98.005 10.055 98.805 ;
        RECT 10.260 98.175 10.955 98.805 ;
        RECT 11.240 98.635 12.195 98.805 ;
        RECT 12.365 99.535 12.765 100.385 ;
        RECT 12.955 99.925 13.235 100.385 ;
        RECT 13.755 100.095 14.080 100.555 ;
        RECT 12.955 99.705 14.080 99.925 ;
        RECT 12.365 98.975 13.460 99.535 ;
        RECT 13.630 99.245 14.080 99.705 ;
        RECT 14.250 99.415 14.635 100.385 ;
        RECT 15.265 100.045 15.565 100.555 ;
        RECT 15.735 99.875 16.065 100.385 ;
        RECT 16.235 100.045 16.865 100.555 ;
        RECT 17.445 100.045 17.825 100.215 ;
        RECT 17.995 100.045 18.295 100.555 ;
        RECT 17.655 99.875 17.825 100.045 ;
        RECT 11.240 98.175 11.525 98.635 ;
        RECT 11.695 98.005 11.965 98.465 ;
        RECT 12.365 98.175 12.765 98.975 ;
        RECT 13.630 98.915 14.185 99.245 ;
        RECT 13.630 98.805 14.080 98.915 ;
        RECT 12.955 98.635 14.080 98.805 ;
        RECT 14.355 98.745 14.635 99.415 ;
        RECT 12.955 98.175 13.235 98.635 ;
        RECT 13.755 98.005 14.080 98.465 ;
        RECT 14.250 98.175 14.635 98.745 ;
        RECT 15.265 99.705 17.485 99.875 ;
        RECT 15.265 98.745 15.435 99.705 ;
        RECT 15.605 99.365 17.145 99.535 ;
        RECT 15.605 98.915 15.850 99.365 ;
        RECT 16.110 98.995 16.805 99.195 ;
        RECT 16.975 99.165 17.145 99.365 ;
        RECT 17.315 99.505 17.485 99.705 ;
        RECT 17.655 99.675 18.315 99.875 ;
        RECT 17.315 99.335 17.975 99.505 ;
        RECT 16.975 98.995 17.575 99.165 ;
        RECT 17.805 98.915 17.975 99.335 ;
        RECT 15.265 98.200 15.730 98.745 ;
        RECT 16.235 98.005 16.405 98.825 ;
        RECT 16.575 98.745 17.485 98.825 ;
        RECT 18.145 98.745 18.315 99.675 ;
        RECT 18.485 99.390 18.775 100.555 ;
        RECT 19.035 99.885 19.205 100.385 ;
        RECT 19.375 100.055 19.705 100.555 ;
        RECT 19.035 99.715 19.700 99.885 ;
        RECT 18.950 98.895 19.300 99.545 ;
        RECT 16.575 98.655 17.825 98.745 ;
        RECT 16.575 98.175 16.905 98.655 ;
        RECT 17.315 98.575 17.825 98.655 ;
        RECT 17.075 98.005 17.425 98.395 ;
        RECT 17.595 98.175 17.825 98.575 ;
        RECT 17.995 98.265 18.315 98.745 ;
        RECT 18.485 98.005 18.775 98.730 ;
        RECT 19.470 98.725 19.700 99.715 ;
        RECT 19.035 98.555 19.700 98.725 ;
        RECT 19.035 98.265 19.205 98.555 ;
        RECT 19.375 98.005 19.705 98.385 ;
        RECT 19.875 98.265 20.060 100.385 ;
        RECT 20.300 100.095 20.565 100.555 ;
        RECT 20.735 99.960 20.985 100.385 ;
        RECT 21.195 100.110 22.300 100.280 ;
        RECT 20.680 99.830 20.985 99.960 ;
        RECT 20.230 98.635 20.510 99.585 ;
        RECT 20.680 98.725 20.850 99.830 ;
        RECT 21.020 99.045 21.260 99.640 ;
        RECT 21.430 99.575 21.960 99.940 ;
        RECT 21.430 98.875 21.600 99.575 ;
        RECT 22.130 99.495 22.300 100.110 ;
        RECT 22.470 99.755 22.640 100.555 ;
        RECT 22.810 100.055 23.060 100.385 ;
        RECT 23.285 100.085 24.170 100.255 ;
        RECT 22.130 99.405 22.640 99.495 ;
        RECT 20.680 98.595 20.905 98.725 ;
        RECT 21.075 98.655 21.600 98.875 ;
        RECT 21.770 99.235 22.640 99.405 ;
        RECT 20.315 98.005 20.565 98.465 ;
        RECT 20.735 98.455 20.905 98.595 ;
        RECT 21.770 98.455 21.940 99.235 ;
        RECT 22.470 99.165 22.640 99.235 ;
        RECT 22.150 98.985 22.350 99.015 ;
        RECT 22.810 98.985 22.980 100.055 ;
        RECT 23.150 99.165 23.340 99.885 ;
        RECT 22.150 98.685 22.980 98.985 ;
        RECT 23.510 98.955 23.830 99.915 ;
        RECT 20.735 98.285 21.070 98.455 ;
        RECT 21.265 98.285 21.940 98.455 ;
        RECT 22.260 98.005 22.630 98.505 ;
        RECT 22.810 98.455 22.980 98.685 ;
        RECT 23.365 98.625 23.830 98.955 ;
        RECT 24.000 99.245 24.170 100.085 ;
        RECT 24.350 100.055 24.665 100.555 ;
        RECT 24.895 99.825 25.235 100.385 ;
        RECT 24.340 99.450 25.235 99.825 ;
        RECT 25.405 99.545 25.575 100.555 ;
        RECT 25.045 99.245 25.235 99.450 ;
        RECT 25.745 99.495 26.075 100.340 ;
        RECT 25.745 99.415 26.135 99.495 ;
        RECT 26.305 99.465 29.815 100.555 ;
        RECT 25.920 99.365 26.135 99.415 ;
        RECT 24.000 98.915 24.875 99.245 ;
        RECT 25.045 98.915 25.795 99.245 ;
        RECT 24.000 98.455 24.170 98.915 ;
        RECT 25.045 98.745 25.245 98.915 ;
        RECT 25.965 98.785 26.135 99.365 ;
        RECT 25.910 98.745 26.135 98.785 ;
        RECT 22.810 98.285 23.215 98.455 ;
        RECT 23.385 98.285 24.170 98.455 ;
        RECT 24.445 98.005 24.655 98.535 ;
        RECT 24.915 98.220 25.245 98.745 ;
        RECT 25.755 98.660 26.135 98.745 ;
        RECT 26.305 98.775 27.955 99.295 ;
        RECT 28.125 98.945 29.815 99.465 ;
        RECT 30.445 99.415 30.705 100.555 ;
        RECT 30.875 99.405 31.205 100.385 ;
        RECT 31.375 99.415 31.655 100.555 ;
        RECT 32.290 99.605 32.555 100.375 ;
        RECT 32.725 99.835 33.055 100.555 ;
        RECT 33.245 100.015 33.505 100.375 ;
        RECT 33.675 100.185 34.005 100.555 ;
        RECT 34.175 100.015 34.435 100.375 ;
        RECT 33.245 99.785 34.435 100.015 ;
        RECT 35.005 99.605 35.295 100.375 ;
        RECT 30.465 98.995 30.800 99.245 ;
        RECT 30.970 98.805 31.140 99.405 ;
        RECT 31.310 98.975 31.645 99.245 ;
        RECT 25.415 98.005 25.585 98.615 ;
        RECT 25.755 98.225 26.085 98.660 ;
        RECT 26.305 98.005 29.815 98.775 ;
        RECT 30.445 98.175 31.140 98.805 ;
        RECT 31.345 98.005 31.655 98.805 ;
        RECT 32.290 98.185 32.625 99.605 ;
        RECT 32.800 99.425 35.295 99.605 ;
        RECT 32.800 98.735 33.025 99.425 ;
        RECT 35.505 99.415 35.795 100.555 ;
        RECT 36.590 100.215 37.955 100.385 ;
        RECT 36.590 100.005 36.920 100.215 ;
        RECT 35.965 99.755 36.920 100.005 ;
        RECT 33.225 98.915 33.505 99.245 ;
        RECT 33.685 98.915 34.260 99.245 ;
        RECT 34.440 98.915 34.875 99.245 ;
        RECT 35.055 98.915 35.325 99.245 ;
        RECT 35.505 98.915 35.780 99.245 ;
        RECT 35.965 98.745 36.135 99.755 ;
        RECT 36.305 98.915 36.660 99.580 ;
        RECT 36.845 98.915 37.120 99.580 ;
        RECT 37.290 99.245 37.615 100.045 ;
        RECT 37.785 99.585 37.955 100.215 ;
        RECT 38.125 99.755 38.415 100.555 ;
        RECT 37.785 99.415 38.460 99.585 ;
        RECT 38.630 99.415 39.015 100.375 ;
        RECT 39.185 99.465 42.695 100.555 ;
        RECT 38.290 99.245 38.460 99.415 ;
        RECT 37.290 98.915 37.635 99.245 ;
        RECT 37.845 98.995 38.095 99.245 ;
        RECT 38.290 98.995 38.655 99.245 ;
        RECT 37.925 98.915 38.095 98.995 ;
        RECT 38.465 98.915 38.655 98.995 ;
        RECT 38.840 98.745 39.015 99.415 ;
        RECT 32.800 98.545 35.285 98.735 ;
        RECT 32.805 98.005 33.550 98.375 ;
        RECT 34.115 98.185 34.370 98.545 ;
        RECT 34.550 98.005 34.880 98.375 ;
        RECT 35.060 98.185 35.285 98.545 ;
        RECT 35.505 98.385 35.795 98.655 ;
        RECT 35.965 98.555 36.390 98.745 ;
        RECT 36.560 98.575 37.960 98.745 ;
        RECT 36.560 98.385 36.890 98.575 ;
        RECT 35.505 98.175 36.890 98.385 ;
        RECT 37.125 98.005 37.455 98.405 ;
        RECT 37.630 98.175 37.960 98.575 ;
        RECT 38.165 98.005 38.335 98.565 ;
        RECT 38.505 98.175 39.015 98.745 ;
        RECT 39.185 98.775 40.835 99.295 ;
        RECT 41.005 98.945 42.695 99.465 ;
        RECT 42.925 99.415 43.135 100.555 ;
        RECT 43.305 99.405 43.635 100.385 ;
        RECT 43.805 99.415 44.035 100.555 ;
        RECT 39.185 98.005 42.695 98.775 ;
        RECT 42.925 98.005 43.135 98.825 ;
        RECT 43.305 98.805 43.555 99.405 ;
        RECT 44.245 99.390 44.535 100.555 ;
        RECT 45.685 99.495 46.015 100.340 ;
        RECT 46.185 99.545 46.355 100.555 ;
        RECT 46.525 99.825 46.865 100.385 ;
        RECT 47.095 100.055 47.410 100.555 ;
        RECT 47.590 100.085 48.475 100.255 ;
        RECT 45.625 99.415 46.015 99.495 ;
        RECT 46.525 99.450 47.420 99.825 ;
        RECT 45.625 99.365 45.840 99.415 ;
        RECT 43.725 98.995 44.055 99.245 ;
        RECT 43.305 98.175 43.635 98.805 ;
        RECT 43.805 98.005 44.035 98.825 ;
        RECT 45.625 98.785 45.795 99.365 ;
        RECT 46.525 99.245 46.715 99.450 ;
        RECT 47.590 99.245 47.760 100.085 ;
        RECT 48.700 100.055 48.950 100.385 ;
        RECT 45.965 98.915 46.715 99.245 ;
        RECT 46.885 98.915 47.760 99.245 ;
        RECT 45.625 98.745 45.850 98.785 ;
        RECT 46.515 98.745 46.715 98.915 ;
        RECT 44.245 98.005 44.535 98.730 ;
        RECT 45.625 98.660 46.005 98.745 ;
        RECT 45.675 98.225 46.005 98.660 ;
        RECT 46.175 98.005 46.345 98.615 ;
        RECT 46.515 98.220 46.845 98.745 ;
        RECT 47.105 98.005 47.315 98.535 ;
        RECT 47.590 98.455 47.760 98.915 ;
        RECT 47.930 98.955 48.250 99.915 ;
        RECT 48.420 99.165 48.610 99.885 ;
        RECT 48.780 98.985 48.950 100.055 ;
        RECT 49.120 99.755 49.290 100.555 ;
        RECT 49.460 100.110 50.565 100.280 ;
        RECT 49.460 99.495 49.630 100.110 ;
        RECT 50.775 99.960 51.025 100.385 ;
        RECT 51.195 100.095 51.460 100.555 ;
        RECT 49.800 99.575 50.330 99.940 ;
        RECT 50.775 99.830 51.080 99.960 ;
        RECT 49.120 99.405 49.630 99.495 ;
        RECT 49.120 99.235 49.990 99.405 ;
        RECT 49.120 99.165 49.290 99.235 ;
        RECT 49.410 98.985 49.610 99.015 ;
        RECT 47.930 98.625 48.395 98.955 ;
        RECT 48.780 98.685 49.610 98.985 ;
        RECT 48.780 98.455 48.950 98.685 ;
        RECT 47.590 98.285 48.375 98.455 ;
        RECT 48.545 98.285 48.950 98.455 ;
        RECT 49.130 98.005 49.500 98.505 ;
        RECT 49.820 98.455 49.990 99.235 ;
        RECT 50.160 98.875 50.330 99.575 ;
        RECT 50.500 99.045 50.740 99.640 ;
        RECT 50.160 98.655 50.685 98.875 ;
        RECT 50.910 98.725 51.080 99.830 ;
        RECT 50.855 98.595 51.080 98.725 ;
        RECT 51.250 98.635 51.530 99.585 ;
        RECT 50.855 98.455 51.025 98.595 ;
        RECT 49.820 98.285 50.495 98.455 ;
        RECT 50.690 98.285 51.025 98.455 ;
        RECT 51.195 98.005 51.445 98.465 ;
        RECT 51.700 98.265 51.885 100.385 ;
        RECT 52.055 100.055 52.385 100.555 ;
        RECT 52.555 99.885 52.725 100.385 ;
        RECT 52.060 99.715 52.725 99.885 ;
        RECT 52.060 98.725 52.290 99.715 ;
        RECT 52.460 98.895 52.810 99.545 ;
        RECT 52.990 99.415 53.325 100.385 ;
        RECT 53.495 99.415 53.665 100.555 ;
        RECT 53.835 100.215 55.865 100.385 ;
        RECT 52.990 98.745 53.160 99.415 ;
        RECT 53.835 99.245 54.005 100.215 ;
        RECT 53.330 98.915 53.585 99.245 ;
        RECT 53.810 98.915 54.005 99.245 ;
        RECT 54.175 99.875 55.300 100.045 ;
        RECT 53.415 98.745 53.585 98.915 ;
        RECT 54.175 98.745 54.345 99.875 ;
        RECT 52.060 98.555 52.725 98.725 ;
        RECT 52.055 98.005 52.385 98.385 ;
        RECT 52.555 98.265 52.725 98.555 ;
        RECT 52.990 98.175 53.245 98.745 ;
        RECT 53.415 98.575 54.345 98.745 ;
        RECT 54.515 99.535 55.525 99.705 ;
        RECT 54.515 98.735 54.685 99.535 ;
        RECT 54.890 98.855 55.165 99.335 ;
        RECT 54.885 98.685 55.165 98.855 ;
        RECT 54.170 98.540 54.345 98.575 ;
        RECT 53.415 98.005 53.745 98.405 ;
        RECT 54.170 98.175 54.700 98.540 ;
        RECT 54.890 98.175 55.165 98.685 ;
        RECT 55.335 98.175 55.525 99.535 ;
        RECT 55.695 99.550 55.865 100.215 ;
        RECT 56.035 99.795 56.205 100.555 ;
        RECT 56.440 99.795 56.955 100.205 ;
        RECT 55.695 99.360 56.445 99.550 ;
        RECT 56.615 98.985 56.955 99.795 ;
        RECT 57.215 99.625 57.385 100.385 ;
        RECT 57.600 99.795 57.930 100.555 ;
        RECT 57.215 99.455 57.930 99.625 ;
        RECT 58.100 99.480 58.355 100.385 ;
        RECT 55.725 98.815 56.955 98.985 ;
        RECT 57.125 98.905 57.480 99.275 ;
        RECT 57.760 99.245 57.930 99.455 ;
        RECT 57.760 98.915 58.015 99.245 ;
        RECT 55.705 98.005 56.215 98.540 ;
        RECT 56.435 98.210 56.680 98.815 ;
        RECT 57.760 98.725 57.930 98.915 ;
        RECT 58.185 98.750 58.355 99.480 ;
        RECT 58.530 99.405 58.790 100.555 ;
        RECT 58.975 99.585 59.305 100.370 ;
        RECT 58.975 99.415 59.655 99.585 ;
        RECT 59.835 99.415 60.165 100.555 ;
        RECT 60.345 99.465 63.855 100.555 ;
        RECT 58.965 98.995 59.315 99.245 ;
        RECT 57.215 98.555 57.930 98.725 ;
        RECT 57.215 98.175 57.385 98.555 ;
        RECT 57.600 98.005 57.930 98.385 ;
        RECT 58.100 98.175 58.355 98.750 ;
        RECT 58.530 98.005 58.790 98.845 ;
        RECT 59.485 98.815 59.655 99.415 ;
        RECT 59.825 98.995 60.175 99.245 ;
        RECT 58.985 98.005 59.225 98.815 ;
        RECT 59.395 98.175 59.725 98.815 ;
        RECT 59.895 98.005 60.165 98.815 ;
        RECT 60.345 98.775 61.995 99.295 ;
        RECT 62.165 98.945 63.855 99.465 ;
        RECT 64.945 99.415 65.205 100.555 ;
        RECT 65.375 99.405 65.705 100.385 ;
        RECT 65.875 99.415 66.155 100.555 ;
        RECT 65.465 99.365 65.640 99.405 ;
        RECT 66.325 99.375 66.645 100.555 ;
        RECT 66.815 99.535 67.015 100.325 ;
        RECT 67.340 99.725 67.725 100.385 ;
        RECT 68.120 99.795 68.905 100.555 ;
        RECT 67.315 99.625 67.725 99.725 ;
        RECT 66.815 99.365 67.145 99.535 ;
        RECT 67.315 99.415 68.925 99.625 ;
        RECT 64.965 98.995 65.300 99.245 ;
        RECT 65.470 98.805 65.640 99.365 ;
        RECT 66.965 99.245 67.145 99.365 ;
        RECT 65.810 98.975 66.145 99.245 ;
        RECT 66.325 98.995 66.790 99.195 ;
        RECT 66.965 98.995 67.295 99.245 ;
        RECT 67.465 99.195 67.930 99.245 ;
        RECT 67.465 99.025 67.935 99.195 ;
        RECT 67.465 98.995 67.930 99.025 ;
        RECT 68.125 98.995 68.480 99.245 ;
        RECT 68.650 98.815 68.925 99.415 ;
        RECT 60.345 98.005 63.855 98.775 ;
        RECT 64.945 98.175 65.640 98.805 ;
        RECT 65.845 98.005 66.155 98.805 ;
        RECT 66.325 98.615 67.505 98.785 ;
        RECT 66.325 98.200 66.665 98.615 ;
        RECT 66.835 98.005 67.005 98.445 ;
        RECT 67.175 98.395 67.505 98.615 ;
        RECT 67.675 98.635 68.925 98.815 ;
        RECT 67.675 98.565 68.040 98.635 ;
        RECT 67.175 98.215 68.425 98.395 ;
        RECT 68.695 98.005 68.865 98.465 ;
        RECT 69.095 98.285 69.375 100.385 ;
        RECT 70.005 99.390 70.295 100.555 ;
        RECT 70.465 99.465 72.135 100.555 ;
        RECT 72.855 99.885 73.025 100.385 ;
        RECT 73.195 100.055 73.525 100.555 ;
        RECT 72.855 99.715 73.520 99.885 ;
        RECT 70.465 98.775 71.215 99.295 ;
        RECT 71.385 98.945 72.135 99.465 ;
        RECT 72.770 98.895 73.120 99.545 ;
        RECT 70.005 98.005 70.295 98.730 ;
        RECT 70.465 98.005 72.135 98.775 ;
        RECT 73.290 98.725 73.520 99.715 ;
        RECT 72.855 98.555 73.520 98.725 ;
        RECT 72.855 98.265 73.025 98.555 ;
        RECT 73.195 98.005 73.525 98.385 ;
        RECT 73.695 98.265 73.880 100.385 ;
        RECT 74.120 100.095 74.385 100.555 ;
        RECT 74.555 99.960 74.805 100.385 ;
        RECT 75.015 100.110 76.120 100.280 ;
        RECT 74.500 99.830 74.805 99.960 ;
        RECT 74.050 98.635 74.330 99.585 ;
        RECT 74.500 98.725 74.670 99.830 ;
        RECT 74.840 99.045 75.080 99.640 ;
        RECT 75.250 99.575 75.780 99.940 ;
        RECT 75.250 98.875 75.420 99.575 ;
        RECT 75.950 99.495 76.120 100.110 ;
        RECT 76.290 99.755 76.460 100.555 ;
        RECT 76.630 100.055 76.880 100.385 ;
        RECT 77.105 100.085 77.990 100.255 ;
        RECT 75.950 99.405 76.460 99.495 ;
        RECT 74.500 98.595 74.725 98.725 ;
        RECT 74.895 98.655 75.420 98.875 ;
        RECT 75.590 99.235 76.460 99.405 ;
        RECT 74.135 98.005 74.385 98.465 ;
        RECT 74.555 98.455 74.725 98.595 ;
        RECT 75.590 98.455 75.760 99.235 ;
        RECT 76.290 99.165 76.460 99.235 ;
        RECT 75.970 98.985 76.170 99.015 ;
        RECT 76.630 98.985 76.800 100.055 ;
        RECT 76.970 99.165 77.160 99.885 ;
        RECT 75.970 98.685 76.800 98.985 ;
        RECT 77.330 98.955 77.650 99.915 ;
        RECT 74.555 98.285 74.890 98.455 ;
        RECT 75.085 98.285 75.760 98.455 ;
        RECT 76.080 98.005 76.450 98.505 ;
        RECT 76.630 98.455 76.800 98.685 ;
        RECT 77.185 98.625 77.650 98.955 ;
        RECT 77.820 99.245 77.990 100.085 ;
        RECT 78.170 100.055 78.485 100.555 ;
        RECT 78.715 99.825 79.055 100.385 ;
        RECT 78.160 99.450 79.055 99.825 ;
        RECT 79.225 99.545 79.395 100.555 ;
        RECT 78.865 99.245 79.055 99.450 ;
        RECT 79.565 99.495 79.895 100.340 ;
        RECT 79.565 99.415 79.955 99.495 ;
        RECT 80.125 99.465 82.715 100.555 ;
        RECT 79.740 99.365 79.955 99.415 ;
        RECT 77.820 98.915 78.695 99.245 ;
        RECT 78.865 98.915 79.615 99.245 ;
        RECT 77.820 98.455 77.990 98.915 ;
        RECT 78.865 98.745 79.065 98.915 ;
        RECT 79.785 98.785 79.955 99.365 ;
        RECT 79.730 98.745 79.955 98.785 ;
        RECT 76.630 98.285 77.035 98.455 ;
        RECT 77.205 98.285 77.990 98.455 ;
        RECT 78.265 98.005 78.475 98.535 ;
        RECT 78.735 98.220 79.065 98.745 ;
        RECT 79.575 98.660 79.955 98.745 ;
        RECT 80.125 98.775 81.335 99.295 ;
        RECT 81.505 98.945 82.715 99.465 ;
        RECT 82.885 99.465 84.095 100.555 ;
        RECT 82.885 98.925 83.405 99.465 ;
        RECT 79.235 98.005 79.405 98.615 ;
        RECT 79.575 98.225 79.905 98.660 ;
        RECT 80.125 98.005 82.715 98.775 ;
        RECT 83.575 98.755 84.095 99.295 ;
        RECT 82.885 98.005 84.095 98.755 ;
        RECT 5.520 97.835 84.180 98.005 ;
        RECT 5.605 97.085 6.815 97.835 ;
        RECT 7.075 97.285 7.245 97.575 ;
        RECT 7.415 97.455 7.745 97.835 ;
        RECT 7.075 97.115 7.740 97.285 ;
        RECT 5.605 96.545 6.125 97.085 ;
        RECT 6.295 96.375 6.815 96.915 ;
        RECT 5.605 95.285 6.815 96.375 ;
        RECT 6.990 96.295 7.340 96.945 ;
        RECT 7.510 96.125 7.740 97.115 ;
        RECT 7.075 95.955 7.740 96.125 ;
        RECT 7.075 95.455 7.245 95.955 ;
        RECT 7.415 95.285 7.745 95.785 ;
        RECT 7.915 95.455 8.100 97.575 ;
        RECT 8.355 97.375 8.605 97.835 ;
        RECT 8.775 97.385 9.110 97.555 ;
        RECT 9.305 97.385 9.980 97.555 ;
        RECT 8.775 97.245 8.945 97.385 ;
        RECT 8.270 96.255 8.550 97.205 ;
        RECT 8.720 97.115 8.945 97.245 ;
        RECT 8.720 96.010 8.890 97.115 ;
        RECT 9.115 96.965 9.640 97.185 ;
        RECT 9.060 96.200 9.300 96.795 ;
        RECT 9.470 96.265 9.640 96.965 ;
        RECT 9.810 96.605 9.980 97.385 ;
        RECT 10.300 97.335 10.670 97.835 ;
        RECT 10.850 97.385 11.255 97.555 ;
        RECT 11.425 97.385 12.210 97.555 ;
        RECT 10.850 97.155 11.020 97.385 ;
        RECT 10.190 96.855 11.020 97.155 ;
        RECT 11.405 96.885 11.870 97.215 ;
        RECT 10.190 96.825 10.390 96.855 ;
        RECT 10.510 96.605 10.680 96.675 ;
        RECT 9.810 96.435 10.680 96.605 ;
        RECT 10.170 96.345 10.680 96.435 ;
        RECT 8.720 95.880 9.025 96.010 ;
        RECT 9.470 95.900 10.000 96.265 ;
        RECT 8.340 95.285 8.605 95.745 ;
        RECT 8.775 95.455 9.025 95.880 ;
        RECT 10.170 95.730 10.340 96.345 ;
        RECT 9.235 95.560 10.340 95.730 ;
        RECT 10.510 95.285 10.680 96.085 ;
        RECT 10.850 95.785 11.020 96.855 ;
        RECT 11.190 95.955 11.380 96.675 ;
        RECT 11.550 95.925 11.870 96.885 ;
        RECT 12.040 96.925 12.210 97.385 ;
        RECT 12.485 97.305 12.695 97.835 ;
        RECT 12.955 97.095 13.285 97.620 ;
        RECT 13.455 97.225 13.625 97.835 ;
        RECT 13.795 97.180 14.125 97.615 ;
        RECT 14.350 97.580 14.685 97.625 ;
        RECT 13.795 97.095 14.175 97.180 ;
        RECT 13.085 96.925 13.285 97.095 ;
        RECT 13.950 97.055 14.175 97.095 ;
        RECT 12.040 96.595 12.915 96.925 ;
        RECT 13.085 96.595 13.835 96.925 ;
        RECT 10.850 95.455 11.100 95.785 ;
        RECT 12.040 95.755 12.210 96.595 ;
        RECT 13.085 96.390 13.275 96.595 ;
        RECT 14.005 96.475 14.175 97.055 ;
        RECT 13.960 96.425 14.175 96.475 ;
        RECT 12.380 96.015 13.275 96.390 ;
        RECT 13.785 96.345 14.175 96.425 ;
        RECT 14.345 97.115 14.685 97.580 ;
        RECT 14.855 97.455 15.185 97.835 ;
        RECT 15.645 97.495 15.915 97.500 ;
        RECT 15.645 97.325 15.955 97.495 ;
        RECT 14.345 96.425 14.515 97.115 ;
        RECT 14.685 96.595 14.945 96.925 ;
        RECT 11.325 95.585 12.210 95.755 ;
        RECT 12.390 95.285 12.705 95.785 ;
        RECT 12.935 95.455 13.275 96.015 ;
        RECT 13.445 95.285 13.615 96.295 ;
        RECT 13.785 95.500 14.115 96.345 ;
        RECT 14.345 95.455 14.605 96.425 ;
        RECT 14.775 96.045 14.945 96.595 ;
        RECT 15.115 96.225 15.455 97.255 ;
        RECT 15.645 96.225 15.915 97.325 ;
        RECT 16.140 96.225 16.420 97.500 ;
        RECT 16.620 97.335 16.850 97.665 ;
        RECT 17.095 97.455 17.425 97.835 ;
        RECT 16.620 96.045 16.790 97.335 ;
        RECT 17.595 97.265 17.770 97.665 ;
        RECT 17.140 97.095 17.770 97.265 ;
        RECT 17.140 96.925 17.310 97.095 ;
        RECT 18.025 97.035 18.335 97.835 ;
        RECT 18.540 97.035 19.235 97.665 ;
        RECT 19.405 97.290 24.750 97.835 ;
        RECT 24.925 97.290 30.270 97.835 ;
        RECT 18.540 96.985 18.715 97.035 ;
        RECT 16.960 96.595 17.310 96.925 ;
        RECT 14.775 95.875 16.790 96.045 ;
        RECT 17.140 96.075 17.310 96.595 ;
        RECT 17.490 96.245 17.855 96.925 ;
        RECT 18.035 96.595 18.370 96.865 ;
        RECT 18.540 96.435 18.710 96.985 ;
        RECT 18.880 96.595 19.215 96.845 ;
        RECT 20.990 96.460 21.330 97.290 ;
        RECT 17.140 95.905 17.770 96.075 ;
        RECT 14.800 95.285 15.130 95.695 ;
        RECT 15.330 95.455 15.500 95.875 ;
        RECT 15.715 95.285 16.385 95.695 ;
        RECT 16.620 95.455 16.790 95.875 ;
        RECT 17.095 95.285 17.425 95.725 ;
        RECT 17.595 95.455 17.770 95.905 ;
        RECT 18.025 95.285 18.305 96.425 ;
        RECT 18.475 95.455 18.805 96.435 ;
        RECT 18.975 95.285 19.235 96.425 ;
        RECT 22.810 95.720 23.160 96.970 ;
        RECT 26.510 96.460 26.850 97.290 ;
        RECT 31.365 97.110 31.655 97.835 ;
        RECT 31.825 97.065 34.415 97.835 ;
        RECT 35.050 97.095 35.305 97.665 ;
        RECT 35.475 97.435 35.805 97.835 ;
        RECT 36.230 97.300 36.760 97.665 ;
        RECT 36.950 97.495 37.225 97.665 ;
        RECT 36.945 97.325 37.225 97.495 ;
        RECT 36.230 97.265 36.405 97.300 ;
        RECT 35.475 97.095 36.405 97.265 ;
        RECT 28.330 95.720 28.680 96.970 ;
        RECT 31.825 96.545 33.035 97.065 ;
        RECT 19.405 95.285 24.750 95.720 ;
        RECT 24.925 95.285 30.270 95.720 ;
        RECT 31.365 95.285 31.655 96.450 ;
        RECT 33.205 96.375 34.415 96.895 ;
        RECT 31.825 95.285 34.415 96.375 ;
        RECT 35.050 96.425 35.220 97.095 ;
        RECT 35.475 96.925 35.645 97.095 ;
        RECT 35.390 96.595 35.645 96.925 ;
        RECT 35.870 96.595 36.065 96.925 ;
        RECT 35.050 95.455 35.385 96.425 ;
        RECT 35.555 95.285 35.725 96.425 ;
        RECT 35.895 95.625 36.065 96.595 ;
        RECT 36.235 95.965 36.405 97.095 ;
        RECT 36.575 96.305 36.745 97.105 ;
        RECT 36.950 96.505 37.225 97.325 ;
        RECT 37.395 96.305 37.585 97.665 ;
        RECT 37.765 97.300 38.275 97.835 ;
        RECT 38.495 97.025 38.740 97.630 ;
        RECT 39.275 97.285 39.445 97.575 ;
        RECT 39.615 97.455 39.945 97.835 ;
        RECT 39.275 97.115 39.940 97.285 ;
        RECT 37.785 96.855 39.015 97.025 ;
        RECT 36.575 96.135 37.585 96.305 ;
        RECT 37.755 96.290 38.505 96.480 ;
        RECT 36.235 95.795 37.360 95.965 ;
        RECT 37.755 95.625 37.925 96.290 ;
        RECT 38.675 96.045 39.015 96.855 ;
        RECT 39.190 96.295 39.540 96.945 ;
        RECT 39.710 96.125 39.940 97.115 ;
        RECT 35.895 95.455 37.925 95.625 ;
        RECT 38.095 95.285 38.265 96.045 ;
        RECT 38.500 95.635 39.015 96.045 ;
        RECT 39.275 95.955 39.940 96.125 ;
        RECT 39.275 95.455 39.445 95.955 ;
        RECT 39.615 95.285 39.945 95.785 ;
        RECT 40.115 95.455 40.300 97.575 ;
        RECT 40.555 97.375 40.805 97.835 ;
        RECT 40.975 97.385 41.310 97.555 ;
        RECT 41.505 97.385 42.180 97.555 ;
        RECT 40.975 97.245 41.145 97.385 ;
        RECT 40.470 96.255 40.750 97.205 ;
        RECT 40.920 97.115 41.145 97.245 ;
        RECT 40.920 96.010 41.090 97.115 ;
        RECT 41.315 96.965 41.840 97.185 ;
        RECT 41.260 96.200 41.500 96.795 ;
        RECT 41.670 96.265 41.840 96.965 ;
        RECT 42.010 96.605 42.180 97.385 ;
        RECT 42.500 97.335 42.870 97.835 ;
        RECT 43.050 97.385 43.455 97.555 ;
        RECT 43.625 97.385 44.410 97.555 ;
        RECT 43.050 97.155 43.220 97.385 ;
        RECT 42.390 96.855 43.220 97.155 ;
        RECT 43.605 96.885 44.070 97.215 ;
        RECT 42.390 96.825 42.590 96.855 ;
        RECT 42.710 96.605 42.880 96.675 ;
        RECT 42.010 96.435 42.880 96.605 ;
        RECT 42.370 96.345 42.880 96.435 ;
        RECT 40.920 95.880 41.225 96.010 ;
        RECT 41.670 95.900 42.200 96.265 ;
        RECT 40.540 95.285 40.805 95.745 ;
        RECT 40.975 95.455 41.225 95.880 ;
        RECT 42.370 95.730 42.540 96.345 ;
        RECT 41.435 95.560 42.540 95.730 ;
        RECT 42.710 95.285 42.880 96.085 ;
        RECT 43.050 95.785 43.220 96.855 ;
        RECT 43.390 95.955 43.580 96.675 ;
        RECT 43.750 95.925 44.070 96.885 ;
        RECT 44.240 96.925 44.410 97.385 ;
        RECT 44.685 97.305 44.895 97.835 ;
        RECT 45.155 97.095 45.485 97.620 ;
        RECT 45.655 97.225 45.825 97.835 ;
        RECT 45.995 97.180 46.325 97.615 ;
        RECT 46.730 97.355 46.900 97.835 ;
        RECT 47.070 97.185 47.400 97.655 ;
        RECT 47.570 97.355 47.740 97.835 ;
        RECT 47.910 97.185 48.240 97.655 ;
        RECT 45.995 97.095 46.375 97.180 ;
        RECT 45.285 96.925 45.485 97.095 ;
        RECT 46.150 97.055 46.375 97.095 ;
        RECT 44.240 96.595 45.115 96.925 ;
        RECT 45.285 96.595 46.035 96.925 ;
        RECT 43.050 95.455 43.300 95.785 ;
        RECT 44.240 95.755 44.410 96.595 ;
        RECT 45.285 96.390 45.475 96.595 ;
        RECT 46.205 96.475 46.375 97.055 ;
        RECT 46.160 96.425 46.375 96.475 ;
        RECT 44.580 96.015 45.475 96.390 ;
        RECT 45.985 96.345 46.375 96.425 ;
        RECT 46.545 97.015 48.240 97.185 ;
        RECT 48.450 97.095 48.620 97.835 ;
        RECT 48.835 97.095 49.165 97.630 ;
        RECT 49.335 97.325 49.575 97.835 ;
        RECT 49.855 97.285 50.025 97.575 ;
        RECT 50.195 97.455 50.525 97.835 ;
        RECT 46.545 96.425 46.890 97.015 ;
        RECT 47.060 96.675 48.270 96.845 ;
        RECT 48.065 96.425 48.270 96.675 ;
        RECT 48.440 96.595 48.815 96.925 ;
        RECT 48.985 96.425 49.165 97.095 ;
        RECT 49.335 96.595 49.590 97.155 ;
        RECT 49.855 97.115 50.520 97.285 ;
        RECT 43.525 95.585 44.410 95.755 ;
        RECT 44.590 95.285 44.905 95.785 ;
        RECT 45.135 95.455 45.475 96.015 ;
        RECT 45.645 95.285 45.815 96.295 ;
        RECT 45.985 95.500 46.315 96.345 ;
        RECT 46.545 96.255 47.400 96.425 ;
        RECT 48.065 96.255 49.525 96.425 ;
        RECT 49.770 96.295 50.120 96.945 ;
        RECT 47.070 96.085 47.400 96.255 ;
        RECT 46.730 95.285 46.900 96.085 ;
        RECT 47.070 95.915 48.240 96.085 ;
        RECT 47.070 95.455 47.400 95.915 ;
        RECT 47.570 95.285 47.740 95.745 ;
        RECT 47.910 95.455 48.240 95.915 ;
        RECT 48.450 95.285 48.620 96.085 ;
        RECT 49.165 95.455 49.525 96.255 ;
        RECT 50.290 96.125 50.520 97.115 ;
        RECT 49.855 95.955 50.520 96.125 ;
        RECT 49.855 95.455 50.025 95.955 ;
        RECT 50.195 95.285 50.525 95.785 ;
        RECT 50.695 95.455 50.880 97.575 ;
        RECT 51.135 97.375 51.385 97.835 ;
        RECT 51.555 97.385 51.890 97.555 ;
        RECT 52.085 97.385 52.760 97.555 ;
        RECT 51.555 97.245 51.725 97.385 ;
        RECT 51.050 96.255 51.330 97.205 ;
        RECT 51.500 97.115 51.725 97.245 ;
        RECT 51.500 96.010 51.670 97.115 ;
        RECT 51.895 96.965 52.420 97.185 ;
        RECT 51.840 96.200 52.080 96.795 ;
        RECT 52.250 96.265 52.420 96.965 ;
        RECT 52.590 96.605 52.760 97.385 ;
        RECT 53.080 97.335 53.450 97.835 ;
        RECT 53.630 97.385 54.035 97.555 ;
        RECT 54.205 97.385 54.990 97.555 ;
        RECT 53.630 97.155 53.800 97.385 ;
        RECT 52.970 96.855 53.800 97.155 ;
        RECT 54.185 96.885 54.650 97.215 ;
        RECT 52.970 96.825 53.170 96.855 ;
        RECT 53.290 96.605 53.460 96.675 ;
        RECT 52.590 96.435 53.460 96.605 ;
        RECT 52.950 96.345 53.460 96.435 ;
        RECT 51.500 95.880 51.805 96.010 ;
        RECT 52.250 95.900 52.780 96.265 ;
        RECT 51.120 95.285 51.385 95.745 ;
        RECT 51.555 95.455 51.805 95.880 ;
        RECT 52.950 95.730 53.120 96.345 ;
        RECT 52.015 95.560 53.120 95.730 ;
        RECT 53.290 95.285 53.460 96.085 ;
        RECT 53.630 95.785 53.800 96.855 ;
        RECT 53.970 95.955 54.160 96.675 ;
        RECT 54.330 95.925 54.650 96.885 ;
        RECT 54.820 96.925 54.990 97.385 ;
        RECT 55.265 97.305 55.475 97.835 ;
        RECT 55.735 97.095 56.065 97.620 ;
        RECT 56.235 97.225 56.405 97.835 ;
        RECT 56.575 97.180 56.905 97.615 ;
        RECT 56.575 97.095 56.955 97.180 ;
        RECT 57.125 97.110 57.415 97.835 ;
        RECT 55.865 96.925 56.065 97.095 ;
        RECT 56.730 97.055 56.955 97.095 ;
        RECT 54.820 96.595 55.695 96.925 ;
        RECT 55.865 96.595 56.615 96.925 ;
        RECT 53.630 95.455 53.880 95.785 ;
        RECT 54.820 95.755 54.990 96.595 ;
        RECT 55.865 96.390 56.055 96.595 ;
        RECT 56.785 96.475 56.955 97.055 ;
        RECT 56.740 96.425 56.955 96.475 ;
        RECT 57.590 97.095 57.845 97.665 ;
        RECT 58.015 97.435 58.345 97.835 ;
        RECT 58.770 97.300 59.300 97.665 ;
        RECT 58.770 97.265 58.945 97.300 ;
        RECT 58.015 97.095 58.945 97.265 ;
        RECT 55.160 96.015 56.055 96.390 ;
        RECT 56.565 96.345 56.955 96.425 ;
        RECT 54.105 95.585 54.990 95.755 ;
        RECT 55.170 95.285 55.485 95.785 ;
        RECT 55.715 95.455 56.055 96.015 ;
        RECT 56.225 95.285 56.395 96.295 ;
        RECT 56.565 95.500 56.895 96.345 ;
        RECT 57.125 95.285 57.415 96.450 ;
        RECT 57.590 96.425 57.760 97.095 ;
        RECT 58.015 96.925 58.185 97.095 ;
        RECT 57.930 96.595 58.185 96.925 ;
        RECT 58.410 96.595 58.605 96.925 ;
        RECT 57.590 95.455 57.925 96.425 ;
        RECT 58.095 95.285 58.265 96.425 ;
        RECT 58.435 95.625 58.605 96.595 ;
        RECT 58.775 95.965 58.945 97.095 ;
        RECT 59.115 96.305 59.285 97.105 ;
        RECT 59.490 96.815 59.765 97.665 ;
        RECT 59.485 96.645 59.765 96.815 ;
        RECT 59.490 96.505 59.765 96.645 ;
        RECT 59.935 96.305 60.125 97.665 ;
        RECT 60.305 97.300 60.815 97.835 ;
        RECT 61.035 97.025 61.280 97.630 ;
        RECT 61.725 97.065 63.395 97.835 ;
        RECT 64.025 97.095 64.515 97.665 ;
        RECT 64.685 97.265 64.915 97.665 ;
        RECT 65.085 97.435 65.505 97.835 ;
        RECT 65.675 97.265 65.845 97.665 ;
        RECT 64.685 97.095 65.845 97.265 ;
        RECT 66.015 97.095 66.465 97.835 ;
        RECT 66.635 97.095 67.075 97.655 ;
        RECT 67.295 97.365 67.585 97.835 ;
        RECT 67.755 97.195 68.085 97.665 ;
        RECT 68.255 97.365 68.425 97.835 ;
        RECT 68.595 97.195 68.925 97.665 ;
        RECT 67.755 97.185 68.925 97.195 ;
        RECT 60.325 96.855 61.555 97.025 ;
        RECT 59.115 96.135 60.125 96.305 ;
        RECT 60.295 96.290 61.045 96.480 ;
        RECT 58.775 95.795 59.900 95.965 ;
        RECT 60.295 95.625 60.465 96.290 ;
        RECT 61.215 96.045 61.555 96.855 ;
        RECT 61.725 96.545 62.475 97.065 ;
        RECT 62.645 96.375 63.395 96.895 ;
        RECT 58.435 95.455 60.465 95.625 ;
        RECT 60.635 95.285 60.805 96.045 ;
        RECT 61.040 95.635 61.555 96.045 ;
        RECT 61.725 95.285 63.395 96.375 ;
        RECT 64.025 96.425 64.195 97.095 ;
        RECT 64.365 96.595 64.770 96.925 ;
        RECT 64.025 96.255 64.795 96.425 ;
        RECT 64.035 95.285 64.365 96.085 ;
        RECT 64.545 95.625 64.795 96.255 ;
        RECT 64.985 95.795 65.235 96.925 ;
        RECT 65.435 96.595 65.680 96.925 ;
        RECT 65.865 96.645 66.255 96.925 ;
        RECT 65.435 95.795 65.635 96.595 ;
        RECT 66.425 96.475 66.595 96.925 ;
        RECT 65.805 96.305 66.595 96.475 ;
        RECT 65.805 95.625 65.975 96.305 ;
        RECT 64.545 95.455 65.975 95.625 ;
        RECT 66.145 95.285 66.460 96.135 ;
        RECT 66.765 96.085 67.075 97.095 ;
        RECT 67.325 97.015 68.925 97.185 ;
        RECT 69.095 97.015 69.370 97.835 ;
        RECT 69.550 97.160 69.825 97.505 ;
        RECT 70.015 97.435 70.395 97.835 ;
        RECT 70.565 97.265 70.735 97.615 ;
        RECT 70.905 97.435 71.235 97.835 ;
        RECT 71.405 97.265 71.660 97.615 ;
        RECT 71.865 97.325 72.105 97.835 ;
        RECT 72.275 97.325 72.565 97.665 ;
        RECT 72.795 97.325 73.110 97.835 ;
        RECT 67.325 96.475 67.540 97.015 ;
        RECT 67.710 96.645 68.480 96.845 ;
        RECT 68.650 96.645 69.370 96.845 ;
        RECT 67.325 96.255 68.085 96.475 ;
        RECT 66.635 95.455 67.075 96.085 ;
        RECT 67.285 95.625 67.585 96.085 ;
        RECT 67.755 95.795 68.085 96.255 ;
        RECT 68.255 96.255 69.370 96.465 ;
        RECT 68.255 95.625 68.425 96.255 ;
        RECT 67.285 95.455 68.425 95.625 ;
        RECT 68.595 95.285 68.925 96.085 ;
        RECT 69.095 95.455 69.370 96.255 ;
        RECT 69.550 96.425 69.720 97.160 ;
        RECT 69.995 97.095 71.660 97.265 ;
        RECT 69.995 96.925 70.165 97.095 ;
        RECT 69.890 96.595 70.165 96.925 ;
        RECT 70.335 96.595 71.160 96.925 ;
        RECT 71.330 96.595 71.675 96.925 ;
        RECT 71.910 96.815 72.105 97.155 ;
        RECT 71.905 96.645 72.105 96.815 ;
        RECT 71.910 96.595 72.105 96.645 ;
        RECT 69.995 96.425 70.165 96.595 ;
        RECT 69.550 95.455 69.825 96.425 ;
        RECT 69.995 96.255 70.655 96.425 ;
        RECT 70.965 96.305 71.160 96.595 ;
        RECT 72.275 96.425 72.455 97.325 ;
        RECT 73.280 97.265 73.450 97.535 ;
        RECT 73.620 97.435 73.950 97.835 ;
        RECT 72.625 96.595 73.035 97.155 ;
        RECT 73.280 97.095 73.975 97.265 ;
        RECT 73.205 96.425 73.375 96.925 ;
        RECT 70.485 96.135 70.655 96.255 ;
        RECT 71.330 96.135 71.655 96.425 ;
        RECT 70.035 95.285 70.315 96.085 ;
        RECT 70.485 95.965 71.655 96.135 ;
        RECT 71.915 96.255 73.375 96.425 ;
        RECT 71.915 96.080 72.275 96.255 ;
        RECT 73.545 96.085 73.975 97.095 ;
        RECT 70.485 95.505 71.675 95.795 ;
        RECT 72.860 95.285 73.030 96.085 ;
        RECT 73.200 95.915 73.975 96.085 ;
        RECT 74.610 97.095 74.865 97.665 ;
        RECT 75.035 97.435 75.365 97.835 ;
        RECT 75.790 97.300 76.320 97.665 ;
        RECT 76.510 97.495 76.785 97.665 ;
        RECT 76.505 97.325 76.785 97.495 ;
        RECT 75.790 97.265 75.965 97.300 ;
        RECT 75.035 97.095 75.965 97.265 ;
        RECT 74.610 96.425 74.780 97.095 ;
        RECT 75.035 96.925 75.205 97.095 ;
        RECT 74.950 96.595 75.205 96.925 ;
        RECT 75.430 96.595 75.625 96.925 ;
        RECT 73.200 95.455 73.530 95.915 ;
        RECT 73.700 95.285 73.870 95.745 ;
        RECT 74.610 95.455 74.945 96.425 ;
        RECT 75.115 95.285 75.285 96.425 ;
        RECT 75.455 95.625 75.625 96.595 ;
        RECT 75.795 95.965 75.965 97.095 ;
        RECT 76.135 96.305 76.305 97.105 ;
        RECT 76.510 96.505 76.785 97.325 ;
        RECT 76.955 96.305 77.145 97.665 ;
        RECT 77.325 97.300 77.835 97.835 ;
        RECT 78.055 97.025 78.300 97.630 ;
        RECT 78.745 97.065 82.255 97.835 ;
        RECT 82.885 97.085 84.095 97.835 ;
        RECT 77.345 96.855 78.575 97.025 ;
        RECT 76.135 96.135 77.145 96.305 ;
        RECT 77.315 96.290 78.065 96.480 ;
        RECT 75.795 95.795 76.920 95.965 ;
        RECT 77.315 95.625 77.485 96.290 ;
        RECT 78.235 96.045 78.575 96.855 ;
        RECT 78.745 96.545 80.395 97.065 ;
        RECT 80.565 96.375 82.255 96.895 ;
        RECT 75.455 95.455 77.485 95.625 ;
        RECT 77.655 95.285 77.825 96.045 ;
        RECT 78.060 95.635 78.575 96.045 ;
        RECT 78.745 95.285 82.255 96.375 ;
        RECT 82.885 96.375 83.405 96.915 ;
        RECT 83.575 96.545 84.095 97.085 ;
        RECT 82.885 95.285 84.095 96.375 ;
        RECT 5.520 95.115 84.180 95.285 ;
        RECT 5.605 94.025 6.815 95.115 ;
        RECT 6.985 94.025 10.495 95.115 ;
        RECT 5.605 93.315 6.125 93.855 ;
        RECT 6.295 93.485 6.815 94.025 ;
        RECT 6.985 93.335 8.635 93.855 ;
        RECT 8.805 93.505 10.495 94.025 ;
        RECT 10.670 93.975 10.990 95.115 ;
        RECT 11.170 93.805 11.365 94.855 ;
        RECT 11.545 94.265 11.875 94.945 ;
        RECT 12.075 94.315 12.330 95.115 ;
        RECT 11.545 93.985 11.895 94.265 ;
        RECT 10.730 93.755 10.990 93.805 ;
        RECT 10.725 93.585 10.990 93.755 ;
        RECT 10.730 93.475 10.990 93.585 ;
        RECT 11.170 93.475 11.555 93.805 ;
        RECT 11.725 93.605 11.895 93.985 ;
        RECT 12.085 93.775 12.330 94.135 ;
        RECT 12.505 93.975 12.890 94.945 ;
        RECT 13.060 94.655 13.385 95.115 ;
        RECT 13.905 94.485 14.185 94.945 ;
        RECT 13.060 94.265 14.185 94.485 ;
        RECT 11.725 93.435 12.245 93.605 ;
        RECT 5.605 92.565 6.815 93.315 ;
        RECT 6.985 92.565 10.495 93.335 ;
        RECT 10.670 93.095 11.885 93.265 ;
        RECT 10.670 92.745 10.960 93.095 ;
        RECT 11.155 92.565 11.485 92.925 ;
        RECT 11.655 92.790 11.885 93.095 ;
        RECT 12.075 92.870 12.245 93.435 ;
        RECT 12.505 93.305 12.785 93.975 ;
        RECT 13.060 93.805 13.510 94.265 ;
        RECT 14.375 94.095 14.775 94.945 ;
        RECT 15.175 94.655 15.445 95.115 ;
        RECT 15.615 94.485 15.900 94.945 ;
        RECT 12.955 93.475 13.510 93.805 ;
        RECT 13.680 93.535 14.775 94.095 ;
        RECT 13.060 93.365 13.510 93.475 ;
        RECT 12.505 92.735 12.890 93.305 ;
        RECT 13.060 93.195 14.185 93.365 ;
        RECT 13.060 92.565 13.385 93.025 ;
        RECT 13.905 92.735 14.185 93.195 ;
        RECT 14.375 92.735 14.775 93.535 ;
        RECT 14.945 94.265 15.900 94.485 ;
        RECT 14.945 93.365 15.155 94.265 ;
        RECT 15.325 93.535 16.015 94.095 ;
        RECT 16.185 94.025 17.855 95.115 ;
        RECT 14.945 93.195 15.900 93.365 ;
        RECT 15.175 92.565 15.445 93.025 ;
        RECT 15.615 92.735 15.900 93.195 ;
        RECT 16.185 93.335 16.935 93.855 ;
        RECT 17.105 93.505 17.855 94.025 ;
        RECT 18.485 93.950 18.775 95.115 ;
        RECT 18.945 94.680 24.290 95.115 ;
        RECT 16.185 92.565 17.855 93.335 ;
        RECT 18.485 92.565 18.775 93.290 ;
        RECT 20.530 93.110 20.870 93.940 ;
        RECT 22.350 93.430 22.700 94.680 ;
        RECT 24.465 94.025 26.135 95.115 ;
        RECT 26.395 94.445 26.565 94.945 ;
        RECT 26.735 94.615 27.065 95.115 ;
        RECT 26.395 94.275 27.060 94.445 ;
        RECT 24.465 93.335 25.215 93.855 ;
        RECT 25.385 93.505 26.135 94.025 ;
        RECT 26.310 93.455 26.660 94.105 ;
        RECT 18.945 92.565 24.290 93.110 ;
        RECT 24.465 92.565 26.135 93.335 ;
        RECT 26.830 93.285 27.060 94.275 ;
        RECT 26.395 93.115 27.060 93.285 ;
        RECT 26.395 92.825 26.565 93.115 ;
        RECT 26.735 92.565 27.065 92.945 ;
        RECT 27.235 92.825 27.420 94.945 ;
        RECT 27.660 94.655 27.925 95.115 ;
        RECT 28.095 94.520 28.345 94.945 ;
        RECT 28.555 94.670 29.660 94.840 ;
        RECT 28.040 94.390 28.345 94.520 ;
        RECT 27.590 93.195 27.870 94.145 ;
        RECT 28.040 93.285 28.210 94.390 ;
        RECT 28.380 93.605 28.620 94.200 ;
        RECT 28.790 94.135 29.320 94.500 ;
        RECT 28.790 93.435 28.960 94.135 ;
        RECT 29.490 94.055 29.660 94.670 ;
        RECT 29.830 94.315 30.000 95.115 ;
        RECT 30.170 94.615 30.420 94.945 ;
        RECT 30.645 94.645 31.530 94.815 ;
        RECT 29.490 93.965 30.000 94.055 ;
        RECT 28.040 93.155 28.265 93.285 ;
        RECT 28.435 93.215 28.960 93.435 ;
        RECT 29.130 93.795 30.000 93.965 ;
        RECT 27.675 92.565 27.925 93.025 ;
        RECT 28.095 93.015 28.265 93.155 ;
        RECT 29.130 93.015 29.300 93.795 ;
        RECT 29.830 93.725 30.000 93.795 ;
        RECT 29.510 93.545 29.710 93.575 ;
        RECT 30.170 93.545 30.340 94.615 ;
        RECT 30.510 93.725 30.700 94.445 ;
        RECT 29.510 93.245 30.340 93.545 ;
        RECT 30.870 93.515 31.190 94.475 ;
        RECT 28.095 92.845 28.430 93.015 ;
        RECT 28.625 92.845 29.300 93.015 ;
        RECT 29.620 92.565 29.990 93.065 ;
        RECT 30.170 93.015 30.340 93.245 ;
        RECT 30.725 93.185 31.190 93.515 ;
        RECT 31.360 93.805 31.530 94.645 ;
        RECT 31.710 94.615 32.025 95.115 ;
        RECT 32.255 94.385 32.595 94.945 ;
        RECT 31.700 94.010 32.595 94.385 ;
        RECT 32.765 94.105 32.935 95.115 ;
        RECT 32.405 93.805 32.595 94.010 ;
        RECT 33.105 94.055 33.435 94.900 ;
        RECT 33.105 93.975 33.495 94.055 ;
        RECT 33.280 93.925 33.495 93.975 ;
        RECT 31.360 93.475 32.235 93.805 ;
        RECT 32.405 93.475 33.155 93.805 ;
        RECT 31.360 93.015 31.530 93.475 ;
        RECT 32.405 93.305 32.605 93.475 ;
        RECT 33.325 93.345 33.495 93.925 ;
        RECT 33.270 93.305 33.495 93.345 ;
        RECT 30.170 92.845 30.575 93.015 ;
        RECT 30.745 92.845 31.530 93.015 ;
        RECT 31.805 92.565 32.015 93.095 ;
        RECT 32.275 92.780 32.605 93.305 ;
        RECT 33.115 93.220 33.495 93.305 ;
        RECT 33.665 93.975 34.050 94.945 ;
        RECT 34.220 94.655 34.545 95.115 ;
        RECT 35.065 94.485 35.345 94.945 ;
        RECT 34.220 94.265 35.345 94.485 ;
        RECT 33.665 93.305 33.945 93.975 ;
        RECT 34.220 93.805 34.670 94.265 ;
        RECT 35.535 94.095 35.935 94.945 ;
        RECT 36.335 94.655 36.605 95.115 ;
        RECT 36.775 94.485 37.060 94.945 ;
        RECT 34.115 93.475 34.670 93.805 ;
        RECT 34.840 93.535 35.935 94.095 ;
        RECT 34.220 93.365 34.670 93.475 ;
        RECT 32.775 92.565 32.945 93.175 ;
        RECT 33.115 92.785 33.445 93.220 ;
        RECT 33.665 92.735 34.050 93.305 ;
        RECT 34.220 93.195 35.345 93.365 ;
        RECT 34.220 92.565 34.545 93.025 ;
        RECT 35.065 92.735 35.345 93.195 ;
        RECT 35.535 92.735 35.935 93.535 ;
        RECT 36.105 94.265 37.060 94.485 ;
        RECT 36.105 93.365 36.315 94.265 ;
        RECT 36.485 93.535 37.175 94.095 ;
        RECT 37.345 94.025 39.935 95.115 ;
        RECT 36.105 93.195 37.060 93.365 ;
        RECT 36.335 92.565 36.605 93.025 ;
        RECT 36.775 92.735 37.060 93.195 ;
        RECT 37.345 93.335 38.555 93.855 ;
        RECT 38.725 93.505 39.935 94.025 ;
        RECT 40.110 93.975 40.445 94.945 ;
        RECT 40.615 93.975 40.785 95.115 ;
        RECT 40.955 94.775 42.985 94.945 ;
        RECT 37.345 92.565 39.935 93.335 ;
        RECT 40.110 93.305 40.280 93.975 ;
        RECT 40.955 93.805 41.125 94.775 ;
        RECT 40.450 93.475 40.705 93.805 ;
        RECT 40.930 93.475 41.125 93.805 ;
        RECT 41.295 94.435 42.420 94.605 ;
        RECT 40.535 93.305 40.705 93.475 ;
        RECT 41.295 93.305 41.465 94.435 ;
        RECT 40.110 92.735 40.365 93.305 ;
        RECT 40.535 93.135 41.465 93.305 ;
        RECT 41.635 94.095 42.645 94.265 ;
        RECT 41.635 93.295 41.805 94.095 ;
        RECT 42.010 93.415 42.285 93.895 ;
        RECT 42.005 93.245 42.285 93.415 ;
        RECT 41.290 93.100 41.465 93.135 ;
        RECT 40.535 92.565 40.865 92.965 ;
        RECT 41.290 92.735 41.820 93.100 ;
        RECT 42.010 92.735 42.285 93.245 ;
        RECT 42.455 92.735 42.645 94.095 ;
        RECT 42.815 94.110 42.985 94.775 ;
        RECT 43.155 94.355 43.325 95.115 ;
        RECT 43.560 94.355 44.075 94.765 ;
        RECT 42.815 93.920 43.565 94.110 ;
        RECT 43.735 93.545 44.075 94.355 ;
        RECT 44.245 93.950 44.535 95.115 ;
        RECT 44.710 93.975 45.045 94.945 ;
        RECT 45.215 93.975 45.385 95.115 ;
        RECT 45.555 94.775 47.585 94.945 ;
        RECT 42.845 93.375 44.075 93.545 ;
        RECT 42.825 92.565 43.335 93.100 ;
        RECT 43.555 92.770 43.800 93.375 ;
        RECT 44.710 93.305 44.880 93.975 ;
        RECT 45.555 93.805 45.725 94.775 ;
        RECT 45.050 93.475 45.305 93.805 ;
        RECT 45.530 93.475 45.725 93.805 ;
        RECT 45.895 94.435 47.020 94.605 ;
        RECT 45.135 93.305 45.305 93.475 ;
        RECT 45.895 93.305 46.065 94.435 ;
        RECT 44.245 92.565 44.535 93.290 ;
        RECT 44.710 92.735 44.965 93.305 ;
        RECT 45.135 93.135 46.065 93.305 ;
        RECT 46.235 94.095 47.245 94.265 ;
        RECT 46.235 93.295 46.405 94.095 ;
        RECT 46.610 93.755 46.885 93.895 ;
        RECT 46.605 93.585 46.885 93.755 ;
        RECT 45.890 93.100 46.065 93.135 ;
        RECT 45.135 92.565 45.465 92.965 ;
        RECT 45.890 92.735 46.420 93.100 ;
        RECT 46.610 92.735 46.885 93.585 ;
        RECT 47.055 92.735 47.245 94.095 ;
        RECT 47.415 94.110 47.585 94.775 ;
        RECT 47.755 94.355 47.925 95.115 ;
        RECT 48.160 94.355 48.675 94.765 ;
        RECT 47.415 93.920 48.165 94.110 ;
        RECT 48.335 93.545 48.675 94.355 ;
        RECT 48.845 94.025 52.355 95.115 ;
        RECT 52.525 94.025 53.735 95.115 ;
        RECT 54.020 94.485 54.305 94.945 ;
        RECT 54.475 94.655 54.745 95.115 ;
        RECT 54.020 94.265 54.975 94.485 ;
        RECT 47.445 93.375 48.675 93.545 ;
        RECT 47.425 92.565 47.935 93.100 ;
        RECT 48.155 92.770 48.400 93.375 ;
        RECT 48.845 93.335 50.495 93.855 ;
        RECT 50.665 93.505 52.355 94.025 ;
        RECT 48.845 92.565 52.355 93.335 ;
        RECT 52.525 93.315 53.045 93.855 ;
        RECT 53.215 93.485 53.735 94.025 ;
        RECT 53.905 93.535 54.595 94.095 ;
        RECT 54.765 93.365 54.975 94.265 ;
        RECT 52.525 92.565 53.735 93.315 ;
        RECT 54.020 93.195 54.975 93.365 ;
        RECT 55.145 94.095 55.545 94.945 ;
        RECT 55.735 94.485 56.015 94.945 ;
        RECT 56.535 94.655 56.860 95.115 ;
        RECT 55.735 94.265 56.860 94.485 ;
        RECT 55.145 93.535 56.240 94.095 ;
        RECT 56.410 93.805 56.860 94.265 ;
        RECT 57.030 93.975 57.415 94.945 ;
        RECT 57.585 94.025 59.255 95.115 ;
        RECT 54.020 92.735 54.305 93.195 ;
        RECT 54.475 92.565 54.745 93.025 ;
        RECT 55.145 92.735 55.545 93.535 ;
        RECT 56.410 93.475 56.965 93.805 ;
        RECT 56.410 93.365 56.860 93.475 ;
        RECT 55.735 93.195 56.860 93.365 ;
        RECT 57.135 93.305 57.415 93.975 ;
        RECT 55.735 92.735 56.015 93.195 ;
        RECT 56.535 92.565 56.860 93.025 ;
        RECT 57.030 92.735 57.415 93.305 ;
        RECT 57.585 93.335 58.335 93.855 ;
        RECT 58.505 93.505 59.255 94.025 ;
        RECT 59.425 94.245 59.700 94.945 ;
        RECT 59.870 94.570 60.125 95.115 ;
        RECT 60.295 94.605 60.775 94.945 ;
        RECT 60.950 94.560 61.555 95.115 ;
        RECT 60.940 94.460 61.555 94.560 ;
        RECT 60.940 94.435 61.125 94.460 ;
        RECT 57.585 92.565 59.255 93.335 ;
        RECT 59.425 93.215 59.595 94.245 ;
        RECT 59.870 94.115 60.625 94.365 ;
        RECT 60.795 94.190 61.125 94.435 ;
        RECT 59.870 94.080 60.640 94.115 ;
        RECT 59.870 94.070 60.655 94.080 ;
        RECT 59.765 94.055 60.660 94.070 ;
        RECT 59.765 94.040 60.680 94.055 ;
        RECT 59.765 94.030 60.700 94.040 ;
        RECT 59.765 94.020 60.725 94.030 ;
        RECT 59.765 93.990 60.795 94.020 ;
        RECT 59.765 93.960 60.815 93.990 ;
        RECT 59.765 93.930 60.835 93.960 ;
        RECT 59.765 93.905 60.865 93.930 ;
        RECT 59.765 93.870 60.900 93.905 ;
        RECT 59.765 93.865 60.930 93.870 ;
        RECT 59.765 93.470 59.995 93.865 ;
        RECT 60.540 93.860 60.930 93.865 ;
        RECT 60.565 93.850 60.930 93.860 ;
        RECT 60.580 93.845 60.930 93.850 ;
        RECT 60.595 93.840 60.930 93.845 ;
        RECT 61.295 93.840 61.555 94.290 ;
        RECT 61.735 94.145 62.065 94.930 ;
        RECT 61.735 93.975 62.415 94.145 ;
        RECT 62.595 93.975 62.925 95.115 ;
        RECT 63.105 94.025 65.695 95.115 ;
        RECT 66.325 94.605 67.515 94.895 ;
        RECT 60.595 93.835 61.555 93.840 ;
        RECT 60.605 93.825 61.555 93.835 ;
        RECT 60.615 93.820 61.555 93.825 ;
        RECT 60.625 93.810 61.555 93.820 ;
        RECT 60.630 93.800 61.555 93.810 ;
        RECT 60.635 93.795 61.555 93.800 ;
        RECT 60.645 93.780 61.555 93.795 ;
        RECT 60.650 93.765 61.555 93.780 ;
        RECT 60.660 93.740 61.555 93.765 ;
        RECT 60.165 93.270 60.495 93.695 ;
        RECT 59.425 92.735 59.685 93.215 ;
        RECT 59.855 92.565 60.105 93.105 ;
        RECT 60.275 92.785 60.495 93.270 ;
        RECT 60.665 93.670 61.555 93.740 ;
        RECT 60.665 92.945 60.835 93.670 ;
        RECT 61.725 93.555 62.075 93.805 ;
        RECT 61.005 93.115 61.555 93.500 ;
        RECT 62.245 93.375 62.415 93.975 ;
        RECT 62.585 93.555 62.935 93.805 ;
        RECT 60.665 92.775 61.555 92.945 ;
        RECT 61.745 92.565 61.985 93.375 ;
        RECT 62.155 92.735 62.485 93.375 ;
        RECT 62.655 92.565 62.925 93.375 ;
        RECT 63.105 93.335 64.315 93.855 ;
        RECT 64.485 93.505 65.695 94.025 ;
        RECT 66.345 94.265 67.515 94.435 ;
        RECT 67.685 94.315 67.965 95.115 ;
        RECT 66.345 93.975 66.670 94.265 ;
        RECT 67.345 94.145 67.515 94.265 ;
        RECT 66.840 93.805 67.035 94.095 ;
        RECT 67.345 93.975 68.005 94.145 ;
        RECT 68.175 93.975 68.450 94.945 ;
        RECT 68.625 94.025 69.835 95.115 ;
        RECT 67.835 93.805 68.005 93.975 ;
        RECT 66.325 93.475 66.670 93.805 ;
        RECT 66.840 93.475 67.665 93.805 ;
        RECT 67.835 93.475 68.110 93.805 ;
        RECT 63.105 92.565 65.695 93.335 ;
        RECT 67.835 93.305 68.005 93.475 ;
        RECT 66.340 93.135 68.005 93.305 ;
        RECT 68.280 93.240 68.450 93.975 ;
        RECT 66.340 92.785 66.595 93.135 ;
        RECT 66.765 92.565 67.095 92.965 ;
        RECT 67.265 92.785 67.435 93.135 ;
        RECT 67.605 92.565 67.985 92.965 ;
        RECT 68.175 92.895 68.450 93.240 ;
        RECT 68.625 93.315 69.145 93.855 ;
        RECT 69.315 93.485 69.835 94.025 ;
        RECT 70.005 93.950 70.295 95.115 ;
        RECT 71.385 94.355 71.900 94.765 ;
        RECT 72.135 94.355 72.305 95.115 ;
        RECT 72.475 94.775 74.505 94.945 ;
        RECT 71.385 93.545 71.725 94.355 ;
        RECT 72.475 94.110 72.645 94.775 ;
        RECT 73.040 94.435 74.165 94.605 ;
        RECT 71.895 93.920 72.645 94.110 ;
        RECT 72.815 94.095 73.825 94.265 ;
        RECT 71.385 93.375 72.615 93.545 ;
        RECT 68.625 92.565 69.835 93.315 ;
        RECT 70.005 92.565 70.295 93.290 ;
        RECT 71.660 92.770 71.905 93.375 ;
        RECT 72.125 92.565 72.635 93.100 ;
        RECT 72.815 92.735 73.005 94.095 ;
        RECT 73.175 93.075 73.450 93.895 ;
        RECT 73.655 93.295 73.825 94.095 ;
        RECT 73.995 93.305 74.165 94.435 ;
        RECT 74.335 93.805 74.505 94.775 ;
        RECT 74.675 93.975 74.845 95.115 ;
        RECT 75.015 93.975 75.350 94.945 ;
        RECT 75.525 94.680 80.870 95.115 ;
        RECT 74.335 93.475 74.530 93.805 ;
        RECT 74.755 93.475 75.010 93.805 ;
        RECT 74.755 93.305 74.925 93.475 ;
        RECT 75.180 93.305 75.350 93.975 ;
        RECT 73.995 93.135 74.925 93.305 ;
        RECT 73.995 93.100 74.170 93.135 ;
        RECT 73.175 92.905 73.455 93.075 ;
        RECT 73.175 92.735 73.450 92.905 ;
        RECT 73.640 92.735 74.170 93.100 ;
        RECT 74.595 92.565 74.925 92.965 ;
        RECT 75.095 92.735 75.350 93.305 ;
        RECT 77.110 93.110 77.450 93.940 ;
        RECT 78.930 93.430 79.280 94.680 ;
        RECT 81.045 94.025 82.715 95.115 ;
        RECT 81.045 93.335 81.795 93.855 ;
        RECT 81.965 93.505 82.715 94.025 ;
        RECT 82.885 94.025 84.095 95.115 ;
        RECT 82.885 93.485 83.405 94.025 ;
        RECT 75.525 92.565 80.870 93.110 ;
        RECT 81.045 92.565 82.715 93.335 ;
        RECT 83.575 93.315 84.095 93.855 ;
        RECT 82.885 92.565 84.095 93.315 ;
        RECT 5.520 92.395 84.180 92.565 ;
        RECT 5.605 91.645 6.815 92.395 ;
        RECT 6.985 91.645 8.195 92.395 ;
        RECT 8.370 91.655 8.625 92.225 ;
        RECT 8.795 91.995 9.125 92.395 ;
        RECT 9.550 91.860 10.080 92.225 ;
        RECT 9.550 91.825 9.725 91.860 ;
        RECT 8.795 91.655 9.725 91.825 ;
        RECT 5.605 91.105 6.125 91.645 ;
        RECT 6.295 90.935 6.815 91.475 ;
        RECT 6.985 91.105 7.505 91.645 ;
        RECT 7.675 90.935 8.195 91.475 ;
        RECT 5.605 89.845 6.815 90.935 ;
        RECT 6.985 89.845 8.195 90.935 ;
        RECT 8.370 90.985 8.540 91.655 ;
        RECT 8.795 91.485 8.965 91.655 ;
        RECT 8.710 91.155 8.965 91.485 ;
        RECT 9.190 91.155 9.385 91.485 ;
        RECT 8.370 90.015 8.705 90.985 ;
        RECT 8.875 89.845 9.045 90.985 ;
        RECT 9.215 90.185 9.385 91.155 ;
        RECT 9.555 90.525 9.725 91.655 ;
        RECT 9.895 90.865 10.065 91.665 ;
        RECT 10.270 91.375 10.545 92.225 ;
        RECT 10.265 91.205 10.545 91.375 ;
        RECT 10.270 91.065 10.545 91.205 ;
        RECT 10.715 90.865 10.905 92.225 ;
        RECT 11.085 91.860 11.595 92.395 ;
        RECT 11.815 91.585 12.060 92.190 ;
        RECT 12.985 91.825 13.240 92.175 ;
        RECT 13.410 91.995 13.740 92.395 ;
        RECT 13.910 91.825 14.080 92.175 ;
        RECT 14.250 91.995 14.630 92.395 ;
        RECT 12.985 91.655 14.650 91.825 ;
        RECT 14.820 91.720 15.095 92.065 ;
        RECT 11.105 91.415 12.335 91.585 ;
        RECT 14.480 91.485 14.650 91.655 ;
        RECT 9.895 90.695 10.905 90.865 ;
        RECT 11.075 90.850 11.825 91.040 ;
        RECT 9.555 90.355 10.680 90.525 ;
        RECT 11.075 90.185 11.245 90.850 ;
        RECT 11.995 90.605 12.335 91.415 ;
        RECT 12.965 91.155 13.315 91.485 ;
        RECT 13.485 91.155 14.310 91.485 ;
        RECT 14.480 91.155 14.755 91.485 ;
        RECT 9.215 90.015 11.245 90.185 ;
        RECT 11.415 89.845 11.585 90.605 ;
        RECT 11.820 90.195 12.335 90.605 ;
        RECT 12.985 90.695 13.315 90.985 ;
        RECT 13.485 90.865 13.710 91.155 ;
        RECT 14.480 90.985 14.650 91.155 ;
        RECT 14.925 90.985 15.095 91.720 ;
        RECT 15.265 91.565 15.555 92.395 ;
        RECT 15.725 91.625 18.315 92.395 ;
        RECT 18.575 91.845 18.745 92.135 ;
        RECT 18.915 92.015 19.245 92.395 ;
        RECT 18.575 91.675 19.240 91.845 ;
        RECT 15.725 91.105 16.935 91.625 ;
        RECT 13.980 90.815 14.650 90.985 ;
        RECT 13.980 90.695 14.150 90.815 ;
        RECT 12.985 90.525 14.150 90.695 ;
        RECT 12.965 90.065 14.160 90.355 ;
        RECT 14.330 89.845 14.610 90.645 ;
        RECT 14.820 90.015 15.095 90.985 ;
        RECT 15.265 89.845 15.555 91.050 ;
        RECT 17.105 90.935 18.315 91.455 ;
        RECT 15.725 89.845 18.315 90.935 ;
        RECT 18.490 90.855 18.840 91.505 ;
        RECT 19.010 90.685 19.240 91.675 ;
        RECT 18.575 90.515 19.240 90.685 ;
        RECT 18.575 90.015 18.745 90.515 ;
        RECT 18.915 89.845 19.245 90.345 ;
        RECT 19.415 90.015 19.600 92.135 ;
        RECT 19.855 91.935 20.105 92.395 ;
        RECT 20.275 91.945 20.610 92.115 ;
        RECT 20.805 91.945 21.480 92.115 ;
        RECT 20.275 91.805 20.445 91.945 ;
        RECT 19.770 90.815 20.050 91.765 ;
        RECT 20.220 91.675 20.445 91.805 ;
        RECT 20.220 90.570 20.390 91.675 ;
        RECT 20.615 91.525 21.140 91.745 ;
        RECT 20.560 90.760 20.800 91.355 ;
        RECT 20.970 90.825 21.140 91.525 ;
        RECT 21.310 91.165 21.480 91.945 ;
        RECT 21.800 91.895 22.170 92.395 ;
        RECT 22.350 91.945 22.755 92.115 ;
        RECT 22.925 91.945 23.710 92.115 ;
        RECT 22.350 91.715 22.520 91.945 ;
        RECT 21.690 91.415 22.520 91.715 ;
        RECT 22.905 91.445 23.370 91.775 ;
        RECT 21.690 91.385 21.890 91.415 ;
        RECT 22.010 91.165 22.180 91.235 ;
        RECT 21.310 90.995 22.180 91.165 ;
        RECT 21.670 90.905 22.180 90.995 ;
        RECT 20.220 90.440 20.525 90.570 ;
        RECT 20.970 90.460 21.500 90.825 ;
        RECT 19.840 89.845 20.105 90.305 ;
        RECT 20.275 90.015 20.525 90.440 ;
        RECT 21.670 90.290 21.840 90.905 ;
        RECT 20.735 90.120 21.840 90.290 ;
        RECT 22.010 89.845 22.180 90.645 ;
        RECT 22.350 90.345 22.520 91.415 ;
        RECT 22.690 90.515 22.880 91.235 ;
        RECT 23.050 90.485 23.370 91.445 ;
        RECT 23.540 91.485 23.710 91.945 ;
        RECT 23.985 91.865 24.195 92.395 ;
        RECT 24.455 91.655 24.785 92.180 ;
        RECT 24.955 91.785 25.125 92.395 ;
        RECT 25.295 91.740 25.625 92.175 ;
        RECT 25.795 91.880 25.965 92.395 ;
        RECT 25.295 91.655 25.675 91.740 ;
        RECT 24.585 91.485 24.785 91.655 ;
        RECT 25.450 91.615 25.675 91.655 ;
        RECT 23.540 91.155 24.415 91.485 ;
        RECT 24.585 91.155 25.335 91.485 ;
        RECT 22.350 90.015 22.600 90.345 ;
        RECT 23.540 90.315 23.710 91.155 ;
        RECT 24.585 90.950 24.775 91.155 ;
        RECT 25.505 91.035 25.675 91.615 ;
        RECT 25.460 90.985 25.675 91.035 ;
        RECT 23.880 90.575 24.775 90.950 ;
        RECT 25.285 90.905 25.675 90.985 ;
        RECT 27.230 91.655 27.485 92.225 ;
        RECT 27.655 91.995 27.985 92.395 ;
        RECT 28.410 91.860 28.940 92.225 ;
        RECT 29.130 92.055 29.405 92.225 ;
        RECT 29.125 91.885 29.405 92.055 ;
        RECT 28.410 91.825 28.585 91.860 ;
        RECT 27.655 91.655 28.585 91.825 ;
        RECT 27.230 90.985 27.400 91.655 ;
        RECT 27.655 91.485 27.825 91.655 ;
        RECT 27.570 91.155 27.825 91.485 ;
        RECT 28.050 91.155 28.245 91.485 ;
        RECT 22.825 90.145 23.710 90.315 ;
        RECT 23.890 89.845 24.205 90.345 ;
        RECT 24.435 90.015 24.775 90.575 ;
        RECT 24.945 89.845 25.115 90.855 ;
        RECT 25.285 90.060 25.615 90.905 ;
        RECT 25.785 89.845 25.955 90.760 ;
        RECT 27.230 90.015 27.565 90.985 ;
        RECT 27.735 89.845 27.905 90.985 ;
        RECT 28.075 90.185 28.245 91.155 ;
        RECT 28.415 90.525 28.585 91.655 ;
        RECT 28.755 90.865 28.925 91.665 ;
        RECT 29.130 91.065 29.405 91.885 ;
        RECT 29.575 90.865 29.765 92.225 ;
        RECT 29.945 91.860 30.455 92.395 ;
        RECT 30.675 91.585 30.920 92.190 ;
        RECT 31.365 91.670 31.655 92.395 ;
        RECT 32.290 91.655 32.545 92.225 ;
        RECT 32.715 91.995 33.045 92.395 ;
        RECT 33.470 91.860 34.000 92.225 ;
        RECT 33.470 91.825 33.645 91.860 ;
        RECT 32.715 91.655 33.645 91.825 ;
        RECT 29.965 91.415 31.195 91.585 ;
        RECT 28.755 90.695 29.765 90.865 ;
        RECT 29.935 90.850 30.685 91.040 ;
        RECT 28.415 90.355 29.540 90.525 ;
        RECT 29.935 90.185 30.105 90.850 ;
        RECT 30.855 90.605 31.195 91.415 ;
        RECT 28.075 90.015 30.105 90.185 ;
        RECT 30.275 89.845 30.445 90.605 ;
        RECT 30.680 90.195 31.195 90.605 ;
        RECT 31.365 89.845 31.655 91.010 ;
        RECT 32.290 90.985 32.460 91.655 ;
        RECT 32.715 91.485 32.885 91.655 ;
        RECT 32.630 91.155 32.885 91.485 ;
        RECT 33.110 91.155 33.305 91.485 ;
        RECT 32.290 90.015 32.625 90.985 ;
        RECT 32.795 89.845 32.965 90.985 ;
        RECT 33.135 90.185 33.305 91.155 ;
        RECT 33.475 90.525 33.645 91.655 ;
        RECT 33.815 90.865 33.985 91.665 ;
        RECT 34.190 91.375 34.465 92.225 ;
        RECT 34.185 91.205 34.465 91.375 ;
        RECT 34.190 91.065 34.465 91.205 ;
        RECT 34.635 90.865 34.825 92.225 ;
        RECT 35.005 91.860 35.515 92.395 ;
        RECT 35.735 91.585 35.980 92.190 ;
        RECT 36.425 92.015 37.315 92.185 ;
        RECT 35.025 91.415 36.255 91.585 ;
        RECT 36.425 91.460 36.975 91.845 ;
        RECT 33.815 90.695 34.825 90.865 ;
        RECT 34.995 90.850 35.745 91.040 ;
        RECT 33.475 90.355 34.600 90.525 ;
        RECT 34.995 90.185 35.165 90.850 ;
        RECT 35.915 90.605 36.255 91.415 ;
        RECT 37.145 91.290 37.315 92.015 ;
        RECT 36.425 91.220 37.315 91.290 ;
        RECT 37.485 91.690 37.705 92.175 ;
        RECT 37.875 91.855 38.125 92.395 ;
        RECT 38.295 91.745 38.555 92.225 ;
        RECT 38.725 91.850 44.070 92.395 ;
        RECT 37.485 91.265 37.815 91.690 ;
        RECT 36.425 91.195 37.320 91.220 ;
        RECT 36.425 91.180 37.330 91.195 ;
        RECT 36.425 91.165 37.335 91.180 ;
        RECT 36.425 91.160 37.345 91.165 ;
        RECT 36.425 91.150 37.350 91.160 ;
        RECT 36.425 91.140 37.355 91.150 ;
        RECT 36.425 91.135 37.365 91.140 ;
        RECT 36.425 91.125 37.375 91.135 ;
        RECT 36.425 91.120 37.385 91.125 ;
        RECT 36.425 90.670 36.685 91.120 ;
        RECT 37.050 91.115 37.385 91.120 ;
        RECT 37.050 91.110 37.400 91.115 ;
        RECT 37.050 91.100 37.415 91.110 ;
        RECT 37.050 91.095 37.440 91.100 ;
        RECT 37.985 91.095 38.215 91.490 ;
        RECT 37.050 91.090 38.215 91.095 ;
        RECT 37.080 91.055 38.215 91.090 ;
        RECT 37.115 91.030 38.215 91.055 ;
        RECT 37.145 91.000 38.215 91.030 ;
        RECT 37.165 90.970 38.215 91.000 ;
        RECT 37.185 90.940 38.215 90.970 ;
        RECT 37.255 90.930 38.215 90.940 ;
        RECT 37.280 90.920 38.215 90.930 ;
        RECT 37.300 90.905 38.215 90.920 ;
        RECT 37.320 90.890 38.215 90.905 ;
        RECT 37.325 90.880 38.110 90.890 ;
        RECT 37.340 90.845 38.110 90.880 ;
        RECT 33.135 90.015 35.165 90.185 ;
        RECT 35.335 89.845 35.505 90.605 ;
        RECT 35.740 90.195 36.255 90.605 ;
        RECT 36.855 90.525 37.185 90.770 ;
        RECT 37.355 90.595 38.110 90.845 ;
        RECT 38.385 90.715 38.555 91.745 ;
        RECT 40.310 91.020 40.650 91.850 ;
        RECT 44.245 91.625 46.835 92.395 ;
        RECT 47.515 91.740 47.845 92.175 ;
        RECT 48.015 91.785 48.185 92.395 ;
        RECT 47.465 91.655 47.845 91.740 ;
        RECT 48.355 91.655 48.685 92.180 ;
        RECT 48.945 91.865 49.155 92.395 ;
        RECT 49.430 91.945 50.215 92.115 ;
        RECT 50.385 91.945 50.790 92.115 ;
        RECT 36.855 90.500 37.040 90.525 ;
        RECT 36.425 90.400 37.040 90.500 ;
        RECT 36.425 89.845 37.030 90.400 ;
        RECT 37.205 90.015 37.685 90.355 ;
        RECT 37.855 89.845 38.110 90.390 ;
        RECT 38.280 90.015 38.555 90.715 ;
        RECT 42.130 90.280 42.480 91.530 ;
        RECT 44.245 91.105 45.455 91.625 ;
        RECT 47.465 91.615 47.690 91.655 ;
        RECT 45.625 90.935 46.835 91.455 ;
        RECT 38.725 89.845 44.070 90.280 ;
        RECT 44.245 89.845 46.835 90.935 ;
        RECT 47.465 91.035 47.635 91.615 ;
        RECT 48.355 91.485 48.555 91.655 ;
        RECT 49.430 91.485 49.600 91.945 ;
        RECT 47.805 91.155 48.555 91.485 ;
        RECT 48.725 91.155 49.600 91.485 ;
        RECT 47.465 90.985 47.680 91.035 ;
        RECT 47.465 90.905 47.855 90.985 ;
        RECT 47.525 90.060 47.855 90.905 ;
        RECT 48.365 90.950 48.555 91.155 ;
        RECT 48.025 89.845 48.195 90.855 ;
        RECT 48.365 90.575 49.260 90.950 ;
        RECT 48.365 90.015 48.705 90.575 ;
        RECT 48.935 89.845 49.250 90.345 ;
        RECT 49.430 90.315 49.600 91.155 ;
        RECT 49.770 91.445 50.235 91.775 ;
        RECT 50.620 91.715 50.790 91.945 ;
        RECT 50.970 91.895 51.340 92.395 ;
        RECT 51.660 91.945 52.335 92.115 ;
        RECT 52.530 91.945 52.865 92.115 ;
        RECT 49.770 90.485 50.090 91.445 ;
        RECT 50.620 91.415 51.450 91.715 ;
        RECT 50.260 90.515 50.450 91.235 ;
        RECT 50.620 90.345 50.790 91.415 ;
        RECT 51.250 91.385 51.450 91.415 ;
        RECT 50.960 91.165 51.130 91.235 ;
        RECT 51.660 91.165 51.830 91.945 ;
        RECT 52.695 91.805 52.865 91.945 ;
        RECT 53.035 91.935 53.285 92.395 ;
        RECT 50.960 90.995 51.830 91.165 ;
        RECT 52.000 91.525 52.525 91.745 ;
        RECT 52.695 91.675 52.920 91.805 ;
        RECT 50.960 90.905 51.470 90.995 ;
        RECT 49.430 90.145 50.315 90.315 ;
        RECT 50.540 90.015 50.790 90.345 ;
        RECT 50.960 89.845 51.130 90.645 ;
        RECT 51.300 90.290 51.470 90.905 ;
        RECT 52.000 90.825 52.170 91.525 ;
        RECT 51.640 90.460 52.170 90.825 ;
        RECT 52.340 90.760 52.580 91.355 ;
        RECT 52.750 90.570 52.920 91.675 ;
        RECT 53.090 90.815 53.370 91.765 ;
        RECT 52.615 90.440 52.920 90.570 ;
        RECT 51.300 90.120 52.405 90.290 ;
        RECT 52.615 90.015 52.865 90.440 ;
        RECT 53.035 89.845 53.300 90.305 ;
        RECT 53.540 90.015 53.725 92.135 ;
        RECT 53.895 92.015 54.225 92.395 ;
        RECT 54.395 91.845 54.565 92.135 ;
        RECT 53.900 91.675 54.565 91.845 ;
        RECT 53.900 90.685 54.130 91.675 ;
        RECT 54.825 91.625 56.495 92.395 ;
        RECT 57.125 91.670 57.415 92.395 ;
        RECT 57.585 91.895 57.845 92.225 ;
        RECT 58.015 92.035 58.345 92.395 ;
        RECT 58.600 92.015 59.900 92.225 ;
        RECT 57.585 91.885 57.815 91.895 ;
        RECT 54.300 90.855 54.650 91.505 ;
        RECT 54.825 91.105 55.575 91.625 ;
        RECT 55.745 90.935 56.495 91.455 ;
        RECT 53.900 90.515 54.565 90.685 ;
        RECT 53.895 89.845 54.225 90.345 ;
        RECT 54.395 90.015 54.565 90.515 ;
        RECT 54.825 89.845 56.495 90.935 ;
        RECT 57.125 89.845 57.415 91.010 ;
        RECT 57.585 90.695 57.755 91.885 ;
        RECT 58.600 91.865 58.770 92.015 ;
        RECT 58.015 91.740 58.770 91.865 ;
        RECT 57.925 91.695 58.770 91.740 ;
        RECT 57.925 91.575 58.195 91.695 ;
        RECT 57.925 91.000 58.095 91.575 ;
        RECT 58.325 91.135 58.735 91.440 ;
        RECT 59.025 91.405 59.235 91.805 ;
        RECT 58.905 91.195 59.235 91.405 ;
        RECT 59.480 91.405 59.700 91.805 ;
        RECT 60.175 91.630 60.630 92.395 ;
        RECT 59.480 91.195 59.955 91.405 ;
        RECT 60.145 91.205 60.635 91.405 ;
        RECT 57.925 90.965 58.125 91.000 ;
        RECT 59.455 90.965 60.630 91.025 ;
        RECT 57.925 90.855 60.630 90.965 ;
        RECT 57.985 90.795 59.785 90.855 ;
        RECT 59.455 90.765 59.785 90.795 ;
        RECT 57.585 90.015 57.845 90.695 ;
        RECT 58.015 89.845 58.265 90.625 ;
        RECT 58.515 90.595 59.350 90.605 ;
        RECT 59.940 90.595 60.125 90.685 ;
        RECT 58.515 90.395 60.125 90.595 ;
        RECT 58.515 90.015 58.765 90.395 ;
        RECT 59.895 90.355 60.125 90.395 ;
        RECT 60.375 90.235 60.630 90.855 ;
        RECT 58.935 89.845 59.290 90.225 ;
        RECT 60.295 90.015 60.630 90.235 ;
        RECT 61.270 90.795 61.605 92.215 ;
        RECT 61.785 92.025 62.530 92.395 ;
        RECT 63.095 91.855 63.350 92.215 ;
        RECT 63.530 92.025 63.860 92.395 ;
        RECT 64.040 91.855 64.265 92.215 ;
        RECT 61.780 91.665 64.265 91.855 ;
        RECT 61.780 90.975 62.005 91.665 ;
        RECT 64.485 91.625 66.155 92.395 ;
        RECT 66.340 91.825 66.595 92.175 ;
        RECT 66.765 91.995 67.095 92.395 ;
        RECT 67.265 91.825 67.435 92.175 ;
        RECT 67.605 91.995 67.985 92.395 ;
        RECT 66.340 91.655 68.005 91.825 ;
        RECT 68.175 91.720 68.450 92.065 ;
        RECT 68.790 91.885 69.030 92.395 ;
        RECT 69.210 91.885 69.490 92.215 ;
        RECT 69.720 91.885 69.935 92.395 ;
        RECT 62.205 91.155 62.485 91.485 ;
        RECT 62.665 91.155 63.240 91.485 ;
        RECT 63.420 91.155 63.855 91.485 ;
        RECT 64.035 91.155 64.305 91.485 ;
        RECT 64.485 91.105 65.235 91.625 ;
        RECT 67.835 91.485 68.005 91.655 ;
        RECT 61.780 90.795 64.275 90.975 ;
        RECT 65.405 90.935 66.155 91.455 ;
        RECT 66.325 91.155 66.670 91.485 ;
        RECT 66.840 91.155 67.665 91.485 ;
        RECT 67.835 91.155 68.110 91.485 ;
        RECT 61.270 90.025 61.535 90.795 ;
        RECT 61.705 89.845 62.035 90.565 ;
        RECT 62.225 90.385 63.415 90.615 ;
        RECT 62.225 90.025 62.485 90.385 ;
        RECT 62.655 89.845 62.985 90.215 ;
        RECT 63.155 90.025 63.415 90.385 ;
        RECT 63.985 90.025 64.275 90.795 ;
        RECT 64.485 89.845 66.155 90.935 ;
        RECT 66.345 90.695 66.670 90.985 ;
        RECT 66.840 90.865 67.035 91.155 ;
        RECT 67.835 90.985 68.005 91.155 ;
        RECT 68.280 90.985 68.450 91.720 ;
        RECT 68.685 91.155 69.040 91.715 ;
        RECT 69.210 90.985 69.380 91.885 ;
        RECT 69.550 91.155 69.815 91.715 ;
        RECT 70.105 91.655 70.720 92.225 ;
        RECT 70.065 90.985 70.235 91.485 ;
        RECT 67.345 90.815 68.005 90.985 ;
        RECT 67.345 90.695 67.515 90.815 ;
        RECT 66.345 90.525 67.515 90.695 ;
        RECT 66.325 90.065 67.515 90.355 ;
        RECT 67.685 89.845 67.965 90.645 ;
        RECT 68.175 90.015 68.450 90.985 ;
        RECT 68.810 90.815 70.235 90.985 ;
        RECT 68.810 90.640 69.200 90.815 ;
        RECT 69.685 89.845 70.015 90.645 ;
        RECT 70.405 90.635 70.720 91.655 ;
        RECT 71.850 91.630 72.305 92.395 ;
        RECT 72.580 92.015 73.880 92.225 ;
        RECT 74.135 92.035 74.465 92.395 ;
        RECT 73.710 91.865 73.880 92.015 ;
        RECT 74.635 91.895 74.895 92.225 ;
        RECT 74.665 91.885 74.895 91.895 ;
        RECT 72.780 91.405 73.000 91.805 ;
        RECT 71.845 91.205 72.335 91.405 ;
        RECT 72.525 91.195 73.000 91.405 ;
        RECT 73.245 91.405 73.455 91.805 ;
        RECT 73.710 91.740 74.465 91.865 ;
        RECT 73.710 91.695 74.555 91.740 ;
        RECT 74.285 91.575 74.555 91.695 ;
        RECT 73.245 91.195 73.575 91.405 ;
        RECT 73.745 91.135 74.155 91.440 ;
        RECT 70.185 90.015 70.720 90.635 ;
        RECT 71.850 90.965 73.025 91.025 ;
        RECT 74.385 91.000 74.555 91.575 ;
        RECT 74.355 90.965 74.555 91.000 ;
        RECT 71.850 90.855 74.555 90.965 ;
        RECT 71.850 90.235 72.105 90.855 ;
        RECT 72.695 90.795 74.495 90.855 ;
        RECT 72.695 90.765 73.025 90.795 ;
        RECT 74.725 90.695 74.895 91.885 ;
        RECT 75.065 91.850 80.410 92.395 ;
        RECT 76.650 91.020 76.990 91.850 ;
        RECT 80.585 91.625 82.255 92.395 ;
        RECT 82.885 91.645 84.095 92.395 ;
        RECT 72.355 90.595 72.540 90.685 ;
        RECT 73.130 90.595 73.965 90.605 ;
        RECT 72.355 90.395 73.965 90.595 ;
        RECT 72.355 90.355 72.585 90.395 ;
        RECT 71.850 90.015 72.185 90.235 ;
        RECT 73.190 89.845 73.545 90.225 ;
        RECT 73.715 90.015 73.965 90.395 ;
        RECT 74.215 89.845 74.465 90.625 ;
        RECT 74.635 90.015 74.895 90.695 ;
        RECT 78.470 90.280 78.820 91.530 ;
        RECT 80.585 91.105 81.335 91.625 ;
        RECT 81.505 90.935 82.255 91.455 ;
        RECT 75.065 89.845 80.410 90.280 ;
        RECT 80.585 89.845 82.255 90.935 ;
        RECT 82.885 90.935 83.405 91.475 ;
        RECT 83.575 91.105 84.095 91.645 ;
        RECT 82.885 89.845 84.095 90.935 ;
        RECT 5.520 89.675 84.180 89.845 ;
        RECT 5.605 88.585 6.815 89.675 ;
        RECT 7.075 89.005 7.245 89.505 ;
        RECT 7.415 89.175 7.745 89.675 ;
        RECT 7.075 88.835 7.740 89.005 ;
        RECT 5.605 87.875 6.125 88.415 ;
        RECT 6.295 88.045 6.815 88.585 ;
        RECT 6.990 88.015 7.340 88.665 ;
        RECT 5.605 87.125 6.815 87.875 ;
        RECT 7.510 87.845 7.740 88.835 ;
        RECT 7.075 87.675 7.740 87.845 ;
        RECT 7.075 87.385 7.245 87.675 ;
        RECT 7.415 87.125 7.745 87.505 ;
        RECT 7.915 87.385 8.100 89.505 ;
        RECT 8.340 89.215 8.605 89.675 ;
        RECT 8.775 89.080 9.025 89.505 ;
        RECT 9.235 89.230 10.340 89.400 ;
        RECT 8.720 88.950 9.025 89.080 ;
        RECT 8.270 87.755 8.550 88.705 ;
        RECT 8.720 87.845 8.890 88.950 ;
        RECT 9.060 88.165 9.300 88.760 ;
        RECT 9.470 88.695 10.000 89.060 ;
        RECT 9.470 87.995 9.640 88.695 ;
        RECT 10.170 88.615 10.340 89.230 ;
        RECT 10.510 88.875 10.680 89.675 ;
        RECT 10.850 89.175 11.100 89.505 ;
        RECT 11.325 89.205 12.210 89.375 ;
        RECT 10.170 88.525 10.680 88.615 ;
        RECT 8.720 87.715 8.945 87.845 ;
        RECT 9.115 87.775 9.640 87.995 ;
        RECT 9.810 88.355 10.680 88.525 ;
        RECT 8.355 87.125 8.605 87.585 ;
        RECT 8.775 87.575 8.945 87.715 ;
        RECT 9.810 87.575 9.980 88.355 ;
        RECT 10.510 88.285 10.680 88.355 ;
        RECT 10.190 88.105 10.390 88.135 ;
        RECT 10.850 88.105 11.020 89.175 ;
        RECT 11.190 88.285 11.380 89.005 ;
        RECT 10.190 87.805 11.020 88.105 ;
        RECT 11.550 88.075 11.870 89.035 ;
        RECT 8.775 87.405 9.110 87.575 ;
        RECT 9.305 87.405 9.980 87.575 ;
        RECT 10.300 87.125 10.670 87.625 ;
        RECT 10.850 87.575 11.020 87.805 ;
        RECT 11.405 87.745 11.870 88.075 ;
        RECT 12.040 88.365 12.210 89.205 ;
        RECT 12.390 89.175 12.705 89.675 ;
        RECT 12.935 88.945 13.275 89.505 ;
        RECT 12.380 88.570 13.275 88.945 ;
        RECT 13.445 88.665 13.615 89.675 ;
        RECT 13.085 88.365 13.275 88.570 ;
        RECT 13.785 88.615 14.115 89.460 ;
        RECT 14.285 88.760 14.455 89.675 ;
        RECT 15.725 89.120 16.330 89.675 ;
        RECT 16.505 89.165 16.985 89.505 ;
        RECT 17.155 89.130 17.410 89.675 ;
        RECT 15.725 89.020 16.340 89.120 ;
        RECT 16.155 88.995 16.340 89.020 ;
        RECT 13.785 88.535 14.175 88.615 ;
        RECT 13.960 88.485 14.175 88.535 ;
        RECT 12.040 88.035 12.915 88.365 ;
        RECT 13.085 88.035 13.835 88.365 ;
        RECT 12.040 87.575 12.210 88.035 ;
        RECT 13.085 87.865 13.285 88.035 ;
        RECT 14.005 87.905 14.175 88.485 ;
        RECT 15.725 88.400 15.985 88.850 ;
        RECT 16.155 88.750 16.485 88.995 ;
        RECT 16.655 88.675 17.410 88.925 ;
        RECT 17.580 88.805 17.855 89.505 ;
        RECT 16.640 88.640 17.410 88.675 ;
        RECT 16.625 88.630 17.410 88.640 ;
        RECT 16.620 88.615 17.515 88.630 ;
        RECT 16.600 88.600 17.515 88.615 ;
        RECT 16.580 88.590 17.515 88.600 ;
        RECT 16.555 88.580 17.515 88.590 ;
        RECT 16.485 88.550 17.515 88.580 ;
        RECT 16.465 88.520 17.515 88.550 ;
        RECT 16.445 88.490 17.515 88.520 ;
        RECT 16.415 88.465 17.515 88.490 ;
        RECT 16.380 88.430 17.515 88.465 ;
        RECT 16.350 88.425 17.515 88.430 ;
        RECT 16.350 88.420 16.740 88.425 ;
        RECT 16.350 88.410 16.715 88.420 ;
        RECT 16.350 88.405 16.700 88.410 ;
        RECT 16.350 88.400 16.685 88.405 ;
        RECT 15.725 88.395 16.685 88.400 ;
        RECT 15.725 88.385 16.675 88.395 ;
        RECT 15.725 88.380 16.665 88.385 ;
        RECT 15.725 88.370 16.655 88.380 ;
        RECT 15.725 88.360 16.650 88.370 ;
        RECT 15.725 88.355 16.645 88.360 ;
        RECT 15.725 88.340 16.635 88.355 ;
        RECT 15.725 88.325 16.630 88.340 ;
        RECT 15.725 88.300 16.620 88.325 ;
        RECT 15.725 88.230 16.615 88.300 ;
        RECT 13.950 87.865 14.175 87.905 ;
        RECT 10.850 87.405 11.255 87.575 ;
        RECT 11.425 87.405 12.210 87.575 ;
        RECT 12.485 87.125 12.695 87.655 ;
        RECT 12.955 87.340 13.285 87.865 ;
        RECT 13.795 87.780 14.175 87.865 ;
        RECT 13.455 87.125 13.625 87.735 ;
        RECT 13.795 87.345 14.125 87.780 ;
        RECT 15.725 87.675 16.275 88.060 ;
        RECT 14.295 87.125 14.465 87.640 ;
        RECT 16.445 87.505 16.615 88.230 ;
        RECT 15.725 87.335 16.615 87.505 ;
        RECT 16.785 87.830 17.115 88.255 ;
        RECT 17.285 88.030 17.515 88.425 ;
        RECT 16.785 87.345 17.005 87.830 ;
        RECT 17.685 87.775 17.855 88.805 ;
        RECT 18.485 88.510 18.775 89.675 ;
        RECT 19.410 88.535 19.745 89.505 ;
        RECT 19.915 88.535 20.085 89.675 ;
        RECT 20.255 89.335 22.285 89.505 ;
        RECT 19.410 87.865 19.580 88.535 ;
        RECT 20.255 88.365 20.425 89.335 ;
        RECT 19.750 88.035 20.005 88.365 ;
        RECT 20.230 88.035 20.425 88.365 ;
        RECT 20.595 88.995 21.720 89.165 ;
        RECT 19.835 87.865 20.005 88.035 ;
        RECT 20.595 87.865 20.765 88.995 ;
        RECT 17.175 87.125 17.425 87.665 ;
        RECT 17.595 87.295 17.855 87.775 ;
        RECT 18.485 87.125 18.775 87.850 ;
        RECT 19.410 87.295 19.665 87.865 ;
        RECT 19.835 87.695 20.765 87.865 ;
        RECT 20.935 88.655 21.945 88.825 ;
        RECT 20.935 87.855 21.105 88.655 ;
        RECT 21.310 87.975 21.585 88.455 ;
        RECT 21.305 87.805 21.585 87.975 ;
        RECT 20.590 87.660 20.765 87.695 ;
        RECT 19.835 87.125 20.165 87.525 ;
        RECT 20.590 87.295 21.120 87.660 ;
        RECT 21.310 87.295 21.585 87.805 ;
        RECT 21.755 87.295 21.945 88.655 ;
        RECT 22.115 88.670 22.285 89.335 ;
        RECT 22.455 88.915 22.625 89.675 ;
        RECT 22.860 88.915 23.375 89.325 ;
        RECT 23.545 89.240 28.890 89.675 ;
        RECT 22.115 88.480 22.865 88.670 ;
        RECT 23.035 88.105 23.375 88.915 ;
        RECT 22.145 87.935 23.375 88.105 ;
        RECT 22.125 87.125 22.635 87.660 ;
        RECT 22.855 87.330 23.100 87.935 ;
        RECT 25.130 87.670 25.470 88.500 ;
        RECT 26.950 87.990 27.300 89.240 ;
        RECT 29.065 88.585 32.575 89.675 ;
        RECT 32.860 89.045 33.145 89.505 ;
        RECT 33.315 89.215 33.585 89.675 ;
        RECT 32.860 88.825 33.815 89.045 ;
        RECT 29.065 87.895 30.715 88.415 ;
        RECT 30.885 88.065 32.575 88.585 ;
        RECT 32.745 88.095 33.435 88.655 ;
        RECT 33.605 87.925 33.815 88.825 ;
        RECT 23.545 87.125 28.890 87.670 ;
        RECT 29.065 87.125 32.575 87.895 ;
        RECT 32.860 87.755 33.815 87.925 ;
        RECT 33.985 88.655 34.385 89.505 ;
        RECT 34.575 89.045 34.855 89.505 ;
        RECT 35.375 89.215 35.700 89.675 ;
        RECT 34.575 88.825 35.700 89.045 ;
        RECT 33.985 88.095 35.080 88.655 ;
        RECT 35.250 88.365 35.700 88.825 ;
        RECT 35.870 88.535 36.255 89.505 ;
        RECT 36.425 88.585 38.095 89.675 ;
        RECT 38.725 88.600 39.065 89.675 ;
        RECT 39.250 89.165 41.300 89.455 ;
        RECT 32.860 87.295 33.145 87.755 ;
        RECT 33.315 87.125 33.585 87.585 ;
        RECT 33.985 87.295 34.385 88.095 ;
        RECT 35.250 88.035 35.805 88.365 ;
        RECT 35.250 87.925 35.700 88.035 ;
        RECT 34.575 87.755 35.700 87.925 ;
        RECT 35.975 87.865 36.255 88.535 ;
        RECT 34.575 87.295 34.855 87.755 ;
        RECT 35.375 87.125 35.700 87.585 ;
        RECT 35.870 87.295 36.255 87.865 ;
        RECT 36.425 87.895 37.175 88.415 ;
        RECT 37.345 88.065 38.095 88.585 ;
        RECT 39.235 88.365 39.475 88.960 ;
        RECT 39.670 88.825 41.300 88.995 ;
        RECT 41.470 88.875 41.750 89.675 ;
        RECT 39.670 88.535 39.990 88.825 ;
        RECT 41.130 88.705 41.300 88.825 ;
        RECT 36.425 87.125 38.095 87.895 ;
        RECT 38.725 87.795 39.065 88.365 ;
        RECT 39.235 88.035 39.890 88.365 ;
        RECT 40.160 88.035 40.900 88.655 ;
        RECT 41.130 88.535 41.790 88.705 ;
        RECT 41.960 88.535 42.235 89.505 ;
        RECT 42.405 88.585 44.075 89.675 ;
        RECT 41.620 88.365 41.790 88.535 ;
        RECT 41.070 88.035 41.450 88.365 ;
        RECT 41.620 88.035 41.895 88.365 ;
        RECT 38.725 87.125 39.065 87.625 ;
        RECT 39.235 87.345 39.480 88.035 ;
        RECT 41.620 87.865 41.790 88.035 ;
        RECT 40.205 87.695 41.790 87.865 ;
        RECT 42.065 87.800 42.235 88.535 ;
        RECT 39.675 87.125 40.005 87.625 ;
        RECT 40.205 87.345 40.375 87.695 ;
        RECT 40.550 87.125 40.880 87.525 ;
        RECT 41.050 87.345 41.220 87.695 ;
        RECT 41.390 87.125 41.770 87.525 ;
        RECT 41.960 87.455 42.235 87.800 ;
        RECT 42.405 87.895 43.155 88.415 ;
        RECT 43.325 88.065 44.075 88.585 ;
        RECT 44.245 88.510 44.535 89.675 ;
        RECT 44.705 89.240 50.050 89.675 ;
        RECT 50.225 89.240 55.570 89.675 ;
        RECT 42.405 87.125 44.075 87.895 ;
        RECT 44.245 87.125 44.535 87.850 ;
        RECT 46.290 87.670 46.630 88.500 ;
        RECT 48.110 87.990 48.460 89.240 ;
        RECT 51.810 87.670 52.150 88.500 ;
        RECT 53.630 87.990 53.980 89.240 ;
        RECT 55.745 88.585 59.255 89.675 ;
        RECT 59.530 88.875 59.785 89.675 ;
        RECT 59.955 88.705 60.285 89.505 ;
        RECT 60.455 88.875 60.625 89.675 ;
        RECT 60.795 88.705 61.125 89.505 ;
        RECT 55.745 87.895 57.395 88.415 ;
        RECT 57.565 88.065 59.255 88.585 ;
        RECT 59.425 88.535 61.125 88.705 ;
        RECT 61.295 88.535 61.555 89.675 ;
        RECT 61.725 88.585 63.395 89.675 ;
        RECT 63.565 89.120 64.170 89.675 ;
        RECT 64.345 89.165 64.825 89.505 ;
        RECT 64.995 89.130 65.250 89.675 ;
        RECT 63.565 89.020 64.180 89.120 ;
        RECT 63.995 88.995 64.180 89.020 ;
        RECT 59.425 87.945 59.705 88.535 ;
        RECT 59.875 88.115 60.625 88.365 ;
        RECT 60.795 88.115 61.555 88.365 ;
        RECT 44.705 87.125 50.050 87.670 ;
        RECT 50.225 87.125 55.570 87.670 ;
        RECT 55.745 87.125 59.255 87.895 ;
        RECT 59.425 87.695 60.285 87.945 ;
        RECT 60.455 87.755 61.555 87.925 ;
        RECT 59.535 87.505 59.865 87.525 ;
        RECT 60.455 87.505 60.705 87.755 ;
        RECT 59.535 87.295 60.705 87.505 ;
        RECT 60.875 87.125 61.045 87.585 ;
        RECT 61.215 87.295 61.555 87.755 ;
        RECT 61.725 87.895 62.475 88.415 ;
        RECT 62.645 88.065 63.395 88.585 ;
        RECT 63.565 88.400 63.825 88.850 ;
        RECT 63.995 88.750 64.325 88.995 ;
        RECT 64.495 88.675 65.250 88.925 ;
        RECT 65.420 88.805 65.695 89.505 ;
        RECT 64.480 88.640 65.250 88.675 ;
        RECT 64.465 88.630 65.250 88.640 ;
        RECT 64.460 88.615 65.355 88.630 ;
        RECT 64.440 88.600 65.355 88.615 ;
        RECT 64.420 88.590 65.355 88.600 ;
        RECT 64.395 88.580 65.355 88.590 ;
        RECT 64.325 88.550 65.355 88.580 ;
        RECT 64.305 88.520 65.355 88.550 ;
        RECT 64.285 88.490 65.355 88.520 ;
        RECT 64.255 88.465 65.355 88.490 ;
        RECT 64.220 88.430 65.355 88.465 ;
        RECT 64.190 88.425 65.355 88.430 ;
        RECT 64.190 88.420 64.580 88.425 ;
        RECT 64.190 88.410 64.555 88.420 ;
        RECT 64.190 88.405 64.540 88.410 ;
        RECT 64.190 88.400 64.525 88.405 ;
        RECT 63.565 88.395 64.525 88.400 ;
        RECT 63.565 88.385 64.515 88.395 ;
        RECT 63.565 88.380 64.505 88.385 ;
        RECT 63.565 88.370 64.495 88.380 ;
        RECT 63.565 88.360 64.490 88.370 ;
        RECT 63.565 88.355 64.485 88.360 ;
        RECT 63.565 88.340 64.475 88.355 ;
        RECT 63.565 88.325 64.470 88.340 ;
        RECT 63.565 88.300 64.460 88.325 ;
        RECT 63.565 88.230 64.455 88.300 ;
        RECT 61.725 87.125 63.395 87.895 ;
        RECT 63.565 87.675 64.115 88.060 ;
        RECT 64.285 87.505 64.455 88.230 ;
        RECT 63.565 87.335 64.455 87.505 ;
        RECT 64.625 87.830 64.955 88.255 ;
        RECT 65.125 88.030 65.355 88.425 ;
        RECT 64.625 87.345 64.845 87.830 ;
        RECT 65.525 87.775 65.695 88.805 ;
        RECT 65.865 88.585 69.375 89.675 ;
        RECT 65.015 87.125 65.265 87.665 ;
        RECT 65.435 87.295 65.695 87.775 ;
        RECT 65.865 87.895 67.515 88.415 ;
        RECT 67.685 88.065 69.375 88.585 ;
        RECT 70.005 88.510 70.295 89.675 ;
        RECT 70.470 88.705 70.745 89.505 ;
        RECT 70.915 88.875 71.245 89.675 ;
        RECT 71.415 89.335 72.555 89.505 ;
        RECT 71.415 88.705 71.585 89.335 ;
        RECT 70.470 88.495 71.585 88.705 ;
        RECT 71.755 88.705 72.085 89.165 ;
        RECT 72.255 88.875 72.555 89.335 ;
        RECT 71.755 88.655 72.515 88.705 ;
        RECT 71.755 88.485 72.535 88.655 ;
        RECT 72.825 88.535 73.035 89.675 ;
        RECT 73.205 88.525 73.535 89.505 ;
        RECT 73.705 88.535 73.935 89.675 ;
        RECT 74.145 88.585 77.655 89.675 ;
        RECT 77.825 88.585 79.035 89.675 ;
        RECT 70.470 88.115 71.190 88.315 ;
        RECT 71.360 88.115 72.130 88.315 ;
        RECT 72.300 87.945 72.515 88.485 ;
        RECT 65.865 87.125 69.375 87.895 ;
        RECT 70.005 87.125 70.295 87.850 ;
        RECT 70.470 87.125 70.745 87.945 ;
        RECT 70.915 87.775 72.515 87.945 ;
        RECT 70.915 87.765 72.085 87.775 ;
        RECT 70.915 87.295 71.245 87.765 ;
        RECT 71.415 87.125 71.585 87.595 ;
        RECT 71.755 87.295 72.085 87.765 ;
        RECT 72.255 87.125 72.545 87.595 ;
        RECT 72.825 87.125 73.035 87.945 ;
        RECT 73.205 87.925 73.455 88.525 ;
        RECT 73.625 88.115 73.955 88.365 ;
        RECT 73.205 87.295 73.535 87.925 ;
        RECT 73.705 87.125 73.935 87.945 ;
        RECT 74.145 87.895 75.795 88.415 ;
        RECT 75.965 88.065 77.655 88.585 ;
        RECT 74.145 87.125 77.655 87.895 ;
        RECT 77.825 87.875 78.345 88.415 ;
        RECT 78.515 88.045 79.035 88.585 ;
        RECT 79.205 88.535 79.590 89.505 ;
        RECT 79.760 89.215 80.085 89.675 ;
        RECT 80.605 89.045 80.885 89.505 ;
        RECT 79.760 88.825 80.885 89.045 ;
        RECT 77.825 87.125 79.035 87.875 ;
        RECT 79.205 87.865 79.485 88.535 ;
        RECT 79.760 88.365 80.210 88.825 ;
        RECT 81.075 88.655 81.475 89.505 ;
        RECT 81.875 89.215 82.145 89.675 ;
        RECT 82.315 89.045 82.600 89.505 ;
        RECT 79.655 88.035 80.210 88.365 ;
        RECT 80.380 88.095 81.475 88.655 ;
        RECT 79.760 87.925 80.210 88.035 ;
        RECT 79.205 87.295 79.590 87.865 ;
        RECT 79.760 87.755 80.885 87.925 ;
        RECT 79.760 87.125 80.085 87.585 ;
        RECT 80.605 87.295 80.885 87.755 ;
        RECT 81.075 87.295 81.475 88.095 ;
        RECT 81.645 88.825 82.600 89.045 ;
        RECT 81.645 87.925 81.855 88.825 ;
        RECT 82.025 88.095 82.715 88.655 ;
        RECT 82.885 88.585 84.095 89.675 ;
        RECT 82.885 88.045 83.405 88.585 ;
        RECT 81.645 87.755 82.600 87.925 ;
        RECT 83.575 87.875 84.095 88.415 ;
        RECT 81.875 87.125 82.145 87.585 ;
        RECT 82.315 87.295 82.600 87.755 ;
        RECT 82.885 87.125 84.095 87.875 ;
        RECT 5.520 86.955 84.180 87.125 ;
        RECT 5.605 86.205 6.815 86.955 ;
        RECT 5.605 85.665 6.125 86.205 ;
        RECT 6.985 86.185 8.655 86.955 ;
        RECT 9.290 86.280 9.565 86.625 ;
        RECT 9.755 86.555 10.135 86.955 ;
        RECT 10.305 86.385 10.475 86.735 ;
        RECT 10.645 86.555 10.975 86.955 ;
        RECT 11.145 86.385 11.400 86.735 ;
        RECT 6.295 85.495 6.815 86.035 ;
        RECT 6.985 85.665 7.735 86.185 ;
        RECT 7.905 85.495 8.655 86.015 ;
        RECT 5.605 84.405 6.815 85.495 ;
        RECT 6.985 84.405 8.655 85.495 ;
        RECT 9.290 85.545 9.460 86.280 ;
        RECT 9.735 86.215 11.400 86.385 ;
        RECT 11.675 86.405 11.845 86.695 ;
        RECT 12.015 86.575 12.345 86.955 ;
        RECT 11.675 86.235 12.340 86.405 ;
        RECT 9.735 86.045 9.905 86.215 ;
        RECT 9.630 85.715 9.905 86.045 ;
        RECT 10.075 85.715 10.900 86.045 ;
        RECT 11.070 85.715 11.415 86.045 ;
        RECT 9.735 85.545 9.905 85.715 ;
        RECT 9.290 84.575 9.565 85.545 ;
        RECT 9.735 85.375 10.395 85.545 ;
        RECT 10.705 85.425 10.900 85.715 ;
        RECT 10.225 85.255 10.395 85.375 ;
        RECT 11.070 85.255 11.395 85.545 ;
        RECT 11.590 85.415 11.940 86.065 ;
        RECT 9.775 84.405 10.055 85.205 ;
        RECT 10.225 85.085 11.395 85.255 ;
        RECT 12.110 85.245 12.340 86.235 ;
        RECT 11.675 85.075 12.340 85.245 ;
        RECT 10.225 84.625 11.415 84.915 ;
        RECT 11.675 84.575 11.845 85.075 ;
        RECT 12.015 84.405 12.345 84.905 ;
        RECT 12.515 84.575 12.700 86.695 ;
        RECT 12.955 86.495 13.205 86.955 ;
        RECT 13.375 86.505 13.710 86.675 ;
        RECT 13.905 86.505 14.580 86.675 ;
        RECT 13.375 86.365 13.545 86.505 ;
        RECT 12.870 85.375 13.150 86.325 ;
        RECT 13.320 86.235 13.545 86.365 ;
        RECT 13.320 85.130 13.490 86.235 ;
        RECT 13.715 86.085 14.240 86.305 ;
        RECT 13.660 85.320 13.900 85.915 ;
        RECT 14.070 85.385 14.240 86.085 ;
        RECT 14.410 85.725 14.580 86.505 ;
        RECT 14.900 86.455 15.270 86.955 ;
        RECT 15.450 86.505 15.855 86.675 ;
        RECT 16.025 86.505 16.810 86.675 ;
        RECT 15.450 86.275 15.620 86.505 ;
        RECT 14.790 85.975 15.620 86.275 ;
        RECT 16.005 86.005 16.470 86.335 ;
        RECT 14.790 85.945 14.990 85.975 ;
        RECT 15.110 85.725 15.280 85.795 ;
        RECT 14.410 85.555 15.280 85.725 ;
        RECT 14.770 85.465 15.280 85.555 ;
        RECT 13.320 85.000 13.625 85.130 ;
        RECT 14.070 85.020 14.600 85.385 ;
        RECT 12.940 84.405 13.205 84.865 ;
        RECT 13.375 84.575 13.625 85.000 ;
        RECT 14.770 84.850 14.940 85.465 ;
        RECT 13.835 84.680 14.940 84.850 ;
        RECT 15.110 84.405 15.280 85.205 ;
        RECT 15.450 84.905 15.620 85.975 ;
        RECT 15.790 85.075 15.980 85.795 ;
        RECT 16.150 85.045 16.470 86.005 ;
        RECT 16.640 86.045 16.810 86.505 ;
        RECT 17.085 86.425 17.295 86.955 ;
        RECT 17.555 86.215 17.885 86.740 ;
        RECT 18.055 86.345 18.225 86.955 ;
        RECT 18.395 86.300 18.725 86.735 ;
        RECT 18.945 86.575 19.835 86.745 ;
        RECT 18.395 86.215 18.775 86.300 ;
        RECT 17.685 86.045 17.885 86.215 ;
        RECT 18.550 86.175 18.775 86.215 ;
        RECT 16.640 85.715 17.515 86.045 ;
        RECT 17.685 85.715 18.435 86.045 ;
        RECT 15.450 84.575 15.700 84.905 ;
        RECT 16.640 84.875 16.810 85.715 ;
        RECT 17.685 85.510 17.875 85.715 ;
        RECT 18.605 85.595 18.775 86.175 ;
        RECT 18.945 86.020 19.495 86.405 ;
        RECT 19.665 85.850 19.835 86.575 ;
        RECT 18.560 85.545 18.775 85.595 ;
        RECT 16.980 85.135 17.875 85.510 ;
        RECT 18.385 85.465 18.775 85.545 ;
        RECT 18.945 85.780 19.835 85.850 ;
        RECT 20.005 86.250 20.225 86.735 ;
        RECT 20.395 86.415 20.645 86.955 ;
        RECT 20.815 86.305 21.075 86.785 ;
        RECT 20.005 85.825 20.335 86.250 ;
        RECT 18.945 85.755 19.840 85.780 ;
        RECT 18.945 85.740 19.850 85.755 ;
        RECT 18.945 85.725 19.855 85.740 ;
        RECT 18.945 85.720 19.865 85.725 ;
        RECT 18.945 85.710 19.870 85.720 ;
        RECT 18.945 85.700 19.875 85.710 ;
        RECT 18.945 85.695 19.885 85.700 ;
        RECT 18.945 85.685 19.895 85.695 ;
        RECT 18.945 85.680 19.905 85.685 ;
        RECT 15.925 84.705 16.810 84.875 ;
        RECT 16.990 84.405 17.305 84.905 ;
        RECT 17.535 84.575 17.875 85.135 ;
        RECT 18.045 84.405 18.215 85.415 ;
        RECT 18.385 84.620 18.715 85.465 ;
        RECT 18.945 85.230 19.205 85.680 ;
        RECT 19.570 85.675 19.905 85.680 ;
        RECT 19.570 85.670 19.920 85.675 ;
        RECT 19.570 85.660 19.935 85.670 ;
        RECT 19.570 85.655 19.960 85.660 ;
        RECT 20.505 85.655 20.735 86.050 ;
        RECT 19.570 85.650 20.735 85.655 ;
        RECT 19.600 85.615 20.735 85.650 ;
        RECT 19.635 85.590 20.735 85.615 ;
        RECT 19.665 85.560 20.735 85.590 ;
        RECT 19.685 85.530 20.735 85.560 ;
        RECT 19.705 85.500 20.735 85.530 ;
        RECT 19.775 85.490 20.735 85.500 ;
        RECT 19.800 85.480 20.735 85.490 ;
        RECT 19.820 85.465 20.735 85.480 ;
        RECT 19.840 85.450 20.735 85.465 ;
        RECT 19.845 85.440 20.630 85.450 ;
        RECT 19.860 85.405 20.630 85.440 ;
        RECT 19.375 85.085 19.705 85.330 ;
        RECT 19.875 85.155 20.630 85.405 ;
        RECT 20.905 85.275 21.075 86.305 ;
        RECT 21.245 86.185 23.835 86.955 ;
        RECT 24.095 86.405 24.265 86.695 ;
        RECT 24.435 86.575 24.765 86.955 ;
        RECT 24.095 86.235 24.760 86.405 ;
        RECT 21.245 85.665 22.455 86.185 ;
        RECT 22.625 85.495 23.835 86.015 ;
        RECT 19.375 85.060 19.560 85.085 ;
        RECT 18.945 84.960 19.560 85.060 ;
        RECT 18.945 84.405 19.550 84.960 ;
        RECT 19.725 84.575 20.205 84.915 ;
        RECT 20.375 84.405 20.630 84.950 ;
        RECT 20.800 84.575 21.075 85.275 ;
        RECT 21.245 84.405 23.835 85.495 ;
        RECT 24.010 85.415 24.360 86.065 ;
        RECT 24.530 85.245 24.760 86.235 ;
        RECT 24.095 85.075 24.760 85.245 ;
        RECT 24.095 84.575 24.265 85.075 ;
        RECT 24.435 84.405 24.765 84.905 ;
        RECT 24.935 84.575 25.120 86.695 ;
        RECT 25.375 86.495 25.625 86.955 ;
        RECT 25.795 86.505 26.130 86.675 ;
        RECT 26.325 86.505 27.000 86.675 ;
        RECT 25.795 86.365 25.965 86.505 ;
        RECT 25.290 85.375 25.570 86.325 ;
        RECT 25.740 86.235 25.965 86.365 ;
        RECT 25.740 85.130 25.910 86.235 ;
        RECT 26.135 86.085 26.660 86.305 ;
        RECT 26.080 85.320 26.320 85.915 ;
        RECT 26.490 85.385 26.660 86.085 ;
        RECT 26.830 85.725 27.000 86.505 ;
        RECT 27.320 86.455 27.690 86.955 ;
        RECT 27.870 86.505 28.275 86.675 ;
        RECT 28.445 86.505 29.230 86.675 ;
        RECT 27.870 86.275 28.040 86.505 ;
        RECT 27.210 85.975 28.040 86.275 ;
        RECT 28.425 86.005 28.890 86.335 ;
        RECT 27.210 85.945 27.410 85.975 ;
        RECT 27.530 85.725 27.700 85.795 ;
        RECT 26.830 85.555 27.700 85.725 ;
        RECT 27.190 85.465 27.700 85.555 ;
        RECT 25.740 85.000 26.045 85.130 ;
        RECT 26.490 85.020 27.020 85.385 ;
        RECT 25.360 84.405 25.625 84.865 ;
        RECT 25.795 84.575 26.045 85.000 ;
        RECT 27.190 84.850 27.360 85.465 ;
        RECT 26.255 84.680 27.360 84.850 ;
        RECT 27.530 84.405 27.700 85.205 ;
        RECT 27.870 84.905 28.040 85.975 ;
        RECT 28.210 85.075 28.400 85.795 ;
        RECT 28.570 85.045 28.890 86.005 ;
        RECT 29.060 86.045 29.230 86.505 ;
        RECT 29.505 86.425 29.715 86.955 ;
        RECT 29.975 86.215 30.305 86.740 ;
        RECT 30.475 86.345 30.645 86.955 ;
        RECT 30.815 86.300 31.145 86.735 ;
        RECT 30.815 86.215 31.195 86.300 ;
        RECT 31.365 86.230 31.655 86.955 ;
        RECT 30.105 86.045 30.305 86.215 ;
        RECT 30.970 86.175 31.195 86.215 ;
        RECT 29.060 85.715 29.935 86.045 ;
        RECT 30.105 85.715 30.855 86.045 ;
        RECT 27.870 84.575 28.120 84.905 ;
        RECT 29.060 84.875 29.230 85.715 ;
        RECT 30.105 85.510 30.295 85.715 ;
        RECT 31.025 85.595 31.195 86.175 ;
        RECT 30.980 85.545 31.195 85.595 ;
        RECT 31.830 86.215 32.085 86.785 ;
        RECT 32.255 86.555 32.585 86.955 ;
        RECT 33.010 86.420 33.540 86.785 ;
        RECT 33.730 86.615 34.005 86.785 ;
        RECT 33.725 86.445 34.005 86.615 ;
        RECT 33.010 86.385 33.185 86.420 ;
        RECT 32.255 86.215 33.185 86.385 ;
        RECT 29.400 85.135 30.295 85.510 ;
        RECT 30.805 85.465 31.195 85.545 ;
        RECT 28.345 84.705 29.230 84.875 ;
        RECT 29.410 84.405 29.725 84.905 ;
        RECT 29.955 84.575 30.295 85.135 ;
        RECT 30.465 84.405 30.635 85.415 ;
        RECT 30.805 84.620 31.135 85.465 ;
        RECT 31.365 84.405 31.655 85.570 ;
        RECT 31.830 85.545 32.000 86.215 ;
        RECT 32.255 86.045 32.425 86.215 ;
        RECT 32.170 85.715 32.425 86.045 ;
        RECT 32.650 85.715 32.845 86.045 ;
        RECT 31.830 84.575 32.165 85.545 ;
        RECT 32.335 84.405 32.505 85.545 ;
        RECT 32.675 84.745 32.845 85.715 ;
        RECT 33.015 85.085 33.185 86.215 ;
        RECT 33.355 85.425 33.525 86.225 ;
        RECT 33.730 85.625 34.005 86.445 ;
        RECT 34.175 85.425 34.365 86.785 ;
        RECT 34.545 86.420 35.055 86.955 ;
        RECT 35.275 86.145 35.520 86.750 ;
        RECT 35.965 86.185 37.635 86.955 ;
        RECT 34.565 85.975 35.795 86.145 ;
        RECT 33.355 85.255 34.365 85.425 ;
        RECT 34.535 85.410 35.285 85.600 ;
        RECT 33.015 84.915 34.140 85.085 ;
        RECT 34.535 84.745 34.705 85.410 ;
        RECT 35.455 85.165 35.795 85.975 ;
        RECT 35.965 85.665 36.715 86.185 ;
        RECT 37.805 86.155 38.145 86.785 ;
        RECT 38.315 86.155 38.565 86.955 ;
        RECT 38.755 86.305 39.085 86.785 ;
        RECT 39.255 86.495 39.480 86.955 ;
        RECT 39.650 86.305 39.980 86.785 ;
        RECT 36.885 85.495 37.635 86.015 ;
        RECT 32.675 84.575 34.705 84.745 ;
        RECT 34.875 84.405 35.045 85.165 ;
        RECT 35.280 84.755 35.795 85.165 ;
        RECT 35.965 84.405 37.635 85.495 ;
        RECT 37.805 85.545 37.980 86.155 ;
        RECT 38.755 86.135 39.980 86.305 ;
        RECT 40.610 86.175 41.110 86.785 ;
        RECT 41.485 86.305 41.745 86.785 ;
        RECT 41.915 86.495 42.245 86.955 ;
        RECT 42.435 86.315 42.635 86.735 ;
        RECT 38.150 85.795 38.845 85.965 ;
        RECT 38.675 85.545 38.845 85.795 ;
        RECT 39.020 85.765 39.440 85.965 ;
        RECT 39.610 85.765 39.940 85.965 ;
        RECT 40.110 85.765 40.440 85.965 ;
        RECT 40.610 85.545 40.780 86.175 ;
        RECT 40.965 85.715 41.315 85.965 ;
        RECT 37.805 84.575 38.145 85.545 ;
        RECT 38.315 84.405 38.485 85.545 ;
        RECT 38.675 85.375 41.110 85.545 ;
        RECT 38.755 84.405 39.005 85.205 ;
        RECT 39.650 84.575 39.980 85.375 ;
        RECT 40.280 84.405 40.610 85.205 ;
        RECT 40.780 84.575 41.110 85.375 ;
        RECT 41.485 85.275 41.655 86.305 ;
        RECT 41.825 85.615 42.055 86.045 ;
        RECT 42.225 85.795 42.635 86.315 ;
        RECT 42.805 86.470 43.595 86.735 ;
        RECT 42.805 85.615 43.060 86.470 ;
        RECT 43.775 86.135 44.105 86.555 ;
        RECT 44.275 86.135 44.535 86.955 ;
        RECT 44.725 86.265 44.965 86.785 ;
        RECT 45.135 86.460 45.530 86.955 ;
        RECT 46.095 86.625 46.265 86.770 ;
        RECT 45.890 86.430 46.265 86.625 ;
        RECT 43.775 86.045 44.025 86.135 ;
        RECT 43.230 85.795 44.025 86.045 ;
        RECT 41.825 85.445 43.615 85.615 ;
        RECT 41.485 84.575 41.760 85.275 ;
        RECT 41.930 85.150 42.645 85.445 ;
        RECT 42.865 85.085 43.195 85.275 ;
        RECT 41.970 84.405 42.185 84.950 ;
        RECT 42.355 84.575 42.830 84.915 ;
        RECT 43.000 84.910 43.195 85.085 ;
        RECT 43.365 85.080 43.615 85.445 ;
        RECT 43.000 84.405 43.615 84.910 ;
        RECT 43.855 84.575 44.025 85.795 ;
        RECT 44.195 85.085 44.535 85.965 ;
        RECT 44.725 85.460 44.900 86.265 ;
        RECT 45.890 86.095 46.060 86.430 ;
        RECT 46.545 86.385 46.785 86.760 ;
        RECT 46.955 86.450 47.290 86.955 ;
        RECT 46.545 86.235 46.765 86.385 ;
        RECT 45.075 85.735 46.060 86.095 ;
        RECT 46.230 85.905 46.765 86.235 ;
        RECT 45.075 85.715 46.360 85.735 ;
        RECT 45.500 85.565 46.360 85.715 ;
        RECT 44.275 84.405 44.535 84.915 ;
        RECT 44.725 84.675 45.030 85.460 ;
        RECT 45.205 85.085 45.900 85.395 ;
        RECT 45.210 84.405 45.895 84.875 ;
        RECT 46.075 84.620 46.360 85.565 ;
        RECT 46.530 85.255 46.765 85.905 ;
        RECT 46.935 85.425 47.235 86.275 ;
        RECT 47.465 86.185 49.135 86.955 ;
        RECT 49.395 86.405 49.565 86.695 ;
        RECT 49.735 86.575 50.065 86.955 ;
        RECT 49.395 86.235 50.060 86.405 ;
        RECT 47.465 85.665 48.215 86.185 ;
        RECT 48.385 85.495 49.135 86.015 ;
        RECT 46.530 85.025 47.205 85.255 ;
        RECT 46.535 84.405 46.865 84.855 ;
        RECT 47.035 84.595 47.205 85.025 ;
        RECT 47.465 84.405 49.135 85.495 ;
        RECT 49.310 85.415 49.660 86.065 ;
        RECT 49.830 85.245 50.060 86.235 ;
        RECT 49.395 85.075 50.060 85.245 ;
        RECT 49.395 84.575 49.565 85.075 ;
        RECT 49.735 84.405 50.065 84.905 ;
        RECT 50.235 84.575 50.420 86.695 ;
        RECT 50.675 86.495 50.925 86.955 ;
        RECT 51.095 86.505 51.430 86.675 ;
        RECT 51.625 86.505 52.300 86.675 ;
        RECT 51.095 86.365 51.265 86.505 ;
        RECT 50.590 85.375 50.870 86.325 ;
        RECT 51.040 86.235 51.265 86.365 ;
        RECT 51.040 85.130 51.210 86.235 ;
        RECT 51.435 86.085 51.960 86.305 ;
        RECT 51.380 85.320 51.620 85.915 ;
        RECT 51.790 85.385 51.960 86.085 ;
        RECT 52.130 85.725 52.300 86.505 ;
        RECT 52.620 86.455 52.990 86.955 ;
        RECT 53.170 86.505 53.575 86.675 ;
        RECT 53.745 86.505 54.530 86.675 ;
        RECT 53.170 86.275 53.340 86.505 ;
        RECT 52.510 85.975 53.340 86.275 ;
        RECT 53.725 86.005 54.190 86.335 ;
        RECT 52.510 85.945 52.710 85.975 ;
        RECT 52.830 85.725 53.000 85.795 ;
        RECT 52.130 85.555 53.000 85.725 ;
        RECT 52.490 85.465 53.000 85.555 ;
        RECT 51.040 85.000 51.345 85.130 ;
        RECT 51.790 85.020 52.320 85.385 ;
        RECT 50.660 84.405 50.925 84.865 ;
        RECT 51.095 84.575 51.345 85.000 ;
        RECT 52.490 84.850 52.660 85.465 ;
        RECT 51.555 84.680 52.660 84.850 ;
        RECT 52.830 84.405 53.000 85.205 ;
        RECT 53.170 84.905 53.340 85.975 ;
        RECT 53.510 85.075 53.700 85.795 ;
        RECT 53.870 85.045 54.190 86.005 ;
        RECT 54.360 86.045 54.530 86.505 ;
        RECT 54.805 86.425 55.015 86.955 ;
        RECT 55.275 86.215 55.605 86.740 ;
        RECT 55.775 86.345 55.945 86.955 ;
        RECT 56.115 86.300 56.445 86.735 ;
        RECT 56.115 86.215 56.495 86.300 ;
        RECT 57.125 86.230 57.415 86.955 ;
        RECT 57.590 86.480 57.925 86.740 ;
        RECT 58.095 86.555 58.425 86.955 ;
        RECT 58.595 86.555 60.210 86.725 ;
        RECT 55.405 86.045 55.605 86.215 ;
        RECT 56.270 86.175 56.495 86.215 ;
        RECT 54.360 85.715 55.235 86.045 ;
        RECT 55.405 85.715 56.155 86.045 ;
        RECT 53.170 84.575 53.420 84.905 ;
        RECT 54.360 84.875 54.530 85.715 ;
        RECT 55.405 85.510 55.595 85.715 ;
        RECT 56.325 85.595 56.495 86.175 ;
        RECT 56.280 85.545 56.495 85.595 ;
        RECT 54.700 85.135 55.595 85.510 ;
        RECT 56.105 85.465 56.495 85.545 ;
        RECT 53.645 84.705 54.530 84.875 ;
        RECT 54.710 84.405 55.025 84.905 ;
        RECT 55.255 84.575 55.595 85.135 ;
        RECT 55.765 84.405 55.935 85.415 ;
        RECT 56.105 84.620 56.435 85.465 ;
        RECT 57.125 84.405 57.415 85.570 ;
        RECT 57.590 85.125 57.845 86.480 ;
        RECT 58.595 86.385 58.765 86.555 ;
        RECT 58.205 86.215 58.765 86.385 ;
        RECT 58.205 86.045 58.375 86.215 ;
        RECT 58.070 85.715 58.375 86.045 ;
        RECT 58.570 85.935 58.820 86.045 ;
        RECT 59.030 85.935 59.300 86.375 ;
        RECT 59.490 86.275 59.780 86.375 ;
        RECT 59.485 86.105 59.780 86.275 ;
        RECT 58.565 85.765 58.820 85.935 ;
        RECT 59.025 85.765 59.300 85.935 ;
        RECT 58.570 85.715 58.820 85.765 ;
        RECT 59.030 85.715 59.300 85.765 ;
        RECT 59.490 85.715 59.780 86.105 ;
        RECT 59.950 85.715 60.370 86.380 ;
        RECT 60.755 86.235 61.085 86.955 ;
        RECT 62.190 86.450 62.525 86.955 ;
        RECT 62.695 86.385 62.935 86.760 ;
        RECT 63.215 86.625 63.385 86.770 ;
        RECT 63.215 86.430 63.590 86.625 ;
        RECT 63.950 86.460 64.345 86.955 ;
        RECT 60.680 85.935 61.030 86.045 ;
        RECT 60.680 85.765 61.035 85.935 ;
        RECT 60.680 85.715 61.030 85.765 ;
        RECT 58.205 85.545 58.375 85.715 ;
        RECT 58.205 85.375 60.575 85.545 ;
        RECT 60.825 85.425 61.030 85.715 ;
        RECT 62.245 85.425 62.545 86.275 ;
        RECT 62.715 86.235 62.935 86.385 ;
        RECT 62.715 85.905 63.250 86.235 ;
        RECT 63.420 86.095 63.590 86.430 ;
        RECT 64.515 86.265 64.755 86.785 ;
        RECT 57.590 84.615 57.925 85.125 ;
        RECT 58.175 84.405 58.505 85.205 ;
        RECT 58.750 84.995 60.175 85.165 ;
        RECT 58.750 84.575 59.035 84.995 ;
        RECT 59.290 84.405 59.620 84.825 ;
        RECT 59.845 84.745 60.175 84.995 ;
        RECT 60.405 84.915 60.575 85.375 ;
        RECT 62.715 85.255 62.950 85.905 ;
        RECT 63.420 85.735 64.405 86.095 ;
        RECT 60.835 84.745 61.005 85.245 ;
        RECT 59.845 84.575 61.005 84.745 ;
        RECT 62.275 85.025 62.950 85.255 ;
        RECT 63.120 85.715 64.405 85.735 ;
        RECT 63.120 85.565 63.980 85.715 ;
        RECT 62.275 84.595 62.445 85.025 ;
        RECT 62.615 84.405 62.945 84.855 ;
        RECT 63.120 84.620 63.405 85.565 ;
        RECT 64.580 85.460 64.755 86.265 ;
        RECT 64.950 86.425 65.240 86.775 ;
        RECT 65.435 86.595 65.765 86.955 ;
        RECT 65.935 86.425 66.165 86.730 ;
        RECT 64.950 86.255 66.165 86.425 ;
        RECT 66.355 86.615 66.525 86.650 ;
        RECT 66.355 86.445 66.555 86.615 ;
        RECT 66.355 86.085 66.525 86.445 ;
        RECT 65.010 85.935 65.270 86.045 ;
        RECT 65.005 85.765 65.270 85.935 ;
        RECT 65.010 85.715 65.270 85.765 ;
        RECT 65.450 85.715 65.835 86.045 ;
        RECT 66.005 85.915 66.525 86.085 ;
        RECT 66.785 86.185 69.375 86.955 ;
        RECT 70.010 86.190 70.465 86.955 ;
        RECT 70.740 86.575 72.040 86.785 ;
        RECT 72.295 86.595 72.625 86.955 ;
        RECT 71.870 86.425 72.040 86.575 ;
        RECT 72.795 86.455 73.055 86.785 ;
        RECT 63.580 85.085 64.275 85.395 ;
        RECT 63.585 84.405 64.270 84.875 ;
        RECT 64.450 84.675 64.755 85.460 ;
        RECT 64.950 84.405 65.270 85.545 ;
        RECT 65.450 84.665 65.645 85.715 ;
        RECT 66.005 85.535 66.175 85.915 ;
        RECT 65.825 85.255 66.175 85.535 ;
        RECT 66.365 85.385 66.610 85.745 ;
        RECT 66.785 85.665 67.995 86.185 ;
        RECT 68.165 85.495 69.375 86.015 ;
        RECT 70.940 85.965 71.160 86.365 ;
        RECT 70.005 85.765 70.495 85.965 ;
        RECT 70.685 85.755 71.160 85.965 ;
        RECT 71.405 85.965 71.615 86.365 ;
        RECT 71.870 86.300 72.625 86.425 ;
        RECT 71.870 86.255 72.715 86.300 ;
        RECT 72.445 86.135 72.715 86.255 ;
        RECT 71.405 85.755 71.735 85.965 ;
        RECT 71.905 85.695 72.315 86.000 ;
        RECT 65.825 84.575 66.155 85.255 ;
        RECT 66.355 84.405 66.610 85.205 ;
        RECT 66.785 84.405 69.375 85.495 ;
        RECT 70.010 85.525 71.185 85.585 ;
        RECT 72.545 85.560 72.715 86.135 ;
        RECT 72.515 85.525 72.715 85.560 ;
        RECT 70.010 85.415 72.715 85.525 ;
        RECT 70.010 84.795 70.265 85.415 ;
        RECT 70.855 85.355 72.655 85.415 ;
        RECT 70.855 85.325 71.185 85.355 ;
        RECT 72.885 85.255 73.055 86.455 ;
        RECT 73.775 86.405 73.945 86.695 ;
        RECT 74.115 86.575 74.445 86.955 ;
        RECT 73.775 86.235 74.440 86.405 ;
        RECT 73.690 85.415 74.040 86.065 ;
        RECT 70.515 85.155 70.700 85.245 ;
        RECT 71.290 85.155 72.125 85.165 ;
        RECT 70.515 84.955 72.125 85.155 ;
        RECT 70.515 84.915 70.745 84.955 ;
        RECT 70.010 84.575 70.345 84.795 ;
        RECT 71.350 84.405 71.705 84.785 ;
        RECT 71.875 84.575 72.125 84.955 ;
        RECT 72.375 84.405 72.625 85.185 ;
        RECT 72.795 84.575 73.055 85.255 ;
        RECT 74.210 85.245 74.440 86.235 ;
        RECT 73.775 85.075 74.440 85.245 ;
        RECT 73.775 84.575 73.945 85.075 ;
        RECT 74.115 84.405 74.445 84.905 ;
        RECT 74.615 84.575 74.800 86.695 ;
        RECT 75.055 86.495 75.305 86.955 ;
        RECT 75.475 86.505 75.810 86.675 ;
        RECT 76.005 86.505 76.680 86.675 ;
        RECT 75.475 86.365 75.645 86.505 ;
        RECT 74.970 85.375 75.250 86.325 ;
        RECT 75.420 86.235 75.645 86.365 ;
        RECT 75.420 85.130 75.590 86.235 ;
        RECT 75.815 86.085 76.340 86.305 ;
        RECT 75.760 85.320 76.000 85.915 ;
        RECT 76.170 85.385 76.340 86.085 ;
        RECT 76.510 85.725 76.680 86.505 ;
        RECT 77.000 86.455 77.370 86.955 ;
        RECT 77.550 86.505 77.955 86.675 ;
        RECT 78.125 86.505 78.910 86.675 ;
        RECT 77.550 86.275 77.720 86.505 ;
        RECT 76.890 85.975 77.720 86.275 ;
        RECT 78.105 86.005 78.570 86.335 ;
        RECT 76.890 85.945 77.090 85.975 ;
        RECT 77.210 85.725 77.380 85.795 ;
        RECT 76.510 85.555 77.380 85.725 ;
        RECT 76.870 85.465 77.380 85.555 ;
        RECT 75.420 85.000 75.725 85.130 ;
        RECT 76.170 85.020 76.700 85.385 ;
        RECT 75.040 84.405 75.305 84.865 ;
        RECT 75.475 84.575 75.725 85.000 ;
        RECT 76.870 84.850 77.040 85.465 ;
        RECT 75.935 84.680 77.040 84.850 ;
        RECT 77.210 84.405 77.380 85.205 ;
        RECT 77.550 84.905 77.720 85.975 ;
        RECT 77.890 85.075 78.080 85.795 ;
        RECT 78.250 85.045 78.570 86.005 ;
        RECT 78.740 86.045 78.910 86.505 ;
        RECT 79.185 86.425 79.395 86.955 ;
        RECT 79.655 86.215 79.985 86.740 ;
        RECT 80.155 86.345 80.325 86.955 ;
        RECT 80.495 86.300 80.825 86.735 ;
        RECT 81.135 86.405 81.305 86.785 ;
        RECT 81.520 86.575 81.850 86.955 ;
        RECT 80.495 86.215 80.875 86.300 ;
        RECT 81.135 86.235 81.850 86.405 ;
        RECT 79.785 86.045 79.985 86.215 ;
        RECT 80.650 86.175 80.875 86.215 ;
        RECT 78.740 85.715 79.615 86.045 ;
        RECT 79.785 85.715 80.535 86.045 ;
        RECT 77.550 84.575 77.800 84.905 ;
        RECT 78.740 84.875 78.910 85.715 ;
        RECT 79.785 85.510 79.975 85.715 ;
        RECT 80.705 85.595 80.875 86.175 ;
        RECT 81.045 85.685 81.400 86.055 ;
        RECT 81.680 86.045 81.850 86.235 ;
        RECT 82.020 86.210 82.275 86.785 ;
        RECT 81.680 85.715 81.935 86.045 ;
        RECT 80.660 85.545 80.875 85.595 ;
        RECT 79.080 85.135 79.975 85.510 ;
        RECT 80.485 85.465 80.875 85.545 ;
        RECT 81.680 85.505 81.850 85.715 ;
        RECT 78.025 84.705 78.910 84.875 ;
        RECT 79.090 84.405 79.405 84.905 ;
        RECT 79.635 84.575 79.975 85.135 ;
        RECT 80.145 84.405 80.315 85.415 ;
        RECT 80.485 84.620 80.815 85.465 ;
        RECT 81.135 85.335 81.850 85.505 ;
        RECT 82.105 85.480 82.275 86.210 ;
        RECT 82.450 86.115 82.710 86.955 ;
        RECT 82.885 86.205 84.095 86.955 ;
        RECT 81.135 84.575 81.305 85.335 ;
        RECT 81.520 84.405 81.850 85.165 ;
        RECT 82.020 84.575 82.275 85.480 ;
        RECT 82.450 84.405 82.710 85.555 ;
        RECT 82.885 85.495 83.405 86.035 ;
        RECT 83.575 85.665 84.095 86.205 ;
        RECT 82.885 84.405 84.095 85.495 ;
        RECT 5.520 84.235 84.180 84.405 ;
        RECT 5.605 83.145 6.815 84.235 ;
        RECT 6.985 83.145 10.495 84.235 ;
        RECT 10.665 83.145 11.875 84.235 ;
        RECT 5.605 82.435 6.125 82.975 ;
        RECT 6.295 82.605 6.815 83.145 ;
        RECT 6.985 82.455 8.635 82.975 ;
        RECT 8.805 82.625 10.495 83.145 ;
        RECT 5.605 81.685 6.815 82.435 ;
        RECT 6.985 81.685 10.495 82.455 ;
        RECT 10.665 82.435 11.185 82.975 ;
        RECT 11.355 82.605 11.875 83.145 ;
        RECT 12.230 83.265 12.620 83.440 ;
        RECT 13.105 83.435 13.435 84.235 ;
        RECT 13.605 83.445 14.140 84.065 ;
        RECT 12.230 83.095 13.655 83.265 ;
        RECT 10.665 81.685 11.875 82.435 ;
        RECT 12.105 82.365 12.460 82.925 ;
        RECT 12.630 82.195 12.800 83.095 ;
        RECT 12.970 82.365 13.235 82.925 ;
        RECT 13.485 82.595 13.655 83.095 ;
        RECT 13.825 82.425 14.140 83.445 ;
        RECT 12.210 81.685 12.450 82.195 ;
        RECT 12.630 81.865 12.910 82.195 ;
        RECT 13.140 81.685 13.355 82.195 ;
        RECT 13.525 81.855 14.140 82.425 ;
        RECT 14.345 83.515 14.805 84.065 ;
        RECT 14.995 83.515 15.325 84.235 ;
        RECT 14.345 82.145 14.595 83.515 ;
        RECT 15.525 83.345 15.825 83.895 ;
        RECT 15.995 83.565 16.275 84.235 ;
        RECT 14.885 83.175 15.825 83.345 ;
        RECT 14.885 82.925 15.055 83.175 ;
        RECT 16.195 82.925 16.460 83.285 ;
        RECT 17.145 83.095 17.375 84.235 ;
        RECT 17.545 83.085 17.875 84.065 ;
        RECT 18.045 83.095 18.255 84.235 ;
        RECT 14.765 82.595 15.055 82.925 ;
        RECT 15.225 82.675 15.565 82.925 ;
        RECT 15.785 82.675 16.460 82.925 ;
        RECT 17.125 82.675 17.455 82.925 ;
        RECT 14.885 82.505 15.055 82.595 ;
        RECT 14.885 82.315 16.275 82.505 ;
        RECT 14.345 81.855 14.905 82.145 ;
        RECT 15.075 81.685 15.325 82.145 ;
        RECT 15.945 81.955 16.275 82.315 ;
        RECT 17.145 81.685 17.375 82.505 ;
        RECT 17.625 82.485 17.875 83.085 ;
        RECT 18.485 83.070 18.775 84.235 ;
        RECT 19.955 83.565 20.125 84.065 ;
        RECT 20.295 83.735 20.625 84.235 ;
        RECT 19.955 83.395 20.620 83.565 ;
        RECT 19.870 82.575 20.220 83.225 ;
        RECT 17.545 81.855 17.875 82.485 ;
        RECT 18.045 81.685 18.255 82.505 ;
        RECT 18.485 81.685 18.775 82.410 ;
        RECT 20.390 82.405 20.620 83.395 ;
        RECT 19.955 82.235 20.620 82.405 ;
        RECT 19.955 81.945 20.125 82.235 ;
        RECT 20.295 81.685 20.625 82.065 ;
        RECT 20.795 81.945 20.980 84.065 ;
        RECT 21.220 83.775 21.485 84.235 ;
        RECT 21.655 83.640 21.905 84.065 ;
        RECT 22.115 83.790 23.220 83.960 ;
        RECT 21.600 83.510 21.905 83.640 ;
        RECT 21.150 82.315 21.430 83.265 ;
        RECT 21.600 82.405 21.770 83.510 ;
        RECT 21.940 82.725 22.180 83.320 ;
        RECT 22.350 83.255 22.880 83.620 ;
        RECT 22.350 82.555 22.520 83.255 ;
        RECT 23.050 83.175 23.220 83.790 ;
        RECT 23.390 83.435 23.560 84.235 ;
        RECT 23.730 83.735 23.980 84.065 ;
        RECT 24.205 83.765 25.090 83.935 ;
        RECT 23.050 83.085 23.560 83.175 ;
        RECT 21.600 82.275 21.825 82.405 ;
        RECT 21.995 82.335 22.520 82.555 ;
        RECT 22.690 82.915 23.560 83.085 ;
        RECT 21.235 81.685 21.485 82.145 ;
        RECT 21.655 82.135 21.825 82.275 ;
        RECT 22.690 82.135 22.860 82.915 ;
        RECT 23.390 82.845 23.560 82.915 ;
        RECT 23.070 82.665 23.270 82.695 ;
        RECT 23.730 82.665 23.900 83.735 ;
        RECT 24.070 82.845 24.260 83.565 ;
        RECT 23.070 82.365 23.900 82.665 ;
        RECT 24.430 82.635 24.750 83.595 ;
        RECT 21.655 81.965 21.990 82.135 ;
        RECT 22.185 81.965 22.860 82.135 ;
        RECT 23.180 81.685 23.550 82.185 ;
        RECT 23.730 82.135 23.900 82.365 ;
        RECT 24.285 82.305 24.750 82.635 ;
        RECT 24.920 82.925 25.090 83.765 ;
        RECT 25.270 83.735 25.585 84.235 ;
        RECT 25.815 83.505 26.155 84.065 ;
        RECT 25.260 83.130 26.155 83.505 ;
        RECT 26.325 83.225 26.495 84.235 ;
        RECT 25.965 82.925 26.155 83.130 ;
        RECT 26.665 83.175 26.995 84.020 ;
        RECT 27.165 83.320 27.335 84.235 ;
        RECT 26.665 83.095 27.055 83.175 ;
        RECT 27.685 83.145 31.195 84.235 ;
        RECT 26.840 83.045 27.055 83.095 ;
        RECT 24.920 82.595 25.795 82.925 ;
        RECT 25.965 82.595 26.715 82.925 ;
        RECT 24.920 82.135 25.090 82.595 ;
        RECT 25.965 82.425 26.165 82.595 ;
        RECT 26.885 82.465 27.055 83.045 ;
        RECT 26.830 82.425 27.055 82.465 ;
        RECT 23.730 81.965 24.135 82.135 ;
        RECT 24.305 81.965 25.090 82.135 ;
        RECT 25.365 81.685 25.575 82.215 ;
        RECT 25.835 81.900 26.165 82.425 ;
        RECT 26.675 82.340 27.055 82.425 ;
        RECT 27.685 82.455 29.335 82.975 ;
        RECT 29.505 82.625 31.195 83.145 ;
        RECT 32.285 83.095 32.670 84.065 ;
        RECT 32.840 83.775 33.165 84.235 ;
        RECT 33.685 83.605 33.965 84.065 ;
        RECT 32.840 83.385 33.965 83.605 ;
        RECT 26.335 81.685 26.505 82.295 ;
        RECT 26.675 81.905 27.005 82.340 ;
        RECT 27.175 81.685 27.345 82.200 ;
        RECT 27.685 81.685 31.195 82.455 ;
        RECT 32.285 82.425 32.565 83.095 ;
        RECT 32.840 82.925 33.290 83.385 ;
        RECT 34.155 83.215 34.555 84.065 ;
        RECT 34.955 83.775 35.225 84.235 ;
        RECT 35.395 83.605 35.680 84.065 ;
        RECT 35.965 83.725 36.225 84.235 ;
        RECT 32.735 82.595 33.290 82.925 ;
        RECT 33.460 82.655 34.555 83.215 ;
        RECT 32.840 82.485 33.290 82.595 ;
        RECT 32.285 81.855 32.670 82.425 ;
        RECT 32.840 82.315 33.965 82.485 ;
        RECT 32.840 81.685 33.165 82.145 ;
        RECT 33.685 81.855 33.965 82.315 ;
        RECT 34.155 81.855 34.555 82.655 ;
        RECT 34.725 83.385 35.680 83.605 ;
        RECT 34.725 82.485 34.935 83.385 ;
        RECT 35.105 82.655 35.795 83.215 ;
        RECT 35.965 82.675 36.305 83.555 ;
        RECT 36.475 82.845 36.645 84.065 ;
        RECT 36.885 83.730 37.500 84.235 ;
        RECT 36.885 83.195 37.135 83.560 ;
        RECT 37.305 83.555 37.500 83.730 ;
        RECT 37.670 83.725 38.145 84.065 ;
        RECT 38.315 83.690 38.530 84.235 ;
        RECT 37.305 83.365 37.635 83.555 ;
        RECT 37.855 83.195 38.570 83.490 ;
        RECT 38.740 83.365 39.015 84.065 ;
        RECT 36.885 83.025 38.675 83.195 ;
        RECT 36.475 82.595 37.270 82.845 ;
        RECT 36.475 82.505 36.725 82.595 ;
        RECT 34.725 82.315 35.680 82.485 ;
        RECT 34.955 81.685 35.225 82.145 ;
        RECT 35.395 81.855 35.680 82.315 ;
        RECT 35.965 81.685 36.225 82.505 ;
        RECT 36.395 82.085 36.725 82.505 ;
        RECT 37.440 82.170 37.695 83.025 ;
        RECT 36.905 81.905 37.695 82.170 ;
        RECT 37.865 82.325 38.275 82.845 ;
        RECT 38.445 82.595 38.675 83.025 ;
        RECT 38.845 82.335 39.015 83.365 ;
        RECT 37.865 81.905 38.065 82.325 ;
        RECT 38.255 81.685 38.585 82.145 ;
        RECT 38.755 81.855 39.015 82.335 ;
        RECT 40.125 83.180 40.430 83.965 ;
        RECT 40.610 83.765 41.295 84.235 ;
        RECT 40.605 83.245 41.300 83.555 ;
        RECT 40.125 82.375 40.300 83.180 ;
        RECT 41.475 83.075 41.760 84.020 ;
        RECT 41.935 83.785 42.265 84.235 ;
        RECT 42.435 83.615 42.605 84.045 ;
        RECT 40.900 82.925 41.760 83.075 ;
        RECT 40.475 82.905 41.760 82.925 ;
        RECT 41.930 83.385 42.605 83.615 ;
        RECT 40.475 82.545 41.460 82.905 ;
        RECT 41.930 82.735 42.165 83.385 ;
        RECT 40.125 81.855 40.365 82.375 ;
        RECT 41.290 82.210 41.460 82.545 ;
        RECT 41.630 82.405 42.165 82.735 ;
        RECT 41.945 82.255 42.165 82.405 ;
        RECT 42.335 82.365 42.635 83.215 ;
        RECT 42.865 83.145 44.075 84.235 ;
        RECT 42.865 82.435 43.385 82.975 ;
        RECT 43.555 82.605 44.075 83.145 ;
        RECT 44.245 83.070 44.535 84.235 ;
        RECT 44.710 83.095 45.045 84.065 ;
        RECT 45.215 83.095 45.385 84.235 ;
        RECT 45.555 83.895 47.585 84.065 ;
        RECT 40.535 81.685 40.930 82.180 ;
        RECT 41.290 82.015 41.665 82.210 ;
        RECT 41.495 81.870 41.665 82.015 ;
        RECT 41.945 81.880 42.185 82.255 ;
        RECT 42.355 81.685 42.690 82.190 ;
        RECT 42.865 81.685 44.075 82.435 ;
        RECT 44.710 82.425 44.880 83.095 ;
        RECT 45.555 82.925 45.725 83.895 ;
        RECT 45.050 82.595 45.305 82.925 ;
        RECT 45.530 82.595 45.725 82.925 ;
        RECT 45.895 83.555 47.020 83.725 ;
        RECT 45.135 82.425 45.305 82.595 ;
        RECT 45.895 82.425 46.065 83.555 ;
        RECT 44.245 81.685 44.535 82.410 ;
        RECT 44.710 81.855 44.965 82.425 ;
        RECT 45.135 82.255 46.065 82.425 ;
        RECT 46.235 83.215 47.245 83.385 ;
        RECT 46.235 82.415 46.405 83.215 ;
        RECT 45.890 82.220 46.065 82.255 ;
        RECT 45.135 81.685 45.465 82.085 ;
        RECT 45.890 81.855 46.420 82.220 ;
        RECT 46.610 82.195 46.885 83.015 ;
        RECT 46.605 82.025 46.885 82.195 ;
        RECT 46.610 81.855 46.885 82.025 ;
        RECT 47.055 81.855 47.245 83.215 ;
        RECT 47.415 83.230 47.585 83.895 ;
        RECT 47.755 83.475 47.925 84.235 ;
        RECT 48.160 83.475 48.675 83.885 ;
        RECT 47.415 83.040 48.165 83.230 ;
        RECT 48.335 82.665 48.675 83.475 ;
        RECT 49.395 83.565 49.565 84.065 ;
        RECT 49.735 83.735 50.065 84.235 ;
        RECT 49.395 83.395 50.060 83.565 ;
        RECT 47.445 82.495 48.675 82.665 ;
        RECT 49.310 82.575 49.660 83.225 ;
        RECT 47.425 81.685 47.935 82.220 ;
        RECT 48.155 81.890 48.400 82.495 ;
        RECT 49.830 82.405 50.060 83.395 ;
        RECT 49.395 82.235 50.060 82.405 ;
        RECT 49.395 81.945 49.565 82.235 ;
        RECT 49.735 81.685 50.065 82.065 ;
        RECT 50.235 81.945 50.420 84.065 ;
        RECT 50.660 83.775 50.925 84.235 ;
        RECT 51.095 83.640 51.345 84.065 ;
        RECT 51.555 83.790 52.660 83.960 ;
        RECT 51.040 83.510 51.345 83.640 ;
        RECT 50.590 82.315 50.870 83.265 ;
        RECT 51.040 82.405 51.210 83.510 ;
        RECT 51.380 82.725 51.620 83.320 ;
        RECT 51.790 83.255 52.320 83.620 ;
        RECT 51.790 82.555 51.960 83.255 ;
        RECT 52.490 83.175 52.660 83.790 ;
        RECT 52.830 83.435 53.000 84.235 ;
        RECT 53.170 83.735 53.420 84.065 ;
        RECT 53.645 83.765 54.530 83.935 ;
        RECT 52.490 83.085 53.000 83.175 ;
        RECT 51.040 82.275 51.265 82.405 ;
        RECT 51.435 82.335 51.960 82.555 ;
        RECT 52.130 82.915 53.000 83.085 ;
        RECT 50.675 81.685 50.925 82.145 ;
        RECT 51.095 82.135 51.265 82.275 ;
        RECT 52.130 82.135 52.300 82.915 ;
        RECT 52.830 82.845 53.000 82.915 ;
        RECT 52.510 82.665 52.710 82.695 ;
        RECT 53.170 82.665 53.340 83.735 ;
        RECT 53.510 82.845 53.700 83.565 ;
        RECT 52.510 82.365 53.340 82.665 ;
        RECT 53.870 82.635 54.190 83.595 ;
        RECT 51.095 81.965 51.430 82.135 ;
        RECT 51.625 81.965 52.300 82.135 ;
        RECT 52.620 81.685 52.990 82.185 ;
        RECT 53.170 82.135 53.340 82.365 ;
        RECT 53.725 82.305 54.190 82.635 ;
        RECT 54.360 82.925 54.530 83.765 ;
        RECT 54.710 83.735 55.025 84.235 ;
        RECT 55.255 83.505 55.595 84.065 ;
        RECT 54.700 83.130 55.595 83.505 ;
        RECT 55.765 83.225 55.935 84.235 ;
        RECT 55.405 82.925 55.595 83.130 ;
        RECT 56.105 83.175 56.435 84.020 ;
        RECT 56.670 83.285 56.935 84.055 ;
        RECT 57.105 83.515 57.435 84.235 ;
        RECT 57.625 83.695 57.885 84.055 ;
        RECT 58.055 83.865 58.385 84.235 ;
        RECT 58.555 83.695 58.815 84.055 ;
        RECT 57.625 83.465 58.815 83.695 ;
        RECT 59.385 83.285 59.675 84.055 ;
        RECT 56.105 83.095 56.495 83.175 ;
        RECT 56.280 83.045 56.495 83.095 ;
        RECT 54.360 82.595 55.235 82.925 ;
        RECT 55.405 82.595 56.155 82.925 ;
        RECT 54.360 82.135 54.530 82.595 ;
        RECT 55.405 82.425 55.605 82.595 ;
        RECT 56.325 82.465 56.495 83.045 ;
        RECT 56.270 82.425 56.495 82.465 ;
        RECT 53.170 81.965 53.575 82.135 ;
        RECT 53.745 81.965 54.530 82.135 ;
        RECT 54.805 81.685 55.015 82.215 ;
        RECT 55.275 81.900 55.605 82.425 ;
        RECT 56.115 82.340 56.495 82.425 ;
        RECT 55.775 81.685 55.945 82.295 ;
        RECT 56.115 81.905 56.445 82.340 ;
        RECT 56.670 81.865 57.005 83.285 ;
        RECT 57.180 83.105 59.675 83.285 ;
        RECT 59.920 83.445 60.455 84.065 ;
        RECT 57.180 82.415 57.405 83.105 ;
        RECT 57.605 82.595 57.885 82.925 ;
        RECT 58.065 82.595 58.640 82.925 ;
        RECT 58.820 82.595 59.255 82.925 ;
        RECT 59.435 82.595 59.705 82.925 ;
        RECT 59.920 82.425 60.235 83.445 ;
        RECT 60.625 83.435 60.955 84.235 ;
        RECT 61.440 83.265 61.830 83.440 ;
        RECT 60.405 83.095 61.830 83.265 ;
        RECT 62.185 83.095 62.445 84.235 ;
        RECT 60.405 82.595 60.575 83.095 ;
        RECT 57.180 82.225 59.665 82.415 ;
        RECT 57.185 81.685 57.930 82.055 ;
        RECT 58.495 81.865 58.750 82.225 ;
        RECT 58.930 81.685 59.260 82.055 ;
        RECT 59.440 81.865 59.665 82.225 ;
        RECT 59.920 81.855 60.535 82.425 ;
        RECT 60.825 82.365 61.090 82.925 ;
        RECT 61.260 82.195 61.430 83.095 ;
        RECT 62.615 83.085 62.945 84.065 ;
        RECT 63.115 83.095 63.395 84.235 ;
        RECT 63.565 83.145 64.775 84.235 ;
        RECT 61.600 82.365 61.955 82.925 ;
        RECT 62.205 82.675 62.540 82.925 ;
        RECT 62.710 82.485 62.880 83.085 ;
        RECT 63.050 82.655 63.385 82.925 ;
        RECT 60.705 81.685 60.920 82.195 ;
        RECT 61.150 81.865 61.430 82.195 ;
        RECT 61.610 81.685 61.850 82.195 ;
        RECT 62.185 81.855 62.880 82.485 ;
        RECT 63.085 81.685 63.395 82.485 ;
        RECT 63.565 82.435 64.085 82.975 ;
        RECT 64.255 82.605 64.775 83.145 ;
        RECT 64.950 83.095 65.270 84.235 ;
        RECT 65.450 82.925 65.645 83.975 ;
        RECT 65.825 83.385 66.155 84.065 ;
        RECT 66.355 83.435 66.610 84.235 ;
        RECT 65.825 83.105 66.175 83.385 ;
        RECT 67.890 83.265 68.280 83.440 ;
        RECT 68.765 83.435 69.095 84.235 ;
        RECT 69.265 83.445 69.800 84.065 ;
        RECT 65.010 82.875 65.270 82.925 ;
        RECT 65.005 82.705 65.270 82.875 ;
        RECT 65.010 82.595 65.270 82.705 ;
        RECT 65.450 82.595 65.835 82.925 ;
        RECT 66.005 82.725 66.175 83.105 ;
        RECT 66.365 82.895 66.610 83.255 ;
        RECT 67.890 83.095 69.315 83.265 ;
        RECT 66.005 82.555 66.525 82.725 ;
        RECT 63.565 81.685 64.775 82.435 ;
        RECT 64.950 82.215 66.165 82.385 ;
        RECT 64.950 81.865 65.240 82.215 ;
        RECT 65.435 81.685 65.765 82.045 ;
        RECT 65.935 81.910 66.165 82.215 ;
        RECT 66.355 82.195 66.525 82.555 ;
        RECT 67.765 82.365 68.120 82.925 ;
        RECT 68.290 82.195 68.460 83.095 ;
        RECT 68.630 82.365 68.895 82.925 ;
        RECT 69.145 82.595 69.315 83.095 ;
        RECT 69.485 82.425 69.800 83.445 ;
        RECT 70.005 83.070 70.295 84.235 ;
        RECT 70.620 83.225 70.920 84.065 ;
        RECT 71.115 83.395 71.365 84.235 ;
        RECT 71.955 83.645 72.760 84.065 ;
        RECT 71.535 83.475 73.100 83.645 ;
        RECT 71.535 83.225 71.705 83.475 ;
        RECT 70.620 83.055 71.705 83.225 ;
        RECT 70.465 82.595 70.795 82.885 ;
        RECT 70.965 82.425 71.135 83.055 ;
        RECT 71.875 82.925 72.195 83.305 ;
        RECT 72.385 83.215 72.760 83.305 ;
        RECT 72.365 83.045 72.760 83.215 ;
        RECT 72.930 83.225 73.100 83.475 ;
        RECT 73.270 83.395 73.600 84.235 ;
        RECT 73.770 83.475 74.435 84.065 ;
        RECT 72.930 83.055 73.850 83.225 ;
        RECT 71.305 82.675 71.635 82.885 ;
        RECT 71.815 82.675 72.195 82.925 ;
        RECT 72.385 82.885 72.760 83.045 ;
        RECT 73.680 82.885 73.850 83.055 ;
        RECT 72.385 82.675 72.870 82.885 ;
        RECT 73.060 82.675 73.510 82.885 ;
        RECT 73.680 82.675 74.015 82.885 ;
        RECT 74.185 82.505 74.435 83.475 ;
        RECT 66.355 82.025 66.555 82.195 ;
        RECT 66.355 81.990 66.525 82.025 ;
        RECT 67.870 81.685 68.110 82.195 ;
        RECT 68.290 81.865 68.570 82.195 ;
        RECT 68.800 81.685 69.015 82.195 ;
        RECT 69.185 81.855 69.800 82.425 ;
        RECT 70.005 81.685 70.295 82.410 ;
        RECT 70.625 82.245 71.135 82.425 ;
        RECT 71.540 82.335 73.240 82.505 ;
        RECT 71.540 82.245 71.925 82.335 ;
        RECT 70.625 81.855 70.955 82.245 ;
        RECT 71.125 81.905 72.310 82.075 ;
        RECT 72.570 81.685 72.740 82.155 ;
        RECT 72.910 81.870 73.240 82.335 ;
        RECT 73.410 81.685 73.580 82.505 ;
        RECT 73.750 81.865 74.435 82.505 ;
        RECT 75.530 83.095 75.865 84.065 ;
        RECT 76.035 83.095 76.205 84.235 ;
        RECT 76.375 83.895 78.405 84.065 ;
        RECT 75.530 82.425 75.700 83.095 ;
        RECT 76.375 82.925 76.545 83.895 ;
        RECT 75.870 82.595 76.125 82.925 ;
        RECT 76.350 82.595 76.545 82.925 ;
        RECT 76.715 83.555 77.840 83.725 ;
        RECT 75.955 82.425 76.125 82.595 ;
        RECT 76.715 82.425 76.885 83.555 ;
        RECT 75.530 81.855 75.785 82.425 ;
        RECT 75.955 82.255 76.885 82.425 ;
        RECT 77.055 83.215 78.065 83.385 ;
        RECT 77.055 82.415 77.225 83.215 ;
        RECT 77.430 82.875 77.705 83.015 ;
        RECT 77.425 82.705 77.705 82.875 ;
        RECT 76.710 82.220 76.885 82.255 ;
        RECT 75.955 81.685 76.285 82.085 ;
        RECT 76.710 81.855 77.240 82.220 ;
        RECT 77.430 81.855 77.705 82.705 ;
        RECT 77.875 81.855 78.065 83.215 ;
        RECT 78.235 83.230 78.405 83.895 ;
        RECT 78.575 83.475 78.745 84.235 ;
        RECT 78.980 83.475 79.495 83.885 ;
        RECT 78.235 83.040 78.985 83.230 ;
        RECT 79.155 82.665 79.495 83.475 ;
        RECT 79.755 83.305 79.925 84.065 ;
        RECT 80.105 83.475 80.435 84.235 ;
        RECT 79.755 83.135 80.420 83.305 ;
        RECT 80.605 83.160 80.875 84.065 ;
        RECT 80.250 82.990 80.420 83.135 ;
        RECT 78.265 82.495 79.495 82.665 ;
        RECT 79.685 82.585 80.015 82.955 ;
        RECT 80.250 82.660 80.535 82.990 ;
        RECT 78.245 81.685 78.755 82.220 ;
        RECT 78.975 81.890 79.220 82.495 ;
        RECT 80.250 82.405 80.420 82.660 ;
        RECT 79.755 82.235 80.420 82.405 ;
        RECT 80.705 82.360 80.875 83.160 ;
        RECT 81.045 83.145 82.715 84.235 ;
        RECT 79.755 81.855 79.925 82.235 ;
        RECT 80.105 81.685 80.435 82.065 ;
        RECT 80.615 81.855 80.875 82.360 ;
        RECT 81.045 82.455 81.795 82.975 ;
        RECT 81.965 82.625 82.715 83.145 ;
        RECT 82.885 83.145 84.095 84.235 ;
        RECT 82.885 82.605 83.405 83.145 ;
        RECT 81.045 81.685 82.715 82.455 ;
        RECT 83.575 82.435 84.095 82.975 ;
        RECT 82.885 81.685 84.095 82.435 ;
        RECT 5.520 81.515 84.180 81.685 ;
        RECT 5.605 80.765 6.815 81.515 ;
        RECT 6.985 80.970 12.330 81.515 ;
        RECT 12.505 80.970 17.850 81.515 ;
        RECT 5.605 80.225 6.125 80.765 ;
        RECT 6.295 80.055 6.815 80.595 ;
        RECT 8.570 80.140 8.910 80.970 ;
        RECT 5.605 78.965 6.815 80.055 ;
        RECT 10.390 79.400 10.740 80.650 ;
        RECT 14.090 80.140 14.430 80.970 ;
        RECT 18.025 80.745 19.695 81.515 ;
        RECT 20.330 80.775 20.585 81.345 ;
        RECT 20.755 81.115 21.085 81.515 ;
        RECT 21.510 80.980 22.040 81.345 ;
        RECT 21.510 80.945 21.685 80.980 ;
        RECT 20.755 80.775 21.685 80.945 ;
        RECT 15.910 79.400 16.260 80.650 ;
        RECT 18.025 80.225 18.775 80.745 ;
        RECT 18.945 80.055 19.695 80.575 ;
        RECT 6.985 78.965 12.330 79.400 ;
        RECT 12.505 78.965 17.850 79.400 ;
        RECT 18.025 78.965 19.695 80.055 ;
        RECT 20.330 80.105 20.500 80.775 ;
        RECT 20.755 80.605 20.925 80.775 ;
        RECT 20.670 80.275 20.925 80.605 ;
        RECT 21.150 80.275 21.345 80.605 ;
        RECT 20.330 79.135 20.665 80.105 ;
        RECT 20.835 78.965 21.005 80.105 ;
        RECT 21.175 79.305 21.345 80.275 ;
        RECT 21.515 79.645 21.685 80.775 ;
        RECT 21.855 79.985 22.025 80.785 ;
        RECT 22.230 80.495 22.505 81.345 ;
        RECT 22.225 80.325 22.505 80.495 ;
        RECT 22.230 80.185 22.505 80.325 ;
        RECT 22.675 79.985 22.865 81.345 ;
        RECT 23.045 80.980 23.555 81.515 ;
        RECT 23.775 80.705 24.020 81.310 ;
        RECT 24.465 80.970 29.810 81.515 ;
        RECT 23.065 80.535 24.295 80.705 ;
        RECT 21.855 79.815 22.865 79.985 ;
        RECT 23.035 79.970 23.785 80.160 ;
        RECT 21.515 79.475 22.640 79.645 ;
        RECT 23.035 79.305 23.205 79.970 ;
        RECT 23.955 79.725 24.295 80.535 ;
        RECT 26.050 80.140 26.390 80.970 ;
        RECT 29.985 80.765 31.195 81.515 ;
        RECT 31.365 80.790 31.655 81.515 ;
        RECT 31.915 80.965 32.085 81.255 ;
        RECT 32.255 81.135 32.585 81.515 ;
        RECT 31.915 80.795 32.580 80.965 ;
        RECT 21.175 79.135 23.205 79.305 ;
        RECT 23.375 78.965 23.545 79.725 ;
        RECT 23.780 79.315 24.295 79.725 ;
        RECT 27.870 79.400 28.220 80.650 ;
        RECT 29.985 80.225 30.505 80.765 ;
        RECT 30.675 80.055 31.195 80.595 ;
        RECT 24.465 78.965 29.810 79.400 ;
        RECT 29.985 78.965 31.195 80.055 ;
        RECT 31.365 78.965 31.655 80.130 ;
        RECT 31.830 79.975 32.180 80.625 ;
        RECT 32.350 79.805 32.580 80.795 ;
        RECT 31.915 79.635 32.580 79.805 ;
        RECT 31.915 79.135 32.085 79.635 ;
        RECT 32.255 78.965 32.585 79.465 ;
        RECT 32.755 79.135 32.940 81.255 ;
        RECT 33.195 81.055 33.445 81.515 ;
        RECT 33.615 81.065 33.950 81.235 ;
        RECT 34.145 81.065 34.820 81.235 ;
        RECT 33.615 80.925 33.785 81.065 ;
        RECT 33.110 79.935 33.390 80.885 ;
        RECT 33.560 80.795 33.785 80.925 ;
        RECT 33.560 79.690 33.730 80.795 ;
        RECT 33.955 80.645 34.480 80.865 ;
        RECT 33.900 79.880 34.140 80.475 ;
        RECT 34.310 79.945 34.480 80.645 ;
        RECT 34.650 80.285 34.820 81.065 ;
        RECT 35.140 81.015 35.510 81.515 ;
        RECT 35.690 81.065 36.095 81.235 ;
        RECT 36.265 81.065 37.050 81.235 ;
        RECT 35.690 80.835 35.860 81.065 ;
        RECT 35.030 80.535 35.860 80.835 ;
        RECT 36.245 80.565 36.710 80.895 ;
        RECT 35.030 80.505 35.230 80.535 ;
        RECT 35.350 80.285 35.520 80.355 ;
        RECT 34.650 80.115 35.520 80.285 ;
        RECT 35.010 80.025 35.520 80.115 ;
        RECT 33.560 79.560 33.865 79.690 ;
        RECT 34.310 79.580 34.840 79.945 ;
        RECT 33.180 78.965 33.445 79.425 ;
        RECT 33.615 79.135 33.865 79.560 ;
        RECT 35.010 79.410 35.180 80.025 ;
        RECT 34.075 79.240 35.180 79.410 ;
        RECT 35.350 78.965 35.520 79.765 ;
        RECT 35.690 79.465 35.860 80.535 ;
        RECT 36.030 79.635 36.220 80.355 ;
        RECT 36.390 79.605 36.710 80.565 ;
        RECT 36.880 80.605 37.050 81.065 ;
        RECT 37.325 80.985 37.535 81.515 ;
        RECT 37.795 80.775 38.125 81.300 ;
        RECT 38.295 80.905 38.465 81.515 ;
        RECT 38.635 80.860 38.965 81.295 ;
        RECT 38.635 80.775 39.015 80.860 ;
        RECT 37.925 80.605 38.125 80.775 ;
        RECT 38.790 80.735 39.015 80.775 ;
        RECT 36.880 80.275 37.755 80.605 ;
        RECT 37.925 80.275 38.675 80.605 ;
        RECT 35.690 79.135 35.940 79.465 ;
        RECT 36.880 79.435 37.050 80.275 ;
        RECT 37.925 80.070 38.115 80.275 ;
        RECT 38.845 80.155 39.015 80.735 ;
        RECT 38.800 80.105 39.015 80.155 ;
        RECT 37.220 79.695 38.115 80.070 ;
        RECT 38.625 80.025 39.015 80.105 ;
        RECT 39.185 80.840 39.455 81.185 ;
        RECT 39.645 81.115 40.025 81.515 ;
        RECT 40.195 80.945 40.365 81.295 ;
        RECT 40.535 81.115 40.865 81.515 ;
        RECT 41.065 80.945 41.235 81.295 ;
        RECT 41.435 81.015 41.765 81.515 ;
        RECT 39.185 80.105 39.355 80.840 ;
        RECT 39.625 80.775 41.235 80.945 ;
        RECT 42.495 80.965 42.665 81.255 ;
        RECT 42.835 81.135 43.165 81.515 ;
        RECT 39.625 80.605 39.795 80.775 ;
        RECT 39.525 80.275 39.795 80.605 ;
        RECT 39.965 80.275 40.370 80.605 ;
        RECT 39.625 80.105 39.795 80.275 ;
        RECT 36.165 79.265 37.050 79.435 ;
        RECT 37.230 78.965 37.545 79.465 ;
        RECT 37.775 79.135 38.115 79.695 ;
        RECT 38.285 78.965 38.455 79.975 ;
        RECT 38.625 79.180 38.955 80.025 ;
        RECT 39.185 79.135 39.455 80.105 ;
        RECT 39.625 79.935 40.350 80.105 ;
        RECT 40.540 79.985 41.250 80.605 ;
        RECT 41.420 80.275 41.770 80.845 ;
        RECT 42.495 80.795 43.160 80.965 ;
        RECT 40.180 79.815 40.350 79.935 ;
        RECT 41.450 79.815 41.770 80.105 ;
        RECT 42.410 79.975 42.760 80.625 ;
        RECT 39.665 78.965 39.945 79.765 ;
        RECT 40.180 79.645 41.770 79.815 ;
        RECT 42.930 79.805 43.160 80.795 ;
        RECT 42.495 79.635 43.160 79.805 ;
        RECT 40.115 79.185 41.770 79.475 ;
        RECT 42.495 79.135 42.665 79.635 ;
        RECT 42.835 78.965 43.165 79.465 ;
        RECT 43.335 79.135 43.520 81.255 ;
        RECT 43.775 81.055 44.025 81.515 ;
        RECT 44.195 81.065 44.530 81.235 ;
        RECT 44.725 81.065 45.400 81.235 ;
        RECT 44.195 80.925 44.365 81.065 ;
        RECT 43.690 79.935 43.970 80.885 ;
        RECT 44.140 80.795 44.365 80.925 ;
        RECT 44.140 79.690 44.310 80.795 ;
        RECT 44.535 80.645 45.060 80.865 ;
        RECT 44.480 79.880 44.720 80.475 ;
        RECT 44.890 79.945 45.060 80.645 ;
        RECT 45.230 80.285 45.400 81.065 ;
        RECT 45.720 81.015 46.090 81.515 ;
        RECT 46.270 81.065 46.675 81.235 ;
        RECT 46.845 81.065 47.630 81.235 ;
        RECT 46.270 80.835 46.440 81.065 ;
        RECT 45.610 80.535 46.440 80.835 ;
        RECT 46.825 80.565 47.290 80.895 ;
        RECT 45.610 80.505 45.810 80.535 ;
        RECT 45.930 80.285 46.100 80.355 ;
        RECT 45.230 80.115 46.100 80.285 ;
        RECT 45.590 80.025 46.100 80.115 ;
        RECT 44.140 79.560 44.445 79.690 ;
        RECT 44.890 79.580 45.420 79.945 ;
        RECT 43.760 78.965 44.025 79.425 ;
        RECT 44.195 79.135 44.445 79.560 ;
        RECT 45.590 79.410 45.760 80.025 ;
        RECT 44.655 79.240 45.760 79.410 ;
        RECT 45.930 78.965 46.100 79.765 ;
        RECT 46.270 79.465 46.440 80.535 ;
        RECT 46.610 79.635 46.800 80.355 ;
        RECT 46.970 79.605 47.290 80.565 ;
        RECT 47.460 80.605 47.630 81.065 ;
        RECT 47.905 80.985 48.115 81.515 ;
        RECT 48.375 80.775 48.705 81.300 ;
        RECT 48.875 80.905 49.045 81.515 ;
        RECT 49.215 80.860 49.545 81.295 ;
        RECT 49.215 80.775 49.595 80.860 ;
        RECT 48.505 80.605 48.705 80.775 ;
        RECT 49.370 80.735 49.595 80.775 ;
        RECT 47.460 80.275 48.335 80.605 ;
        RECT 48.505 80.275 49.255 80.605 ;
        RECT 46.270 79.135 46.520 79.465 ;
        RECT 47.460 79.435 47.630 80.275 ;
        RECT 48.505 80.070 48.695 80.275 ;
        RECT 49.425 80.155 49.595 80.735 ;
        RECT 49.380 80.105 49.595 80.155 ;
        RECT 47.800 79.695 48.695 80.070 ;
        RECT 49.205 80.025 49.595 80.105 ;
        RECT 49.765 80.775 50.150 81.345 ;
        RECT 50.320 81.055 50.645 81.515 ;
        RECT 51.165 80.885 51.445 81.345 ;
        RECT 49.765 80.105 50.045 80.775 ;
        RECT 50.320 80.715 51.445 80.885 ;
        RECT 50.320 80.605 50.770 80.715 ;
        RECT 50.215 80.275 50.770 80.605 ;
        RECT 51.635 80.545 52.035 81.345 ;
        RECT 52.435 81.055 52.705 81.515 ;
        RECT 52.875 80.885 53.160 81.345 ;
        RECT 46.745 79.265 47.630 79.435 ;
        RECT 47.810 78.965 48.125 79.465 ;
        RECT 48.355 79.135 48.695 79.695 ;
        RECT 48.865 78.965 49.035 79.975 ;
        RECT 49.205 79.180 49.535 80.025 ;
        RECT 49.765 79.135 50.150 80.105 ;
        RECT 50.320 79.815 50.770 80.275 ;
        RECT 50.940 79.985 52.035 80.545 ;
        RECT 50.320 79.595 51.445 79.815 ;
        RECT 50.320 78.965 50.645 79.425 ;
        RECT 51.165 79.135 51.445 79.595 ;
        RECT 51.635 79.135 52.035 79.985 ;
        RECT 52.205 80.715 53.160 80.885 ;
        RECT 53.445 80.745 56.955 81.515 ;
        RECT 57.125 80.790 57.415 81.515 ;
        RECT 52.205 79.815 52.415 80.715 ;
        RECT 52.585 79.985 53.275 80.545 ;
        RECT 53.445 80.225 55.095 80.745 ;
        RECT 58.505 80.695 58.765 81.515 ;
        RECT 58.935 80.695 59.265 81.115 ;
        RECT 59.445 81.030 60.235 81.295 ;
        RECT 59.015 80.605 59.265 80.695 ;
        RECT 55.265 80.055 56.955 80.575 ;
        RECT 52.205 79.595 53.160 79.815 ;
        RECT 52.435 78.965 52.705 79.425 ;
        RECT 52.875 79.135 53.160 79.595 ;
        RECT 53.445 78.965 56.955 80.055 ;
        RECT 57.125 78.965 57.415 80.130 ;
        RECT 58.505 79.645 58.845 80.525 ;
        RECT 59.015 80.355 59.810 80.605 ;
        RECT 58.505 78.965 58.765 79.475 ;
        RECT 59.015 79.135 59.185 80.355 ;
        RECT 59.980 80.175 60.235 81.030 ;
        RECT 60.405 80.875 60.605 81.295 ;
        RECT 60.795 81.055 61.125 81.515 ;
        RECT 60.405 80.355 60.815 80.875 ;
        RECT 61.295 80.865 61.555 81.345 ;
        RECT 60.985 80.175 61.215 80.605 ;
        RECT 59.425 80.005 61.215 80.175 ;
        RECT 59.425 79.640 59.675 80.005 ;
        RECT 59.845 79.645 60.175 79.835 ;
        RECT 60.395 79.710 61.110 80.005 ;
        RECT 61.385 79.835 61.555 80.865 ;
        RECT 59.845 79.470 60.040 79.645 ;
        RECT 59.425 78.965 60.040 79.470 ;
        RECT 60.210 79.135 60.685 79.475 ;
        RECT 60.855 78.965 61.070 79.510 ;
        RECT 61.280 79.135 61.555 79.835 ;
        RECT 61.745 80.825 61.985 81.345 ;
        RECT 62.155 81.020 62.550 81.515 ;
        RECT 63.115 81.185 63.285 81.330 ;
        RECT 62.910 80.990 63.285 81.185 ;
        RECT 61.745 80.020 61.920 80.825 ;
        RECT 62.910 80.655 63.080 80.990 ;
        RECT 63.565 80.945 63.805 81.320 ;
        RECT 63.975 81.010 64.310 81.515 ;
        RECT 63.565 80.795 63.785 80.945 ;
        RECT 62.095 80.295 63.080 80.655 ;
        RECT 63.250 80.465 63.785 80.795 ;
        RECT 62.095 80.275 63.380 80.295 ;
        RECT 62.520 80.125 63.380 80.275 ;
        RECT 61.745 79.235 62.050 80.020 ;
        RECT 62.225 79.645 62.920 79.955 ;
        RECT 62.230 78.965 62.915 79.435 ;
        RECT 63.095 79.180 63.380 80.125 ;
        RECT 63.550 79.815 63.785 80.465 ;
        RECT 63.955 79.985 64.255 80.835 ;
        RECT 64.485 80.745 67.075 81.515 ;
        RECT 67.245 80.865 67.505 81.345 ;
        RECT 67.675 80.975 67.925 81.515 ;
        RECT 64.485 80.225 65.695 80.745 ;
        RECT 65.865 80.055 67.075 80.575 ;
        RECT 63.550 79.585 64.225 79.815 ;
        RECT 63.555 78.965 63.885 79.415 ;
        RECT 64.055 79.155 64.225 79.585 ;
        RECT 64.485 78.965 67.075 80.055 ;
        RECT 67.245 79.835 67.415 80.865 ;
        RECT 68.095 80.810 68.315 81.295 ;
        RECT 67.585 80.215 67.815 80.610 ;
        RECT 67.985 80.385 68.315 80.810 ;
        RECT 68.485 81.135 69.375 81.305 ;
        RECT 68.485 80.410 68.655 81.135 ;
        RECT 69.545 80.970 74.890 81.515 ;
        RECT 68.825 80.580 69.375 80.965 ;
        RECT 68.485 80.340 69.375 80.410 ;
        RECT 68.480 80.315 69.375 80.340 ;
        RECT 68.470 80.300 69.375 80.315 ;
        RECT 68.465 80.285 69.375 80.300 ;
        RECT 68.455 80.280 69.375 80.285 ;
        RECT 68.450 80.270 69.375 80.280 ;
        RECT 68.445 80.260 69.375 80.270 ;
        RECT 68.435 80.255 69.375 80.260 ;
        RECT 68.425 80.245 69.375 80.255 ;
        RECT 68.415 80.240 69.375 80.245 ;
        RECT 68.415 80.235 68.750 80.240 ;
        RECT 68.400 80.230 68.750 80.235 ;
        RECT 68.385 80.220 68.750 80.230 ;
        RECT 68.360 80.215 68.750 80.220 ;
        RECT 67.585 80.210 68.750 80.215 ;
        RECT 67.585 80.175 68.720 80.210 ;
        RECT 67.585 80.150 68.685 80.175 ;
        RECT 67.585 80.120 68.655 80.150 ;
        RECT 67.585 80.090 68.635 80.120 ;
        RECT 67.585 80.060 68.615 80.090 ;
        RECT 67.585 80.050 68.545 80.060 ;
        RECT 67.585 80.040 68.520 80.050 ;
        RECT 67.585 80.025 68.500 80.040 ;
        RECT 67.585 80.010 68.480 80.025 ;
        RECT 67.690 80.000 68.475 80.010 ;
        RECT 67.690 79.965 68.460 80.000 ;
        RECT 67.245 79.135 67.520 79.835 ;
        RECT 67.690 79.715 68.445 79.965 ;
        RECT 68.615 79.645 68.945 79.890 ;
        RECT 69.115 79.790 69.375 80.240 ;
        RECT 71.130 80.140 71.470 80.970 ;
        RECT 75.065 80.745 77.655 81.515 ;
        RECT 77.915 80.965 78.085 81.345 ;
        RECT 78.265 81.135 78.595 81.515 ;
        RECT 77.915 80.795 78.580 80.965 ;
        RECT 78.775 80.840 79.035 81.345 ;
        RECT 68.760 79.620 68.945 79.645 ;
        RECT 68.760 79.520 69.375 79.620 ;
        RECT 67.690 78.965 67.945 79.510 ;
        RECT 68.115 79.135 68.595 79.475 ;
        RECT 68.770 78.965 69.375 79.520 ;
        RECT 72.950 79.400 73.300 80.650 ;
        RECT 75.065 80.225 76.275 80.745 ;
        RECT 76.445 80.055 77.655 80.575 ;
        RECT 77.845 80.245 78.175 80.615 ;
        RECT 78.410 80.540 78.580 80.795 ;
        RECT 78.410 80.210 78.695 80.540 ;
        RECT 78.410 80.065 78.580 80.210 ;
        RECT 69.545 78.965 74.890 79.400 ;
        RECT 75.065 78.965 77.655 80.055 ;
        RECT 77.915 79.895 78.580 80.065 ;
        RECT 78.865 80.040 79.035 80.840 ;
        RECT 77.915 79.135 78.085 79.895 ;
        RECT 78.265 78.965 78.595 79.725 ;
        RECT 78.765 79.135 79.035 80.040 ;
        RECT 79.205 80.775 79.590 81.345 ;
        RECT 79.760 81.055 80.085 81.515 ;
        RECT 80.605 80.885 80.885 81.345 ;
        RECT 79.205 80.105 79.485 80.775 ;
        RECT 79.760 80.715 80.885 80.885 ;
        RECT 79.760 80.605 80.210 80.715 ;
        RECT 79.655 80.275 80.210 80.605 ;
        RECT 81.075 80.545 81.475 81.345 ;
        RECT 81.875 81.055 82.145 81.515 ;
        RECT 82.315 80.885 82.600 81.345 ;
        RECT 79.205 79.135 79.590 80.105 ;
        RECT 79.760 79.815 80.210 80.275 ;
        RECT 80.380 79.985 81.475 80.545 ;
        RECT 79.760 79.595 80.885 79.815 ;
        RECT 79.760 78.965 80.085 79.425 ;
        RECT 80.605 79.135 80.885 79.595 ;
        RECT 81.075 79.135 81.475 79.985 ;
        RECT 81.645 80.715 82.600 80.885 ;
        RECT 82.885 80.765 84.095 81.515 ;
        RECT 81.645 79.815 81.855 80.715 ;
        RECT 82.025 79.985 82.715 80.545 ;
        RECT 82.885 80.055 83.405 80.595 ;
        RECT 83.575 80.225 84.095 80.765 ;
        RECT 81.645 79.595 82.600 79.815 ;
        RECT 81.875 78.965 82.145 79.425 ;
        RECT 82.315 79.135 82.600 79.595 ;
        RECT 82.885 78.965 84.095 80.055 ;
        RECT 5.520 78.795 84.180 78.965 ;
        RECT 5.605 77.705 6.815 78.795 ;
        RECT 6.985 77.705 8.655 78.795 ;
        RECT 5.605 76.995 6.125 77.535 ;
        RECT 6.295 77.165 6.815 77.705 ;
        RECT 6.985 77.015 7.735 77.535 ;
        RECT 7.905 77.185 8.655 77.705 ;
        RECT 9.285 78.075 9.745 78.625 ;
        RECT 9.935 78.075 10.265 78.795 ;
        RECT 5.605 76.245 6.815 76.995 ;
        RECT 6.985 76.245 8.655 77.015 ;
        RECT 9.285 76.705 9.535 78.075 ;
        RECT 10.465 77.905 10.765 78.455 ;
        RECT 10.935 78.125 11.215 78.795 ;
        RECT 9.825 77.735 10.765 77.905 ;
        RECT 9.825 77.485 9.995 77.735 ;
        RECT 11.135 77.485 11.400 77.845 ;
        RECT 11.585 77.655 11.845 78.795 ;
        RECT 12.015 77.645 12.345 78.625 ;
        RECT 12.515 77.655 12.795 78.795 ;
        RECT 12.975 77.825 13.305 78.610 ;
        RECT 12.975 77.655 13.655 77.825 ;
        RECT 13.835 77.655 14.165 78.795 ;
        RECT 15.265 77.655 15.525 78.795 ;
        RECT 15.765 78.285 17.380 78.615 ;
        RECT 12.105 77.605 12.280 77.645 ;
        RECT 9.705 77.155 9.995 77.485 ;
        RECT 10.165 77.235 10.505 77.485 ;
        RECT 10.725 77.235 11.400 77.485 ;
        RECT 11.605 77.235 11.940 77.485 ;
        RECT 9.825 77.065 9.995 77.155 ;
        RECT 9.825 76.875 11.215 77.065 ;
        RECT 12.110 77.045 12.280 77.605 ;
        RECT 12.450 77.215 12.785 77.485 ;
        RECT 12.965 77.235 13.315 77.485 ;
        RECT 13.485 77.055 13.655 77.655 ;
        RECT 15.775 77.485 15.945 78.045 ;
        RECT 16.205 77.945 17.380 78.115 ;
        RECT 17.550 77.995 17.830 78.795 ;
        RECT 16.205 77.655 16.535 77.945 ;
        RECT 17.210 77.825 17.380 77.945 ;
        RECT 16.705 77.485 16.950 77.775 ;
        RECT 17.210 77.655 17.870 77.825 ;
        RECT 18.040 77.655 18.315 78.625 ;
        RECT 17.700 77.485 17.870 77.655 ;
        RECT 13.825 77.235 14.175 77.485 ;
        RECT 15.270 77.235 15.605 77.485 ;
        RECT 15.775 77.155 16.490 77.485 ;
        RECT 16.705 77.155 17.530 77.485 ;
        RECT 17.700 77.155 17.975 77.485 ;
        RECT 15.775 77.065 16.025 77.155 ;
        RECT 9.285 76.415 9.845 76.705 ;
        RECT 10.015 76.245 10.265 76.705 ;
        RECT 10.885 76.515 11.215 76.875 ;
        RECT 11.585 76.415 12.280 77.045 ;
        RECT 12.485 76.245 12.795 77.045 ;
        RECT 12.985 76.245 13.225 77.055 ;
        RECT 13.395 76.415 13.725 77.055 ;
        RECT 13.895 76.245 14.165 77.055 ;
        RECT 15.265 76.245 15.525 77.065 ;
        RECT 15.695 76.645 16.025 77.065 ;
        RECT 17.700 76.985 17.870 77.155 ;
        RECT 16.205 76.815 17.870 76.985 ;
        RECT 18.145 76.920 18.315 77.655 ;
        RECT 18.485 77.630 18.775 78.795 ;
        RECT 18.945 77.705 20.155 78.795 ;
        RECT 18.945 76.995 19.465 77.535 ;
        RECT 19.635 77.165 20.155 77.705 ;
        RECT 20.330 77.655 20.665 78.625 ;
        RECT 20.835 77.655 21.005 78.795 ;
        RECT 21.175 78.455 23.205 78.625 ;
        RECT 16.205 76.415 16.465 76.815 ;
        RECT 16.635 76.245 16.965 76.645 ;
        RECT 17.135 76.465 17.305 76.815 ;
        RECT 17.475 76.245 17.850 76.645 ;
        RECT 18.040 76.575 18.315 76.920 ;
        RECT 18.485 76.245 18.775 76.970 ;
        RECT 18.945 76.245 20.155 76.995 ;
        RECT 20.330 76.985 20.500 77.655 ;
        RECT 21.175 77.485 21.345 78.455 ;
        RECT 20.670 77.155 20.925 77.485 ;
        RECT 21.150 77.155 21.345 77.485 ;
        RECT 21.515 78.115 22.640 78.285 ;
        RECT 20.755 76.985 20.925 77.155 ;
        RECT 21.515 76.985 21.685 78.115 ;
        RECT 20.330 76.415 20.585 76.985 ;
        RECT 20.755 76.815 21.685 76.985 ;
        RECT 21.855 77.775 22.865 77.945 ;
        RECT 21.855 76.975 22.025 77.775 ;
        RECT 22.230 77.435 22.505 77.575 ;
        RECT 22.225 77.265 22.505 77.435 ;
        RECT 21.510 76.780 21.685 76.815 ;
        RECT 20.755 76.245 21.085 76.645 ;
        RECT 21.510 76.415 22.040 76.780 ;
        RECT 22.230 76.415 22.505 77.265 ;
        RECT 22.675 76.415 22.865 77.775 ;
        RECT 23.035 77.790 23.205 78.455 ;
        RECT 23.375 78.035 23.545 78.795 ;
        RECT 23.780 78.035 24.295 78.445 ;
        RECT 24.465 78.360 29.810 78.795 ;
        RECT 23.035 77.600 23.785 77.790 ;
        RECT 23.955 77.225 24.295 78.035 ;
        RECT 23.065 77.055 24.295 77.225 ;
        RECT 23.045 76.245 23.555 76.780 ;
        RECT 23.775 76.450 24.020 77.055 ;
        RECT 26.050 76.790 26.390 77.620 ;
        RECT 27.870 77.110 28.220 78.360 ;
        RECT 30.905 78.035 31.420 78.445 ;
        RECT 31.655 78.035 31.825 78.795 ;
        RECT 31.995 78.455 34.025 78.625 ;
        RECT 30.905 77.225 31.245 78.035 ;
        RECT 31.995 77.790 32.165 78.455 ;
        RECT 32.560 78.115 33.685 78.285 ;
        RECT 31.415 77.600 32.165 77.790 ;
        RECT 32.335 77.775 33.345 77.945 ;
        RECT 30.905 77.055 32.135 77.225 ;
        RECT 24.465 76.245 29.810 76.790 ;
        RECT 31.180 76.450 31.425 77.055 ;
        RECT 31.645 76.245 32.155 76.780 ;
        RECT 32.335 76.415 32.525 77.775 ;
        RECT 32.695 76.755 32.970 77.575 ;
        RECT 33.175 76.975 33.345 77.775 ;
        RECT 33.515 76.985 33.685 78.115 ;
        RECT 33.855 77.485 34.025 78.455 ;
        RECT 34.195 77.655 34.365 78.795 ;
        RECT 34.535 77.655 34.870 78.625 ;
        RECT 35.045 77.705 36.715 78.795 ;
        RECT 33.855 77.155 34.050 77.485 ;
        RECT 34.275 77.155 34.530 77.485 ;
        RECT 34.275 76.985 34.445 77.155 ;
        RECT 34.700 76.985 34.870 77.655 ;
        RECT 33.515 76.815 34.445 76.985 ;
        RECT 33.515 76.780 33.690 76.815 ;
        RECT 32.695 76.585 32.975 76.755 ;
        RECT 32.695 76.415 32.970 76.585 ;
        RECT 33.160 76.415 33.690 76.780 ;
        RECT 34.115 76.245 34.445 76.645 ;
        RECT 34.615 76.415 34.870 76.985 ;
        RECT 35.045 77.015 35.795 77.535 ;
        RECT 35.965 77.185 36.715 77.705 ;
        RECT 36.885 77.655 37.270 78.625 ;
        RECT 37.440 78.335 37.765 78.795 ;
        RECT 38.285 78.165 38.565 78.625 ;
        RECT 37.440 77.945 38.565 78.165 ;
        RECT 35.045 76.245 36.715 77.015 ;
        RECT 36.885 76.985 37.165 77.655 ;
        RECT 37.440 77.485 37.890 77.945 ;
        RECT 38.755 77.775 39.155 78.625 ;
        RECT 39.555 78.335 39.825 78.795 ;
        RECT 39.995 78.165 40.280 78.625 ;
        RECT 37.335 77.155 37.890 77.485 ;
        RECT 38.060 77.215 39.155 77.775 ;
        RECT 37.440 77.045 37.890 77.155 ;
        RECT 36.885 76.415 37.270 76.985 ;
        RECT 37.440 76.875 38.565 77.045 ;
        RECT 37.440 76.245 37.765 76.705 ;
        RECT 38.285 76.415 38.565 76.875 ;
        RECT 38.755 76.415 39.155 77.215 ;
        RECT 39.325 77.945 40.280 78.165 ;
        RECT 40.680 78.165 40.965 78.625 ;
        RECT 41.135 78.335 41.405 78.795 ;
        RECT 40.680 77.945 41.635 78.165 ;
        RECT 39.325 77.045 39.535 77.945 ;
        RECT 39.705 77.215 40.395 77.775 ;
        RECT 40.565 77.215 41.255 77.775 ;
        RECT 41.425 77.045 41.635 77.945 ;
        RECT 39.325 76.875 40.280 77.045 ;
        RECT 39.555 76.245 39.825 76.705 ;
        RECT 39.995 76.415 40.280 76.875 ;
        RECT 40.680 76.875 41.635 77.045 ;
        RECT 41.805 77.775 42.205 78.625 ;
        RECT 42.395 78.165 42.675 78.625 ;
        RECT 43.195 78.335 43.520 78.795 ;
        RECT 42.395 77.945 43.520 78.165 ;
        RECT 41.805 77.215 42.900 77.775 ;
        RECT 43.070 77.485 43.520 77.945 ;
        RECT 43.690 77.655 44.075 78.625 ;
        RECT 40.680 76.415 40.965 76.875 ;
        RECT 41.135 76.245 41.405 76.705 ;
        RECT 41.805 76.415 42.205 77.215 ;
        RECT 43.070 77.155 43.625 77.485 ;
        RECT 43.070 77.045 43.520 77.155 ;
        RECT 42.395 76.875 43.520 77.045 ;
        RECT 43.795 76.985 44.075 77.655 ;
        RECT 44.245 77.630 44.535 78.795 ;
        RECT 44.705 77.925 44.980 78.625 ;
        RECT 45.150 78.250 45.405 78.795 ;
        RECT 45.575 78.285 46.055 78.625 ;
        RECT 46.230 78.240 46.835 78.795 ;
        RECT 46.220 78.140 46.835 78.240 ;
        RECT 46.220 78.115 46.405 78.140 ;
        RECT 42.395 76.415 42.675 76.875 ;
        RECT 43.195 76.245 43.520 76.705 ;
        RECT 43.690 76.415 44.075 76.985 ;
        RECT 44.245 76.245 44.535 76.970 ;
        RECT 44.705 76.895 44.875 77.925 ;
        RECT 45.150 77.795 45.905 78.045 ;
        RECT 46.075 77.870 46.405 78.115 ;
        RECT 45.150 77.760 45.920 77.795 ;
        RECT 45.150 77.750 45.935 77.760 ;
        RECT 45.045 77.735 45.940 77.750 ;
        RECT 45.045 77.720 45.960 77.735 ;
        RECT 45.045 77.710 45.980 77.720 ;
        RECT 45.045 77.700 46.005 77.710 ;
        RECT 45.045 77.670 46.075 77.700 ;
        RECT 45.045 77.640 46.095 77.670 ;
        RECT 45.045 77.610 46.115 77.640 ;
        RECT 45.045 77.585 46.145 77.610 ;
        RECT 45.045 77.550 46.180 77.585 ;
        RECT 45.045 77.545 46.210 77.550 ;
        RECT 45.045 77.150 45.275 77.545 ;
        RECT 45.820 77.540 46.210 77.545 ;
        RECT 45.845 77.530 46.210 77.540 ;
        RECT 45.860 77.525 46.210 77.530 ;
        RECT 45.875 77.520 46.210 77.525 ;
        RECT 46.575 77.520 46.835 77.970 ;
        RECT 45.875 77.515 46.835 77.520 ;
        RECT 45.885 77.505 46.835 77.515 ;
        RECT 45.895 77.500 46.835 77.505 ;
        RECT 45.905 77.490 46.835 77.500 ;
        RECT 45.910 77.480 46.835 77.490 ;
        RECT 45.915 77.475 46.835 77.480 ;
        RECT 45.925 77.460 46.835 77.475 ;
        RECT 45.930 77.445 46.835 77.460 ;
        RECT 45.940 77.420 46.835 77.445 ;
        RECT 45.445 76.950 45.775 77.375 ;
        RECT 44.705 76.415 44.965 76.895 ;
        RECT 45.135 76.245 45.385 76.785 ;
        RECT 45.555 76.465 45.775 76.950 ;
        RECT 45.945 77.350 46.835 77.420 ;
        RECT 47.010 77.655 47.345 78.625 ;
        RECT 47.515 77.655 47.685 78.795 ;
        RECT 47.855 78.455 49.885 78.625 ;
        RECT 45.945 76.625 46.115 77.350 ;
        RECT 46.285 76.795 46.835 77.180 ;
        RECT 47.010 76.985 47.180 77.655 ;
        RECT 47.855 77.485 48.025 78.455 ;
        RECT 47.350 77.155 47.605 77.485 ;
        RECT 47.830 77.155 48.025 77.485 ;
        RECT 48.195 78.115 49.320 78.285 ;
        RECT 47.435 76.985 47.605 77.155 ;
        RECT 48.195 76.985 48.365 78.115 ;
        RECT 45.945 76.455 46.835 76.625 ;
        RECT 47.010 76.415 47.265 76.985 ;
        RECT 47.435 76.815 48.365 76.985 ;
        RECT 48.535 77.775 49.545 77.945 ;
        RECT 48.535 76.975 48.705 77.775 ;
        RECT 48.190 76.780 48.365 76.815 ;
        RECT 47.435 76.245 47.765 76.645 ;
        RECT 48.190 76.415 48.720 76.780 ;
        RECT 48.910 76.755 49.185 77.575 ;
        RECT 48.905 76.585 49.185 76.755 ;
        RECT 48.910 76.415 49.185 76.585 ;
        RECT 49.355 76.415 49.545 77.775 ;
        RECT 49.715 77.790 49.885 78.455 ;
        RECT 50.055 78.035 50.225 78.795 ;
        RECT 50.460 78.035 50.975 78.445 ;
        RECT 51.145 78.360 56.490 78.795 ;
        RECT 49.715 77.600 50.465 77.790 ;
        RECT 50.635 77.225 50.975 78.035 ;
        RECT 49.745 77.055 50.975 77.225 ;
        RECT 49.725 76.245 50.235 76.780 ;
        RECT 50.455 76.450 50.700 77.055 ;
        RECT 52.730 76.790 53.070 77.620 ;
        RECT 54.550 77.110 54.900 78.360 ;
        RECT 56.780 78.165 57.065 78.625 ;
        RECT 57.235 78.335 57.505 78.795 ;
        RECT 56.780 77.945 57.735 78.165 ;
        RECT 56.665 77.215 57.355 77.775 ;
        RECT 57.525 77.045 57.735 77.945 ;
        RECT 56.780 76.875 57.735 77.045 ;
        RECT 57.905 77.775 58.305 78.625 ;
        RECT 58.495 78.165 58.775 78.625 ;
        RECT 59.295 78.335 59.620 78.795 ;
        RECT 58.495 77.945 59.620 78.165 ;
        RECT 57.905 77.215 59.000 77.775 ;
        RECT 59.170 77.485 59.620 77.945 ;
        RECT 59.790 77.655 60.175 78.625 ;
        RECT 60.345 78.240 60.950 78.795 ;
        RECT 61.125 78.285 61.605 78.625 ;
        RECT 61.775 78.250 62.030 78.795 ;
        RECT 60.345 78.140 60.960 78.240 ;
        RECT 60.775 78.115 60.960 78.140 ;
        RECT 51.145 76.245 56.490 76.790 ;
        RECT 56.780 76.415 57.065 76.875 ;
        RECT 57.235 76.245 57.505 76.705 ;
        RECT 57.905 76.415 58.305 77.215 ;
        RECT 59.170 77.155 59.725 77.485 ;
        RECT 59.170 77.045 59.620 77.155 ;
        RECT 58.495 76.875 59.620 77.045 ;
        RECT 59.895 76.985 60.175 77.655 ;
        RECT 60.345 77.520 60.605 77.970 ;
        RECT 60.775 77.870 61.105 78.115 ;
        RECT 61.275 77.795 62.030 78.045 ;
        RECT 62.200 77.925 62.475 78.625 ;
        RECT 61.260 77.760 62.030 77.795 ;
        RECT 61.245 77.750 62.030 77.760 ;
        RECT 61.240 77.735 62.135 77.750 ;
        RECT 61.220 77.720 62.135 77.735 ;
        RECT 61.200 77.710 62.135 77.720 ;
        RECT 61.175 77.700 62.135 77.710 ;
        RECT 61.105 77.670 62.135 77.700 ;
        RECT 61.085 77.640 62.135 77.670 ;
        RECT 61.065 77.610 62.135 77.640 ;
        RECT 61.035 77.585 62.135 77.610 ;
        RECT 61.000 77.550 62.135 77.585 ;
        RECT 60.970 77.545 62.135 77.550 ;
        RECT 60.970 77.540 61.360 77.545 ;
        RECT 60.970 77.530 61.335 77.540 ;
        RECT 60.970 77.525 61.320 77.530 ;
        RECT 60.970 77.520 61.305 77.525 ;
        RECT 60.345 77.515 61.305 77.520 ;
        RECT 60.345 77.505 61.295 77.515 ;
        RECT 60.345 77.500 61.285 77.505 ;
        RECT 60.345 77.490 61.275 77.500 ;
        RECT 60.345 77.480 61.270 77.490 ;
        RECT 60.345 77.475 61.265 77.480 ;
        RECT 60.345 77.460 61.255 77.475 ;
        RECT 60.345 77.445 61.250 77.460 ;
        RECT 60.345 77.420 61.240 77.445 ;
        RECT 60.345 77.350 61.235 77.420 ;
        RECT 58.495 76.415 58.775 76.875 ;
        RECT 59.295 76.245 59.620 76.705 ;
        RECT 59.790 76.415 60.175 76.985 ;
        RECT 60.345 76.795 60.895 77.180 ;
        RECT 61.065 76.625 61.235 77.350 ;
        RECT 60.345 76.455 61.235 76.625 ;
        RECT 61.405 76.950 61.735 77.375 ;
        RECT 61.905 77.150 62.135 77.545 ;
        RECT 61.405 76.465 61.625 76.950 ;
        RECT 62.305 76.895 62.475 77.925 ;
        RECT 62.645 77.705 65.235 78.795 ;
        RECT 61.795 76.245 62.045 76.785 ;
        RECT 62.215 76.415 62.475 76.895 ;
        RECT 62.645 77.015 63.855 77.535 ;
        RECT 64.025 77.185 65.235 77.705 ;
        RECT 66.020 77.785 66.320 78.625 ;
        RECT 66.515 77.955 66.765 78.795 ;
        RECT 67.355 78.205 68.160 78.625 ;
        RECT 66.935 78.035 68.500 78.205 ;
        RECT 66.935 77.785 67.105 78.035 ;
        RECT 66.020 77.615 67.105 77.785 ;
        RECT 65.865 77.155 66.195 77.445 ;
        RECT 62.645 76.245 65.235 77.015 ;
        RECT 66.365 76.985 66.535 77.615 ;
        RECT 67.275 77.485 67.595 77.865 ;
        RECT 66.705 77.235 67.035 77.445 ;
        RECT 67.215 77.235 67.595 77.485 ;
        RECT 67.785 77.445 68.160 77.865 ;
        RECT 68.330 77.785 68.500 78.035 ;
        RECT 68.670 77.955 69.000 78.795 ;
        RECT 69.170 78.035 69.835 78.625 ;
        RECT 68.330 77.615 69.250 77.785 ;
        RECT 69.080 77.445 69.250 77.615 ;
        RECT 67.785 77.435 68.270 77.445 ;
        RECT 67.765 77.265 68.270 77.435 ;
        RECT 67.785 77.235 68.270 77.265 ;
        RECT 68.460 77.235 68.910 77.445 ;
        RECT 69.080 77.235 69.415 77.445 ;
        RECT 69.585 77.065 69.835 78.035 ;
        RECT 70.005 77.630 70.295 78.795 ;
        RECT 70.470 78.405 70.805 78.625 ;
        RECT 71.810 78.415 72.165 78.795 ;
        RECT 70.470 77.785 70.725 78.405 ;
        RECT 70.975 78.245 71.205 78.285 ;
        RECT 72.335 78.245 72.585 78.625 ;
        RECT 70.975 78.045 72.585 78.245 ;
        RECT 70.975 77.955 71.160 78.045 ;
        RECT 71.750 78.035 72.585 78.045 ;
        RECT 72.835 78.015 73.085 78.795 ;
        RECT 73.255 77.945 73.515 78.625 ;
        RECT 73.775 78.125 73.945 78.625 ;
        RECT 74.115 78.295 74.445 78.795 ;
        RECT 73.775 77.955 74.440 78.125 ;
        RECT 71.315 77.845 71.645 77.875 ;
        RECT 71.315 77.785 73.115 77.845 ;
        RECT 70.470 77.675 73.175 77.785 ;
        RECT 70.470 77.615 71.645 77.675 ;
        RECT 72.975 77.640 73.175 77.675 ;
        RECT 70.465 77.235 70.955 77.435 ;
        RECT 71.145 77.235 71.620 77.445 ;
        RECT 66.025 76.805 66.535 76.985 ;
        RECT 66.940 76.895 68.640 77.065 ;
        RECT 66.940 76.805 67.325 76.895 ;
        RECT 66.025 76.415 66.355 76.805 ;
        RECT 66.525 76.465 67.710 76.635 ;
        RECT 67.970 76.245 68.140 76.715 ;
        RECT 68.310 76.430 68.640 76.895 ;
        RECT 68.810 76.245 68.980 77.065 ;
        RECT 69.150 76.425 69.835 77.065 ;
        RECT 70.005 76.245 70.295 76.970 ;
        RECT 70.470 76.245 70.925 77.010 ;
        RECT 71.400 76.835 71.620 77.235 ;
        RECT 71.865 77.235 72.195 77.445 ;
        RECT 71.865 76.835 72.075 77.235 ;
        RECT 72.365 77.200 72.775 77.505 ;
        RECT 73.005 77.065 73.175 77.640 ;
        RECT 72.905 76.945 73.175 77.065 ;
        RECT 72.330 76.900 73.175 76.945 ;
        RECT 72.330 76.775 73.085 76.900 ;
        RECT 72.330 76.625 72.500 76.775 ;
        RECT 73.345 76.755 73.515 77.945 ;
        RECT 73.690 77.135 74.040 77.785 ;
        RECT 74.210 76.965 74.440 77.955 ;
        RECT 73.285 76.745 73.515 76.755 ;
        RECT 71.200 76.415 72.500 76.625 ;
        RECT 72.755 76.245 73.085 76.605 ;
        RECT 73.255 76.415 73.515 76.745 ;
        RECT 73.775 76.795 74.440 76.965 ;
        RECT 73.775 76.505 73.945 76.795 ;
        RECT 74.115 76.245 74.445 76.625 ;
        RECT 74.615 76.505 74.800 78.625 ;
        RECT 75.040 78.335 75.305 78.795 ;
        RECT 75.475 78.200 75.725 78.625 ;
        RECT 75.935 78.350 77.040 78.520 ;
        RECT 75.420 78.070 75.725 78.200 ;
        RECT 74.970 76.875 75.250 77.825 ;
        RECT 75.420 76.965 75.590 78.070 ;
        RECT 75.760 77.285 76.000 77.880 ;
        RECT 76.170 77.815 76.700 78.180 ;
        RECT 76.170 77.115 76.340 77.815 ;
        RECT 76.870 77.735 77.040 78.350 ;
        RECT 77.210 77.995 77.380 78.795 ;
        RECT 77.550 78.295 77.800 78.625 ;
        RECT 78.025 78.325 78.910 78.495 ;
        RECT 76.870 77.645 77.380 77.735 ;
        RECT 75.420 76.835 75.645 76.965 ;
        RECT 75.815 76.895 76.340 77.115 ;
        RECT 76.510 77.475 77.380 77.645 ;
        RECT 75.055 76.245 75.305 76.705 ;
        RECT 75.475 76.695 75.645 76.835 ;
        RECT 76.510 76.695 76.680 77.475 ;
        RECT 77.210 77.405 77.380 77.475 ;
        RECT 76.890 77.225 77.090 77.255 ;
        RECT 77.550 77.225 77.720 78.295 ;
        RECT 77.890 77.405 78.080 78.125 ;
        RECT 76.890 76.925 77.720 77.225 ;
        RECT 78.250 77.195 78.570 78.155 ;
        RECT 75.475 76.525 75.810 76.695 ;
        RECT 76.005 76.525 76.680 76.695 ;
        RECT 77.000 76.245 77.370 76.745 ;
        RECT 77.550 76.695 77.720 76.925 ;
        RECT 78.105 76.865 78.570 77.195 ;
        RECT 78.740 77.485 78.910 78.325 ;
        RECT 79.090 78.295 79.405 78.795 ;
        RECT 79.635 78.065 79.975 78.625 ;
        RECT 79.080 77.690 79.975 78.065 ;
        RECT 80.145 77.785 80.315 78.795 ;
        RECT 79.785 77.485 79.975 77.690 ;
        RECT 80.485 77.735 80.815 78.580 ;
        RECT 81.135 77.865 81.305 78.625 ;
        RECT 81.520 78.035 81.850 78.795 ;
        RECT 80.485 77.655 80.875 77.735 ;
        RECT 81.135 77.695 81.850 77.865 ;
        RECT 82.020 77.720 82.275 78.625 ;
        RECT 80.660 77.605 80.875 77.655 ;
        RECT 78.740 77.155 79.615 77.485 ;
        RECT 79.785 77.155 80.535 77.485 ;
        RECT 78.740 76.695 78.910 77.155 ;
        RECT 79.785 76.985 79.985 77.155 ;
        RECT 80.705 77.025 80.875 77.605 ;
        RECT 81.045 77.145 81.400 77.515 ;
        RECT 81.680 77.485 81.850 77.695 ;
        RECT 81.680 77.155 81.935 77.485 ;
        RECT 80.650 76.985 80.875 77.025 ;
        RECT 77.550 76.525 77.955 76.695 ;
        RECT 78.125 76.525 78.910 76.695 ;
        RECT 79.185 76.245 79.395 76.775 ;
        RECT 79.655 76.460 79.985 76.985 ;
        RECT 80.495 76.900 80.875 76.985 ;
        RECT 81.680 76.965 81.850 77.155 ;
        RECT 82.105 76.990 82.275 77.720 ;
        RECT 82.450 77.645 82.710 78.795 ;
        RECT 82.885 77.705 84.095 78.795 ;
        RECT 82.885 77.165 83.405 77.705 ;
        RECT 80.155 76.245 80.325 76.855 ;
        RECT 80.495 76.465 80.825 76.900 ;
        RECT 81.135 76.795 81.850 76.965 ;
        RECT 81.135 76.415 81.305 76.795 ;
        RECT 81.520 76.245 81.850 76.625 ;
        RECT 82.020 76.415 82.275 76.990 ;
        RECT 82.450 76.245 82.710 77.085 ;
        RECT 83.575 76.995 84.095 77.535 ;
        RECT 82.885 76.245 84.095 76.995 ;
        RECT 5.520 76.075 84.180 76.245 ;
        RECT 5.605 75.325 6.815 76.075 ;
        RECT 7.995 75.525 8.165 75.815 ;
        RECT 8.335 75.695 8.665 76.075 ;
        RECT 7.995 75.355 8.660 75.525 ;
        RECT 5.605 74.785 6.125 75.325 ;
        RECT 6.295 74.615 6.815 75.155 ;
        RECT 5.605 73.525 6.815 74.615 ;
        RECT 7.910 74.535 8.260 75.185 ;
        RECT 8.430 74.365 8.660 75.355 ;
        RECT 7.995 74.195 8.660 74.365 ;
        RECT 7.995 73.695 8.165 74.195 ;
        RECT 8.335 73.525 8.665 74.025 ;
        RECT 8.835 73.695 9.020 75.815 ;
        RECT 9.275 75.615 9.525 76.075 ;
        RECT 9.695 75.625 10.030 75.795 ;
        RECT 10.225 75.625 10.900 75.795 ;
        RECT 9.695 75.485 9.865 75.625 ;
        RECT 9.190 74.495 9.470 75.445 ;
        RECT 9.640 75.355 9.865 75.485 ;
        RECT 9.640 74.250 9.810 75.355 ;
        RECT 10.035 75.205 10.560 75.425 ;
        RECT 9.980 74.440 10.220 75.035 ;
        RECT 10.390 74.505 10.560 75.205 ;
        RECT 10.730 74.845 10.900 75.625 ;
        RECT 11.220 75.575 11.590 76.075 ;
        RECT 11.770 75.625 12.175 75.795 ;
        RECT 12.345 75.625 13.130 75.795 ;
        RECT 11.770 75.395 11.940 75.625 ;
        RECT 11.110 75.095 11.940 75.395 ;
        RECT 12.325 75.125 12.790 75.455 ;
        RECT 11.110 75.065 11.310 75.095 ;
        RECT 11.430 74.845 11.600 74.915 ;
        RECT 10.730 74.675 11.600 74.845 ;
        RECT 11.090 74.585 11.600 74.675 ;
        RECT 9.640 74.120 9.945 74.250 ;
        RECT 10.390 74.140 10.920 74.505 ;
        RECT 9.260 73.525 9.525 73.985 ;
        RECT 9.695 73.695 9.945 74.120 ;
        RECT 11.090 73.970 11.260 74.585 ;
        RECT 10.155 73.800 11.260 73.970 ;
        RECT 11.430 73.525 11.600 74.325 ;
        RECT 11.770 74.025 11.940 75.095 ;
        RECT 12.110 74.195 12.300 74.915 ;
        RECT 12.470 74.165 12.790 75.125 ;
        RECT 12.960 75.165 13.130 75.625 ;
        RECT 13.405 75.545 13.615 76.075 ;
        RECT 13.875 75.335 14.205 75.860 ;
        RECT 14.375 75.465 14.545 76.075 ;
        RECT 14.715 75.420 15.045 75.855 ;
        RECT 14.715 75.335 15.095 75.420 ;
        RECT 14.005 75.165 14.205 75.335 ;
        RECT 14.870 75.295 15.095 75.335 ;
        RECT 12.960 74.835 13.835 75.165 ;
        RECT 14.005 74.835 14.755 75.165 ;
        RECT 11.770 73.695 12.020 74.025 ;
        RECT 12.960 73.995 13.130 74.835 ;
        RECT 14.005 74.630 14.195 74.835 ;
        RECT 14.925 74.715 15.095 75.295 ;
        RECT 15.265 75.305 16.935 76.075 ;
        RECT 15.265 74.785 16.015 75.305 ;
        RECT 17.105 75.255 17.365 76.075 ;
        RECT 17.535 75.255 17.865 75.675 ;
        RECT 18.045 75.505 18.305 75.905 ;
        RECT 18.475 75.675 18.805 76.075 ;
        RECT 18.975 75.505 19.145 75.855 ;
        RECT 19.315 75.675 19.690 76.075 ;
        RECT 18.045 75.335 19.710 75.505 ;
        RECT 19.880 75.400 20.155 75.745 ;
        RECT 17.615 75.165 17.865 75.255 ;
        RECT 19.540 75.165 19.710 75.335 ;
        RECT 14.880 74.665 15.095 74.715 ;
        RECT 13.300 74.255 14.195 74.630 ;
        RECT 14.705 74.585 15.095 74.665 ;
        RECT 16.185 74.615 16.935 75.135 ;
        RECT 17.110 74.835 17.445 75.085 ;
        RECT 17.615 74.835 18.330 75.165 ;
        RECT 18.545 74.835 19.370 75.165 ;
        RECT 19.540 74.835 19.815 75.165 ;
        RECT 12.245 73.825 13.130 73.995 ;
        RECT 13.310 73.525 13.625 74.025 ;
        RECT 13.855 73.695 14.195 74.255 ;
        RECT 14.365 73.525 14.535 74.535 ;
        RECT 14.705 73.740 15.035 74.585 ;
        RECT 15.265 73.525 16.935 74.615 ;
        RECT 17.105 73.525 17.365 74.665 ;
        RECT 17.615 74.275 17.785 74.835 ;
        RECT 18.045 74.375 18.375 74.665 ;
        RECT 18.545 74.545 18.790 74.835 ;
        RECT 19.540 74.665 19.710 74.835 ;
        RECT 19.985 74.665 20.155 75.400 ;
        RECT 20.875 75.525 21.045 75.815 ;
        RECT 21.215 75.695 21.545 76.075 ;
        RECT 20.875 75.355 21.540 75.525 ;
        RECT 19.050 74.495 19.710 74.665 ;
        RECT 19.050 74.375 19.220 74.495 ;
        RECT 18.045 74.205 19.220 74.375 ;
        RECT 17.605 73.705 19.220 74.035 ;
        RECT 19.390 73.525 19.670 74.325 ;
        RECT 19.880 73.695 20.155 74.665 ;
        RECT 20.790 74.535 21.140 75.185 ;
        RECT 21.310 74.365 21.540 75.355 ;
        RECT 20.875 74.195 21.540 74.365 ;
        RECT 20.875 73.695 21.045 74.195 ;
        RECT 21.215 73.525 21.545 74.025 ;
        RECT 21.715 73.695 21.900 75.815 ;
        RECT 22.155 75.615 22.405 76.075 ;
        RECT 22.575 75.625 22.910 75.795 ;
        RECT 23.105 75.625 23.780 75.795 ;
        RECT 22.575 75.485 22.745 75.625 ;
        RECT 22.070 74.495 22.350 75.445 ;
        RECT 22.520 75.355 22.745 75.485 ;
        RECT 22.520 74.250 22.690 75.355 ;
        RECT 22.915 75.205 23.440 75.425 ;
        RECT 22.860 74.440 23.100 75.035 ;
        RECT 23.270 74.505 23.440 75.205 ;
        RECT 23.610 74.845 23.780 75.625 ;
        RECT 24.100 75.575 24.470 76.075 ;
        RECT 24.650 75.625 25.055 75.795 ;
        RECT 25.225 75.625 26.010 75.795 ;
        RECT 24.650 75.395 24.820 75.625 ;
        RECT 23.990 75.095 24.820 75.395 ;
        RECT 25.205 75.125 25.670 75.455 ;
        RECT 23.990 75.065 24.190 75.095 ;
        RECT 24.310 74.845 24.480 74.915 ;
        RECT 23.610 74.675 24.480 74.845 ;
        RECT 23.970 74.585 24.480 74.675 ;
        RECT 22.520 74.120 22.825 74.250 ;
        RECT 23.270 74.140 23.800 74.505 ;
        RECT 22.140 73.525 22.405 73.985 ;
        RECT 22.575 73.695 22.825 74.120 ;
        RECT 23.970 73.970 24.140 74.585 ;
        RECT 23.035 73.800 24.140 73.970 ;
        RECT 24.310 73.525 24.480 74.325 ;
        RECT 24.650 74.025 24.820 75.095 ;
        RECT 24.990 74.195 25.180 74.915 ;
        RECT 25.350 74.165 25.670 75.125 ;
        RECT 25.840 75.165 26.010 75.625 ;
        RECT 26.285 75.545 26.495 76.075 ;
        RECT 26.755 75.335 27.085 75.860 ;
        RECT 27.255 75.465 27.425 76.075 ;
        RECT 27.595 75.420 27.925 75.855 ;
        RECT 28.095 75.560 28.265 76.075 ;
        RECT 27.595 75.335 27.975 75.420 ;
        RECT 26.885 75.165 27.085 75.335 ;
        RECT 27.750 75.295 27.975 75.335 ;
        RECT 25.840 74.835 26.715 75.165 ;
        RECT 26.885 74.835 27.635 75.165 ;
        RECT 24.650 73.695 24.900 74.025 ;
        RECT 25.840 73.995 26.010 74.835 ;
        RECT 26.885 74.630 27.075 74.835 ;
        RECT 27.805 74.715 27.975 75.295 ;
        RECT 28.605 75.305 31.195 76.075 ;
        RECT 31.365 75.350 31.655 76.075 ;
        RECT 31.915 75.525 32.085 75.815 ;
        RECT 32.255 75.695 32.585 76.075 ;
        RECT 31.915 75.355 32.580 75.525 ;
        RECT 28.605 74.785 29.815 75.305 ;
        RECT 27.760 74.665 27.975 74.715 ;
        RECT 26.180 74.255 27.075 74.630 ;
        RECT 27.585 74.585 27.975 74.665 ;
        RECT 29.985 74.615 31.195 75.135 ;
        RECT 25.125 73.825 26.010 73.995 ;
        RECT 26.190 73.525 26.505 74.025 ;
        RECT 26.735 73.695 27.075 74.255 ;
        RECT 27.245 73.525 27.415 74.535 ;
        RECT 27.585 73.740 27.915 74.585 ;
        RECT 28.085 73.525 28.255 74.440 ;
        RECT 28.605 73.525 31.195 74.615 ;
        RECT 31.365 73.525 31.655 74.690 ;
        RECT 31.830 74.535 32.180 75.185 ;
        RECT 32.350 74.365 32.580 75.355 ;
        RECT 31.915 74.195 32.580 74.365 ;
        RECT 31.915 73.695 32.085 74.195 ;
        RECT 32.255 73.525 32.585 74.025 ;
        RECT 32.755 73.695 32.940 75.815 ;
        RECT 33.195 75.615 33.445 76.075 ;
        RECT 33.615 75.625 33.950 75.795 ;
        RECT 34.145 75.625 34.820 75.795 ;
        RECT 33.615 75.485 33.785 75.625 ;
        RECT 33.110 74.495 33.390 75.445 ;
        RECT 33.560 75.355 33.785 75.485 ;
        RECT 33.560 74.250 33.730 75.355 ;
        RECT 33.955 75.205 34.480 75.425 ;
        RECT 33.900 74.440 34.140 75.035 ;
        RECT 34.310 74.505 34.480 75.205 ;
        RECT 34.650 74.845 34.820 75.625 ;
        RECT 35.140 75.575 35.510 76.075 ;
        RECT 35.690 75.625 36.095 75.795 ;
        RECT 36.265 75.625 37.050 75.795 ;
        RECT 35.690 75.395 35.860 75.625 ;
        RECT 35.030 75.095 35.860 75.395 ;
        RECT 36.245 75.125 36.710 75.455 ;
        RECT 35.030 75.065 35.230 75.095 ;
        RECT 35.350 74.845 35.520 74.915 ;
        RECT 34.650 74.675 35.520 74.845 ;
        RECT 35.010 74.585 35.520 74.675 ;
        RECT 33.560 74.120 33.865 74.250 ;
        RECT 34.310 74.140 34.840 74.505 ;
        RECT 33.180 73.525 33.445 73.985 ;
        RECT 33.615 73.695 33.865 74.120 ;
        RECT 35.010 73.970 35.180 74.585 ;
        RECT 34.075 73.800 35.180 73.970 ;
        RECT 35.350 73.525 35.520 74.325 ;
        RECT 35.690 74.025 35.860 75.095 ;
        RECT 36.030 74.195 36.220 74.915 ;
        RECT 36.390 74.165 36.710 75.125 ;
        RECT 36.880 75.165 37.050 75.625 ;
        RECT 37.325 75.545 37.535 76.075 ;
        RECT 37.795 75.335 38.125 75.860 ;
        RECT 38.295 75.465 38.465 76.075 ;
        RECT 38.635 75.420 38.965 75.855 ;
        RECT 39.695 75.420 40.025 75.855 ;
        RECT 40.195 75.465 40.365 76.075 ;
        RECT 38.635 75.335 39.015 75.420 ;
        RECT 37.925 75.165 38.125 75.335 ;
        RECT 38.790 75.295 39.015 75.335 ;
        RECT 36.880 74.835 37.755 75.165 ;
        RECT 37.925 74.835 38.675 75.165 ;
        RECT 35.690 73.695 35.940 74.025 ;
        RECT 36.880 73.995 37.050 74.835 ;
        RECT 37.925 74.630 38.115 74.835 ;
        RECT 38.845 74.715 39.015 75.295 ;
        RECT 38.800 74.665 39.015 74.715 ;
        RECT 37.220 74.255 38.115 74.630 ;
        RECT 38.625 74.585 39.015 74.665 ;
        RECT 39.645 75.335 40.025 75.420 ;
        RECT 40.535 75.335 40.865 75.860 ;
        RECT 41.125 75.545 41.335 76.075 ;
        RECT 41.610 75.625 42.395 75.795 ;
        RECT 42.565 75.625 42.970 75.795 ;
        RECT 39.645 75.295 39.870 75.335 ;
        RECT 39.645 74.715 39.815 75.295 ;
        RECT 40.535 75.165 40.735 75.335 ;
        RECT 41.610 75.165 41.780 75.625 ;
        RECT 39.985 74.835 40.735 75.165 ;
        RECT 40.905 74.835 41.780 75.165 ;
        RECT 39.645 74.665 39.860 74.715 ;
        RECT 39.645 74.585 40.035 74.665 ;
        RECT 36.165 73.825 37.050 73.995 ;
        RECT 37.230 73.525 37.545 74.025 ;
        RECT 37.775 73.695 38.115 74.255 ;
        RECT 38.285 73.525 38.455 74.535 ;
        RECT 38.625 73.740 38.955 74.585 ;
        RECT 39.705 73.740 40.035 74.585 ;
        RECT 40.545 74.630 40.735 74.835 ;
        RECT 40.205 73.525 40.375 74.535 ;
        RECT 40.545 74.255 41.440 74.630 ;
        RECT 40.545 73.695 40.885 74.255 ;
        RECT 41.115 73.525 41.430 74.025 ;
        RECT 41.610 73.995 41.780 74.835 ;
        RECT 41.950 75.125 42.415 75.455 ;
        RECT 42.800 75.395 42.970 75.625 ;
        RECT 43.150 75.575 43.520 76.075 ;
        RECT 43.840 75.625 44.515 75.795 ;
        RECT 44.710 75.625 45.045 75.795 ;
        RECT 41.950 74.165 42.270 75.125 ;
        RECT 42.800 75.095 43.630 75.395 ;
        RECT 42.440 74.195 42.630 74.915 ;
        RECT 42.800 74.025 42.970 75.095 ;
        RECT 43.430 75.065 43.630 75.095 ;
        RECT 43.140 74.845 43.310 74.915 ;
        RECT 43.840 74.845 44.010 75.625 ;
        RECT 44.875 75.485 45.045 75.625 ;
        RECT 45.215 75.615 45.465 76.075 ;
        RECT 43.140 74.675 44.010 74.845 ;
        RECT 44.180 75.205 44.705 75.425 ;
        RECT 44.875 75.355 45.100 75.485 ;
        RECT 43.140 74.585 43.650 74.675 ;
        RECT 41.610 73.825 42.495 73.995 ;
        RECT 42.720 73.695 42.970 74.025 ;
        RECT 43.140 73.525 43.310 74.325 ;
        RECT 43.480 73.970 43.650 74.585 ;
        RECT 44.180 74.505 44.350 75.205 ;
        RECT 43.820 74.140 44.350 74.505 ;
        RECT 44.520 74.440 44.760 75.035 ;
        RECT 44.930 74.250 45.100 75.355 ;
        RECT 45.270 74.495 45.550 75.445 ;
        RECT 44.795 74.120 45.100 74.250 ;
        RECT 43.480 73.800 44.585 73.970 ;
        RECT 44.795 73.695 45.045 74.120 ;
        RECT 45.215 73.525 45.480 73.985 ;
        RECT 45.720 73.695 45.905 75.815 ;
        RECT 46.075 75.695 46.405 76.075 ;
        RECT 46.575 75.525 46.745 75.815 ;
        RECT 46.080 75.355 46.745 75.525 ;
        RECT 46.080 74.365 46.310 75.355 ;
        RECT 47.005 75.305 49.595 76.075 ;
        RECT 49.815 75.420 50.145 75.855 ;
        RECT 50.315 75.465 50.485 76.075 ;
        RECT 49.765 75.335 50.145 75.420 ;
        RECT 50.655 75.335 50.985 75.860 ;
        RECT 51.245 75.545 51.455 76.075 ;
        RECT 51.730 75.625 52.515 75.795 ;
        RECT 52.685 75.625 53.090 75.795 ;
        RECT 46.480 74.535 46.830 75.185 ;
        RECT 47.005 74.785 48.215 75.305 ;
        RECT 49.765 75.295 49.990 75.335 ;
        RECT 48.385 74.615 49.595 75.135 ;
        RECT 46.080 74.195 46.745 74.365 ;
        RECT 46.075 73.525 46.405 74.025 ;
        RECT 46.575 73.695 46.745 74.195 ;
        RECT 47.005 73.525 49.595 74.615 ;
        RECT 49.765 74.715 49.935 75.295 ;
        RECT 50.655 75.165 50.855 75.335 ;
        RECT 51.730 75.165 51.900 75.625 ;
        RECT 50.105 74.835 50.855 75.165 ;
        RECT 51.025 74.835 51.900 75.165 ;
        RECT 49.765 74.665 49.980 74.715 ;
        RECT 49.765 74.585 50.155 74.665 ;
        RECT 49.825 73.740 50.155 74.585 ;
        RECT 50.665 74.630 50.855 74.835 ;
        RECT 50.325 73.525 50.495 74.535 ;
        RECT 50.665 74.255 51.560 74.630 ;
        RECT 50.665 73.695 51.005 74.255 ;
        RECT 51.235 73.525 51.550 74.025 ;
        RECT 51.730 73.995 51.900 74.835 ;
        RECT 52.070 75.125 52.535 75.455 ;
        RECT 52.920 75.395 53.090 75.625 ;
        RECT 53.270 75.575 53.640 76.075 ;
        RECT 53.960 75.625 54.635 75.795 ;
        RECT 54.830 75.625 55.165 75.795 ;
        RECT 52.070 74.165 52.390 75.125 ;
        RECT 52.920 75.095 53.750 75.395 ;
        RECT 52.560 74.195 52.750 74.915 ;
        RECT 52.920 74.025 53.090 75.095 ;
        RECT 53.550 75.065 53.750 75.095 ;
        RECT 53.260 74.845 53.430 74.915 ;
        RECT 53.960 74.845 54.130 75.625 ;
        RECT 54.995 75.485 55.165 75.625 ;
        RECT 55.335 75.615 55.585 76.075 ;
        RECT 53.260 74.675 54.130 74.845 ;
        RECT 54.300 75.205 54.825 75.425 ;
        RECT 54.995 75.355 55.220 75.485 ;
        RECT 53.260 74.585 53.770 74.675 ;
        RECT 51.730 73.825 52.615 73.995 ;
        RECT 52.840 73.695 53.090 74.025 ;
        RECT 53.260 73.525 53.430 74.325 ;
        RECT 53.600 73.970 53.770 74.585 ;
        RECT 54.300 74.505 54.470 75.205 ;
        RECT 53.940 74.140 54.470 74.505 ;
        RECT 54.640 74.440 54.880 75.035 ;
        RECT 55.050 74.250 55.220 75.355 ;
        RECT 55.390 74.495 55.670 75.445 ;
        RECT 54.915 74.120 55.220 74.250 ;
        RECT 53.600 73.800 54.705 73.970 ;
        RECT 54.915 73.695 55.165 74.120 ;
        RECT 55.335 73.525 55.600 73.985 ;
        RECT 55.840 73.695 56.025 75.815 ;
        RECT 56.195 75.695 56.525 76.075 ;
        RECT 56.695 75.525 56.865 75.815 ;
        RECT 56.200 75.355 56.865 75.525 ;
        RECT 56.200 74.365 56.430 75.355 ;
        RECT 57.125 75.350 57.415 76.075 ;
        RECT 57.585 75.335 58.025 75.895 ;
        RECT 58.195 75.335 58.645 76.075 ;
        RECT 58.815 75.505 58.985 75.905 ;
        RECT 59.155 75.675 59.575 76.075 ;
        RECT 59.745 75.505 59.975 75.905 ;
        RECT 58.815 75.335 59.975 75.505 ;
        RECT 60.145 75.335 60.635 75.905 ;
        RECT 56.600 74.535 56.950 75.185 ;
        RECT 56.200 74.195 56.865 74.365 ;
        RECT 56.195 73.525 56.525 74.025 ;
        RECT 56.695 73.695 56.865 74.195 ;
        RECT 57.125 73.525 57.415 74.690 ;
        RECT 57.585 74.325 57.895 75.335 ;
        RECT 58.065 74.715 58.235 75.165 ;
        RECT 58.405 74.885 58.795 75.165 ;
        RECT 58.980 74.835 59.225 75.165 ;
        RECT 58.065 74.545 58.855 74.715 ;
        RECT 57.585 73.695 58.025 74.325 ;
        RECT 58.200 73.525 58.515 74.375 ;
        RECT 58.685 73.865 58.855 74.545 ;
        RECT 59.025 74.035 59.225 74.835 ;
        RECT 59.425 74.035 59.675 75.165 ;
        RECT 59.890 74.835 60.295 75.165 ;
        RECT 60.465 74.665 60.635 75.335 ;
        RECT 59.865 74.495 60.635 74.665 ;
        RECT 60.815 75.350 61.145 75.860 ;
        RECT 61.315 75.675 61.645 76.075 ;
        RECT 62.695 75.505 63.025 75.845 ;
        RECT 63.195 75.675 63.525 76.075 ;
        RECT 60.815 74.715 61.005 75.350 ;
        RECT 61.315 75.335 63.680 75.505 ;
        RECT 64.965 75.345 65.255 76.075 ;
        RECT 61.315 75.165 61.485 75.335 ;
        RECT 61.175 74.835 61.485 75.165 ;
        RECT 61.655 74.835 61.960 75.165 ;
        RECT 60.815 74.585 61.035 74.715 ;
        RECT 59.865 73.865 60.115 74.495 ;
        RECT 58.685 73.695 60.115 73.865 ;
        RECT 60.295 73.525 60.625 74.325 ;
        RECT 60.815 73.735 61.145 74.585 ;
        RECT 61.315 73.525 61.565 74.665 ;
        RECT 61.745 74.505 61.960 74.835 ;
        RECT 62.135 74.505 62.420 75.165 ;
        RECT 62.615 74.505 62.880 75.165 ;
        RECT 63.095 74.505 63.340 75.165 ;
        RECT 63.510 74.335 63.680 75.335 ;
        RECT 64.955 74.835 65.255 75.165 ;
        RECT 65.435 75.145 65.665 75.785 ;
        RECT 65.845 75.525 66.155 75.895 ;
        RECT 66.335 75.705 67.005 76.075 ;
        RECT 65.845 75.325 67.075 75.525 ;
        RECT 65.435 74.835 65.960 75.145 ;
        RECT 66.140 74.835 66.605 75.145 ;
        RECT 66.785 74.655 67.075 75.325 ;
        RECT 61.755 74.165 63.045 74.335 ;
        RECT 61.755 73.745 62.005 74.165 ;
        RECT 62.235 73.525 62.565 73.995 ;
        RECT 62.795 73.745 63.045 74.165 ;
        RECT 63.225 74.165 63.680 74.335 ;
        RECT 64.965 74.415 66.125 74.655 ;
        RECT 63.225 73.735 63.555 74.165 ;
        RECT 64.965 73.705 65.225 74.415 ;
        RECT 65.395 73.525 65.725 74.235 ;
        RECT 65.895 73.705 66.125 74.415 ;
        RECT 66.305 74.435 67.075 74.655 ;
        RECT 66.305 73.705 66.575 74.435 ;
        RECT 66.755 73.525 67.095 74.255 ;
        RECT 67.265 73.705 67.525 75.895 ;
        RECT 67.725 75.345 68.015 76.075 ;
        RECT 67.715 74.835 68.015 75.165 ;
        RECT 68.195 75.145 68.425 75.785 ;
        RECT 68.605 75.525 68.915 75.895 ;
        RECT 69.095 75.705 69.765 76.075 ;
        RECT 68.605 75.325 69.835 75.525 ;
        RECT 68.195 74.835 68.720 75.145 ;
        RECT 68.900 74.835 69.365 75.145 ;
        RECT 69.545 74.655 69.835 75.325 ;
        RECT 67.725 74.415 68.885 74.655 ;
        RECT 67.725 73.705 67.985 74.415 ;
        RECT 68.155 73.525 68.485 74.235 ;
        RECT 68.655 73.705 68.885 74.415 ;
        RECT 69.065 74.435 69.835 74.655 ;
        RECT 69.065 73.705 69.335 74.435 ;
        RECT 69.515 73.525 69.855 74.255 ;
        RECT 70.025 73.705 70.285 75.895 ;
        RECT 70.465 75.305 73.975 76.075 ;
        RECT 74.145 75.325 75.355 76.075 ;
        RECT 75.530 75.335 75.785 75.905 ;
        RECT 75.955 75.675 76.285 76.075 ;
        RECT 76.710 75.540 77.240 75.905 ;
        RECT 77.430 75.735 77.705 75.905 ;
        RECT 77.425 75.565 77.705 75.735 ;
        RECT 76.710 75.505 76.885 75.540 ;
        RECT 75.955 75.335 76.885 75.505 ;
        RECT 70.465 74.785 72.115 75.305 ;
        RECT 72.285 74.615 73.975 75.135 ;
        RECT 74.145 74.785 74.665 75.325 ;
        RECT 74.835 74.615 75.355 75.155 ;
        RECT 70.465 73.525 73.975 74.615 ;
        RECT 74.145 73.525 75.355 74.615 ;
        RECT 75.530 74.665 75.700 75.335 ;
        RECT 75.955 75.165 76.125 75.335 ;
        RECT 75.870 74.835 76.125 75.165 ;
        RECT 76.350 74.835 76.545 75.165 ;
        RECT 75.530 73.695 75.865 74.665 ;
        RECT 76.035 73.525 76.205 74.665 ;
        RECT 76.375 73.865 76.545 74.835 ;
        RECT 76.715 74.205 76.885 75.335 ;
        RECT 77.055 74.545 77.225 75.345 ;
        RECT 77.430 74.745 77.705 75.565 ;
        RECT 77.875 74.545 78.065 75.905 ;
        RECT 78.245 75.540 78.755 76.075 ;
        RECT 78.975 75.265 79.220 75.870 ;
        RECT 79.755 75.525 79.925 75.905 ;
        RECT 80.105 75.695 80.435 76.075 ;
        RECT 79.755 75.355 80.420 75.525 ;
        RECT 80.615 75.400 80.875 75.905 ;
        RECT 78.265 75.095 79.495 75.265 ;
        RECT 77.055 74.375 78.065 74.545 ;
        RECT 78.235 74.530 78.985 74.720 ;
        RECT 76.715 74.035 77.840 74.205 ;
        RECT 78.235 73.865 78.405 74.530 ;
        RECT 79.155 74.285 79.495 75.095 ;
        RECT 79.685 74.805 80.015 75.175 ;
        RECT 80.250 75.100 80.420 75.355 ;
        RECT 80.250 74.770 80.535 75.100 ;
        RECT 80.250 74.625 80.420 74.770 ;
        RECT 76.375 73.695 78.405 73.865 ;
        RECT 78.575 73.525 78.745 74.285 ;
        RECT 78.980 73.875 79.495 74.285 ;
        RECT 79.755 74.455 80.420 74.625 ;
        RECT 80.705 74.600 80.875 75.400 ;
        RECT 81.045 75.305 82.715 76.075 ;
        RECT 82.885 75.325 84.095 76.075 ;
        RECT 81.045 74.785 81.795 75.305 ;
        RECT 81.965 74.615 82.715 75.135 ;
        RECT 79.755 73.695 79.925 74.455 ;
        RECT 80.105 73.525 80.435 74.285 ;
        RECT 80.605 73.695 80.875 74.600 ;
        RECT 81.045 73.525 82.715 74.615 ;
        RECT 82.885 74.615 83.405 75.155 ;
        RECT 83.575 74.785 84.095 75.325 ;
        RECT 82.885 73.525 84.095 74.615 ;
        RECT 5.520 73.355 84.180 73.525 ;
        RECT 5.605 72.265 6.815 73.355 ;
        RECT 6.985 72.265 8.655 73.355 ;
        RECT 5.605 71.555 6.125 72.095 ;
        RECT 6.295 71.725 6.815 72.265 ;
        RECT 6.985 71.575 7.735 72.095 ;
        RECT 7.905 71.745 8.655 72.265 ;
        RECT 8.860 72.565 9.395 73.185 ;
        RECT 5.605 70.805 6.815 71.555 ;
        RECT 6.985 70.805 8.655 71.575 ;
        RECT 8.860 71.545 9.175 72.565 ;
        RECT 9.565 72.555 9.895 73.355 ;
        RECT 11.585 72.845 11.845 73.355 ;
        RECT 10.380 72.385 10.770 72.560 ;
        RECT 9.345 72.215 10.770 72.385 ;
        RECT 9.345 71.715 9.515 72.215 ;
        RECT 8.860 70.975 9.475 71.545 ;
        RECT 9.765 71.485 10.030 72.045 ;
        RECT 10.200 71.315 10.370 72.215 ;
        RECT 10.540 71.485 10.895 72.045 ;
        RECT 11.585 71.795 11.925 72.675 ;
        RECT 12.095 71.965 12.265 73.185 ;
        RECT 12.505 72.850 13.120 73.355 ;
        RECT 12.505 72.315 12.755 72.680 ;
        RECT 12.925 72.675 13.120 72.850 ;
        RECT 13.290 72.845 13.765 73.185 ;
        RECT 13.935 72.810 14.150 73.355 ;
        RECT 12.925 72.485 13.255 72.675 ;
        RECT 13.475 72.315 14.190 72.610 ;
        RECT 14.360 72.485 14.635 73.185 ;
        RECT 12.505 72.145 14.295 72.315 ;
        RECT 12.095 71.715 12.890 71.965 ;
        RECT 12.095 71.625 12.345 71.715 ;
        RECT 9.645 70.805 9.860 71.315 ;
        RECT 10.090 70.985 10.370 71.315 ;
        RECT 10.550 70.805 10.790 71.315 ;
        RECT 11.585 70.805 11.845 71.625 ;
        RECT 12.015 71.205 12.345 71.625 ;
        RECT 13.060 71.290 13.315 72.145 ;
        RECT 12.525 71.025 13.315 71.290 ;
        RECT 13.485 71.445 13.895 71.965 ;
        RECT 14.065 71.715 14.295 72.145 ;
        RECT 14.465 71.455 14.635 72.485 ;
        RECT 15.265 72.215 15.525 73.355 ;
        RECT 15.765 72.845 17.380 73.175 ;
        RECT 15.775 72.045 15.945 72.605 ;
        RECT 16.205 72.505 17.380 72.675 ;
        RECT 17.550 72.555 17.830 73.355 ;
        RECT 16.205 72.215 16.535 72.505 ;
        RECT 17.210 72.385 17.380 72.505 ;
        RECT 16.705 72.045 16.950 72.335 ;
        RECT 17.210 72.215 17.870 72.385 ;
        RECT 18.040 72.215 18.315 73.185 ;
        RECT 17.700 72.045 17.870 72.215 ;
        RECT 15.270 71.795 15.605 72.045 ;
        RECT 15.775 71.715 16.490 72.045 ;
        RECT 16.705 71.715 17.530 72.045 ;
        RECT 17.700 71.715 17.975 72.045 ;
        RECT 15.775 71.625 16.025 71.715 ;
        RECT 13.485 71.025 13.685 71.445 ;
        RECT 13.875 70.805 14.205 71.265 ;
        RECT 14.375 70.975 14.635 71.455 ;
        RECT 15.265 70.805 15.525 71.625 ;
        RECT 15.695 71.205 16.025 71.625 ;
        RECT 17.700 71.545 17.870 71.715 ;
        RECT 16.205 71.375 17.870 71.545 ;
        RECT 18.145 71.480 18.315 72.215 ;
        RECT 18.485 72.190 18.775 73.355 ;
        RECT 18.945 72.265 20.615 73.355 ;
        RECT 21.335 72.685 21.505 73.185 ;
        RECT 21.675 72.855 22.005 73.355 ;
        RECT 21.335 72.515 22.000 72.685 ;
        RECT 18.945 71.575 19.695 72.095 ;
        RECT 19.865 71.745 20.615 72.265 ;
        RECT 21.250 71.695 21.600 72.345 ;
        RECT 16.205 70.975 16.465 71.375 ;
        RECT 16.635 70.805 16.965 71.205 ;
        RECT 17.135 71.025 17.305 71.375 ;
        RECT 17.475 70.805 17.850 71.205 ;
        RECT 18.040 71.135 18.315 71.480 ;
        RECT 18.485 70.805 18.775 71.530 ;
        RECT 18.945 70.805 20.615 71.575 ;
        RECT 21.770 71.525 22.000 72.515 ;
        RECT 21.335 71.355 22.000 71.525 ;
        RECT 21.335 71.065 21.505 71.355 ;
        RECT 21.675 70.805 22.005 71.185 ;
        RECT 22.175 71.065 22.360 73.185 ;
        RECT 22.600 72.895 22.865 73.355 ;
        RECT 23.035 72.760 23.285 73.185 ;
        RECT 23.495 72.910 24.600 73.080 ;
        RECT 22.980 72.630 23.285 72.760 ;
        RECT 22.530 71.435 22.810 72.385 ;
        RECT 22.980 71.525 23.150 72.630 ;
        RECT 23.320 71.845 23.560 72.440 ;
        RECT 23.730 72.375 24.260 72.740 ;
        RECT 23.730 71.675 23.900 72.375 ;
        RECT 24.430 72.295 24.600 72.910 ;
        RECT 24.770 72.555 24.940 73.355 ;
        RECT 25.110 72.855 25.360 73.185 ;
        RECT 25.585 72.885 26.470 73.055 ;
        RECT 24.430 72.205 24.940 72.295 ;
        RECT 22.980 71.395 23.205 71.525 ;
        RECT 23.375 71.455 23.900 71.675 ;
        RECT 24.070 72.035 24.940 72.205 ;
        RECT 22.615 70.805 22.865 71.265 ;
        RECT 23.035 71.255 23.205 71.395 ;
        RECT 24.070 71.255 24.240 72.035 ;
        RECT 24.770 71.965 24.940 72.035 ;
        RECT 24.450 71.785 24.650 71.815 ;
        RECT 25.110 71.785 25.280 72.855 ;
        RECT 25.450 71.965 25.640 72.685 ;
        RECT 24.450 71.485 25.280 71.785 ;
        RECT 25.810 71.755 26.130 72.715 ;
        RECT 23.035 71.085 23.370 71.255 ;
        RECT 23.565 71.085 24.240 71.255 ;
        RECT 24.560 70.805 24.930 71.305 ;
        RECT 25.110 71.255 25.280 71.485 ;
        RECT 25.665 71.425 26.130 71.755 ;
        RECT 26.300 72.045 26.470 72.885 ;
        RECT 26.650 72.855 26.965 73.355 ;
        RECT 27.195 72.625 27.535 73.185 ;
        RECT 26.640 72.250 27.535 72.625 ;
        RECT 27.705 72.345 27.875 73.355 ;
        RECT 27.345 72.045 27.535 72.250 ;
        RECT 28.045 72.295 28.375 73.140 ;
        RECT 28.545 72.440 28.715 73.355 ;
        RECT 28.045 72.215 28.435 72.295 ;
        RECT 29.065 72.265 32.575 73.355 ;
        RECT 28.220 72.165 28.435 72.215 ;
        RECT 26.300 71.715 27.175 72.045 ;
        RECT 27.345 71.715 28.095 72.045 ;
        RECT 26.300 71.255 26.470 71.715 ;
        RECT 27.345 71.545 27.545 71.715 ;
        RECT 28.265 71.585 28.435 72.165 ;
        RECT 28.210 71.545 28.435 71.585 ;
        RECT 25.110 71.085 25.515 71.255 ;
        RECT 25.685 71.085 26.470 71.255 ;
        RECT 26.745 70.805 26.955 71.335 ;
        RECT 27.215 71.020 27.545 71.545 ;
        RECT 28.055 71.460 28.435 71.545 ;
        RECT 29.065 71.575 30.715 72.095 ;
        RECT 30.885 71.745 32.575 72.265 ;
        RECT 32.815 72.350 33.070 73.155 ;
        RECT 33.240 72.520 33.500 73.355 ;
        RECT 33.670 72.350 33.930 73.155 ;
        RECT 34.100 72.520 34.355 73.355 ;
        RECT 32.815 72.180 34.415 72.350 ;
        RECT 32.745 71.785 33.965 72.010 ;
        RECT 34.135 71.615 34.415 72.180 ;
        RECT 27.715 70.805 27.885 71.415 ;
        RECT 28.055 71.025 28.385 71.460 ;
        RECT 28.555 70.805 28.725 71.320 ;
        RECT 29.065 70.805 32.575 71.575 ;
        RECT 33.685 71.445 34.415 71.615 ;
        RECT 34.590 72.215 34.925 73.185 ;
        RECT 35.095 72.215 35.265 73.355 ;
        RECT 35.435 73.015 37.465 73.185 ;
        RECT 34.590 71.545 34.760 72.215 ;
        RECT 35.435 72.045 35.605 73.015 ;
        RECT 34.930 71.715 35.185 72.045 ;
        RECT 35.410 71.715 35.605 72.045 ;
        RECT 35.775 72.675 36.900 72.845 ;
        RECT 35.015 71.545 35.185 71.715 ;
        RECT 35.775 71.545 35.945 72.675 ;
        RECT 33.220 70.805 33.515 71.330 ;
        RECT 33.685 71.000 33.910 71.445 ;
        RECT 34.080 70.805 34.410 71.275 ;
        RECT 34.590 70.975 34.845 71.545 ;
        RECT 35.015 71.375 35.945 71.545 ;
        RECT 36.115 72.335 37.125 72.505 ;
        RECT 36.115 71.535 36.285 72.335 ;
        RECT 35.770 71.340 35.945 71.375 ;
        RECT 35.015 70.805 35.345 71.205 ;
        RECT 35.770 70.975 36.300 71.340 ;
        RECT 36.490 71.315 36.765 72.135 ;
        RECT 36.485 71.145 36.765 71.315 ;
        RECT 36.490 70.975 36.765 71.145 ;
        RECT 36.935 70.975 37.125 72.335 ;
        RECT 37.295 72.350 37.465 73.015 ;
        RECT 37.635 72.595 37.805 73.355 ;
        RECT 38.040 72.595 38.555 73.005 ;
        RECT 37.295 72.160 38.045 72.350 ;
        RECT 38.215 71.785 38.555 72.595 ;
        RECT 37.325 71.615 38.555 71.785 ;
        RECT 38.730 72.215 39.065 73.185 ;
        RECT 39.235 72.215 39.405 73.355 ;
        RECT 39.575 73.015 41.605 73.185 ;
        RECT 37.305 70.805 37.815 71.340 ;
        RECT 38.035 71.010 38.280 71.615 ;
        RECT 38.730 71.545 38.900 72.215 ;
        RECT 39.575 72.045 39.745 73.015 ;
        RECT 39.070 71.715 39.325 72.045 ;
        RECT 39.550 71.715 39.745 72.045 ;
        RECT 39.915 72.675 41.040 72.845 ;
        RECT 39.155 71.545 39.325 71.715 ;
        RECT 39.915 71.545 40.085 72.675 ;
        RECT 38.730 70.975 38.985 71.545 ;
        RECT 39.155 71.375 40.085 71.545 ;
        RECT 40.255 72.335 41.265 72.505 ;
        RECT 40.255 71.535 40.425 72.335 ;
        RECT 39.910 71.340 40.085 71.375 ;
        RECT 39.155 70.805 39.485 71.205 ;
        RECT 39.910 70.975 40.440 71.340 ;
        RECT 40.630 71.315 40.905 72.135 ;
        RECT 40.625 71.145 40.905 71.315 ;
        RECT 40.630 70.975 40.905 71.145 ;
        RECT 41.075 70.975 41.265 72.335 ;
        RECT 41.435 72.350 41.605 73.015 ;
        RECT 41.775 72.595 41.945 73.355 ;
        RECT 42.180 72.595 42.695 73.005 ;
        RECT 41.435 72.160 42.185 72.350 ;
        RECT 42.355 71.785 42.695 72.595 ;
        RECT 42.865 72.265 44.075 73.355 ;
        RECT 41.465 71.615 42.695 71.785 ;
        RECT 41.445 70.805 41.955 71.340 ;
        RECT 42.175 71.010 42.420 71.615 ;
        RECT 42.865 71.555 43.385 72.095 ;
        RECT 43.555 71.725 44.075 72.265 ;
        RECT 44.245 72.190 44.535 73.355 ;
        RECT 44.710 72.215 45.045 73.185 ;
        RECT 45.215 72.215 45.385 73.355 ;
        RECT 45.555 73.015 47.585 73.185 ;
        RECT 42.865 70.805 44.075 71.555 ;
        RECT 44.710 71.545 44.880 72.215 ;
        RECT 45.555 72.045 45.725 73.015 ;
        RECT 45.050 71.715 45.305 72.045 ;
        RECT 45.530 71.715 45.725 72.045 ;
        RECT 45.895 72.675 47.020 72.845 ;
        RECT 45.135 71.545 45.305 71.715 ;
        RECT 45.895 71.545 46.065 72.675 ;
        RECT 44.245 70.805 44.535 71.530 ;
        RECT 44.710 70.975 44.965 71.545 ;
        RECT 45.135 71.375 46.065 71.545 ;
        RECT 46.235 72.335 47.245 72.505 ;
        RECT 46.235 71.535 46.405 72.335 ;
        RECT 45.890 71.340 46.065 71.375 ;
        RECT 45.135 70.805 45.465 71.205 ;
        RECT 45.890 70.975 46.420 71.340 ;
        RECT 46.610 71.315 46.885 72.135 ;
        RECT 46.605 71.145 46.885 71.315 ;
        RECT 46.610 70.975 46.885 71.145 ;
        RECT 47.055 70.975 47.245 72.335 ;
        RECT 47.415 72.350 47.585 73.015 ;
        RECT 47.755 72.595 47.925 73.355 ;
        RECT 48.160 72.595 48.675 73.005 ;
        RECT 47.415 72.160 48.165 72.350 ;
        RECT 48.335 71.785 48.675 72.595 ;
        RECT 49.365 72.295 49.695 73.140 ;
        RECT 49.865 72.345 50.035 73.355 ;
        RECT 50.205 72.625 50.545 73.185 ;
        RECT 50.775 72.855 51.090 73.355 ;
        RECT 51.270 72.885 52.155 73.055 ;
        RECT 47.445 71.615 48.675 71.785 ;
        RECT 49.305 72.215 49.695 72.295 ;
        RECT 50.205 72.250 51.100 72.625 ;
        RECT 49.305 72.165 49.520 72.215 ;
        RECT 47.425 70.805 47.935 71.340 ;
        RECT 48.155 71.010 48.400 71.615 ;
        RECT 49.305 71.585 49.475 72.165 ;
        RECT 50.205 72.045 50.395 72.250 ;
        RECT 51.270 72.045 51.440 72.885 ;
        RECT 52.380 72.855 52.630 73.185 ;
        RECT 49.645 71.715 50.395 72.045 ;
        RECT 50.565 71.715 51.440 72.045 ;
        RECT 49.305 71.545 49.530 71.585 ;
        RECT 50.195 71.545 50.395 71.715 ;
        RECT 49.305 71.460 49.685 71.545 ;
        RECT 49.355 71.025 49.685 71.460 ;
        RECT 49.855 70.805 50.025 71.415 ;
        RECT 50.195 71.020 50.525 71.545 ;
        RECT 50.785 70.805 50.995 71.335 ;
        RECT 51.270 71.255 51.440 71.715 ;
        RECT 51.610 71.755 51.930 72.715 ;
        RECT 52.100 71.965 52.290 72.685 ;
        RECT 52.460 71.785 52.630 72.855 ;
        RECT 52.800 72.555 52.970 73.355 ;
        RECT 53.140 72.910 54.245 73.080 ;
        RECT 53.140 72.295 53.310 72.910 ;
        RECT 54.455 72.760 54.705 73.185 ;
        RECT 54.875 72.895 55.140 73.355 ;
        RECT 53.480 72.375 54.010 72.740 ;
        RECT 54.455 72.630 54.760 72.760 ;
        RECT 52.800 72.205 53.310 72.295 ;
        RECT 52.800 72.035 53.670 72.205 ;
        RECT 52.800 71.965 52.970 72.035 ;
        RECT 53.090 71.785 53.290 71.815 ;
        RECT 51.610 71.425 52.075 71.755 ;
        RECT 52.460 71.485 53.290 71.785 ;
        RECT 52.460 71.255 52.630 71.485 ;
        RECT 51.270 71.085 52.055 71.255 ;
        RECT 52.225 71.085 52.630 71.255 ;
        RECT 52.810 70.805 53.180 71.305 ;
        RECT 53.500 71.255 53.670 72.035 ;
        RECT 53.840 71.675 54.010 72.375 ;
        RECT 54.180 71.845 54.420 72.440 ;
        RECT 53.840 71.455 54.365 71.675 ;
        RECT 54.590 71.525 54.760 72.630 ;
        RECT 54.535 71.395 54.760 71.525 ;
        RECT 54.930 71.435 55.210 72.385 ;
        RECT 54.535 71.255 54.705 71.395 ;
        RECT 53.500 71.085 54.175 71.255 ;
        RECT 54.370 71.085 54.705 71.255 ;
        RECT 54.875 70.805 55.125 71.265 ;
        RECT 55.380 71.065 55.565 73.185 ;
        RECT 55.735 72.855 56.065 73.355 ;
        RECT 56.235 72.685 56.405 73.185 ;
        RECT 55.740 72.515 56.405 72.685 ;
        RECT 56.780 72.725 57.065 73.185 ;
        RECT 57.235 72.895 57.505 73.355 ;
        RECT 55.740 71.525 55.970 72.515 ;
        RECT 56.780 72.505 57.735 72.725 ;
        RECT 56.140 71.695 56.490 72.345 ;
        RECT 56.665 71.775 57.355 72.335 ;
        RECT 57.525 71.605 57.735 72.505 ;
        RECT 55.740 71.355 56.405 71.525 ;
        RECT 55.735 70.805 56.065 71.185 ;
        RECT 56.235 71.065 56.405 71.355 ;
        RECT 56.780 71.435 57.735 71.605 ;
        RECT 57.905 72.335 58.305 73.185 ;
        RECT 58.495 72.725 58.775 73.185 ;
        RECT 59.295 72.895 59.620 73.355 ;
        RECT 58.495 72.505 59.620 72.725 ;
        RECT 57.905 71.775 59.000 72.335 ;
        RECT 59.170 72.045 59.620 72.505 ;
        RECT 59.790 72.215 60.175 73.185 ;
        RECT 56.780 70.975 57.065 71.435 ;
        RECT 57.235 70.805 57.505 71.265 ;
        RECT 57.905 70.975 58.305 71.775 ;
        RECT 59.170 71.715 59.725 72.045 ;
        RECT 59.170 71.605 59.620 71.715 ;
        RECT 58.495 71.435 59.620 71.605 ;
        RECT 59.895 71.545 60.175 72.215 ;
        RECT 58.495 70.975 58.775 71.435 ;
        RECT 59.295 70.805 59.620 71.265 ;
        RECT 59.790 70.975 60.175 71.545 ;
        RECT 60.345 71.085 60.625 73.185 ;
        RECT 60.815 72.595 61.600 73.355 ;
        RECT 61.995 72.525 62.380 73.185 ;
        RECT 61.995 72.425 62.405 72.525 ;
        RECT 60.795 72.215 62.405 72.425 ;
        RECT 62.705 72.335 62.905 73.125 ;
        RECT 60.795 71.615 61.070 72.215 ;
        RECT 62.575 72.165 62.905 72.335 ;
        RECT 63.075 72.175 63.395 73.355 ;
        RECT 63.765 72.685 64.045 73.355 ;
        RECT 64.215 72.465 64.515 73.015 ;
        RECT 64.715 72.635 65.045 73.355 ;
        RECT 65.235 72.635 65.695 73.185 ;
        RECT 62.575 72.045 62.755 72.165 ;
        RECT 61.240 71.795 61.595 72.045 ;
        RECT 61.790 71.995 62.255 72.045 ;
        RECT 61.785 71.825 62.255 71.995 ;
        RECT 61.790 71.795 62.255 71.825 ;
        RECT 62.425 71.795 62.755 72.045 ;
        RECT 63.580 72.045 63.845 72.405 ;
        RECT 64.215 72.295 65.155 72.465 ;
        RECT 64.985 72.045 65.155 72.295 ;
        RECT 62.930 71.795 63.395 71.995 ;
        RECT 63.580 71.795 64.255 72.045 ;
        RECT 64.475 71.795 64.815 72.045 ;
        RECT 64.985 71.715 65.275 72.045 ;
        RECT 64.985 71.625 65.155 71.715 ;
        RECT 60.795 71.435 62.045 71.615 ;
        RECT 61.680 71.365 62.045 71.435 ;
        RECT 62.215 71.415 63.395 71.585 ;
        RECT 60.855 70.805 61.025 71.265 ;
        RECT 62.215 71.195 62.545 71.415 ;
        RECT 61.295 71.015 62.545 71.195 ;
        RECT 62.715 70.805 62.885 71.245 ;
        RECT 63.055 71.000 63.395 71.415 ;
        RECT 63.765 71.435 65.155 71.625 ;
        RECT 63.765 71.075 64.095 71.435 ;
        RECT 65.445 71.265 65.695 72.635 ;
        RECT 65.865 72.215 66.125 73.355 ;
        RECT 66.295 72.205 66.625 73.185 ;
        RECT 66.795 72.215 67.075 73.355 ;
        RECT 67.795 72.425 67.965 73.185 ;
        RECT 68.180 72.595 68.510 73.355 ;
        RECT 67.795 72.255 68.510 72.425 ;
        RECT 68.680 72.280 68.935 73.185 ;
        RECT 65.885 71.795 66.220 72.045 ;
        RECT 66.390 71.605 66.560 72.205 ;
        RECT 66.730 71.775 67.065 72.045 ;
        RECT 67.705 71.705 68.060 72.075 ;
        RECT 68.340 72.045 68.510 72.255 ;
        RECT 68.340 71.715 68.595 72.045 ;
        RECT 64.715 70.805 64.965 71.265 ;
        RECT 65.135 70.975 65.695 71.265 ;
        RECT 65.865 70.975 66.560 71.605 ;
        RECT 66.765 70.805 67.075 71.605 ;
        RECT 68.340 71.525 68.510 71.715 ;
        RECT 68.765 71.550 68.935 72.280 ;
        RECT 69.110 72.205 69.370 73.355 ;
        RECT 70.005 72.190 70.295 73.355 ;
        RECT 70.465 72.265 73.055 73.355 ;
        RECT 73.775 72.685 73.945 73.185 ;
        RECT 74.115 72.855 74.445 73.355 ;
        RECT 73.775 72.515 74.440 72.685 ;
        RECT 67.795 71.355 68.510 71.525 ;
        RECT 67.795 70.975 67.965 71.355 ;
        RECT 68.180 70.805 68.510 71.185 ;
        RECT 68.680 70.975 68.935 71.550 ;
        RECT 69.110 70.805 69.370 71.645 ;
        RECT 70.465 71.575 71.675 72.095 ;
        RECT 71.845 71.745 73.055 72.265 ;
        RECT 73.690 71.695 74.040 72.345 ;
        RECT 70.005 70.805 70.295 71.530 ;
        RECT 70.465 70.805 73.055 71.575 ;
        RECT 74.210 71.525 74.440 72.515 ;
        RECT 73.775 71.355 74.440 71.525 ;
        RECT 73.775 71.065 73.945 71.355 ;
        RECT 74.115 70.805 74.445 71.185 ;
        RECT 74.615 71.065 74.800 73.185 ;
        RECT 75.040 72.895 75.305 73.355 ;
        RECT 75.475 72.760 75.725 73.185 ;
        RECT 75.935 72.910 77.040 73.080 ;
        RECT 75.420 72.630 75.725 72.760 ;
        RECT 74.970 71.435 75.250 72.385 ;
        RECT 75.420 71.525 75.590 72.630 ;
        RECT 75.760 71.845 76.000 72.440 ;
        RECT 76.170 72.375 76.700 72.740 ;
        RECT 76.170 71.675 76.340 72.375 ;
        RECT 76.870 72.295 77.040 72.910 ;
        RECT 77.210 72.555 77.380 73.355 ;
        RECT 77.550 72.855 77.800 73.185 ;
        RECT 78.025 72.885 78.910 73.055 ;
        RECT 76.870 72.205 77.380 72.295 ;
        RECT 75.420 71.395 75.645 71.525 ;
        RECT 75.815 71.455 76.340 71.675 ;
        RECT 76.510 72.035 77.380 72.205 ;
        RECT 75.055 70.805 75.305 71.265 ;
        RECT 75.475 71.255 75.645 71.395 ;
        RECT 76.510 71.255 76.680 72.035 ;
        RECT 77.210 71.965 77.380 72.035 ;
        RECT 76.890 71.785 77.090 71.815 ;
        RECT 77.550 71.785 77.720 72.855 ;
        RECT 77.890 71.965 78.080 72.685 ;
        RECT 76.890 71.485 77.720 71.785 ;
        RECT 78.250 71.755 78.570 72.715 ;
        RECT 75.475 71.085 75.810 71.255 ;
        RECT 76.005 71.085 76.680 71.255 ;
        RECT 77.000 70.805 77.370 71.305 ;
        RECT 77.550 71.255 77.720 71.485 ;
        RECT 78.105 71.425 78.570 71.755 ;
        RECT 78.740 72.045 78.910 72.885 ;
        RECT 79.090 72.855 79.405 73.355 ;
        RECT 79.635 72.625 79.975 73.185 ;
        RECT 79.080 72.250 79.975 72.625 ;
        RECT 80.145 72.345 80.315 73.355 ;
        RECT 79.785 72.045 79.975 72.250 ;
        RECT 80.485 72.295 80.815 73.140 ;
        RECT 81.135 72.425 81.305 73.185 ;
        RECT 81.520 72.595 81.850 73.355 ;
        RECT 80.485 72.215 80.875 72.295 ;
        RECT 81.135 72.255 81.850 72.425 ;
        RECT 82.020 72.280 82.275 73.185 ;
        RECT 80.660 72.165 80.875 72.215 ;
        RECT 78.740 71.715 79.615 72.045 ;
        RECT 79.785 71.715 80.535 72.045 ;
        RECT 78.740 71.255 78.910 71.715 ;
        RECT 79.785 71.545 79.985 71.715 ;
        RECT 80.705 71.585 80.875 72.165 ;
        RECT 81.045 71.705 81.400 72.075 ;
        RECT 81.680 72.045 81.850 72.255 ;
        RECT 81.680 71.715 81.935 72.045 ;
        RECT 80.650 71.545 80.875 71.585 ;
        RECT 77.550 71.085 77.955 71.255 ;
        RECT 78.125 71.085 78.910 71.255 ;
        RECT 79.185 70.805 79.395 71.335 ;
        RECT 79.655 71.020 79.985 71.545 ;
        RECT 80.495 71.460 80.875 71.545 ;
        RECT 81.680 71.525 81.850 71.715 ;
        RECT 82.105 71.550 82.275 72.280 ;
        RECT 82.450 72.205 82.710 73.355 ;
        RECT 82.885 72.265 84.095 73.355 ;
        RECT 82.885 71.725 83.405 72.265 ;
        RECT 80.155 70.805 80.325 71.415 ;
        RECT 80.495 71.025 80.825 71.460 ;
        RECT 81.135 71.355 81.850 71.525 ;
        RECT 81.135 70.975 81.305 71.355 ;
        RECT 81.520 70.805 81.850 71.185 ;
        RECT 82.020 70.975 82.275 71.550 ;
        RECT 82.450 70.805 82.710 71.645 ;
        RECT 83.575 71.555 84.095 72.095 ;
        RECT 82.885 70.805 84.095 71.555 ;
        RECT 5.520 70.635 84.180 70.805 ;
        RECT 5.605 69.885 6.815 70.635 ;
        RECT 7.450 69.895 7.705 70.465 ;
        RECT 7.875 70.235 8.205 70.635 ;
        RECT 8.630 70.100 9.160 70.465 ;
        RECT 8.630 70.065 8.805 70.100 ;
        RECT 7.875 69.895 8.805 70.065 ;
        RECT 5.605 69.345 6.125 69.885 ;
        RECT 6.295 69.175 6.815 69.715 ;
        RECT 5.605 68.085 6.815 69.175 ;
        RECT 7.450 69.225 7.620 69.895 ;
        RECT 7.875 69.725 8.045 69.895 ;
        RECT 7.790 69.395 8.045 69.725 ;
        RECT 8.270 69.395 8.465 69.725 ;
        RECT 7.450 68.255 7.785 69.225 ;
        RECT 7.955 68.085 8.125 69.225 ;
        RECT 8.295 68.425 8.465 69.395 ;
        RECT 8.635 68.765 8.805 69.895 ;
        RECT 8.975 69.105 9.145 69.905 ;
        RECT 9.350 69.615 9.625 70.465 ;
        RECT 9.345 69.445 9.625 69.615 ;
        RECT 9.350 69.305 9.625 69.445 ;
        RECT 9.795 69.105 9.985 70.465 ;
        RECT 10.165 70.100 10.675 70.635 ;
        RECT 10.895 69.825 11.140 70.430 ;
        RECT 11.590 69.895 11.845 70.465 ;
        RECT 12.015 70.235 12.345 70.635 ;
        RECT 12.770 70.100 13.300 70.465 ;
        RECT 12.770 70.065 12.945 70.100 ;
        RECT 12.015 69.895 12.945 70.065 ;
        RECT 10.185 69.655 11.415 69.825 ;
        RECT 8.975 68.935 9.985 69.105 ;
        RECT 10.155 69.090 10.905 69.280 ;
        RECT 8.635 68.595 9.760 68.765 ;
        RECT 10.155 68.425 10.325 69.090 ;
        RECT 11.075 68.845 11.415 69.655 ;
        RECT 8.295 68.255 10.325 68.425 ;
        RECT 10.495 68.085 10.665 68.845 ;
        RECT 10.900 68.435 11.415 68.845 ;
        RECT 11.590 69.225 11.760 69.895 ;
        RECT 12.015 69.725 12.185 69.895 ;
        RECT 11.930 69.395 12.185 69.725 ;
        RECT 12.410 69.395 12.605 69.725 ;
        RECT 11.590 68.255 11.925 69.225 ;
        RECT 12.095 68.085 12.265 69.225 ;
        RECT 12.435 68.425 12.605 69.395 ;
        RECT 12.775 68.765 12.945 69.895 ;
        RECT 13.115 69.105 13.285 69.905 ;
        RECT 13.490 69.615 13.765 70.465 ;
        RECT 13.485 69.445 13.765 69.615 ;
        RECT 13.490 69.305 13.765 69.445 ;
        RECT 13.935 69.105 14.125 70.465 ;
        RECT 14.305 70.100 14.815 70.635 ;
        RECT 15.035 69.825 15.280 70.430 ;
        RECT 16.920 69.825 17.165 70.430 ;
        RECT 17.385 70.100 17.895 70.635 ;
        RECT 14.325 69.655 15.555 69.825 ;
        RECT 13.115 68.935 14.125 69.105 ;
        RECT 14.295 69.090 15.045 69.280 ;
        RECT 12.775 68.595 13.900 68.765 ;
        RECT 14.295 68.425 14.465 69.090 ;
        RECT 15.215 68.845 15.555 69.655 ;
        RECT 12.435 68.255 14.465 68.425 ;
        RECT 14.635 68.085 14.805 68.845 ;
        RECT 15.040 68.435 15.555 68.845 ;
        RECT 16.645 69.655 17.875 69.825 ;
        RECT 16.645 68.845 16.985 69.655 ;
        RECT 17.155 69.090 17.905 69.280 ;
        RECT 16.645 68.435 17.160 68.845 ;
        RECT 17.395 68.085 17.565 68.845 ;
        RECT 17.735 68.425 17.905 69.090 ;
        RECT 18.075 69.105 18.265 70.465 ;
        RECT 18.435 70.295 18.710 70.465 ;
        RECT 18.435 70.125 18.715 70.295 ;
        RECT 18.435 69.305 18.710 70.125 ;
        RECT 18.900 70.100 19.430 70.465 ;
        RECT 19.855 70.235 20.185 70.635 ;
        RECT 19.255 70.065 19.430 70.100 ;
        RECT 18.915 69.105 19.085 69.905 ;
        RECT 18.075 68.935 19.085 69.105 ;
        RECT 19.255 69.895 20.185 70.065 ;
        RECT 20.355 69.895 20.610 70.465 ;
        RECT 20.845 70.175 21.090 70.635 ;
        RECT 19.255 68.765 19.425 69.895 ;
        RECT 20.015 69.725 20.185 69.895 ;
        RECT 18.300 68.595 19.425 68.765 ;
        RECT 19.595 69.395 19.790 69.725 ;
        RECT 20.015 69.395 20.270 69.725 ;
        RECT 19.595 68.425 19.765 69.395 ;
        RECT 20.440 69.225 20.610 69.895 ;
        RECT 20.785 69.395 21.100 70.005 ;
        RECT 21.270 69.645 21.520 70.455 ;
        RECT 21.690 70.110 21.950 70.635 ;
        RECT 22.120 69.985 22.380 70.440 ;
        RECT 22.550 70.155 22.810 70.635 ;
        RECT 22.980 69.985 23.240 70.440 ;
        RECT 23.410 70.155 23.670 70.635 ;
        RECT 23.840 69.985 24.100 70.440 ;
        RECT 24.270 70.155 24.530 70.635 ;
        RECT 24.700 69.985 24.960 70.440 ;
        RECT 25.130 70.155 25.430 70.635 ;
        RECT 25.845 70.090 31.190 70.635 ;
        RECT 22.120 69.815 25.430 69.985 ;
        RECT 21.270 69.395 24.290 69.645 ;
        RECT 17.735 68.255 19.765 68.425 ;
        RECT 19.935 68.085 20.105 69.225 ;
        RECT 20.275 68.255 20.610 69.225 ;
        RECT 20.795 68.085 21.090 69.195 ;
        RECT 21.270 68.260 21.520 69.395 ;
        RECT 24.460 69.225 25.430 69.815 ;
        RECT 27.430 69.260 27.770 70.090 ;
        RECT 31.365 69.910 31.655 70.635 ;
        RECT 32.805 70.175 33.050 70.635 ;
        RECT 21.690 68.085 21.950 69.195 ;
        RECT 22.120 68.985 25.430 69.225 ;
        RECT 22.120 68.260 22.380 68.985 ;
        RECT 22.550 68.085 22.810 68.815 ;
        RECT 22.980 68.260 23.240 68.985 ;
        RECT 23.410 68.085 23.670 68.815 ;
        RECT 23.840 68.260 24.100 68.985 ;
        RECT 24.270 68.085 24.530 68.815 ;
        RECT 24.700 68.260 24.960 68.985 ;
        RECT 25.130 68.085 25.425 68.815 ;
        RECT 29.250 68.520 29.600 69.770 ;
        RECT 32.745 69.395 33.060 70.005 ;
        RECT 33.230 69.645 33.480 70.455 ;
        RECT 33.650 70.110 33.910 70.635 ;
        RECT 34.080 69.985 34.340 70.440 ;
        RECT 34.510 70.155 34.770 70.635 ;
        RECT 34.940 69.985 35.200 70.440 ;
        RECT 35.370 70.155 35.630 70.635 ;
        RECT 35.800 69.985 36.060 70.440 ;
        RECT 36.230 70.155 36.490 70.635 ;
        RECT 36.660 69.985 36.920 70.440 ;
        RECT 37.090 70.155 37.390 70.635 ;
        RECT 34.080 69.815 37.390 69.985 ;
        RECT 33.230 69.395 36.250 69.645 ;
        RECT 25.845 68.085 31.190 68.520 ;
        RECT 31.365 68.085 31.655 69.250 ;
        RECT 32.755 68.085 33.050 69.195 ;
        RECT 33.230 68.260 33.480 69.395 ;
        RECT 36.420 69.225 37.390 69.815 ;
        RECT 37.805 69.865 40.395 70.635 ;
        RECT 40.655 70.085 40.825 70.375 ;
        RECT 40.995 70.255 41.325 70.635 ;
        RECT 40.655 69.915 41.320 70.085 ;
        RECT 37.805 69.345 39.015 69.865 ;
        RECT 33.650 68.085 33.910 69.195 ;
        RECT 34.080 68.985 37.390 69.225 ;
        RECT 39.185 69.175 40.395 69.695 ;
        RECT 34.080 68.260 34.340 68.985 ;
        RECT 34.510 68.085 34.770 68.815 ;
        RECT 34.940 68.260 35.200 68.985 ;
        RECT 35.370 68.085 35.630 68.815 ;
        RECT 35.800 68.260 36.060 68.985 ;
        RECT 36.230 68.085 36.490 68.815 ;
        RECT 36.660 68.260 36.920 68.985 ;
        RECT 37.090 68.085 37.385 68.815 ;
        RECT 37.805 68.085 40.395 69.175 ;
        RECT 40.570 69.095 40.920 69.745 ;
        RECT 41.090 68.925 41.320 69.915 ;
        RECT 40.655 68.755 41.320 68.925 ;
        RECT 40.655 68.255 40.825 68.755 ;
        RECT 40.995 68.085 41.325 68.585 ;
        RECT 41.495 68.255 41.680 70.375 ;
        RECT 41.935 70.175 42.185 70.635 ;
        RECT 42.355 70.185 42.690 70.355 ;
        RECT 42.885 70.185 43.560 70.355 ;
        RECT 42.355 70.045 42.525 70.185 ;
        RECT 41.850 69.055 42.130 70.005 ;
        RECT 42.300 69.915 42.525 70.045 ;
        RECT 42.300 68.810 42.470 69.915 ;
        RECT 42.695 69.765 43.220 69.985 ;
        RECT 42.640 69.000 42.880 69.595 ;
        RECT 43.050 69.065 43.220 69.765 ;
        RECT 43.390 69.405 43.560 70.185 ;
        RECT 43.880 70.135 44.250 70.635 ;
        RECT 44.430 70.185 44.835 70.355 ;
        RECT 45.005 70.185 45.790 70.355 ;
        RECT 44.430 69.955 44.600 70.185 ;
        RECT 43.770 69.655 44.600 69.955 ;
        RECT 44.985 69.685 45.450 70.015 ;
        RECT 43.770 69.625 43.970 69.655 ;
        RECT 44.090 69.405 44.260 69.475 ;
        RECT 43.390 69.235 44.260 69.405 ;
        RECT 43.750 69.145 44.260 69.235 ;
        RECT 42.300 68.680 42.605 68.810 ;
        RECT 43.050 68.700 43.580 69.065 ;
        RECT 41.920 68.085 42.185 68.545 ;
        RECT 42.355 68.255 42.605 68.680 ;
        RECT 43.750 68.530 43.920 69.145 ;
        RECT 42.815 68.360 43.920 68.530 ;
        RECT 44.090 68.085 44.260 68.885 ;
        RECT 44.430 68.585 44.600 69.655 ;
        RECT 44.770 68.755 44.960 69.475 ;
        RECT 45.130 68.725 45.450 69.685 ;
        RECT 45.620 69.725 45.790 70.185 ;
        RECT 46.065 70.105 46.275 70.635 ;
        RECT 46.535 69.895 46.865 70.420 ;
        RECT 47.035 70.025 47.205 70.635 ;
        RECT 47.375 69.980 47.705 70.415 ;
        RECT 47.375 69.895 47.755 69.980 ;
        RECT 46.665 69.725 46.865 69.895 ;
        RECT 47.530 69.855 47.755 69.895 ;
        RECT 45.620 69.395 46.495 69.725 ;
        RECT 46.665 69.395 47.415 69.725 ;
        RECT 44.430 68.255 44.680 68.585 ;
        RECT 45.620 68.555 45.790 69.395 ;
        RECT 46.665 69.190 46.855 69.395 ;
        RECT 47.585 69.275 47.755 69.855 ;
        RECT 47.540 69.225 47.755 69.275 ;
        RECT 45.960 68.815 46.855 69.190 ;
        RECT 47.365 69.145 47.755 69.225 ;
        RECT 47.930 69.895 48.185 70.465 ;
        RECT 48.355 70.235 48.685 70.635 ;
        RECT 49.110 70.100 49.640 70.465 ;
        RECT 49.110 70.065 49.285 70.100 ;
        RECT 48.355 69.895 49.285 70.065 ;
        RECT 47.930 69.225 48.100 69.895 ;
        RECT 48.355 69.725 48.525 69.895 ;
        RECT 48.270 69.395 48.525 69.725 ;
        RECT 48.750 69.395 48.945 69.725 ;
        RECT 44.905 68.385 45.790 68.555 ;
        RECT 45.970 68.085 46.285 68.585 ;
        RECT 46.515 68.255 46.855 68.815 ;
        RECT 47.025 68.085 47.195 69.095 ;
        RECT 47.365 68.300 47.695 69.145 ;
        RECT 47.930 68.255 48.265 69.225 ;
        RECT 48.435 68.085 48.605 69.225 ;
        RECT 48.775 68.425 48.945 69.395 ;
        RECT 49.115 68.765 49.285 69.895 ;
        RECT 49.455 69.105 49.625 69.905 ;
        RECT 49.830 69.615 50.105 70.465 ;
        RECT 49.825 69.445 50.105 69.615 ;
        RECT 49.830 69.305 50.105 69.445 ;
        RECT 50.275 69.105 50.465 70.465 ;
        RECT 50.645 70.100 51.155 70.635 ;
        RECT 51.375 69.825 51.620 70.430 ;
        RECT 52.065 69.895 52.450 70.465 ;
        RECT 52.620 70.175 52.945 70.635 ;
        RECT 53.465 70.005 53.745 70.465 ;
        RECT 50.665 69.655 51.895 69.825 ;
        RECT 49.455 68.935 50.465 69.105 ;
        RECT 50.635 69.090 51.385 69.280 ;
        RECT 49.115 68.595 50.240 68.765 ;
        RECT 50.635 68.425 50.805 69.090 ;
        RECT 51.555 68.845 51.895 69.655 ;
        RECT 48.775 68.255 50.805 68.425 ;
        RECT 50.975 68.085 51.145 68.845 ;
        RECT 51.380 68.435 51.895 68.845 ;
        RECT 52.065 69.225 52.345 69.895 ;
        RECT 52.620 69.835 53.745 70.005 ;
        RECT 52.620 69.725 53.070 69.835 ;
        RECT 52.515 69.395 53.070 69.725 ;
        RECT 53.935 69.665 54.335 70.465 ;
        RECT 54.735 70.175 55.005 70.635 ;
        RECT 55.175 70.005 55.460 70.465 ;
        RECT 52.065 68.255 52.450 69.225 ;
        RECT 52.620 68.935 53.070 69.395 ;
        RECT 53.240 69.105 54.335 69.665 ;
        RECT 52.620 68.715 53.745 68.935 ;
        RECT 52.620 68.085 52.945 68.545 ;
        RECT 53.465 68.255 53.745 68.715 ;
        RECT 53.935 68.255 54.335 69.105 ;
        RECT 54.505 69.835 55.460 70.005 ;
        RECT 55.745 69.885 56.955 70.635 ;
        RECT 57.125 69.910 57.415 70.635 ;
        RECT 58.065 70.165 58.360 70.635 ;
        RECT 58.530 69.995 58.790 70.440 ;
        RECT 58.960 70.165 59.220 70.635 ;
        RECT 59.390 69.995 59.645 70.440 ;
        RECT 59.815 70.165 60.115 70.635 ;
        RECT 54.505 68.935 54.715 69.835 ;
        RECT 54.885 69.105 55.575 69.665 ;
        RECT 55.745 69.345 56.265 69.885 ;
        RECT 57.605 69.825 60.635 69.995 ;
        RECT 60.805 69.835 61.500 70.465 ;
        RECT 61.705 69.835 62.015 70.635 ;
        RECT 62.185 69.835 62.880 70.465 ;
        RECT 63.085 69.835 63.395 70.635 ;
        RECT 56.435 69.175 56.955 69.715 ;
        RECT 57.605 69.260 57.775 69.825 ;
        RECT 57.945 69.430 60.160 69.655 ;
        RECT 60.335 69.260 60.635 69.825 ;
        RECT 60.825 69.395 61.160 69.645 ;
        RECT 54.505 68.715 55.460 68.935 ;
        RECT 54.735 68.085 55.005 68.545 ;
        RECT 55.175 68.255 55.460 68.715 ;
        RECT 55.745 68.085 56.955 69.175 ;
        RECT 57.125 68.085 57.415 69.250 ;
        RECT 57.605 69.090 60.635 69.260 ;
        RECT 61.330 69.235 61.500 69.835 ;
        RECT 61.670 69.395 62.005 69.665 ;
        RECT 62.205 69.395 62.540 69.645 ;
        RECT 62.710 69.235 62.880 69.835 ;
        RECT 63.575 69.825 63.845 70.635 ;
        RECT 64.015 69.825 64.345 70.465 ;
        RECT 64.515 69.825 64.755 70.635 ;
        RECT 65.870 69.870 66.325 70.635 ;
        RECT 66.600 70.255 67.900 70.465 ;
        RECT 68.155 70.275 68.485 70.635 ;
        RECT 67.730 70.105 67.900 70.255 ;
        RECT 68.655 70.135 68.915 70.465 ;
        RECT 68.685 70.125 68.915 70.135 ;
        RECT 63.050 69.395 63.385 69.665 ;
        RECT 63.565 69.395 63.915 69.645 ;
        RECT 57.585 68.085 57.930 68.920 ;
        RECT 58.105 68.285 58.360 69.090 ;
        RECT 58.530 68.085 58.790 68.920 ;
        RECT 58.965 68.285 59.220 69.090 ;
        RECT 59.390 68.085 59.650 68.920 ;
        RECT 59.820 68.285 60.080 69.090 ;
        RECT 60.250 68.085 60.635 68.920 ;
        RECT 60.805 68.085 61.065 69.225 ;
        RECT 61.235 68.255 61.565 69.235 ;
        RECT 61.735 68.085 62.015 69.225 ;
        RECT 62.185 68.085 62.445 69.225 ;
        RECT 62.615 68.255 62.945 69.235 ;
        RECT 64.085 69.225 64.255 69.825 ;
        RECT 66.800 69.645 67.020 70.045 ;
        RECT 64.425 69.395 64.775 69.645 ;
        RECT 65.865 69.445 66.355 69.645 ;
        RECT 66.545 69.435 67.020 69.645 ;
        RECT 67.265 69.645 67.475 70.045 ;
        RECT 67.730 69.980 68.485 70.105 ;
        RECT 67.730 69.935 68.575 69.980 ;
        RECT 68.305 69.815 68.575 69.935 ;
        RECT 67.265 69.435 67.595 69.645 ;
        RECT 67.765 69.375 68.175 69.680 ;
        RECT 63.115 68.085 63.395 69.225 ;
        RECT 63.575 68.085 63.905 69.225 ;
        RECT 64.085 69.055 64.765 69.225 ;
        RECT 64.435 68.270 64.765 69.055 ;
        RECT 65.870 69.205 67.045 69.265 ;
        RECT 68.405 69.240 68.575 69.815 ;
        RECT 68.375 69.205 68.575 69.240 ;
        RECT 65.870 69.095 68.575 69.205 ;
        RECT 65.870 68.475 66.125 69.095 ;
        RECT 66.715 69.035 68.515 69.095 ;
        RECT 66.715 69.005 67.045 69.035 ;
        RECT 68.745 68.935 68.915 70.125 ;
        RECT 69.290 69.855 69.790 70.465 ;
        RECT 69.085 69.395 69.435 69.645 ;
        RECT 69.620 69.225 69.790 69.855 ;
        RECT 70.420 69.985 70.750 70.465 ;
        RECT 70.920 70.175 71.145 70.635 ;
        RECT 71.315 69.985 71.645 70.465 ;
        RECT 70.420 69.815 71.645 69.985 ;
        RECT 71.835 69.835 72.085 70.635 ;
        RECT 72.255 69.835 72.595 70.465 ;
        RECT 69.960 69.445 70.290 69.645 ;
        RECT 70.460 69.445 70.790 69.645 ;
        RECT 70.960 69.445 71.380 69.645 ;
        RECT 71.555 69.475 72.250 69.645 ;
        RECT 71.555 69.225 71.725 69.475 ;
        RECT 72.420 69.225 72.595 69.835 ;
        RECT 72.765 69.865 74.435 70.635 ;
        RECT 75.070 69.895 75.325 70.465 ;
        RECT 75.495 70.235 75.825 70.635 ;
        RECT 76.250 70.100 76.780 70.465 ;
        RECT 76.250 70.065 76.425 70.100 ;
        RECT 75.495 69.895 76.425 70.065 ;
        RECT 72.765 69.345 73.515 69.865 ;
        RECT 66.375 68.835 66.560 68.925 ;
        RECT 67.150 68.835 67.985 68.845 ;
        RECT 66.375 68.635 67.985 68.835 ;
        RECT 66.375 68.595 66.605 68.635 ;
        RECT 65.870 68.255 66.205 68.475 ;
        RECT 67.210 68.085 67.565 68.465 ;
        RECT 67.735 68.255 67.985 68.635 ;
        RECT 68.235 68.085 68.485 68.865 ;
        RECT 68.655 68.255 68.915 68.935 ;
        RECT 69.290 69.055 71.725 69.225 ;
        RECT 69.290 68.255 69.620 69.055 ;
        RECT 69.790 68.085 70.120 68.885 ;
        RECT 70.420 68.255 70.750 69.055 ;
        RECT 71.395 68.085 71.645 68.885 ;
        RECT 71.915 68.085 72.085 69.225 ;
        RECT 72.255 68.255 72.595 69.225 ;
        RECT 73.685 69.175 74.435 69.695 ;
        RECT 72.765 68.085 74.435 69.175 ;
        RECT 75.070 69.225 75.240 69.895 ;
        RECT 75.495 69.725 75.665 69.895 ;
        RECT 75.410 69.395 75.665 69.725 ;
        RECT 75.890 69.395 76.085 69.725 ;
        RECT 75.070 68.255 75.405 69.225 ;
        RECT 75.575 68.085 75.745 69.225 ;
        RECT 75.915 68.425 76.085 69.395 ;
        RECT 76.255 68.765 76.425 69.895 ;
        RECT 76.595 69.105 76.765 69.905 ;
        RECT 76.970 69.615 77.245 70.465 ;
        RECT 76.965 69.445 77.245 69.615 ;
        RECT 76.970 69.305 77.245 69.445 ;
        RECT 77.415 69.105 77.605 70.465 ;
        RECT 77.785 70.100 78.295 70.635 ;
        RECT 78.515 69.825 78.760 70.430 ;
        RECT 79.205 69.895 79.590 70.465 ;
        RECT 79.760 70.175 80.085 70.635 ;
        RECT 80.605 70.005 80.885 70.465 ;
        RECT 77.805 69.655 79.035 69.825 ;
        RECT 76.595 68.935 77.605 69.105 ;
        RECT 77.775 69.090 78.525 69.280 ;
        RECT 76.255 68.595 77.380 68.765 ;
        RECT 77.775 68.425 77.945 69.090 ;
        RECT 78.695 68.845 79.035 69.655 ;
        RECT 75.915 68.255 77.945 68.425 ;
        RECT 78.115 68.085 78.285 68.845 ;
        RECT 78.520 68.435 79.035 68.845 ;
        RECT 79.205 69.225 79.485 69.895 ;
        RECT 79.760 69.835 80.885 70.005 ;
        RECT 79.760 69.725 80.210 69.835 ;
        RECT 79.655 69.395 80.210 69.725 ;
        RECT 81.075 69.665 81.475 70.465 ;
        RECT 81.875 70.175 82.145 70.635 ;
        RECT 82.315 70.005 82.600 70.465 ;
        RECT 79.205 68.255 79.590 69.225 ;
        RECT 79.760 68.935 80.210 69.395 ;
        RECT 80.380 69.105 81.475 69.665 ;
        RECT 79.760 68.715 80.885 68.935 ;
        RECT 79.760 68.085 80.085 68.545 ;
        RECT 80.605 68.255 80.885 68.715 ;
        RECT 81.075 68.255 81.475 69.105 ;
        RECT 81.645 69.835 82.600 70.005 ;
        RECT 82.885 69.885 84.095 70.635 ;
        RECT 81.645 68.935 81.855 69.835 ;
        RECT 82.025 69.105 82.715 69.665 ;
        RECT 82.885 69.175 83.405 69.715 ;
        RECT 83.575 69.345 84.095 69.885 ;
        RECT 81.645 68.715 82.600 68.935 ;
        RECT 81.875 68.085 82.145 68.545 ;
        RECT 82.315 68.255 82.600 68.715 ;
        RECT 82.885 68.085 84.095 69.175 ;
        RECT 5.520 67.915 84.180 68.085 ;
        RECT 5.605 66.825 6.815 67.915 ;
        RECT 7.075 67.245 7.245 67.745 ;
        RECT 7.415 67.415 7.745 67.915 ;
        RECT 7.075 67.075 7.740 67.245 ;
        RECT 5.605 66.115 6.125 66.655 ;
        RECT 6.295 66.285 6.815 66.825 ;
        RECT 6.990 66.255 7.340 66.905 ;
        RECT 5.605 65.365 6.815 66.115 ;
        RECT 7.510 66.085 7.740 67.075 ;
        RECT 7.075 65.915 7.740 66.085 ;
        RECT 7.075 65.625 7.245 65.915 ;
        RECT 7.415 65.365 7.745 65.745 ;
        RECT 7.915 65.625 8.100 67.745 ;
        RECT 8.340 67.455 8.605 67.915 ;
        RECT 8.775 67.320 9.025 67.745 ;
        RECT 9.235 67.470 10.340 67.640 ;
        RECT 8.720 67.190 9.025 67.320 ;
        RECT 8.270 65.995 8.550 66.945 ;
        RECT 8.720 66.085 8.890 67.190 ;
        RECT 9.060 66.405 9.300 67.000 ;
        RECT 9.470 66.935 10.000 67.300 ;
        RECT 9.470 66.235 9.640 66.935 ;
        RECT 10.170 66.855 10.340 67.470 ;
        RECT 10.510 67.115 10.680 67.915 ;
        RECT 10.850 67.415 11.100 67.745 ;
        RECT 11.325 67.445 12.210 67.615 ;
        RECT 10.170 66.765 10.680 66.855 ;
        RECT 8.720 65.955 8.945 66.085 ;
        RECT 9.115 66.015 9.640 66.235 ;
        RECT 9.810 66.595 10.680 66.765 ;
        RECT 8.355 65.365 8.605 65.825 ;
        RECT 8.775 65.815 8.945 65.955 ;
        RECT 9.810 65.815 9.980 66.595 ;
        RECT 10.510 66.525 10.680 66.595 ;
        RECT 10.190 66.345 10.390 66.375 ;
        RECT 10.850 66.345 11.020 67.415 ;
        RECT 11.190 66.525 11.380 67.245 ;
        RECT 10.190 66.045 11.020 66.345 ;
        RECT 11.550 66.315 11.870 67.275 ;
        RECT 8.775 65.645 9.110 65.815 ;
        RECT 9.305 65.645 9.980 65.815 ;
        RECT 10.300 65.365 10.670 65.865 ;
        RECT 10.850 65.815 11.020 66.045 ;
        RECT 11.405 65.985 11.870 66.315 ;
        RECT 12.040 66.605 12.210 67.445 ;
        RECT 12.390 67.415 12.705 67.915 ;
        RECT 12.935 67.185 13.275 67.745 ;
        RECT 12.380 66.810 13.275 67.185 ;
        RECT 13.445 66.905 13.615 67.915 ;
        RECT 13.085 66.605 13.275 66.810 ;
        RECT 13.785 66.855 14.115 67.700 ;
        RECT 14.285 67.000 14.455 67.915 ;
        RECT 13.785 66.775 14.175 66.855 ;
        RECT 14.805 66.825 18.315 67.915 ;
        RECT 13.960 66.725 14.175 66.775 ;
        RECT 12.040 66.275 12.915 66.605 ;
        RECT 13.085 66.275 13.835 66.605 ;
        RECT 12.040 65.815 12.210 66.275 ;
        RECT 13.085 66.105 13.285 66.275 ;
        RECT 14.005 66.145 14.175 66.725 ;
        RECT 13.950 66.105 14.175 66.145 ;
        RECT 10.850 65.645 11.255 65.815 ;
        RECT 11.425 65.645 12.210 65.815 ;
        RECT 12.485 65.365 12.695 65.895 ;
        RECT 12.955 65.580 13.285 66.105 ;
        RECT 13.795 66.020 14.175 66.105 ;
        RECT 14.805 66.135 16.455 66.655 ;
        RECT 16.625 66.305 18.315 66.825 ;
        RECT 18.485 66.750 18.775 67.915 ;
        RECT 19.035 67.245 19.205 67.745 ;
        RECT 19.375 67.415 19.705 67.915 ;
        RECT 19.035 67.075 19.700 67.245 ;
        RECT 18.950 66.255 19.300 66.905 ;
        RECT 13.455 65.365 13.625 65.975 ;
        RECT 13.795 65.585 14.125 66.020 ;
        RECT 14.295 65.365 14.465 65.880 ;
        RECT 14.805 65.365 18.315 66.135 ;
        RECT 18.485 65.365 18.775 66.090 ;
        RECT 19.470 66.085 19.700 67.075 ;
        RECT 19.035 65.915 19.700 66.085 ;
        RECT 19.035 65.625 19.205 65.915 ;
        RECT 19.375 65.365 19.705 65.745 ;
        RECT 19.875 65.625 20.060 67.745 ;
        RECT 20.300 67.455 20.565 67.915 ;
        RECT 20.735 67.320 20.985 67.745 ;
        RECT 21.195 67.470 22.300 67.640 ;
        RECT 20.680 67.190 20.985 67.320 ;
        RECT 20.230 65.995 20.510 66.945 ;
        RECT 20.680 66.085 20.850 67.190 ;
        RECT 21.020 66.405 21.260 67.000 ;
        RECT 21.430 66.935 21.960 67.300 ;
        RECT 21.430 66.235 21.600 66.935 ;
        RECT 22.130 66.855 22.300 67.470 ;
        RECT 22.470 67.115 22.640 67.915 ;
        RECT 22.810 67.415 23.060 67.745 ;
        RECT 23.285 67.445 24.170 67.615 ;
        RECT 22.130 66.765 22.640 66.855 ;
        RECT 20.680 65.955 20.905 66.085 ;
        RECT 21.075 66.015 21.600 66.235 ;
        RECT 21.770 66.595 22.640 66.765 ;
        RECT 20.315 65.365 20.565 65.825 ;
        RECT 20.735 65.815 20.905 65.955 ;
        RECT 21.770 65.815 21.940 66.595 ;
        RECT 22.470 66.525 22.640 66.595 ;
        RECT 22.150 66.345 22.350 66.375 ;
        RECT 22.810 66.345 22.980 67.415 ;
        RECT 23.150 66.525 23.340 67.245 ;
        RECT 22.150 66.045 22.980 66.345 ;
        RECT 23.510 66.315 23.830 67.275 ;
        RECT 20.735 65.645 21.070 65.815 ;
        RECT 21.265 65.645 21.940 65.815 ;
        RECT 22.260 65.365 22.630 65.865 ;
        RECT 22.810 65.815 22.980 66.045 ;
        RECT 23.365 65.985 23.830 66.315 ;
        RECT 24.000 66.605 24.170 67.445 ;
        RECT 24.350 67.415 24.665 67.915 ;
        RECT 24.895 67.185 25.235 67.745 ;
        RECT 24.340 66.810 25.235 67.185 ;
        RECT 25.405 66.905 25.575 67.915 ;
        RECT 25.045 66.605 25.235 66.810 ;
        RECT 25.745 66.855 26.075 67.700 ;
        RECT 26.245 67.000 26.415 67.915 ;
        RECT 25.745 66.775 26.135 66.855 ;
        RECT 26.765 66.825 28.435 67.915 ;
        RECT 25.920 66.725 26.135 66.775 ;
        RECT 24.000 66.275 24.875 66.605 ;
        RECT 25.045 66.275 25.795 66.605 ;
        RECT 24.000 65.815 24.170 66.275 ;
        RECT 25.045 66.105 25.245 66.275 ;
        RECT 25.965 66.145 26.135 66.725 ;
        RECT 25.910 66.105 26.135 66.145 ;
        RECT 22.810 65.645 23.215 65.815 ;
        RECT 23.385 65.645 24.170 65.815 ;
        RECT 24.445 65.365 24.655 65.895 ;
        RECT 24.915 65.580 25.245 66.105 ;
        RECT 25.755 66.020 26.135 66.105 ;
        RECT 26.765 66.135 27.515 66.655 ;
        RECT 27.685 66.305 28.435 66.825 ;
        RECT 28.610 66.775 28.945 67.745 ;
        RECT 29.115 66.775 29.285 67.915 ;
        RECT 29.455 67.575 31.485 67.745 ;
        RECT 25.415 65.365 25.585 65.975 ;
        RECT 25.755 65.585 26.085 66.020 ;
        RECT 26.255 65.365 26.425 65.880 ;
        RECT 26.765 65.365 28.435 66.135 ;
        RECT 28.610 66.105 28.780 66.775 ;
        RECT 29.455 66.605 29.625 67.575 ;
        RECT 28.950 66.275 29.205 66.605 ;
        RECT 29.430 66.275 29.625 66.605 ;
        RECT 29.795 67.235 30.920 67.405 ;
        RECT 29.035 66.105 29.205 66.275 ;
        RECT 29.795 66.105 29.965 67.235 ;
        RECT 28.610 65.535 28.865 66.105 ;
        RECT 29.035 65.935 29.965 66.105 ;
        RECT 30.135 66.895 31.145 67.065 ;
        RECT 30.135 66.095 30.305 66.895 ;
        RECT 29.790 65.900 29.965 65.935 ;
        RECT 29.035 65.365 29.365 65.765 ;
        RECT 29.790 65.535 30.320 65.900 ;
        RECT 30.510 65.875 30.785 66.695 ;
        RECT 30.505 65.705 30.785 65.875 ;
        RECT 30.510 65.535 30.785 65.705 ;
        RECT 30.955 65.535 31.145 66.895 ;
        RECT 31.315 66.910 31.485 67.575 ;
        RECT 31.655 67.155 31.825 67.915 ;
        RECT 32.060 67.155 32.575 67.565 ;
        RECT 31.315 66.720 32.065 66.910 ;
        RECT 32.235 66.345 32.575 67.155 ;
        RECT 32.835 67.245 33.005 67.745 ;
        RECT 33.175 67.415 33.505 67.915 ;
        RECT 32.835 67.075 33.500 67.245 ;
        RECT 31.345 66.175 32.575 66.345 ;
        RECT 32.750 66.255 33.100 66.905 ;
        RECT 31.325 65.365 31.835 65.900 ;
        RECT 32.055 65.570 32.300 66.175 ;
        RECT 33.270 66.085 33.500 67.075 ;
        RECT 32.835 65.915 33.500 66.085 ;
        RECT 32.835 65.625 33.005 65.915 ;
        RECT 33.175 65.365 33.505 65.745 ;
        RECT 33.675 65.625 33.860 67.745 ;
        RECT 34.100 67.455 34.365 67.915 ;
        RECT 34.535 67.320 34.785 67.745 ;
        RECT 34.995 67.470 36.100 67.640 ;
        RECT 34.480 67.190 34.785 67.320 ;
        RECT 34.030 65.995 34.310 66.945 ;
        RECT 34.480 66.085 34.650 67.190 ;
        RECT 34.820 66.405 35.060 67.000 ;
        RECT 35.230 66.935 35.760 67.300 ;
        RECT 35.230 66.235 35.400 66.935 ;
        RECT 35.930 66.855 36.100 67.470 ;
        RECT 36.270 67.115 36.440 67.915 ;
        RECT 36.610 67.415 36.860 67.745 ;
        RECT 37.085 67.445 37.970 67.615 ;
        RECT 35.930 66.765 36.440 66.855 ;
        RECT 34.480 65.955 34.705 66.085 ;
        RECT 34.875 66.015 35.400 66.235 ;
        RECT 35.570 66.595 36.440 66.765 ;
        RECT 34.115 65.365 34.365 65.825 ;
        RECT 34.535 65.815 34.705 65.955 ;
        RECT 35.570 65.815 35.740 66.595 ;
        RECT 36.270 66.525 36.440 66.595 ;
        RECT 35.950 66.345 36.150 66.375 ;
        RECT 36.610 66.345 36.780 67.415 ;
        RECT 36.950 66.525 37.140 67.245 ;
        RECT 35.950 66.045 36.780 66.345 ;
        RECT 37.310 66.315 37.630 67.275 ;
        RECT 34.535 65.645 34.870 65.815 ;
        RECT 35.065 65.645 35.740 65.815 ;
        RECT 36.060 65.365 36.430 65.865 ;
        RECT 36.610 65.815 36.780 66.045 ;
        RECT 37.165 65.985 37.630 66.315 ;
        RECT 37.800 66.605 37.970 67.445 ;
        RECT 38.150 67.415 38.465 67.915 ;
        RECT 38.695 67.185 39.035 67.745 ;
        RECT 38.140 66.810 39.035 67.185 ;
        RECT 39.205 66.905 39.375 67.915 ;
        RECT 38.845 66.605 39.035 66.810 ;
        RECT 39.545 66.855 39.875 67.700 ;
        RECT 39.545 66.775 39.935 66.855 ;
        RECT 39.720 66.725 39.935 66.775 ;
        RECT 37.800 66.275 38.675 66.605 ;
        RECT 38.845 66.275 39.595 66.605 ;
        RECT 37.800 65.815 37.970 66.275 ;
        RECT 38.845 66.105 39.045 66.275 ;
        RECT 39.765 66.145 39.935 66.725 ;
        RECT 39.710 66.105 39.935 66.145 ;
        RECT 36.610 65.645 37.015 65.815 ;
        RECT 37.185 65.645 37.970 65.815 ;
        RECT 38.245 65.365 38.455 65.895 ;
        RECT 38.715 65.580 39.045 66.105 ;
        RECT 39.555 66.020 39.935 66.105 ;
        RECT 40.110 66.775 40.445 67.745 ;
        RECT 40.615 66.775 40.785 67.915 ;
        RECT 40.955 67.575 42.985 67.745 ;
        RECT 40.110 66.105 40.280 66.775 ;
        RECT 40.955 66.605 41.125 67.575 ;
        RECT 40.450 66.275 40.705 66.605 ;
        RECT 40.930 66.275 41.125 66.605 ;
        RECT 41.295 67.235 42.420 67.405 ;
        RECT 40.535 66.105 40.705 66.275 ;
        RECT 41.295 66.105 41.465 67.235 ;
        RECT 39.215 65.365 39.385 65.975 ;
        RECT 39.555 65.585 39.885 66.020 ;
        RECT 40.110 65.535 40.365 66.105 ;
        RECT 40.535 65.935 41.465 66.105 ;
        RECT 41.635 66.895 42.645 67.065 ;
        RECT 41.635 66.095 41.805 66.895 ;
        RECT 41.290 65.900 41.465 65.935 ;
        RECT 40.535 65.365 40.865 65.765 ;
        RECT 41.290 65.535 41.820 65.900 ;
        RECT 42.010 65.875 42.285 66.695 ;
        RECT 42.005 65.705 42.285 65.875 ;
        RECT 42.010 65.535 42.285 65.705 ;
        RECT 42.455 65.535 42.645 66.895 ;
        RECT 42.815 66.910 42.985 67.575 ;
        RECT 43.155 67.155 43.325 67.915 ;
        RECT 43.560 67.155 44.075 67.565 ;
        RECT 42.815 66.720 43.565 66.910 ;
        RECT 43.735 66.345 44.075 67.155 ;
        RECT 44.245 66.750 44.535 67.915 ;
        RECT 44.705 66.775 45.090 67.745 ;
        RECT 45.260 67.455 45.585 67.915 ;
        RECT 46.105 67.285 46.385 67.745 ;
        RECT 45.260 67.065 46.385 67.285 ;
        RECT 42.845 66.175 44.075 66.345 ;
        RECT 42.825 65.365 43.335 65.900 ;
        RECT 43.555 65.570 43.800 66.175 ;
        RECT 44.705 66.105 44.985 66.775 ;
        RECT 45.260 66.605 45.710 67.065 ;
        RECT 46.575 66.895 46.975 67.745 ;
        RECT 47.375 67.455 47.645 67.915 ;
        RECT 47.815 67.285 48.100 67.745 ;
        RECT 45.155 66.275 45.710 66.605 ;
        RECT 45.880 66.335 46.975 66.895 ;
        RECT 45.260 66.165 45.710 66.275 ;
        RECT 44.245 65.365 44.535 66.090 ;
        RECT 44.705 65.535 45.090 66.105 ;
        RECT 45.260 65.995 46.385 66.165 ;
        RECT 45.260 65.365 45.585 65.825 ;
        RECT 46.105 65.535 46.385 65.995 ;
        RECT 46.575 65.535 46.975 66.335 ;
        RECT 47.145 67.065 48.100 67.285 ;
        RECT 47.145 66.165 47.355 67.065 ;
        RECT 47.525 66.335 48.215 66.895 ;
        RECT 48.385 66.825 51.895 67.915 ;
        RECT 47.145 65.995 48.100 66.165 ;
        RECT 47.375 65.365 47.645 65.825 ;
        RECT 47.815 65.535 48.100 65.995 ;
        RECT 48.385 66.135 50.035 66.655 ;
        RECT 50.205 66.305 51.895 66.825 ;
        RECT 52.995 66.805 53.290 67.915 ;
        RECT 53.470 66.605 53.720 67.740 ;
        RECT 53.890 66.805 54.150 67.915 ;
        RECT 54.320 67.015 54.580 67.740 ;
        RECT 54.750 67.185 55.010 67.915 ;
        RECT 55.180 67.015 55.440 67.740 ;
        RECT 55.610 67.185 55.870 67.915 ;
        RECT 56.040 67.015 56.300 67.740 ;
        RECT 56.470 67.185 56.730 67.915 ;
        RECT 56.900 67.015 57.160 67.740 ;
        RECT 57.330 67.185 57.625 67.915 ;
        RECT 58.160 67.285 58.445 67.745 ;
        RECT 58.615 67.455 58.885 67.915 ;
        RECT 58.160 67.065 59.115 67.285 ;
        RECT 54.320 66.775 57.630 67.015 ;
        RECT 48.385 65.365 51.895 66.135 ;
        RECT 52.985 65.995 53.300 66.605 ;
        RECT 53.470 66.355 56.490 66.605 ;
        RECT 53.045 65.365 53.290 65.825 ;
        RECT 53.470 65.545 53.720 66.355 ;
        RECT 56.660 66.185 57.630 66.775 ;
        RECT 58.045 66.335 58.735 66.895 ;
        RECT 54.320 66.015 57.630 66.185 ;
        RECT 58.905 66.165 59.115 67.065 ;
        RECT 53.890 65.365 54.150 65.890 ;
        RECT 54.320 65.560 54.580 66.015 ;
        RECT 54.750 65.365 55.010 65.845 ;
        RECT 55.180 65.560 55.440 66.015 ;
        RECT 55.610 65.365 55.870 65.845 ;
        RECT 56.040 65.560 56.300 66.015 ;
        RECT 56.470 65.365 56.730 65.845 ;
        RECT 56.900 65.560 57.160 66.015 ;
        RECT 58.160 65.995 59.115 66.165 ;
        RECT 59.285 66.895 59.685 67.745 ;
        RECT 59.875 67.285 60.155 67.745 ;
        RECT 60.675 67.455 61.000 67.915 ;
        RECT 59.875 67.065 61.000 67.285 ;
        RECT 59.285 66.335 60.380 66.895 ;
        RECT 60.550 66.605 61.000 67.065 ;
        RECT 61.170 66.775 61.555 67.745 ;
        RECT 57.330 65.365 57.630 65.845 ;
        RECT 58.160 65.535 58.445 65.995 ;
        RECT 58.615 65.365 58.885 65.825 ;
        RECT 59.285 65.535 59.685 66.335 ;
        RECT 60.550 66.275 61.105 66.605 ;
        RECT 60.550 66.165 61.000 66.275 ;
        RECT 59.875 65.995 61.000 66.165 ;
        RECT 61.275 66.105 61.555 66.775 ;
        RECT 59.875 65.535 60.155 65.995 ;
        RECT 60.675 65.365 61.000 65.825 ;
        RECT 61.170 65.535 61.555 66.105 ;
        RECT 61.725 67.195 62.185 67.745 ;
        RECT 62.375 67.195 62.705 67.915 ;
        RECT 61.725 65.825 61.975 67.195 ;
        RECT 62.905 67.025 63.205 67.575 ;
        RECT 63.375 67.245 63.655 67.915 ;
        RECT 62.265 66.855 63.205 67.025 ;
        RECT 62.265 66.605 62.435 66.855 ;
        RECT 63.575 66.605 63.840 66.965 ;
        RECT 64.085 66.775 64.295 67.915 ;
        RECT 62.145 66.275 62.435 66.605 ;
        RECT 62.605 66.355 62.945 66.605 ;
        RECT 63.165 66.355 63.840 66.605 ;
        RECT 64.465 66.765 64.795 67.745 ;
        RECT 64.965 66.775 65.195 67.915 ;
        RECT 65.405 66.775 65.685 67.915 ;
        RECT 65.855 66.765 66.185 67.745 ;
        RECT 66.355 66.775 66.615 67.915 ;
        RECT 66.785 67.405 67.975 67.695 ;
        RECT 66.805 67.065 67.975 67.235 ;
        RECT 68.145 67.115 68.425 67.915 ;
        RECT 66.805 66.775 67.130 67.065 ;
        RECT 67.805 66.945 67.975 67.065 ;
        RECT 62.265 66.185 62.435 66.275 ;
        RECT 62.265 65.995 63.655 66.185 ;
        RECT 61.725 65.535 62.285 65.825 ;
        RECT 62.455 65.365 62.705 65.825 ;
        RECT 63.325 65.635 63.655 65.995 ;
        RECT 64.085 65.365 64.295 66.185 ;
        RECT 64.465 66.165 64.715 66.765 ;
        RECT 64.885 66.355 65.215 66.605 ;
        RECT 65.415 66.335 65.750 66.605 ;
        RECT 64.465 65.535 64.795 66.165 ;
        RECT 64.965 65.365 65.195 66.185 ;
        RECT 65.920 66.165 66.090 66.765 ;
        RECT 67.300 66.605 67.495 66.895 ;
        RECT 67.805 66.775 68.465 66.945 ;
        RECT 68.635 66.775 68.910 67.745 ;
        RECT 68.295 66.605 68.465 66.775 ;
        RECT 66.260 66.355 66.595 66.605 ;
        RECT 66.785 66.275 67.130 66.605 ;
        RECT 67.300 66.275 68.125 66.605 ;
        RECT 68.295 66.275 68.570 66.605 ;
        RECT 65.405 65.365 65.715 66.165 ;
        RECT 65.920 65.535 66.615 66.165 ;
        RECT 68.295 66.105 68.465 66.275 ;
        RECT 66.800 65.935 68.465 66.105 ;
        RECT 68.740 66.040 68.910 66.775 ;
        RECT 70.005 66.750 70.295 67.915 ;
        RECT 71.390 67.525 71.725 67.745 ;
        RECT 72.730 67.535 73.085 67.915 ;
        RECT 71.390 66.905 71.645 67.525 ;
        RECT 71.895 67.365 72.125 67.405 ;
        RECT 73.255 67.365 73.505 67.745 ;
        RECT 71.895 67.165 73.505 67.365 ;
        RECT 71.895 67.075 72.080 67.165 ;
        RECT 72.670 67.155 73.505 67.165 ;
        RECT 73.755 67.135 74.005 67.915 ;
        RECT 74.175 67.065 74.435 67.745 ;
        RECT 72.235 66.965 72.565 66.995 ;
        RECT 72.235 66.905 74.035 66.965 ;
        RECT 71.390 66.795 74.095 66.905 ;
        RECT 71.390 66.735 72.565 66.795 ;
        RECT 73.895 66.760 74.095 66.795 ;
        RECT 71.385 66.355 71.875 66.555 ;
        RECT 72.065 66.355 72.540 66.565 ;
        RECT 66.800 65.585 67.055 65.935 ;
        RECT 67.225 65.365 67.555 65.765 ;
        RECT 67.725 65.585 67.895 65.935 ;
        RECT 68.065 65.365 68.445 65.765 ;
        RECT 68.635 65.695 68.910 66.040 ;
        RECT 70.005 65.365 70.295 66.090 ;
        RECT 71.390 65.365 71.845 66.130 ;
        RECT 72.320 65.955 72.540 66.355 ;
        RECT 72.785 66.355 73.115 66.565 ;
        RECT 72.785 65.955 72.995 66.355 ;
        RECT 73.285 66.320 73.695 66.625 ;
        RECT 73.925 66.185 74.095 66.760 ;
        RECT 73.825 66.065 74.095 66.185 ;
        RECT 73.250 66.020 74.095 66.065 ;
        RECT 73.250 65.895 74.005 66.020 ;
        RECT 73.250 65.745 73.420 65.895 ;
        RECT 74.265 65.875 74.435 67.065 ;
        RECT 74.605 66.825 77.195 67.915 ;
        RECT 74.205 65.865 74.435 65.875 ;
        RECT 72.120 65.535 73.420 65.745 ;
        RECT 73.675 65.365 74.005 65.725 ;
        RECT 74.175 65.535 74.435 65.865 ;
        RECT 74.605 66.135 75.815 66.655 ;
        RECT 75.985 66.305 77.195 66.825 ;
        RECT 77.370 66.765 77.630 67.915 ;
        RECT 77.805 66.840 78.060 67.745 ;
        RECT 78.230 67.155 78.560 67.915 ;
        RECT 78.775 66.985 78.945 67.745 ;
        RECT 74.605 65.365 77.195 66.135 ;
        RECT 77.370 65.365 77.630 66.205 ;
        RECT 77.805 66.110 77.975 66.840 ;
        RECT 78.230 66.815 78.945 66.985 ;
        RECT 78.230 66.605 78.400 66.815 ;
        RECT 79.205 66.775 79.590 67.745 ;
        RECT 79.760 67.455 80.085 67.915 ;
        RECT 80.605 67.285 80.885 67.745 ;
        RECT 79.760 67.065 80.885 67.285 ;
        RECT 78.145 66.275 78.400 66.605 ;
        RECT 77.805 65.535 78.060 66.110 ;
        RECT 78.230 66.085 78.400 66.275 ;
        RECT 78.680 66.265 79.035 66.635 ;
        RECT 79.205 66.105 79.485 66.775 ;
        RECT 79.760 66.605 80.210 67.065 ;
        RECT 81.075 66.895 81.475 67.745 ;
        RECT 81.875 67.455 82.145 67.915 ;
        RECT 82.315 67.285 82.600 67.745 ;
        RECT 79.655 66.275 80.210 66.605 ;
        RECT 80.380 66.335 81.475 66.895 ;
        RECT 79.760 66.165 80.210 66.275 ;
        RECT 78.230 65.915 78.945 66.085 ;
        RECT 78.230 65.365 78.560 65.745 ;
        RECT 78.775 65.535 78.945 65.915 ;
        RECT 79.205 65.535 79.590 66.105 ;
        RECT 79.760 65.995 80.885 66.165 ;
        RECT 79.760 65.365 80.085 65.825 ;
        RECT 80.605 65.535 80.885 65.995 ;
        RECT 81.075 65.535 81.475 66.335 ;
        RECT 81.645 67.065 82.600 67.285 ;
        RECT 81.645 66.165 81.855 67.065 ;
        RECT 82.025 66.335 82.715 66.895 ;
        RECT 82.885 66.825 84.095 67.915 ;
        RECT 82.885 66.285 83.405 66.825 ;
        RECT 81.645 65.995 82.600 66.165 ;
        RECT 83.575 66.115 84.095 66.655 ;
        RECT 81.875 65.365 82.145 65.825 ;
        RECT 82.315 65.535 82.600 65.995 ;
        RECT 82.885 65.365 84.095 66.115 ;
        RECT 5.520 65.195 84.180 65.365 ;
        RECT 5.605 64.445 6.815 65.195 ;
        RECT 5.605 63.905 6.125 64.445 ;
        RECT 6.990 64.355 7.250 65.195 ;
        RECT 7.425 64.450 7.680 65.025 ;
        RECT 7.850 64.815 8.180 65.195 ;
        RECT 8.395 64.645 8.565 65.025 ;
        RECT 7.850 64.475 8.565 64.645 ;
        RECT 9.835 64.645 10.005 64.935 ;
        RECT 10.175 64.815 10.505 65.195 ;
        RECT 9.835 64.475 10.500 64.645 ;
        RECT 6.295 63.735 6.815 64.275 ;
        RECT 5.605 62.645 6.815 63.735 ;
        RECT 6.990 62.645 7.250 63.795 ;
        RECT 7.425 63.720 7.595 64.450 ;
        RECT 7.850 64.285 8.020 64.475 ;
        RECT 7.765 63.955 8.020 64.285 ;
        RECT 7.850 63.745 8.020 63.955 ;
        RECT 8.300 63.925 8.655 64.295 ;
        RECT 7.425 62.815 7.680 63.720 ;
        RECT 7.850 63.575 8.565 63.745 ;
        RECT 9.750 63.655 10.100 64.305 ;
        RECT 7.850 62.645 8.180 63.405 ;
        RECT 8.395 62.815 8.565 63.575 ;
        RECT 10.270 63.485 10.500 64.475 ;
        RECT 9.835 63.315 10.500 63.485 ;
        RECT 9.835 62.815 10.005 63.315 ;
        RECT 10.175 62.645 10.505 63.145 ;
        RECT 10.675 62.815 10.860 64.935 ;
        RECT 11.115 64.735 11.365 65.195 ;
        RECT 11.535 64.745 11.870 64.915 ;
        RECT 12.065 64.745 12.740 64.915 ;
        RECT 11.535 64.605 11.705 64.745 ;
        RECT 11.030 63.615 11.310 64.565 ;
        RECT 11.480 64.475 11.705 64.605 ;
        RECT 11.480 63.370 11.650 64.475 ;
        RECT 11.875 64.325 12.400 64.545 ;
        RECT 11.820 63.560 12.060 64.155 ;
        RECT 12.230 63.625 12.400 64.325 ;
        RECT 12.570 63.965 12.740 64.745 ;
        RECT 13.060 64.695 13.430 65.195 ;
        RECT 13.610 64.745 14.015 64.915 ;
        RECT 14.185 64.745 14.970 64.915 ;
        RECT 13.610 64.515 13.780 64.745 ;
        RECT 12.950 64.215 13.780 64.515 ;
        RECT 14.165 64.245 14.630 64.575 ;
        RECT 12.950 64.185 13.150 64.215 ;
        RECT 13.270 63.965 13.440 64.035 ;
        RECT 12.570 63.795 13.440 63.965 ;
        RECT 12.930 63.705 13.440 63.795 ;
        RECT 11.480 63.240 11.785 63.370 ;
        RECT 12.230 63.260 12.760 63.625 ;
        RECT 11.100 62.645 11.365 63.105 ;
        RECT 11.535 62.815 11.785 63.240 ;
        RECT 12.930 63.090 13.100 63.705 ;
        RECT 11.995 62.920 13.100 63.090 ;
        RECT 13.270 62.645 13.440 63.445 ;
        RECT 13.610 63.145 13.780 64.215 ;
        RECT 13.950 63.315 14.140 64.035 ;
        RECT 14.310 63.285 14.630 64.245 ;
        RECT 14.800 64.285 14.970 64.745 ;
        RECT 15.245 64.665 15.455 65.195 ;
        RECT 15.715 64.455 16.045 64.980 ;
        RECT 16.215 64.585 16.385 65.195 ;
        RECT 16.555 64.540 16.885 64.975 ;
        RECT 17.055 64.680 17.225 65.195 ;
        RECT 16.555 64.455 16.935 64.540 ;
        RECT 15.845 64.285 16.045 64.455 ;
        RECT 16.710 64.415 16.935 64.455 ;
        RECT 14.800 63.955 15.675 64.285 ;
        RECT 15.845 63.955 16.595 64.285 ;
        RECT 13.610 62.815 13.860 63.145 ;
        RECT 14.800 63.115 14.970 63.955 ;
        RECT 15.845 63.750 16.035 63.955 ;
        RECT 16.765 63.835 16.935 64.415 ;
        RECT 17.840 64.385 18.085 64.990 ;
        RECT 18.305 64.660 18.815 65.195 ;
        RECT 16.720 63.785 16.935 63.835 ;
        RECT 15.140 63.375 16.035 63.750 ;
        RECT 16.545 63.705 16.935 63.785 ;
        RECT 17.565 64.215 18.795 64.385 ;
        RECT 14.085 62.945 14.970 63.115 ;
        RECT 15.150 62.645 15.465 63.145 ;
        RECT 15.695 62.815 16.035 63.375 ;
        RECT 16.205 62.645 16.375 63.655 ;
        RECT 16.545 62.860 16.875 63.705 ;
        RECT 17.045 62.645 17.215 63.560 ;
        RECT 17.565 63.405 17.905 64.215 ;
        RECT 18.075 63.650 18.825 63.840 ;
        RECT 17.565 62.995 18.080 63.405 ;
        RECT 18.315 62.645 18.485 63.405 ;
        RECT 18.655 62.985 18.825 63.650 ;
        RECT 18.995 63.665 19.185 65.025 ;
        RECT 19.355 64.855 19.630 65.025 ;
        RECT 19.355 64.685 19.635 64.855 ;
        RECT 19.355 63.865 19.630 64.685 ;
        RECT 19.820 64.660 20.350 65.025 ;
        RECT 20.775 64.795 21.105 65.195 ;
        RECT 20.175 64.625 20.350 64.660 ;
        RECT 19.835 63.665 20.005 64.465 ;
        RECT 18.995 63.495 20.005 63.665 ;
        RECT 20.175 64.455 21.105 64.625 ;
        RECT 21.275 64.455 21.530 65.025 ;
        RECT 21.705 64.650 27.050 65.195 ;
        RECT 20.175 63.325 20.345 64.455 ;
        RECT 20.935 64.285 21.105 64.455 ;
        RECT 19.220 63.155 20.345 63.325 ;
        RECT 20.515 63.955 20.710 64.285 ;
        RECT 20.935 63.955 21.190 64.285 ;
        RECT 20.515 62.985 20.685 63.955 ;
        RECT 21.360 63.785 21.530 64.455 ;
        RECT 23.290 63.820 23.630 64.650 ;
        RECT 27.225 64.425 30.735 65.195 ;
        RECT 31.365 64.470 31.655 65.195 ;
        RECT 32.285 64.455 32.670 65.025 ;
        RECT 32.840 64.735 33.165 65.195 ;
        RECT 33.685 64.565 33.965 65.025 ;
        RECT 18.655 62.815 20.685 62.985 ;
        RECT 20.855 62.645 21.025 63.785 ;
        RECT 21.195 62.815 21.530 63.785 ;
        RECT 25.110 63.080 25.460 64.330 ;
        RECT 27.225 63.905 28.875 64.425 ;
        RECT 29.045 63.735 30.735 64.255 ;
        RECT 21.705 62.645 27.050 63.080 ;
        RECT 27.225 62.645 30.735 63.735 ;
        RECT 31.365 62.645 31.655 63.810 ;
        RECT 32.285 63.785 32.565 64.455 ;
        RECT 32.840 64.395 33.965 64.565 ;
        RECT 32.840 64.285 33.290 64.395 ;
        RECT 32.735 63.955 33.290 64.285 ;
        RECT 34.155 64.225 34.555 65.025 ;
        RECT 34.955 64.735 35.225 65.195 ;
        RECT 35.395 64.565 35.680 65.025 ;
        RECT 32.285 62.815 32.670 63.785 ;
        RECT 32.840 63.495 33.290 63.955 ;
        RECT 33.460 63.665 34.555 64.225 ;
        RECT 32.840 63.275 33.965 63.495 ;
        RECT 32.840 62.645 33.165 63.105 ;
        RECT 33.685 62.815 33.965 63.275 ;
        RECT 34.155 62.815 34.555 63.665 ;
        RECT 34.725 64.395 35.680 64.565 ;
        RECT 36.015 64.655 36.240 65.015 ;
        RECT 36.420 64.825 36.750 65.195 ;
        RECT 36.930 64.655 37.185 65.015 ;
        RECT 37.750 64.825 38.495 65.195 ;
        RECT 36.015 64.465 38.500 64.655 ;
        RECT 34.725 63.495 34.935 64.395 ;
        RECT 35.105 63.665 35.795 64.225 ;
        RECT 35.975 63.955 36.245 64.285 ;
        RECT 36.425 63.955 36.860 64.285 ;
        RECT 37.040 63.955 37.615 64.285 ;
        RECT 37.795 63.955 38.075 64.285 ;
        RECT 38.275 63.775 38.500 64.465 ;
        RECT 36.005 63.595 38.500 63.775 ;
        RECT 38.675 63.595 39.010 65.015 ;
        RECT 39.185 64.445 40.395 65.195 ;
        RECT 40.565 64.455 40.950 65.025 ;
        RECT 41.120 64.735 41.445 65.195 ;
        RECT 41.965 64.565 42.245 65.025 ;
        RECT 39.185 63.905 39.705 64.445 ;
        RECT 39.875 63.735 40.395 64.275 ;
        RECT 34.725 63.275 35.680 63.495 ;
        RECT 34.955 62.645 35.225 63.105 ;
        RECT 35.395 62.815 35.680 63.275 ;
        RECT 36.005 62.825 36.295 63.595 ;
        RECT 36.865 63.185 38.055 63.415 ;
        RECT 36.865 62.825 37.125 63.185 ;
        RECT 37.295 62.645 37.625 63.015 ;
        RECT 37.795 62.825 38.055 63.185 ;
        RECT 38.245 62.645 38.575 63.365 ;
        RECT 38.745 62.825 39.010 63.595 ;
        RECT 39.185 62.645 40.395 63.735 ;
        RECT 40.565 63.785 40.845 64.455 ;
        RECT 41.120 64.395 42.245 64.565 ;
        RECT 41.120 64.285 41.570 64.395 ;
        RECT 41.015 63.955 41.570 64.285 ;
        RECT 42.435 64.225 42.835 65.025 ;
        RECT 43.235 64.735 43.505 65.195 ;
        RECT 43.675 64.565 43.960 65.025 ;
        RECT 40.565 62.815 40.950 63.785 ;
        RECT 41.120 63.495 41.570 63.955 ;
        RECT 41.740 63.665 42.835 64.225 ;
        RECT 41.120 63.275 42.245 63.495 ;
        RECT 41.120 62.645 41.445 63.105 ;
        RECT 41.965 62.815 42.245 63.275 ;
        RECT 42.435 62.815 42.835 63.665 ;
        RECT 43.005 64.395 43.960 64.565 ;
        RECT 45.170 64.455 45.425 65.025 ;
        RECT 45.595 64.795 45.925 65.195 ;
        RECT 46.350 64.660 46.880 65.025 ;
        RECT 46.350 64.625 46.525 64.660 ;
        RECT 45.595 64.455 46.525 64.625 ;
        RECT 43.005 63.495 43.215 64.395 ;
        RECT 43.385 63.665 44.075 64.225 ;
        RECT 45.170 63.785 45.340 64.455 ;
        RECT 45.595 64.285 45.765 64.455 ;
        RECT 45.510 63.955 45.765 64.285 ;
        RECT 45.990 63.955 46.185 64.285 ;
        RECT 43.005 63.275 43.960 63.495 ;
        RECT 43.235 62.645 43.505 63.105 ;
        RECT 43.675 62.815 43.960 63.275 ;
        RECT 45.170 62.815 45.505 63.785 ;
        RECT 45.675 62.645 45.845 63.785 ;
        RECT 46.015 62.985 46.185 63.955 ;
        RECT 46.355 63.325 46.525 64.455 ;
        RECT 46.695 63.665 46.865 64.465 ;
        RECT 47.070 64.175 47.345 65.025 ;
        RECT 47.065 64.005 47.345 64.175 ;
        RECT 47.070 63.865 47.345 64.005 ;
        RECT 47.515 63.665 47.705 65.025 ;
        RECT 47.885 64.660 48.395 65.195 ;
        RECT 48.615 64.385 48.860 64.990 ;
        RECT 49.355 64.540 49.685 64.975 ;
        RECT 49.855 64.585 50.025 65.195 ;
        RECT 49.305 64.455 49.685 64.540 ;
        RECT 50.195 64.455 50.525 64.980 ;
        RECT 50.785 64.665 50.995 65.195 ;
        RECT 51.270 64.745 52.055 64.915 ;
        RECT 52.225 64.745 52.630 64.915 ;
        RECT 49.305 64.415 49.530 64.455 ;
        RECT 47.905 64.215 49.135 64.385 ;
        RECT 46.695 63.495 47.705 63.665 ;
        RECT 47.875 63.650 48.625 63.840 ;
        RECT 46.355 63.155 47.480 63.325 ;
        RECT 47.875 62.985 48.045 63.650 ;
        RECT 48.795 63.405 49.135 64.215 ;
        RECT 49.305 63.835 49.475 64.415 ;
        RECT 50.195 64.285 50.395 64.455 ;
        RECT 51.270 64.285 51.440 64.745 ;
        RECT 49.645 63.955 50.395 64.285 ;
        RECT 50.565 63.955 51.440 64.285 ;
        RECT 49.305 63.785 49.520 63.835 ;
        RECT 49.305 63.705 49.695 63.785 ;
        RECT 46.015 62.815 48.045 62.985 ;
        RECT 48.215 62.645 48.385 63.405 ;
        RECT 48.620 62.995 49.135 63.405 ;
        RECT 49.365 62.860 49.695 63.705 ;
        RECT 50.205 63.750 50.395 63.955 ;
        RECT 49.865 62.645 50.035 63.655 ;
        RECT 50.205 63.375 51.100 63.750 ;
        RECT 50.205 62.815 50.545 63.375 ;
        RECT 50.775 62.645 51.090 63.145 ;
        RECT 51.270 63.115 51.440 63.955 ;
        RECT 51.610 64.245 52.075 64.575 ;
        RECT 52.460 64.515 52.630 64.745 ;
        RECT 52.810 64.695 53.180 65.195 ;
        RECT 53.500 64.745 54.175 64.915 ;
        RECT 54.370 64.745 54.705 64.915 ;
        RECT 51.610 63.285 51.930 64.245 ;
        RECT 52.460 64.215 53.290 64.515 ;
        RECT 52.100 63.315 52.290 64.035 ;
        RECT 52.460 63.145 52.630 64.215 ;
        RECT 53.090 64.185 53.290 64.215 ;
        RECT 52.800 63.965 52.970 64.035 ;
        RECT 53.500 63.965 53.670 64.745 ;
        RECT 54.535 64.605 54.705 64.745 ;
        RECT 54.875 64.735 55.125 65.195 ;
        RECT 52.800 63.795 53.670 63.965 ;
        RECT 53.840 64.325 54.365 64.545 ;
        RECT 54.535 64.475 54.760 64.605 ;
        RECT 52.800 63.705 53.310 63.795 ;
        RECT 51.270 62.945 52.155 63.115 ;
        RECT 52.380 62.815 52.630 63.145 ;
        RECT 52.800 62.645 52.970 63.445 ;
        RECT 53.140 63.090 53.310 63.705 ;
        RECT 53.840 63.625 54.010 64.325 ;
        RECT 53.480 63.260 54.010 63.625 ;
        RECT 54.180 63.560 54.420 64.155 ;
        RECT 54.590 63.370 54.760 64.475 ;
        RECT 54.930 63.615 55.210 64.565 ;
        RECT 54.455 63.240 54.760 63.370 ;
        RECT 53.140 62.920 54.245 63.090 ;
        RECT 54.455 62.815 54.705 63.240 ;
        RECT 54.875 62.645 55.140 63.105 ;
        RECT 55.380 62.815 55.565 64.935 ;
        RECT 55.735 64.815 56.065 65.195 ;
        RECT 56.235 64.645 56.405 64.935 ;
        RECT 55.740 64.475 56.405 64.645 ;
        RECT 55.740 63.485 55.970 64.475 ;
        RECT 57.125 64.470 57.415 65.195 ;
        RECT 57.590 64.455 57.845 65.025 ;
        RECT 58.015 64.795 58.345 65.195 ;
        RECT 58.770 64.660 59.300 65.025 ;
        RECT 59.490 64.855 59.765 65.025 ;
        RECT 59.485 64.685 59.765 64.855 ;
        RECT 58.770 64.625 58.945 64.660 ;
        RECT 58.015 64.455 58.945 64.625 ;
        RECT 56.140 63.655 56.490 64.305 ;
        RECT 55.740 63.315 56.405 63.485 ;
        RECT 55.735 62.645 56.065 63.145 ;
        RECT 56.235 62.815 56.405 63.315 ;
        RECT 57.125 62.645 57.415 63.810 ;
        RECT 57.590 63.785 57.760 64.455 ;
        RECT 58.015 64.285 58.185 64.455 ;
        RECT 57.930 63.955 58.185 64.285 ;
        RECT 58.410 63.955 58.605 64.285 ;
        RECT 57.590 62.815 57.925 63.785 ;
        RECT 58.095 62.645 58.265 63.785 ;
        RECT 58.435 62.985 58.605 63.955 ;
        RECT 58.775 63.325 58.945 64.455 ;
        RECT 59.115 63.665 59.285 64.465 ;
        RECT 59.490 63.865 59.765 64.685 ;
        RECT 59.935 63.665 60.125 65.025 ;
        RECT 60.305 64.660 60.815 65.195 ;
        RECT 61.035 64.385 61.280 64.990 ;
        RECT 61.725 64.425 64.315 65.195 ;
        RECT 64.960 64.625 65.215 64.975 ;
        RECT 65.385 64.795 65.715 65.195 ;
        RECT 65.885 64.625 66.055 64.975 ;
        RECT 66.225 64.795 66.605 65.195 ;
        RECT 64.960 64.455 66.625 64.625 ;
        RECT 66.795 64.520 67.070 64.865 ;
        RECT 60.325 64.215 61.555 64.385 ;
        RECT 59.115 63.495 60.125 63.665 ;
        RECT 60.295 63.650 61.045 63.840 ;
        RECT 58.775 63.155 59.900 63.325 ;
        RECT 60.295 62.985 60.465 63.650 ;
        RECT 61.215 63.405 61.555 64.215 ;
        RECT 61.725 63.905 62.935 64.425 ;
        RECT 66.455 64.285 66.625 64.455 ;
        RECT 63.105 63.735 64.315 64.255 ;
        RECT 64.945 63.955 65.290 64.285 ;
        RECT 65.460 63.955 66.285 64.285 ;
        RECT 66.455 63.955 66.730 64.285 ;
        RECT 58.435 62.815 60.465 62.985 ;
        RECT 60.635 62.645 60.805 63.405 ;
        RECT 61.040 62.995 61.555 63.405 ;
        RECT 61.725 62.645 64.315 63.735 ;
        RECT 64.965 63.495 65.290 63.785 ;
        RECT 65.460 63.665 65.655 63.955 ;
        RECT 66.455 63.785 66.625 63.955 ;
        RECT 66.900 63.785 67.070 64.520 ;
        RECT 67.450 64.415 67.950 65.025 ;
        RECT 67.245 63.955 67.595 64.205 ;
        RECT 67.780 63.785 67.950 64.415 ;
        RECT 68.580 64.545 68.910 65.025 ;
        RECT 69.080 64.735 69.305 65.195 ;
        RECT 69.475 64.545 69.805 65.025 ;
        RECT 68.580 64.375 69.805 64.545 ;
        RECT 69.995 64.395 70.245 65.195 ;
        RECT 70.415 64.395 70.755 65.025 ;
        RECT 70.930 64.430 71.385 65.195 ;
        RECT 71.660 64.815 72.960 65.025 ;
        RECT 73.215 64.835 73.545 65.195 ;
        RECT 72.790 64.665 72.960 64.815 ;
        RECT 73.715 64.695 73.975 65.025 ;
        RECT 68.120 64.005 68.450 64.205 ;
        RECT 68.620 64.005 68.950 64.205 ;
        RECT 69.120 64.005 69.540 64.205 ;
        RECT 69.715 64.035 70.410 64.205 ;
        RECT 69.715 63.785 69.885 64.035 ;
        RECT 70.580 63.785 70.755 64.395 ;
        RECT 71.860 64.205 72.080 64.605 ;
        RECT 70.925 64.005 71.415 64.205 ;
        RECT 71.605 63.995 72.080 64.205 ;
        RECT 72.325 64.205 72.535 64.605 ;
        RECT 72.790 64.540 73.545 64.665 ;
        RECT 72.790 64.495 73.635 64.540 ;
        RECT 73.365 64.375 73.635 64.495 ;
        RECT 72.325 63.995 72.655 64.205 ;
        RECT 72.825 63.935 73.235 64.240 ;
        RECT 65.965 63.615 66.625 63.785 ;
        RECT 65.965 63.495 66.135 63.615 ;
        RECT 64.965 63.325 66.135 63.495 ;
        RECT 64.945 62.865 66.135 63.155 ;
        RECT 66.305 62.645 66.585 63.445 ;
        RECT 66.795 62.815 67.070 63.785 ;
        RECT 67.450 63.615 69.885 63.785 ;
        RECT 67.450 62.815 67.780 63.615 ;
        RECT 67.950 62.645 68.280 63.445 ;
        RECT 68.580 62.815 68.910 63.615 ;
        RECT 69.555 62.645 69.805 63.445 ;
        RECT 70.075 62.645 70.245 63.785 ;
        RECT 70.415 62.815 70.755 63.785 ;
        RECT 70.930 63.765 72.105 63.825 ;
        RECT 73.465 63.800 73.635 64.375 ;
        RECT 73.435 63.765 73.635 63.800 ;
        RECT 70.930 63.655 73.635 63.765 ;
        RECT 70.930 63.035 71.185 63.655 ;
        RECT 71.775 63.595 73.575 63.655 ;
        RECT 71.775 63.565 72.105 63.595 ;
        RECT 73.805 63.495 73.975 64.695 ;
        RECT 74.235 64.645 74.405 64.935 ;
        RECT 74.575 64.815 74.905 65.195 ;
        RECT 74.235 64.475 74.900 64.645 ;
        RECT 74.150 63.655 74.500 64.305 ;
        RECT 71.435 63.395 71.620 63.485 ;
        RECT 72.210 63.395 73.045 63.405 ;
        RECT 71.435 63.195 73.045 63.395 ;
        RECT 71.435 63.155 71.665 63.195 ;
        RECT 70.930 62.815 71.265 63.035 ;
        RECT 72.270 62.645 72.625 63.025 ;
        RECT 72.795 62.815 73.045 63.195 ;
        RECT 73.295 62.645 73.545 63.425 ;
        RECT 73.715 62.815 73.975 63.495 ;
        RECT 74.670 63.485 74.900 64.475 ;
        RECT 74.235 63.315 74.900 63.485 ;
        RECT 74.235 62.815 74.405 63.315 ;
        RECT 74.575 62.645 74.905 63.145 ;
        RECT 75.075 62.815 75.260 64.935 ;
        RECT 75.515 64.735 75.765 65.195 ;
        RECT 75.935 64.745 76.270 64.915 ;
        RECT 76.465 64.745 77.140 64.915 ;
        RECT 75.935 64.605 76.105 64.745 ;
        RECT 75.430 63.615 75.710 64.565 ;
        RECT 75.880 64.475 76.105 64.605 ;
        RECT 75.880 63.370 76.050 64.475 ;
        RECT 76.275 64.325 76.800 64.545 ;
        RECT 76.220 63.560 76.460 64.155 ;
        RECT 76.630 63.625 76.800 64.325 ;
        RECT 76.970 63.965 77.140 64.745 ;
        RECT 77.460 64.695 77.830 65.195 ;
        RECT 78.010 64.745 78.415 64.915 ;
        RECT 78.585 64.745 79.370 64.915 ;
        RECT 78.010 64.515 78.180 64.745 ;
        RECT 77.350 64.215 78.180 64.515 ;
        RECT 78.565 64.245 79.030 64.575 ;
        RECT 77.350 64.185 77.550 64.215 ;
        RECT 77.670 63.965 77.840 64.035 ;
        RECT 76.970 63.795 77.840 63.965 ;
        RECT 77.330 63.705 77.840 63.795 ;
        RECT 75.880 63.240 76.185 63.370 ;
        RECT 76.630 63.260 77.160 63.625 ;
        RECT 75.500 62.645 75.765 63.105 ;
        RECT 75.935 62.815 76.185 63.240 ;
        RECT 77.330 63.090 77.500 63.705 ;
        RECT 76.395 62.920 77.500 63.090 ;
        RECT 77.670 62.645 77.840 63.445 ;
        RECT 78.010 63.145 78.180 64.215 ;
        RECT 78.350 63.315 78.540 64.035 ;
        RECT 78.710 63.285 79.030 64.245 ;
        RECT 79.200 64.285 79.370 64.745 ;
        RECT 79.645 64.665 79.855 65.195 ;
        RECT 80.115 64.455 80.445 64.980 ;
        RECT 80.615 64.585 80.785 65.195 ;
        RECT 80.955 64.540 81.285 64.975 ;
        RECT 80.955 64.455 81.335 64.540 ;
        RECT 80.245 64.285 80.445 64.455 ;
        RECT 81.110 64.415 81.335 64.455 ;
        RECT 79.200 63.955 80.075 64.285 ;
        RECT 80.245 63.955 80.995 64.285 ;
        RECT 78.010 62.815 78.260 63.145 ;
        RECT 79.200 63.115 79.370 63.955 ;
        RECT 80.245 63.750 80.435 63.955 ;
        RECT 81.165 63.835 81.335 64.415 ;
        RECT 81.120 63.785 81.335 63.835 ;
        RECT 79.540 63.375 80.435 63.750 ;
        RECT 80.945 63.705 81.335 63.785 ;
        RECT 81.505 64.520 81.765 65.025 ;
        RECT 81.945 64.815 82.275 65.195 ;
        RECT 82.455 64.645 82.625 65.025 ;
        RECT 81.505 63.720 81.675 64.520 ;
        RECT 81.960 64.475 82.625 64.645 ;
        RECT 81.960 64.220 82.130 64.475 ;
        RECT 82.885 64.445 84.095 65.195 ;
        RECT 81.845 63.890 82.130 64.220 ;
        RECT 82.365 63.925 82.695 64.295 ;
        RECT 81.960 63.745 82.130 63.890 ;
        RECT 78.485 62.945 79.370 63.115 ;
        RECT 79.550 62.645 79.865 63.145 ;
        RECT 80.095 62.815 80.435 63.375 ;
        RECT 80.605 62.645 80.775 63.655 ;
        RECT 80.945 62.860 81.275 63.705 ;
        RECT 81.505 62.815 81.775 63.720 ;
        RECT 81.960 63.575 82.625 63.745 ;
        RECT 81.945 62.645 82.275 63.405 ;
        RECT 82.455 62.815 82.625 63.575 ;
        RECT 82.885 63.735 83.405 64.275 ;
        RECT 83.575 63.905 84.095 64.445 ;
        RECT 82.885 62.645 84.095 63.735 ;
        RECT 5.520 62.475 84.180 62.645 ;
        RECT 5.605 61.385 6.815 62.475 ;
        RECT 5.605 60.675 6.125 61.215 ;
        RECT 6.295 60.845 6.815 61.385 ;
        RECT 6.990 61.325 7.250 62.475 ;
        RECT 7.425 61.400 7.680 62.305 ;
        RECT 7.850 61.715 8.180 62.475 ;
        RECT 8.395 61.545 8.565 62.305 ;
        RECT 5.605 59.925 6.815 60.675 ;
        RECT 6.990 59.925 7.250 60.765 ;
        RECT 7.425 60.670 7.595 61.400 ;
        RECT 7.850 61.375 8.565 61.545 ;
        RECT 7.850 61.165 8.020 61.375 ;
        RECT 8.830 61.325 9.090 62.475 ;
        RECT 9.265 61.400 9.520 62.305 ;
        RECT 9.690 61.715 10.020 62.475 ;
        RECT 10.235 61.545 10.405 62.305 ;
        RECT 7.765 60.835 8.020 61.165 ;
        RECT 7.425 60.095 7.680 60.670 ;
        RECT 7.850 60.645 8.020 60.835 ;
        RECT 8.300 60.825 8.655 61.195 ;
        RECT 7.850 60.475 8.565 60.645 ;
        RECT 7.850 59.925 8.180 60.305 ;
        RECT 8.395 60.095 8.565 60.475 ;
        RECT 8.830 59.925 9.090 60.765 ;
        RECT 9.265 60.670 9.435 61.400 ;
        RECT 9.690 61.375 10.405 61.545 ;
        RECT 10.665 61.385 11.875 62.475 ;
        RECT 9.690 61.165 9.860 61.375 ;
        RECT 9.605 60.835 9.860 61.165 ;
        RECT 9.265 60.095 9.520 60.670 ;
        RECT 9.690 60.645 9.860 60.835 ;
        RECT 10.140 60.825 10.495 61.195 ;
        RECT 10.665 60.675 11.185 61.215 ;
        RECT 11.355 60.845 11.875 61.385 ;
        RECT 12.050 61.325 12.310 62.475 ;
        RECT 12.485 61.400 12.740 62.305 ;
        RECT 12.910 61.715 13.240 62.475 ;
        RECT 13.455 61.545 13.625 62.305 ;
        RECT 9.690 60.475 10.405 60.645 ;
        RECT 9.690 59.925 10.020 60.305 ;
        RECT 10.235 60.095 10.405 60.475 ;
        RECT 10.665 59.925 11.875 60.675 ;
        RECT 12.050 59.925 12.310 60.765 ;
        RECT 12.485 60.670 12.655 61.400 ;
        RECT 12.910 61.375 13.625 61.545 ;
        RECT 13.885 61.385 17.395 62.475 ;
        RECT 12.910 61.165 13.080 61.375 ;
        RECT 12.825 60.835 13.080 61.165 ;
        RECT 12.485 60.095 12.740 60.670 ;
        RECT 12.910 60.645 13.080 60.835 ;
        RECT 13.360 60.825 13.715 61.195 ;
        RECT 13.885 60.695 15.535 61.215 ;
        RECT 15.705 60.865 17.395 61.385 ;
        RECT 18.485 61.310 18.775 62.475 ;
        RECT 18.945 61.335 19.285 62.305 ;
        RECT 19.455 61.335 19.625 62.475 ;
        RECT 19.895 61.675 20.145 62.475 ;
        RECT 20.790 61.505 21.120 62.305 ;
        RECT 21.420 61.675 21.750 62.475 ;
        RECT 21.920 61.505 22.250 62.305 ;
        RECT 19.815 61.335 22.250 61.505 ;
        RECT 22.810 61.505 23.200 61.680 ;
        RECT 23.685 61.675 24.015 62.475 ;
        RECT 24.185 61.685 24.720 62.305 ;
        RECT 22.810 61.335 24.235 61.505 ;
        RECT 18.945 60.725 19.120 61.335 ;
        RECT 19.815 61.085 19.985 61.335 ;
        RECT 19.290 60.915 19.985 61.085 ;
        RECT 20.160 60.915 20.580 61.115 ;
        RECT 20.750 60.915 21.080 61.115 ;
        RECT 21.250 60.915 21.580 61.115 ;
        RECT 12.910 60.475 13.625 60.645 ;
        RECT 12.910 59.925 13.240 60.305 ;
        RECT 13.455 60.095 13.625 60.475 ;
        RECT 13.885 59.925 17.395 60.695 ;
        RECT 18.485 59.925 18.775 60.650 ;
        RECT 18.945 60.095 19.285 60.725 ;
        RECT 19.455 59.925 19.705 60.725 ;
        RECT 19.895 60.575 21.120 60.745 ;
        RECT 19.895 60.095 20.225 60.575 ;
        RECT 20.395 59.925 20.620 60.385 ;
        RECT 20.790 60.095 21.120 60.575 ;
        RECT 21.750 60.705 21.920 61.335 ;
        RECT 22.105 60.915 22.455 61.165 ;
        RECT 21.750 60.095 22.250 60.705 ;
        RECT 22.685 60.605 23.040 61.165 ;
        RECT 23.210 60.435 23.380 61.335 ;
        RECT 23.550 60.605 23.815 61.165 ;
        RECT 24.065 60.835 24.235 61.335 ;
        RECT 24.405 60.665 24.720 61.685 ;
        RECT 24.925 61.385 26.595 62.475 ;
        RECT 26.855 61.805 27.025 62.305 ;
        RECT 27.195 61.975 27.525 62.475 ;
        RECT 26.855 61.635 27.520 61.805 ;
        RECT 22.790 59.925 23.030 60.435 ;
        RECT 23.210 60.105 23.490 60.435 ;
        RECT 23.720 59.925 23.935 60.435 ;
        RECT 24.105 60.095 24.720 60.665 ;
        RECT 24.925 60.695 25.675 61.215 ;
        RECT 25.845 60.865 26.595 61.385 ;
        RECT 26.770 60.815 27.120 61.465 ;
        RECT 24.925 59.925 26.595 60.695 ;
        RECT 27.290 60.645 27.520 61.635 ;
        RECT 26.855 60.475 27.520 60.645 ;
        RECT 26.855 60.185 27.025 60.475 ;
        RECT 27.195 59.925 27.525 60.305 ;
        RECT 27.695 60.185 27.880 62.305 ;
        RECT 28.120 62.015 28.385 62.475 ;
        RECT 28.555 61.880 28.805 62.305 ;
        RECT 29.015 62.030 30.120 62.200 ;
        RECT 28.500 61.750 28.805 61.880 ;
        RECT 28.050 60.555 28.330 61.505 ;
        RECT 28.500 60.645 28.670 61.750 ;
        RECT 28.840 60.965 29.080 61.560 ;
        RECT 29.250 61.495 29.780 61.860 ;
        RECT 29.250 60.795 29.420 61.495 ;
        RECT 29.950 61.415 30.120 62.030 ;
        RECT 30.290 61.675 30.460 62.475 ;
        RECT 30.630 61.975 30.880 62.305 ;
        RECT 31.105 62.005 31.990 62.175 ;
        RECT 29.950 61.325 30.460 61.415 ;
        RECT 28.500 60.515 28.725 60.645 ;
        RECT 28.895 60.575 29.420 60.795 ;
        RECT 29.590 61.155 30.460 61.325 ;
        RECT 28.135 59.925 28.385 60.385 ;
        RECT 28.555 60.375 28.725 60.515 ;
        RECT 29.590 60.375 29.760 61.155 ;
        RECT 30.290 61.085 30.460 61.155 ;
        RECT 29.970 60.905 30.170 60.935 ;
        RECT 30.630 60.905 30.800 61.975 ;
        RECT 30.970 61.085 31.160 61.805 ;
        RECT 29.970 60.605 30.800 60.905 ;
        RECT 31.330 60.875 31.650 61.835 ;
        RECT 28.555 60.205 28.890 60.375 ;
        RECT 29.085 60.205 29.760 60.375 ;
        RECT 30.080 59.925 30.450 60.425 ;
        RECT 30.630 60.375 30.800 60.605 ;
        RECT 31.185 60.545 31.650 60.875 ;
        RECT 31.820 61.165 31.990 62.005 ;
        RECT 32.170 61.975 32.485 62.475 ;
        RECT 32.715 61.745 33.055 62.305 ;
        RECT 32.160 61.370 33.055 61.745 ;
        RECT 33.225 61.465 33.395 62.475 ;
        RECT 32.865 61.165 33.055 61.370 ;
        RECT 33.565 61.415 33.895 62.260 ;
        RECT 33.565 61.335 33.955 61.415 ;
        RECT 34.125 61.385 36.715 62.475 ;
        RECT 33.740 61.285 33.955 61.335 ;
        RECT 31.820 60.835 32.695 61.165 ;
        RECT 32.865 60.835 33.615 61.165 ;
        RECT 31.820 60.375 31.990 60.835 ;
        RECT 32.865 60.665 33.065 60.835 ;
        RECT 33.785 60.705 33.955 61.285 ;
        RECT 33.730 60.665 33.955 60.705 ;
        RECT 30.630 60.205 31.035 60.375 ;
        RECT 31.205 60.205 31.990 60.375 ;
        RECT 32.265 59.925 32.475 60.455 ;
        RECT 32.735 60.140 33.065 60.665 ;
        RECT 33.575 60.580 33.955 60.665 ;
        RECT 34.125 60.695 35.335 61.215 ;
        RECT 35.505 60.865 36.715 61.385 ;
        RECT 36.890 61.335 37.225 62.305 ;
        RECT 37.395 61.335 37.565 62.475 ;
        RECT 37.735 62.135 39.765 62.305 ;
        RECT 33.235 59.925 33.405 60.535 ;
        RECT 33.575 60.145 33.905 60.580 ;
        RECT 34.125 59.925 36.715 60.695 ;
        RECT 36.890 60.665 37.060 61.335 ;
        RECT 37.735 61.165 37.905 62.135 ;
        RECT 37.230 60.835 37.485 61.165 ;
        RECT 37.710 60.835 37.905 61.165 ;
        RECT 38.075 61.795 39.200 61.965 ;
        RECT 37.315 60.665 37.485 60.835 ;
        RECT 38.075 60.665 38.245 61.795 ;
        RECT 36.890 60.095 37.145 60.665 ;
        RECT 37.315 60.495 38.245 60.665 ;
        RECT 38.415 61.455 39.425 61.625 ;
        RECT 38.415 60.655 38.585 61.455 ;
        RECT 38.790 61.115 39.065 61.255 ;
        RECT 38.785 60.945 39.065 61.115 ;
        RECT 38.070 60.460 38.245 60.495 ;
        RECT 37.315 59.925 37.645 60.325 ;
        RECT 38.070 60.095 38.600 60.460 ;
        RECT 38.790 60.095 39.065 60.945 ;
        RECT 39.235 60.095 39.425 61.455 ;
        RECT 39.595 61.470 39.765 62.135 ;
        RECT 39.935 61.715 40.105 62.475 ;
        RECT 40.340 61.715 40.855 62.125 ;
        RECT 39.595 61.280 40.345 61.470 ;
        RECT 40.515 60.905 40.855 61.715 ;
        RECT 41.540 61.605 41.825 62.475 ;
        RECT 41.995 61.845 42.255 62.305 ;
        RECT 42.430 62.015 42.685 62.475 ;
        RECT 42.855 61.845 43.115 62.305 ;
        RECT 41.995 61.675 43.115 61.845 ;
        RECT 43.285 61.675 43.595 62.475 ;
        RECT 41.995 61.425 42.255 61.675 ;
        RECT 43.765 61.505 44.075 62.305 ;
        RECT 39.625 60.735 40.855 60.905 ;
        RECT 41.500 61.255 42.255 61.425 ;
        RECT 43.045 61.335 44.075 61.505 ;
        RECT 41.500 60.745 41.905 61.255 ;
        RECT 43.045 61.085 43.215 61.335 ;
        RECT 42.075 60.915 43.215 61.085 ;
        RECT 39.605 59.925 40.115 60.460 ;
        RECT 40.335 60.130 40.580 60.735 ;
        RECT 41.500 60.575 43.150 60.745 ;
        RECT 43.385 60.595 43.735 61.165 ;
        RECT 41.545 59.925 41.825 60.405 ;
        RECT 41.995 60.185 42.255 60.575 ;
        RECT 42.430 59.925 42.685 60.405 ;
        RECT 42.855 60.185 43.150 60.575 ;
        RECT 43.905 60.425 44.075 61.335 ;
        RECT 44.245 61.310 44.535 62.475 ;
        RECT 44.795 61.805 44.965 62.305 ;
        RECT 45.135 61.975 45.465 62.475 ;
        RECT 44.795 61.635 45.460 61.805 ;
        RECT 44.710 60.815 45.060 61.465 ;
        RECT 43.330 59.925 43.605 60.405 ;
        RECT 43.775 60.095 44.075 60.425 ;
        RECT 44.245 59.925 44.535 60.650 ;
        RECT 45.230 60.645 45.460 61.635 ;
        RECT 44.795 60.475 45.460 60.645 ;
        RECT 44.795 60.185 44.965 60.475 ;
        RECT 45.135 59.925 45.465 60.305 ;
        RECT 45.635 60.185 45.820 62.305 ;
        RECT 46.060 62.015 46.325 62.475 ;
        RECT 46.495 61.880 46.745 62.305 ;
        RECT 46.955 62.030 48.060 62.200 ;
        RECT 46.440 61.750 46.745 61.880 ;
        RECT 45.990 60.555 46.270 61.505 ;
        RECT 46.440 60.645 46.610 61.750 ;
        RECT 46.780 60.965 47.020 61.560 ;
        RECT 47.190 61.495 47.720 61.860 ;
        RECT 47.190 60.795 47.360 61.495 ;
        RECT 47.890 61.415 48.060 62.030 ;
        RECT 48.230 61.675 48.400 62.475 ;
        RECT 48.570 61.975 48.820 62.305 ;
        RECT 49.045 62.005 49.930 62.175 ;
        RECT 47.890 61.325 48.400 61.415 ;
        RECT 46.440 60.515 46.665 60.645 ;
        RECT 46.835 60.575 47.360 60.795 ;
        RECT 47.530 61.155 48.400 61.325 ;
        RECT 46.075 59.925 46.325 60.385 ;
        RECT 46.495 60.375 46.665 60.515 ;
        RECT 47.530 60.375 47.700 61.155 ;
        RECT 48.230 61.085 48.400 61.155 ;
        RECT 47.910 60.905 48.110 60.935 ;
        RECT 48.570 60.905 48.740 61.975 ;
        RECT 48.910 61.085 49.100 61.805 ;
        RECT 47.910 60.605 48.740 60.905 ;
        RECT 49.270 60.875 49.590 61.835 ;
        RECT 46.495 60.205 46.830 60.375 ;
        RECT 47.025 60.205 47.700 60.375 ;
        RECT 48.020 59.925 48.390 60.425 ;
        RECT 48.570 60.375 48.740 60.605 ;
        RECT 49.125 60.545 49.590 60.875 ;
        RECT 49.760 61.165 49.930 62.005 ;
        RECT 50.110 61.975 50.425 62.475 ;
        RECT 50.655 61.745 50.995 62.305 ;
        RECT 50.100 61.370 50.995 61.745 ;
        RECT 51.165 61.465 51.335 62.475 ;
        RECT 50.805 61.165 50.995 61.370 ;
        RECT 51.505 61.415 51.835 62.260 ;
        RECT 51.505 61.335 51.895 61.415 ;
        RECT 51.680 61.285 51.895 61.335 ;
        RECT 49.760 60.835 50.635 61.165 ;
        RECT 50.805 60.835 51.555 61.165 ;
        RECT 49.760 60.375 49.930 60.835 ;
        RECT 50.805 60.665 51.005 60.835 ;
        RECT 51.725 60.705 51.895 61.285 ;
        RECT 51.670 60.665 51.895 60.705 ;
        RECT 48.570 60.205 48.975 60.375 ;
        RECT 49.145 60.205 49.930 60.375 ;
        RECT 50.205 59.925 50.415 60.455 ;
        RECT 50.675 60.140 51.005 60.665 ;
        RECT 51.515 60.580 51.895 60.665 ;
        RECT 52.065 61.335 52.450 62.305 ;
        RECT 52.620 62.015 52.945 62.475 ;
        RECT 53.465 61.845 53.745 62.305 ;
        RECT 52.620 61.625 53.745 61.845 ;
        RECT 52.065 60.665 52.345 61.335 ;
        RECT 52.620 61.165 53.070 61.625 ;
        RECT 53.935 61.455 54.335 62.305 ;
        RECT 54.735 62.015 55.005 62.475 ;
        RECT 55.175 61.845 55.460 62.305 ;
        RECT 52.515 60.835 53.070 61.165 ;
        RECT 53.240 60.895 54.335 61.455 ;
        RECT 52.620 60.725 53.070 60.835 ;
        RECT 51.175 59.925 51.345 60.535 ;
        RECT 51.515 60.145 51.845 60.580 ;
        RECT 52.065 60.095 52.450 60.665 ;
        RECT 52.620 60.555 53.745 60.725 ;
        RECT 52.620 59.925 52.945 60.385 ;
        RECT 53.465 60.095 53.745 60.555 ;
        RECT 53.935 60.095 54.335 60.895 ;
        RECT 54.505 61.625 55.460 61.845 ;
        RECT 55.860 61.845 56.145 62.305 ;
        RECT 56.315 62.015 56.585 62.475 ;
        RECT 55.860 61.625 56.815 61.845 ;
        RECT 54.505 60.725 54.715 61.625 ;
        RECT 54.885 60.895 55.575 61.455 ;
        RECT 55.745 60.895 56.435 61.455 ;
        RECT 56.605 60.725 56.815 61.625 ;
        RECT 54.505 60.555 55.460 60.725 ;
        RECT 54.735 59.925 55.005 60.385 ;
        RECT 55.175 60.095 55.460 60.555 ;
        RECT 55.860 60.555 56.815 60.725 ;
        RECT 56.985 61.455 57.385 62.305 ;
        RECT 57.575 61.845 57.855 62.305 ;
        RECT 58.375 62.015 58.700 62.475 ;
        RECT 57.575 61.625 58.700 61.845 ;
        RECT 56.985 60.895 58.080 61.455 ;
        RECT 58.250 61.165 58.700 61.625 ;
        RECT 58.870 61.335 59.255 62.305 ;
        RECT 59.430 61.675 59.685 62.475 ;
        RECT 59.885 61.625 60.215 62.305 ;
        RECT 55.860 60.095 56.145 60.555 ;
        RECT 56.315 59.925 56.585 60.385 ;
        RECT 56.985 60.095 57.385 60.895 ;
        RECT 58.250 60.835 58.805 61.165 ;
        RECT 58.250 60.725 58.700 60.835 ;
        RECT 57.575 60.555 58.700 60.725 ;
        RECT 58.975 60.665 59.255 61.335 ;
        RECT 59.430 61.135 59.675 61.495 ;
        RECT 59.865 61.345 60.215 61.625 ;
        RECT 59.865 60.965 60.035 61.345 ;
        RECT 60.395 61.165 60.590 62.215 ;
        RECT 60.770 61.335 61.090 62.475 ;
        RECT 62.195 61.365 62.490 62.475 ;
        RECT 62.670 61.165 62.920 62.300 ;
        RECT 63.090 61.365 63.350 62.475 ;
        RECT 63.520 61.575 63.780 62.300 ;
        RECT 63.950 61.745 64.210 62.475 ;
        RECT 64.380 61.575 64.640 62.300 ;
        RECT 64.810 61.745 65.070 62.475 ;
        RECT 65.240 61.575 65.500 62.300 ;
        RECT 65.670 61.745 65.930 62.475 ;
        RECT 66.100 61.575 66.360 62.300 ;
        RECT 66.530 61.745 66.825 62.475 ;
        RECT 63.520 61.335 66.830 61.575 ;
        RECT 67.890 61.505 68.280 61.680 ;
        RECT 68.765 61.675 69.095 62.475 ;
        RECT 69.265 61.685 69.800 62.305 ;
        RECT 67.890 61.335 69.315 61.505 ;
        RECT 57.575 60.095 57.855 60.555 ;
        RECT 58.375 59.925 58.700 60.385 ;
        RECT 58.870 60.095 59.255 60.665 ;
        RECT 59.515 60.795 60.035 60.965 ;
        RECT 60.205 60.835 60.590 61.165 ;
        RECT 60.770 61.115 61.030 61.165 ;
        RECT 60.770 60.945 61.035 61.115 ;
        RECT 60.770 60.835 61.030 60.945 ;
        RECT 59.515 60.435 59.685 60.795 ;
        RECT 59.485 60.265 59.685 60.435 ;
        RECT 59.515 60.230 59.685 60.265 ;
        RECT 59.875 60.455 61.090 60.625 ;
        RECT 62.185 60.555 62.500 61.165 ;
        RECT 62.670 60.915 65.690 61.165 ;
        RECT 59.875 60.150 60.105 60.455 ;
        RECT 60.275 59.925 60.605 60.285 ;
        RECT 60.800 60.105 61.090 60.455 ;
        RECT 62.245 59.925 62.490 60.385 ;
        RECT 62.670 60.105 62.920 60.915 ;
        RECT 65.860 60.745 66.830 61.335 ;
        RECT 63.520 60.575 66.830 60.745 ;
        RECT 67.765 60.605 68.120 61.165 ;
        RECT 63.090 59.925 63.350 60.450 ;
        RECT 63.520 60.120 63.780 60.575 ;
        RECT 63.950 59.925 64.210 60.405 ;
        RECT 64.380 60.120 64.640 60.575 ;
        RECT 64.810 59.925 65.070 60.405 ;
        RECT 65.240 60.120 65.500 60.575 ;
        RECT 65.670 59.925 65.930 60.405 ;
        RECT 66.100 60.120 66.360 60.575 ;
        RECT 68.290 60.435 68.460 61.335 ;
        RECT 68.630 60.605 68.895 61.165 ;
        RECT 69.145 60.835 69.315 61.335 ;
        RECT 69.485 60.665 69.800 61.685 ;
        RECT 70.005 61.310 70.295 62.475 ;
        RECT 70.465 61.385 72.135 62.475 ;
        RECT 72.420 61.845 72.705 62.305 ;
        RECT 72.875 62.015 73.145 62.475 ;
        RECT 72.420 61.625 73.375 61.845 ;
        RECT 66.530 59.925 66.830 60.405 ;
        RECT 67.870 59.925 68.110 60.435 ;
        RECT 68.290 60.105 68.570 60.435 ;
        RECT 68.800 59.925 69.015 60.435 ;
        RECT 69.185 60.095 69.800 60.665 ;
        RECT 70.465 60.695 71.215 61.215 ;
        RECT 71.385 60.865 72.135 61.385 ;
        RECT 72.305 60.895 72.995 61.455 ;
        RECT 73.165 60.725 73.375 61.625 ;
        RECT 70.005 59.925 70.295 60.650 ;
        RECT 70.465 59.925 72.135 60.695 ;
        RECT 72.420 60.555 73.375 60.725 ;
        RECT 73.545 61.455 73.945 62.305 ;
        RECT 74.135 61.845 74.415 62.305 ;
        RECT 74.935 62.015 75.260 62.475 ;
        RECT 74.135 61.625 75.260 61.845 ;
        RECT 73.545 60.895 74.640 61.455 ;
        RECT 74.810 61.165 75.260 61.625 ;
        RECT 75.430 61.335 75.815 62.305 ;
        RECT 72.420 60.095 72.705 60.555 ;
        RECT 72.875 59.925 73.145 60.385 ;
        RECT 73.545 60.095 73.945 60.895 ;
        RECT 74.810 60.835 75.365 61.165 ;
        RECT 74.810 60.725 75.260 60.835 ;
        RECT 74.135 60.555 75.260 60.725 ;
        RECT 75.535 60.665 75.815 61.335 ;
        RECT 74.135 60.095 74.415 60.555 ;
        RECT 74.935 59.925 75.260 60.385 ;
        RECT 75.430 60.095 75.815 60.665 ;
        RECT 75.990 61.335 76.325 62.305 ;
        RECT 76.495 61.335 76.665 62.475 ;
        RECT 76.835 62.135 78.865 62.305 ;
        RECT 75.990 60.665 76.160 61.335 ;
        RECT 76.835 61.165 77.005 62.135 ;
        RECT 76.330 60.835 76.585 61.165 ;
        RECT 76.810 60.835 77.005 61.165 ;
        RECT 77.175 61.795 78.300 61.965 ;
        RECT 76.415 60.665 76.585 60.835 ;
        RECT 77.175 60.665 77.345 61.795 ;
        RECT 75.990 60.095 76.245 60.665 ;
        RECT 76.415 60.495 77.345 60.665 ;
        RECT 77.515 61.455 78.525 61.625 ;
        RECT 77.515 60.655 77.685 61.455 ;
        RECT 77.890 60.775 78.165 61.255 ;
        RECT 77.885 60.605 78.165 60.775 ;
        RECT 77.170 60.460 77.345 60.495 ;
        RECT 76.415 59.925 76.745 60.325 ;
        RECT 77.170 60.095 77.700 60.460 ;
        RECT 77.890 60.095 78.165 60.605 ;
        RECT 78.335 60.095 78.525 61.455 ;
        RECT 78.695 61.470 78.865 62.135 ;
        RECT 79.035 61.715 79.205 62.475 ;
        RECT 79.440 61.715 79.955 62.125 ;
        RECT 78.695 61.280 79.445 61.470 ;
        RECT 79.615 60.905 79.955 61.715 ;
        RECT 81.135 61.545 81.305 62.305 ;
        RECT 81.520 61.715 81.850 62.475 ;
        RECT 81.135 61.375 81.850 61.545 ;
        RECT 82.020 61.400 82.275 62.305 ;
        RECT 78.725 60.735 79.955 60.905 ;
        RECT 81.045 60.825 81.400 61.195 ;
        RECT 81.680 61.165 81.850 61.375 ;
        RECT 81.680 60.835 81.935 61.165 ;
        RECT 78.705 59.925 79.215 60.460 ;
        RECT 79.435 60.130 79.680 60.735 ;
        RECT 81.680 60.645 81.850 60.835 ;
        RECT 82.105 60.670 82.275 61.400 ;
        RECT 82.450 61.325 82.710 62.475 ;
        RECT 82.885 61.385 84.095 62.475 ;
        RECT 82.885 60.845 83.405 61.385 ;
        RECT 81.135 60.475 81.850 60.645 ;
        RECT 81.135 60.095 81.305 60.475 ;
        RECT 81.520 59.925 81.850 60.305 ;
        RECT 82.020 60.095 82.275 60.670 ;
        RECT 82.450 59.925 82.710 60.765 ;
        RECT 83.575 60.675 84.095 61.215 ;
        RECT 82.885 59.925 84.095 60.675 ;
        RECT 5.520 59.755 84.180 59.925 ;
        RECT 5.605 59.005 6.815 59.755 ;
        RECT 6.985 59.005 8.195 59.755 ;
        RECT 8.530 59.245 8.770 59.755 ;
        RECT 8.950 59.245 9.230 59.575 ;
        RECT 9.460 59.245 9.675 59.755 ;
        RECT 5.605 58.465 6.125 59.005 ;
        RECT 6.295 58.295 6.815 58.835 ;
        RECT 6.985 58.465 7.505 59.005 ;
        RECT 7.675 58.295 8.195 58.835 ;
        RECT 8.425 58.515 8.780 59.075 ;
        RECT 8.950 58.345 9.120 59.245 ;
        RECT 9.290 58.515 9.555 59.075 ;
        RECT 9.845 59.015 10.460 59.585 ;
        RECT 9.805 58.345 9.975 58.845 ;
        RECT 5.605 57.205 6.815 58.295 ;
        RECT 6.985 57.205 8.195 58.295 ;
        RECT 8.550 58.175 9.975 58.345 ;
        RECT 8.550 58.000 8.940 58.175 ;
        RECT 9.425 57.205 9.755 58.005 ;
        RECT 10.145 57.995 10.460 59.015 ;
        RECT 10.665 59.005 11.875 59.755 ;
        RECT 12.045 59.015 12.305 59.585 ;
        RECT 12.475 59.355 12.860 59.755 ;
        RECT 13.030 59.185 13.285 59.585 ;
        RECT 12.475 59.015 13.285 59.185 ;
        RECT 13.475 59.015 13.720 59.585 ;
        RECT 13.890 59.355 14.275 59.755 ;
        RECT 14.445 59.185 14.700 59.585 ;
        RECT 13.890 59.015 14.700 59.185 ;
        RECT 14.890 59.015 15.315 59.585 ;
        RECT 15.485 59.355 15.870 59.755 ;
        RECT 16.040 59.185 16.475 59.585 ;
        RECT 15.485 59.015 16.475 59.185 ;
        RECT 16.735 59.205 16.905 59.495 ;
        RECT 17.075 59.375 17.405 59.755 ;
        RECT 16.735 59.035 17.400 59.205 ;
        RECT 10.665 58.465 11.185 59.005 ;
        RECT 11.355 58.295 11.875 58.835 ;
        RECT 9.925 57.375 10.460 57.995 ;
        RECT 10.665 57.205 11.875 58.295 ;
        RECT 12.045 58.345 12.230 59.015 ;
        RECT 12.475 58.845 12.825 59.015 ;
        RECT 13.475 58.845 13.645 59.015 ;
        RECT 13.890 58.845 14.240 59.015 ;
        RECT 14.890 58.845 15.240 59.015 ;
        RECT 15.485 58.845 15.820 59.015 ;
        RECT 12.400 58.515 12.825 58.845 ;
        RECT 12.045 57.375 12.305 58.345 ;
        RECT 12.475 57.995 12.825 58.515 ;
        RECT 12.995 58.345 13.645 58.845 ;
        RECT 13.815 58.515 14.240 58.845 ;
        RECT 12.995 58.165 13.720 58.345 ;
        RECT 12.475 57.800 13.285 57.995 ;
        RECT 12.475 57.205 12.860 57.630 ;
        RECT 13.030 57.375 13.285 57.800 ;
        RECT 13.475 57.375 13.720 58.165 ;
        RECT 13.890 57.995 14.240 58.515 ;
        RECT 14.410 58.345 15.240 58.845 ;
        RECT 15.410 58.515 15.820 58.845 ;
        RECT 14.410 58.165 15.315 58.345 ;
        RECT 13.890 57.800 14.720 57.995 ;
        RECT 13.890 57.205 14.275 57.630 ;
        RECT 14.445 57.375 14.720 57.800 ;
        RECT 14.890 57.375 15.315 58.165 ;
        RECT 15.485 57.970 15.820 58.515 ;
        RECT 15.990 58.140 16.475 58.845 ;
        RECT 16.650 58.215 17.000 58.865 ;
        RECT 17.170 58.045 17.400 59.035 ;
        RECT 15.485 57.800 16.475 57.970 ;
        RECT 15.485 57.205 15.870 57.630 ;
        RECT 16.040 57.375 16.475 57.800 ;
        RECT 16.735 57.875 17.400 58.045 ;
        RECT 16.735 57.375 16.905 57.875 ;
        RECT 17.075 57.205 17.405 57.705 ;
        RECT 17.575 57.375 17.760 59.495 ;
        RECT 18.015 59.295 18.265 59.755 ;
        RECT 18.435 59.305 18.770 59.475 ;
        RECT 18.965 59.305 19.640 59.475 ;
        RECT 18.435 59.165 18.605 59.305 ;
        RECT 17.930 58.175 18.210 59.125 ;
        RECT 18.380 59.035 18.605 59.165 ;
        RECT 18.380 57.930 18.550 59.035 ;
        RECT 18.775 58.885 19.300 59.105 ;
        RECT 18.720 58.120 18.960 58.715 ;
        RECT 19.130 58.185 19.300 58.885 ;
        RECT 19.470 58.525 19.640 59.305 ;
        RECT 19.960 59.255 20.330 59.755 ;
        RECT 20.510 59.305 20.915 59.475 ;
        RECT 21.085 59.305 21.870 59.475 ;
        RECT 20.510 59.075 20.680 59.305 ;
        RECT 19.850 58.775 20.680 59.075 ;
        RECT 21.065 58.805 21.530 59.135 ;
        RECT 19.850 58.745 20.050 58.775 ;
        RECT 20.170 58.525 20.340 58.595 ;
        RECT 19.470 58.355 20.340 58.525 ;
        RECT 19.830 58.265 20.340 58.355 ;
        RECT 18.380 57.800 18.685 57.930 ;
        RECT 19.130 57.820 19.660 58.185 ;
        RECT 18.000 57.205 18.265 57.665 ;
        RECT 18.435 57.375 18.685 57.800 ;
        RECT 19.830 57.650 20.000 58.265 ;
        RECT 18.895 57.480 20.000 57.650 ;
        RECT 20.170 57.205 20.340 58.005 ;
        RECT 20.510 57.705 20.680 58.775 ;
        RECT 20.850 57.875 21.040 58.595 ;
        RECT 21.210 57.845 21.530 58.805 ;
        RECT 21.700 58.845 21.870 59.305 ;
        RECT 22.145 59.225 22.355 59.755 ;
        RECT 22.615 59.015 22.945 59.540 ;
        RECT 23.115 59.145 23.285 59.755 ;
        RECT 23.455 59.100 23.785 59.535 ;
        RECT 24.095 59.205 24.265 59.495 ;
        RECT 24.435 59.375 24.765 59.755 ;
        RECT 23.455 59.015 23.835 59.100 ;
        RECT 24.095 59.035 24.760 59.205 ;
        RECT 22.745 58.845 22.945 59.015 ;
        RECT 23.610 58.975 23.835 59.015 ;
        RECT 21.700 58.515 22.575 58.845 ;
        RECT 22.745 58.515 23.495 58.845 ;
        RECT 20.510 57.375 20.760 57.705 ;
        RECT 21.700 57.675 21.870 58.515 ;
        RECT 22.745 58.310 22.935 58.515 ;
        RECT 23.665 58.395 23.835 58.975 ;
        RECT 23.620 58.345 23.835 58.395 ;
        RECT 22.040 57.935 22.935 58.310 ;
        RECT 23.445 58.265 23.835 58.345 ;
        RECT 20.985 57.505 21.870 57.675 ;
        RECT 22.050 57.205 22.365 57.705 ;
        RECT 22.595 57.375 22.935 57.935 ;
        RECT 23.105 57.205 23.275 58.215 ;
        RECT 23.445 57.420 23.775 58.265 ;
        RECT 24.010 58.215 24.360 58.865 ;
        RECT 24.530 58.045 24.760 59.035 ;
        RECT 24.095 57.875 24.760 58.045 ;
        RECT 24.095 57.375 24.265 57.875 ;
        RECT 24.435 57.205 24.765 57.705 ;
        RECT 24.935 57.375 25.120 59.495 ;
        RECT 25.375 59.295 25.625 59.755 ;
        RECT 25.795 59.305 26.130 59.475 ;
        RECT 26.325 59.305 27.000 59.475 ;
        RECT 25.795 59.165 25.965 59.305 ;
        RECT 25.290 58.175 25.570 59.125 ;
        RECT 25.740 59.035 25.965 59.165 ;
        RECT 25.740 57.930 25.910 59.035 ;
        RECT 26.135 58.885 26.660 59.105 ;
        RECT 26.080 58.120 26.320 58.715 ;
        RECT 26.490 58.185 26.660 58.885 ;
        RECT 26.830 58.525 27.000 59.305 ;
        RECT 27.320 59.255 27.690 59.755 ;
        RECT 27.870 59.305 28.275 59.475 ;
        RECT 28.445 59.305 29.230 59.475 ;
        RECT 27.870 59.075 28.040 59.305 ;
        RECT 27.210 58.775 28.040 59.075 ;
        RECT 28.425 58.805 28.890 59.135 ;
        RECT 27.210 58.745 27.410 58.775 ;
        RECT 27.530 58.525 27.700 58.595 ;
        RECT 26.830 58.355 27.700 58.525 ;
        RECT 27.190 58.265 27.700 58.355 ;
        RECT 25.740 57.800 26.045 57.930 ;
        RECT 26.490 57.820 27.020 58.185 ;
        RECT 25.360 57.205 25.625 57.665 ;
        RECT 25.795 57.375 26.045 57.800 ;
        RECT 27.190 57.650 27.360 58.265 ;
        RECT 26.255 57.480 27.360 57.650 ;
        RECT 27.530 57.205 27.700 58.005 ;
        RECT 27.870 57.705 28.040 58.775 ;
        RECT 28.210 57.875 28.400 58.595 ;
        RECT 28.570 57.845 28.890 58.805 ;
        RECT 29.060 58.845 29.230 59.305 ;
        RECT 29.505 59.225 29.715 59.755 ;
        RECT 29.975 59.015 30.305 59.540 ;
        RECT 30.475 59.145 30.645 59.755 ;
        RECT 30.815 59.100 31.145 59.535 ;
        RECT 30.815 59.015 31.195 59.100 ;
        RECT 31.365 59.030 31.655 59.755 ;
        RECT 30.105 58.845 30.305 59.015 ;
        RECT 30.970 58.975 31.195 59.015 ;
        RECT 29.060 58.515 29.935 58.845 ;
        RECT 30.105 58.515 30.855 58.845 ;
        RECT 27.870 57.375 28.120 57.705 ;
        RECT 29.060 57.675 29.230 58.515 ;
        RECT 30.105 58.310 30.295 58.515 ;
        RECT 31.025 58.395 31.195 58.975 ;
        RECT 31.825 58.985 34.415 59.755 ;
        RECT 34.675 59.205 34.845 59.495 ;
        RECT 35.015 59.375 35.345 59.755 ;
        RECT 34.675 59.035 35.340 59.205 ;
        RECT 31.825 58.465 33.035 58.985 ;
        RECT 30.980 58.345 31.195 58.395 ;
        RECT 29.400 57.935 30.295 58.310 ;
        RECT 30.805 58.265 31.195 58.345 ;
        RECT 28.345 57.505 29.230 57.675 ;
        RECT 29.410 57.205 29.725 57.705 ;
        RECT 29.955 57.375 30.295 57.935 ;
        RECT 30.465 57.205 30.635 58.215 ;
        RECT 30.805 57.420 31.135 58.265 ;
        RECT 31.365 57.205 31.655 58.370 ;
        RECT 33.205 58.295 34.415 58.815 ;
        RECT 31.825 57.205 34.415 58.295 ;
        RECT 34.590 58.215 34.940 58.865 ;
        RECT 35.110 58.045 35.340 59.035 ;
        RECT 34.675 57.875 35.340 58.045 ;
        RECT 34.675 57.375 34.845 57.875 ;
        RECT 35.015 57.205 35.345 57.705 ;
        RECT 35.515 57.375 35.700 59.495 ;
        RECT 35.955 59.295 36.205 59.755 ;
        RECT 36.375 59.305 36.710 59.475 ;
        RECT 36.905 59.305 37.580 59.475 ;
        RECT 36.375 59.165 36.545 59.305 ;
        RECT 35.870 58.175 36.150 59.125 ;
        RECT 36.320 59.035 36.545 59.165 ;
        RECT 36.320 57.930 36.490 59.035 ;
        RECT 36.715 58.885 37.240 59.105 ;
        RECT 36.660 58.120 36.900 58.715 ;
        RECT 37.070 58.185 37.240 58.885 ;
        RECT 37.410 58.525 37.580 59.305 ;
        RECT 37.900 59.255 38.270 59.755 ;
        RECT 38.450 59.305 38.855 59.475 ;
        RECT 39.025 59.305 39.810 59.475 ;
        RECT 38.450 59.075 38.620 59.305 ;
        RECT 37.790 58.775 38.620 59.075 ;
        RECT 39.005 58.805 39.470 59.135 ;
        RECT 37.790 58.745 37.990 58.775 ;
        RECT 38.110 58.525 38.280 58.595 ;
        RECT 37.410 58.355 38.280 58.525 ;
        RECT 37.770 58.265 38.280 58.355 ;
        RECT 36.320 57.800 36.625 57.930 ;
        RECT 37.070 57.820 37.600 58.185 ;
        RECT 35.940 57.205 36.205 57.665 ;
        RECT 36.375 57.375 36.625 57.800 ;
        RECT 37.770 57.650 37.940 58.265 ;
        RECT 36.835 57.480 37.940 57.650 ;
        RECT 38.110 57.205 38.280 58.005 ;
        RECT 38.450 57.705 38.620 58.775 ;
        RECT 38.790 57.875 38.980 58.595 ;
        RECT 39.150 57.845 39.470 58.805 ;
        RECT 39.640 58.845 39.810 59.305 ;
        RECT 40.085 59.225 40.295 59.755 ;
        RECT 40.555 59.015 40.885 59.540 ;
        RECT 41.055 59.145 41.225 59.755 ;
        RECT 41.395 59.100 41.725 59.535 ;
        RECT 41.395 59.015 41.775 59.100 ;
        RECT 40.685 58.845 40.885 59.015 ;
        RECT 41.550 58.975 41.775 59.015 ;
        RECT 39.640 58.515 40.515 58.845 ;
        RECT 40.685 58.515 41.435 58.845 ;
        RECT 38.450 57.375 38.700 57.705 ;
        RECT 39.640 57.675 39.810 58.515 ;
        RECT 40.685 58.310 40.875 58.515 ;
        RECT 41.605 58.395 41.775 58.975 ;
        RECT 41.945 58.985 43.615 59.755 ;
        RECT 41.945 58.465 42.695 58.985 ;
        RECT 44.060 58.945 44.305 59.550 ;
        RECT 44.525 59.220 45.035 59.755 ;
        RECT 41.560 58.345 41.775 58.395 ;
        RECT 39.980 57.935 40.875 58.310 ;
        RECT 41.385 58.265 41.775 58.345 ;
        RECT 42.865 58.295 43.615 58.815 ;
        RECT 38.925 57.505 39.810 57.675 ;
        RECT 39.990 57.205 40.305 57.705 ;
        RECT 40.535 57.375 40.875 57.935 ;
        RECT 41.045 57.205 41.215 58.215 ;
        RECT 41.385 57.420 41.715 58.265 ;
        RECT 41.945 57.205 43.615 58.295 ;
        RECT 43.785 58.775 45.015 58.945 ;
        RECT 43.785 57.965 44.125 58.775 ;
        RECT 44.295 58.210 45.045 58.400 ;
        RECT 43.785 57.555 44.300 57.965 ;
        RECT 44.535 57.205 44.705 57.965 ;
        RECT 44.875 57.545 45.045 58.210 ;
        RECT 45.215 58.225 45.405 59.585 ;
        RECT 45.575 59.075 45.850 59.585 ;
        RECT 46.040 59.220 46.570 59.585 ;
        RECT 46.995 59.355 47.325 59.755 ;
        RECT 46.395 59.185 46.570 59.220 ;
        RECT 45.575 58.905 45.855 59.075 ;
        RECT 45.575 58.425 45.850 58.905 ;
        RECT 46.055 58.225 46.225 59.025 ;
        RECT 45.215 58.055 46.225 58.225 ;
        RECT 46.395 59.015 47.325 59.185 ;
        RECT 47.495 59.015 47.750 59.585 ;
        RECT 46.395 57.885 46.565 59.015 ;
        RECT 47.155 58.845 47.325 59.015 ;
        RECT 45.440 57.715 46.565 57.885 ;
        RECT 46.735 58.515 46.930 58.845 ;
        RECT 47.155 58.515 47.410 58.845 ;
        RECT 46.735 57.545 46.905 58.515 ;
        RECT 47.580 58.345 47.750 59.015 ;
        RECT 47.925 58.985 49.595 59.755 ;
        RECT 49.815 59.100 50.145 59.535 ;
        RECT 50.315 59.145 50.485 59.755 ;
        RECT 49.765 59.015 50.145 59.100 ;
        RECT 50.655 59.015 50.985 59.540 ;
        RECT 51.245 59.225 51.455 59.755 ;
        RECT 51.730 59.305 52.515 59.475 ;
        RECT 52.685 59.305 53.090 59.475 ;
        RECT 47.925 58.465 48.675 58.985 ;
        RECT 49.765 58.975 49.990 59.015 ;
        RECT 44.875 57.375 46.905 57.545 ;
        RECT 47.075 57.205 47.245 58.345 ;
        RECT 47.415 57.375 47.750 58.345 ;
        RECT 48.845 58.295 49.595 58.815 ;
        RECT 47.925 57.205 49.595 58.295 ;
        RECT 49.765 58.395 49.935 58.975 ;
        RECT 50.655 58.845 50.855 59.015 ;
        RECT 51.730 58.845 51.900 59.305 ;
        RECT 50.105 58.515 50.855 58.845 ;
        RECT 51.025 58.515 51.900 58.845 ;
        RECT 49.765 58.345 49.980 58.395 ;
        RECT 49.765 58.265 50.155 58.345 ;
        RECT 49.825 57.420 50.155 58.265 ;
        RECT 50.665 58.310 50.855 58.515 ;
        RECT 50.325 57.205 50.495 58.215 ;
        RECT 50.665 57.935 51.560 58.310 ;
        RECT 50.665 57.375 51.005 57.935 ;
        RECT 51.235 57.205 51.550 57.705 ;
        RECT 51.730 57.675 51.900 58.515 ;
        RECT 52.070 58.805 52.535 59.135 ;
        RECT 52.920 59.075 53.090 59.305 ;
        RECT 53.270 59.255 53.640 59.755 ;
        RECT 53.960 59.305 54.635 59.475 ;
        RECT 54.830 59.305 55.165 59.475 ;
        RECT 52.070 57.845 52.390 58.805 ;
        RECT 52.920 58.775 53.750 59.075 ;
        RECT 52.560 57.875 52.750 58.595 ;
        RECT 52.920 57.705 53.090 58.775 ;
        RECT 53.550 58.745 53.750 58.775 ;
        RECT 53.260 58.525 53.430 58.595 ;
        RECT 53.960 58.525 54.130 59.305 ;
        RECT 54.995 59.165 55.165 59.305 ;
        RECT 55.335 59.295 55.585 59.755 ;
        RECT 53.260 58.355 54.130 58.525 ;
        RECT 54.300 58.885 54.825 59.105 ;
        RECT 54.995 59.035 55.220 59.165 ;
        RECT 53.260 58.265 53.770 58.355 ;
        RECT 51.730 57.505 52.615 57.675 ;
        RECT 52.840 57.375 53.090 57.705 ;
        RECT 53.260 57.205 53.430 58.005 ;
        RECT 53.600 57.650 53.770 58.265 ;
        RECT 54.300 58.185 54.470 58.885 ;
        RECT 53.940 57.820 54.470 58.185 ;
        RECT 54.640 58.120 54.880 58.715 ;
        RECT 55.050 57.930 55.220 59.035 ;
        RECT 55.390 58.175 55.670 59.125 ;
        RECT 54.915 57.800 55.220 57.930 ;
        RECT 53.600 57.480 54.705 57.650 ;
        RECT 54.915 57.375 55.165 57.800 ;
        RECT 55.335 57.205 55.600 57.665 ;
        RECT 55.840 57.375 56.025 59.495 ;
        RECT 56.195 59.375 56.525 59.755 ;
        RECT 56.695 59.205 56.865 59.495 ;
        RECT 56.200 59.035 56.865 59.205 ;
        RECT 56.200 58.045 56.430 59.035 ;
        RECT 57.125 59.030 57.415 59.755 ;
        RECT 57.585 59.255 57.845 59.585 ;
        RECT 58.015 59.395 58.345 59.755 ;
        RECT 58.600 59.375 59.900 59.585 ;
        RECT 57.585 59.245 57.815 59.255 ;
        RECT 56.600 58.215 56.950 58.865 ;
        RECT 56.200 57.875 56.865 58.045 ;
        RECT 56.195 57.205 56.525 57.705 ;
        RECT 56.695 57.375 56.865 57.875 ;
        RECT 57.125 57.205 57.415 58.370 ;
        RECT 57.585 58.055 57.755 59.245 ;
        RECT 58.600 59.225 58.770 59.375 ;
        RECT 58.015 59.100 58.770 59.225 ;
        RECT 57.925 59.055 58.770 59.100 ;
        RECT 57.925 58.935 58.195 59.055 ;
        RECT 57.925 58.360 58.095 58.935 ;
        RECT 58.325 58.495 58.735 58.800 ;
        RECT 59.025 58.765 59.235 59.165 ;
        RECT 58.905 58.555 59.235 58.765 ;
        RECT 59.480 58.765 59.700 59.165 ;
        RECT 60.175 58.990 60.630 59.755 ;
        RECT 60.805 58.955 61.500 59.585 ;
        RECT 61.705 58.955 62.015 59.755 ;
        RECT 62.195 59.105 62.525 59.580 ;
        RECT 62.695 59.275 62.865 59.755 ;
        RECT 63.035 59.105 63.365 59.580 ;
        RECT 63.535 59.275 63.705 59.755 ;
        RECT 63.875 59.105 64.205 59.580 ;
        RECT 64.375 59.275 64.545 59.755 ;
        RECT 64.715 59.105 65.045 59.580 ;
        RECT 65.215 59.275 65.385 59.755 ;
        RECT 65.555 59.105 65.885 59.580 ;
        RECT 66.055 59.275 66.225 59.755 ;
        RECT 66.395 59.580 66.645 59.585 ;
        RECT 66.395 59.105 66.725 59.580 ;
        RECT 66.895 59.275 67.065 59.755 ;
        RECT 67.315 59.580 67.485 59.585 ;
        RECT 67.235 59.105 67.565 59.580 ;
        RECT 67.735 59.275 67.905 59.755 ;
        RECT 68.155 59.580 68.325 59.585 ;
        RECT 68.075 59.105 68.405 59.580 ;
        RECT 68.575 59.275 68.745 59.755 ;
        RECT 68.915 59.105 69.245 59.580 ;
        RECT 69.415 59.275 69.585 59.755 ;
        RECT 69.755 59.105 70.085 59.580 ;
        RECT 70.255 59.275 70.425 59.755 ;
        RECT 70.595 59.105 70.925 59.580 ;
        RECT 71.095 59.275 71.265 59.755 ;
        RECT 71.435 59.105 71.765 59.580 ;
        RECT 71.935 59.275 72.105 59.755 ;
        RECT 72.275 59.105 72.605 59.580 ;
        RECT 72.775 59.275 72.945 59.755 ;
        RECT 59.480 58.555 59.955 58.765 ;
        RECT 60.145 58.565 60.635 58.765 ;
        RECT 60.825 58.515 61.160 58.765 ;
        RECT 57.925 58.325 58.125 58.360 ;
        RECT 59.455 58.325 60.630 58.385 ;
        RECT 61.330 58.355 61.500 58.955 ;
        RECT 62.195 58.935 63.705 59.105 ;
        RECT 63.875 58.935 66.225 59.105 ;
        RECT 66.395 58.935 73.055 59.105 ;
        RECT 73.225 58.955 73.535 59.755 ;
        RECT 73.740 58.955 74.435 59.585 ;
        RECT 75.530 59.015 75.785 59.585 ;
        RECT 75.955 59.355 76.285 59.755 ;
        RECT 76.710 59.220 77.240 59.585 ;
        RECT 77.430 59.415 77.705 59.585 ;
        RECT 77.425 59.245 77.705 59.415 ;
        RECT 76.710 59.185 76.885 59.220 ;
        RECT 75.955 59.015 76.885 59.185 ;
        RECT 61.670 58.515 62.005 58.785 ;
        RECT 63.535 58.765 63.705 58.935 ;
        RECT 66.050 58.765 66.225 58.935 ;
        RECT 62.190 58.565 63.365 58.765 ;
        RECT 63.535 58.565 65.845 58.765 ;
        RECT 66.050 58.565 72.610 58.765 ;
        RECT 63.535 58.395 63.705 58.565 ;
        RECT 66.050 58.395 66.225 58.565 ;
        RECT 72.780 58.395 73.055 58.935 ;
        RECT 73.235 58.515 73.570 58.785 ;
        RECT 57.925 58.215 60.630 58.325 ;
        RECT 57.985 58.155 59.785 58.215 ;
        RECT 59.455 58.125 59.785 58.155 ;
        RECT 57.585 57.375 57.845 58.055 ;
        RECT 58.015 57.205 58.265 57.985 ;
        RECT 58.515 57.955 59.350 57.965 ;
        RECT 59.940 57.955 60.125 58.045 ;
        RECT 58.515 57.755 60.125 57.955 ;
        RECT 58.515 57.375 58.765 57.755 ;
        RECT 59.895 57.715 60.125 57.755 ;
        RECT 60.375 57.595 60.630 58.215 ;
        RECT 58.935 57.205 59.290 57.585 ;
        RECT 60.295 57.375 60.630 57.595 ;
        RECT 60.805 57.205 61.065 58.345 ;
        RECT 61.235 57.375 61.565 58.355 ;
        RECT 61.735 57.205 62.015 58.345 ;
        RECT 62.195 58.225 63.705 58.395 ;
        RECT 63.875 58.225 66.225 58.395 ;
        RECT 66.395 58.225 73.055 58.395 ;
        RECT 73.740 58.355 73.910 58.955 ;
        RECT 74.080 58.515 74.415 58.765 ;
        RECT 62.195 57.375 62.525 58.225 ;
        RECT 62.695 57.205 62.865 58.055 ;
        RECT 63.035 57.375 63.365 58.225 ;
        RECT 63.535 57.205 63.705 58.055 ;
        RECT 63.875 57.375 64.205 58.225 ;
        RECT 64.375 57.205 64.545 58.005 ;
        RECT 64.715 57.375 65.045 58.225 ;
        RECT 65.215 57.205 65.385 58.005 ;
        RECT 65.555 57.375 65.885 58.225 ;
        RECT 66.055 57.205 66.225 58.005 ;
        RECT 66.395 57.375 66.725 58.225 ;
        RECT 66.895 57.205 67.065 58.005 ;
        RECT 67.235 57.375 67.565 58.225 ;
        RECT 67.735 57.205 67.905 58.005 ;
        RECT 68.075 57.375 68.405 58.225 ;
        RECT 68.575 57.205 68.745 58.005 ;
        RECT 68.915 57.375 69.245 58.225 ;
        RECT 69.415 57.205 69.585 58.005 ;
        RECT 69.755 57.375 70.085 58.225 ;
        RECT 70.255 57.205 70.425 58.005 ;
        RECT 70.595 57.375 70.925 58.225 ;
        RECT 71.095 57.205 71.265 58.005 ;
        RECT 71.435 57.375 71.765 58.225 ;
        RECT 71.935 57.205 72.105 58.005 ;
        RECT 72.275 57.375 72.605 58.225 ;
        RECT 72.775 57.205 72.945 58.005 ;
        RECT 73.225 57.205 73.505 58.345 ;
        RECT 73.675 57.375 74.005 58.355 ;
        RECT 75.530 58.345 75.700 59.015 ;
        RECT 75.955 58.845 76.125 59.015 ;
        RECT 75.870 58.515 76.125 58.845 ;
        RECT 76.350 58.515 76.545 58.845 ;
        RECT 74.175 57.205 74.435 58.345 ;
        RECT 75.530 57.375 75.865 58.345 ;
        RECT 76.035 57.205 76.205 58.345 ;
        RECT 76.375 57.545 76.545 58.515 ;
        RECT 76.715 57.885 76.885 59.015 ;
        RECT 77.055 58.225 77.225 59.025 ;
        RECT 77.430 58.425 77.705 59.245 ;
        RECT 77.875 58.225 78.065 59.585 ;
        RECT 78.245 59.220 78.755 59.755 ;
        RECT 78.975 58.945 79.220 59.550 ;
        RECT 79.665 59.080 79.925 59.585 ;
        RECT 80.105 59.375 80.435 59.755 ;
        RECT 80.615 59.205 80.785 59.585 ;
        RECT 78.265 58.775 79.495 58.945 ;
        RECT 77.055 58.055 78.065 58.225 ;
        RECT 78.235 58.210 78.985 58.400 ;
        RECT 76.715 57.715 77.840 57.885 ;
        RECT 78.235 57.545 78.405 58.210 ;
        RECT 79.155 57.965 79.495 58.775 ;
        RECT 76.375 57.375 78.405 57.545 ;
        RECT 78.575 57.205 78.745 57.965 ;
        RECT 78.980 57.555 79.495 57.965 ;
        RECT 79.665 58.280 79.835 59.080 ;
        RECT 80.120 59.035 80.785 59.205 ;
        RECT 81.135 59.205 81.305 59.585 ;
        RECT 81.520 59.375 81.850 59.755 ;
        RECT 81.135 59.035 81.850 59.205 ;
        RECT 80.120 58.780 80.290 59.035 ;
        RECT 80.005 58.450 80.290 58.780 ;
        RECT 80.525 58.485 80.855 58.855 ;
        RECT 81.045 58.485 81.400 58.855 ;
        RECT 81.680 58.845 81.850 59.035 ;
        RECT 82.020 59.010 82.275 59.585 ;
        RECT 81.680 58.515 81.935 58.845 ;
        RECT 80.120 58.305 80.290 58.450 ;
        RECT 81.680 58.305 81.850 58.515 ;
        RECT 79.665 57.375 79.935 58.280 ;
        RECT 80.120 58.135 80.785 58.305 ;
        RECT 80.105 57.205 80.435 57.965 ;
        RECT 80.615 57.375 80.785 58.135 ;
        RECT 81.135 58.135 81.850 58.305 ;
        RECT 82.105 58.280 82.275 59.010 ;
        RECT 82.450 58.915 82.710 59.755 ;
        RECT 82.885 59.005 84.095 59.755 ;
        RECT 81.135 57.375 81.305 58.135 ;
        RECT 81.520 57.205 81.850 57.965 ;
        RECT 82.020 57.375 82.275 58.280 ;
        RECT 82.450 57.205 82.710 58.355 ;
        RECT 82.885 58.295 83.405 58.835 ;
        RECT 83.575 58.465 84.095 59.005 ;
        RECT 82.885 57.205 84.095 58.295 ;
        RECT 5.520 57.035 84.180 57.205 ;
        RECT 5.605 55.945 6.815 57.035 ;
        RECT 5.605 55.235 6.125 55.775 ;
        RECT 6.295 55.405 6.815 55.945 ;
        RECT 6.990 55.885 7.250 57.035 ;
        RECT 7.425 55.960 7.680 56.865 ;
        RECT 7.850 56.275 8.180 57.035 ;
        RECT 8.395 56.105 8.565 56.865 ;
        RECT 8.915 56.365 9.085 56.865 ;
        RECT 9.255 56.535 9.585 57.035 ;
        RECT 8.915 56.195 9.580 56.365 ;
        RECT 5.605 54.485 6.815 55.235 ;
        RECT 6.990 54.485 7.250 55.325 ;
        RECT 7.425 55.230 7.595 55.960 ;
        RECT 7.850 55.935 8.565 56.105 ;
        RECT 7.850 55.725 8.020 55.935 ;
        RECT 7.765 55.395 8.020 55.725 ;
        RECT 7.425 54.655 7.680 55.230 ;
        RECT 7.850 55.205 8.020 55.395 ;
        RECT 8.300 55.385 8.655 55.755 ;
        RECT 8.830 55.375 9.180 56.025 ;
        RECT 9.350 55.205 9.580 56.195 ;
        RECT 7.850 55.035 8.565 55.205 ;
        RECT 7.850 54.485 8.180 54.865 ;
        RECT 8.395 54.655 8.565 55.035 ;
        RECT 8.915 55.035 9.580 55.205 ;
        RECT 8.915 54.745 9.085 55.035 ;
        RECT 9.255 54.485 9.585 54.865 ;
        RECT 9.755 54.745 9.940 56.865 ;
        RECT 10.180 56.575 10.445 57.035 ;
        RECT 10.615 56.440 10.865 56.865 ;
        RECT 11.075 56.590 12.180 56.760 ;
        RECT 10.560 56.310 10.865 56.440 ;
        RECT 10.110 55.115 10.390 56.065 ;
        RECT 10.560 55.205 10.730 56.310 ;
        RECT 10.900 55.525 11.140 56.120 ;
        RECT 11.310 56.055 11.840 56.420 ;
        RECT 11.310 55.355 11.480 56.055 ;
        RECT 12.010 55.975 12.180 56.590 ;
        RECT 12.350 56.235 12.520 57.035 ;
        RECT 12.690 56.535 12.940 56.865 ;
        RECT 13.165 56.565 14.050 56.735 ;
        RECT 12.010 55.885 12.520 55.975 ;
        RECT 10.560 55.075 10.785 55.205 ;
        RECT 10.955 55.135 11.480 55.355 ;
        RECT 11.650 55.715 12.520 55.885 ;
        RECT 10.195 54.485 10.445 54.945 ;
        RECT 10.615 54.935 10.785 55.075 ;
        RECT 11.650 54.935 11.820 55.715 ;
        RECT 12.350 55.645 12.520 55.715 ;
        RECT 12.030 55.465 12.230 55.495 ;
        RECT 12.690 55.465 12.860 56.535 ;
        RECT 13.030 55.645 13.220 56.365 ;
        RECT 12.030 55.165 12.860 55.465 ;
        RECT 13.390 55.435 13.710 56.395 ;
        RECT 10.615 54.765 10.950 54.935 ;
        RECT 11.145 54.765 11.820 54.935 ;
        RECT 12.140 54.485 12.510 54.985 ;
        RECT 12.690 54.935 12.860 55.165 ;
        RECT 13.245 55.105 13.710 55.435 ;
        RECT 13.880 55.725 14.050 56.565 ;
        RECT 14.230 56.535 14.545 57.035 ;
        RECT 14.775 56.305 15.115 56.865 ;
        RECT 14.220 55.930 15.115 56.305 ;
        RECT 15.285 56.025 15.455 57.035 ;
        RECT 14.925 55.725 15.115 55.930 ;
        RECT 15.625 55.975 15.955 56.820 ;
        RECT 15.625 55.895 16.015 55.975 ;
        RECT 16.185 55.945 17.855 57.035 ;
        RECT 15.800 55.845 16.015 55.895 ;
        RECT 13.880 55.395 14.755 55.725 ;
        RECT 14.925 55.395 15.675 55.725 ;
        RECT 13.880 54.935 14.050 55.395 ;
        RECT 14.925 55.225 15.125 55.395 ;
        RECT 15.845 55.265 16.015 55.845 ;
        RECT 15.790 55.225 16.015 55.265 ;
        RECT 12.690 54.765 13.095 54.935 ;
        RECT 13.265 54.765 14.050 54.935 ;
        RECT 14.325 54.485 14.535 55.015 ;
        RECT 14.795 54.700 15.125 55.225 ;
        RECT 15.635 55.140 16.015 55.225 ;
        RECT 16.185 55.255 16.935 55.775 ;
        RECT 17.105 55.425 17.855 55.945 ;
        RECT 18.485 55.870 18.775 57.035 ;
        RECT 19.130 56.065 19.520 56.240 ;
        RECT 20.005 56.235 20.335 57.035 ;
        RECT 20.505 56.245 21.040 56.865 ;
        RECT 19.130 55.895 20.555 56.065 ;
        RECT 15.295 54.485 15.465 55.095 ;
        RECT 15.635 54.705 15.965 55.140 ;
        RECT 16.185 54.485 17.855 55.255 ;
        RECT 18.485 54.485 18.775 55.210 ;
        RECT 19.005 55.165 19.360 55.725 ;
        RECT 19.530 54.995 19.700 55.895 ;
        RECT 19.870 55.165 20.135 55.725 ;
        RECT 20.385 55.395 20.555 55.895 ;
        RECT 20.725 55.225 21.040 56.245 ;
        RECT 21.910 56.065 22.240 56.865 ;
        RECT 22.410 56.235 22.740 57.035 ;
        RECT 23.040 56.065 23.370 56.865 ;
        RECT 24.015 56.235 24.265 57.035 ;
        RECT 21.910 55.895 24.345 56.065 ;
        RECT 24.535 55.895 24.705 57.035 ;
        RECT 24.875 55.895 25.215 56.865 ;
        RECT 25.385 55.945 27.055 57.035 ;
        RECT 27.315 56.365 27.485 56.865 ;
        RECT 27.655 56.535 27.985 57.035 ;
        RECT 27.315 56.195 27.980 56.365 ;
        RECT 21.705 55.475 22.055 55.725 ;
        RECT 22.240 55.265 22.410 55.895 ;
        RECT 22.580 55.475 22.910 55.675 ;
        RECT 23.080 55.475 23.410 55.675 ;
        RECT 23.580 55.475 24.000 55.675 ;
        RECT 24.175 55.645 24.345 55.895 ;
        RECT 24.175 55.475 24.870 55.645 ;
        RECT 19.110 54.485 19.350 54.995 ;
        RECT 19.530 54.665 19.810 54.995 ;
        RECT 20.040 54.485 20.255 54.995 ;
        RECT 20.425 54.655 21.040 55.225 ;
        RECT 21.910 54.655 22.410 55.265 ;
        RECT 23.040 55.135 24.265 55.305 ;
        RECT 25.040 55.285 25.215 55.895 ;
        RECT 23.040 54.655 23.370 55.135 ;
        RECT 23.540 54.485 23.765 54.945 ;
        RECT 23.935 54.655 24.265 55.135 ;
        RECT 24.455 54.485 24.705 55.285 ;
        RECT 24.875 54.655 25.215 55.285 ;
        RECT 25.385 55.255 26.135 55.775 ;
        RECT 26.305 55.425 27.055 55.945 ;
        RECT 27.230 55.375 27.580 56.025 ;
        RECT 25.385 54.485 27.055 55.255 ;
        RECT 27.750 55.205 27.980 56.195 ;
        RECT 27.315 55.035 27.980 55.205 ;
        RECT 27.315 54.745 27.485 55.035 ;
        RECT 27.655 54.485 27.985 54.865 ;
        RECT 28.155 54.745 28.340 56.865 ;
        RECT 28.580 56.575 28.845 57.035 ;
        RECT 29.015 56.440 29.265 56.865 ;
        RECT 29.475 56.590 30.580 56.760 ;
        RECT 28.960 56.310 29.265 56.440 ;
        RECT 28.510 55.115 28.790 56.065 ;
        RECT 28.960 55.205 29.130 56.310 ;
        RECT 29.300 55.525 29.540 56.120 ;
        RECT 29.710 56.055 30.240 56.420 ;
        RECT 29.710 55.355 29.880 56.055 ;
        RECT 30.410 55.975 30.580 56.590 ;
        RECT 30.750 56.235 30.920 57.035 ;
        RECT 31.090 56.535 31.340 56.865 ;
        RECT 31.565 56.565 32.450 56.735 ;
        RECT 30.410 55.885 30.920 55.975 ;
        RECT 28.960 55.075 29.185 55.205 ;
        RECT 29.355 55.135 29.880 55.355 ;
        RECT 30.050 55.715 30.920 55.885 ;
        RECT 28.595 54.485 28.845 54.945 ;
        RECT 29.015 54.935 29.185 55.075 ;
        RECT 30.050 54.935 30.220 55.715 ;
        RECT 30.750 55.645 30.920 55.715 ;
        RECT 30.430 55.465 30.630 55.495 ;
        RECT 31.090 55.465 31.260 56.535 ;
        RECT 31.430 55.645 31.620 56.365 ;
        RECT 30.430 55.165 31.260 55.465 ;
        RECT 31.790 55.435 32.110 56.395 ;
        RECT 29.015 54.765 29.350 54.935 ;
        RECT 29.545 54.765 30.220 54.935 ;
        RECT 30.540 54.485 30.910 54.985 ;
        RECT 31.090 54.935 31.260 55.165 ;
        RECT 31.645 55.105 32.110 55.435 ;
        RECT 32.280 55.725 32.450 56.565 ;
        RECT 32.630 56.535 32.945 57.035 ;
        RECT 33.175 56.305 33.515 56.865 ;
        RECT 32.620 55.930 33.515 56.305 ;
        RECT 33.685 56.025 33.855 57.035 ;
        RECT 33.325 55.725 33.515 55.930 ;
        RECT 34.025 55.975 34.355 56.820 ;
        RECT 34.025 55.895 34.415 55.975 ;
        RECT 34.200 55.845 34.415 55.895 ;
        RECT 32.280 55.395 33.155 55.725 ;
        RECT 33.325 55.395 34.075 55.725 ;
        RECT 32.280 54.935 32.450 55.395 ;
        RECT 33.325 55.225 33.525 55.395 ;
        RECT 34.245 55.265 34.415 55.845 ;
        RECT 34.190 55.225 34.415 55.265 ;
        RECT 31.090 54.765 31.495 54.935 ;
        RECT 31.665 54.765 32.450 54.935 ;
        RECT 32.725 54.485 32.935 55.015 ;
        RECT 33.195 54.700 33.525 55.225 ;
        RECT 34.035 55.140 34.415 55.225 ;
        RECT 34.590 55.895 34.925 56.865 ;
        RECT 35.095 55.895 35.265 57.035 ;
        RECT 35.435 56.695 37.465 56.865 ;
        RECT 34.590 55.225 34.760 55.895 ;
        RECT 35.435 55.725 35.605 56.695 ;
        RECT 34.930 55.395 35.185 55.725 ;
        RECT 35.410 55.395 35.605 55.725 ;
        RECT 35.775 56.355 36.900 56.525 ;
        RECT 35.015 55.225 35.185 55.395 ;
        RECT 35.775 55.225 35.945 56.355 ;
        RECT 33.695 54.485 33.865 55.095 ;
        RECT 34.035 54.705 34.365 55.140 ;
        RECT 34.590 54.655 34.845 55.225 ;
        RECT 35.015 55.055 35.945 55.225 ;
        RECT 36.115 56.015 37.125 56.185 ;
        RECT 36.115 55.215 36.285 56.015 ;
        RECT 35.770 55.020 35.945 55.055 ;
        RECT 35.015 54.485 35.345 54.885 ;
        RECT 35.770 54.655 36.300 55.020 ;
        RECT 36.490 54.995 36.765 55.815 ;
        RECT 36.485 54.825 36.765 54.995 ;
        RECT 36.490 54.655 36.765 54.825 ;
        RECT 36.935 54.655 37.125 56.015 ;
        RECT 37.295 56.030 37.465 56.695 ;
        RECT 37.635 56.275 37.805 57.035 ;
        RECT 38.040 56.275 38.555 56.685 ;
        RECT 37.295 55.840 38.045 56.030 ;
        RECT 38.215 55.465 38.555 56.275 ;
        RECT 37.325 55.295 38.555 55.465 ;
        RECT 39.185 56.275 39.700 56.685 ;
        RECT 39.935 56.275 40.105 57.035 ;
        RECT 40.275 56.695 42.305 56.865 ;
        RECT 39.185 55.465 39.525 56.275 ;
        RECT 40.275 56.030 40.445 56.695 ;
        RECT 40.840 56.355 41.965 56.525 ;
        RECT 39.695 55.840 40.445 56.030 ;
        RECT 40.615 56.015 41.625 56.185 ;
        RECT 39.185 55.295 40.415 55.465 ;
        RECT 37.305 54.485 37.815 55.020 ;
        RECT 38.035 54.690 38.280 55.295 ;
        RECT 39.460 54.690 39.705 55.295 ;
        RECT 39.925 54.485 40.435 55.020 ;
        RECT 40.615 54.655 40.805 56.015 ;
        RECT 40.975 55.675 41.250 55.815 ;
        RECT 40.975 55.505 41.255 55.675 ;
        RECT 40.975 54.655 41.250 55.505 ;
        RECT 41.455 55.215 41.625 56.015 ;
        RECT 41.795 55.225 41.965 56.355 ;
        RECT 42.135 55.725 42.305 56.695 ;
        RECT 42.475 55.895 42.645 57.035 ;
        RECT 42.815 55.895 43.150 56.865 ;
        RECT 42.135 55.395 42.330 55.725 ;
        RECT 42.555 55.395 42.810 55.725 ;
        RECT 42.555 55.225 42.725 55.395 ;
        RECT 42.980 55.225 43.150 55.895 ;
        RECT 44.245 55.870 44.535 57.035 ;
        RECT 44.705 55.945 48.215 57.035 ;
        RECT 41.795 55.055 42.725 55.225 ;
        RECT 41.795 55.020 41.970 55.055 ;
        RECT 41.440 54.655 41.970 55.020 ;
        RECT 42.395 54.485 42.725 54.885 ;
        RECT 42.895 54.655 43.150 55.225 ;
        RECT 44.705 55.255 46.355 55.775 ;
        RECT 46.525 55.425 48.215 55.945 ;
        RECT 48.390 55.895 48.725 56.865 ;
        RECT 48.895 55.895 49.065 57.035 ;
        RECT 49.235 56.695 51.265 56.865 ;
        RECT 44.245 54.485 44.535 55.210 ;
        RECT 44.705 54.485 48.215 55.255 ;
        RECT 48.390 55.225 48.560 55.895 ;
        RECT 49.235 55.725 49.405 56.695 ;
        RECT 48.730 55.395 48.985 55.725 ;
        RECT 49.210 55.395 49.405 55.725 ;
        RECT 49.575 56.355 50.700 56.525 ;
        RECT 48.815 55.225 48.985 55.395 ;
        RECT 49.575 55.225 49.745 56.355 ;
        RECT 48.390 54.655 48.645 55.225 ;
        RECT 48.815 55.055 49.745 55.225 ;
        RECT 49.915 56.015 50.925 56.185 ;
        RECT 49.915 55.215 50.085 56.015 ;
        RECT 49.570 55.020 49.745 55.055 ;
        RECT 48.815 54.485 49.145 54.885 ;
        RECT 49.570 54.655 50.100 55.020 ;
        RECT 50.290 54.995 50.565 55.815 ;
        RECT 50.285 54.825 50.565 54.995 ;
        RECT 50.290 54.655 50.565 54.825 ;
        RECT 50.735 54.655 50.925 56.015 ;
        RECT 51.095 56.030 51.265 56.695 ;
        RECT 51.435 56.275 51.605 57.035 ;
        RECT 51.840 56.275 52.355 56.685 ;
        RECT 52.525 56.600 57.870 57.035 ;
        RECT 51.095 55.840 51.845 56.030 ;
        RECT 52.015 55.465 52.355 56.275 ;
        RECT 51.125 55.295 52.355 55.465 ;
        RECT 51.105 54.485 51.615 55.020 ;
        RECT 51.835 54.690 52.080 55.295 ;
        RECT 54.110 55.030 54.450 55.860 ;
        RECT 55.930 55.350 56.280 56.600 ;
        RECT 58.045 56.185 58.305 56.865 ;
        RECT 58.475 56.255 58.725 57.035 ;
        RECT 58.975 56.485 59.225 56.865 ;
        RECT 59.395 56.655 59.750 57.035 ;
        RECT 60.755 56.645 61.090 56.865 ;
        RECT 60.355 56.485 60.585 56.525 ;
        RECT 58.975 56.285 60.585 56.485 ;
        RECT 58.975 56.275 59.810 56.285 ;
        RECT 60.400 56.195 60.585 56.285 ;
        RECT 52.525 54.485 57.870 55.030 ;
        RECT 58.045 54.995 58.215 56.185 ;
        RECT 59.915 56.085 60.245 56.115 ;
        RECT 58.445 56.025 60.245 56.085 ;
        RECT 60.835 56.025 61.090 56.645 ;
        RECT 58.385 55.915 61.090 56.025 ;
        RECT 58.385 55.880 58.585 55.915 ;
        RECT 58.385 55.305 58.555 55.880 ;
        RECT 59.915 55.855 61.090 55.915 ;
        RECT 61.265 55.895 61.545 57.035 ;
        RECT 61.715 55.885 62.045 56.865 ;
        RECT 62.215 55.895 62.475 57.035 ;
        RECT 62.655 55.975 62.985 56.825 ;
        RECT 61.780 55.845 61.955 55.885 ;
        RECT 58.785 55.440 59.195 55.745 ;
        RECT 59.365 55.475 59.695 55.685 ;
        RECT 58.385 55.185 58.655 55.305 ;
        RECT 58.385 55.140 59.230 55.185 ;
        RECT 58.475 55.015 59.230 55.140 ;
        RECT 59.485 55.075 59.695 55.475 ;
        RECT 59.940 55.475 60.415 55.685 ;
        RECT 60.605 55.475 61.095 55.675 ;
        RECT 59.940 55.075 60.160 55.475 ;
        RECT 61.275 55.455 61.610 55.725 ;
        RECT 61.780 55.285 61.950 55.845 ;
        RECT 62.120 55.475 62.455 55.725 ;
        RECT 58.045 54.985 58.275 54.995 ;
        RECT 58.045 54.655 58.305 54.985 ;
        RECT 59.060 54.865 59.230 55.015 ;
        RECT 58.475 54.485 58.805 54.845 ;
        RECT 59.060 54.655 60.360 54.865 ;
        RECT 60.635 54.485 61.090 55.250 ;
        RECT 61.265 54.485 61.575 55.285 ;
        RECT 61.780 54.655 62.475 55.285 ;
        RECT 62.655 55.210 62.845 55.975 ;
        RECT 63.155 55.895 63.405 57.035 ;
        RECT 63.595 56.395 63.845 56.815 ;
        RECT 64.075 56.565 64.405 57.035 ;
        RECT 64.635 56.395 64.885 56.815 ;
        RECT 63.595 56.225 64.885 56.395 ;
        RECT 65.065 56.395 65.395 56.825 ;
        RECT 65.065 56.225 65.520 56.395 ;
        RECT 63.585 55.725 63.800 56.055 ;
        RECT 63.015 55.395 63.325 55.725 ;
        RECT 63.495 55.395 63.800 55.725 ;
        RECT 63.975 55.395 64.260 56.055 ;
        RECT 64.455 55.395 64.720 56.055 ;
        RECT 64.935 55.395 65.180 56.055 ;
        RECT 63.155 55.225 63.325 55.395 ;
        RECT 65.350 55.225 65.520 56.225 ;
        RECT 66.020 56.025 66.320 56.865 ;
        RECT 66.515 56.195 66.765 57.035 ;
        RECT 67.355 56.445 68.160 56.865 ;
        RECT 66.935 56.275 68.500 56.445 ;
        RECT 66.935 56.025 67.105 56.275 ;
        RECT 66.020 55.855 67.105 56.025 ;
        RECT 65.865 55.395 66.195 55.685 ;
        RECT 66.365 55.225 66.535 55.855 ;
        RECT 67.275 55.725 67.595 56.105 ;
        RECT 67.785 56.015 68.160 56.105 ;
        RECT 67.765 55.845 68.160 56.015 ;
        RECT 68.330 56.025 68.500 56.275 ;
        RECT 68.670 56.195 69.000 57.035 ;
        RECT 69.170 56.275 69.835 56.865 ;
        RECT 68.330 55.855 69.250 56.025 ;
        RECT 66.705 55.475 67.035 55.685 ;
        RECT 67.215 55.475 67.595 55.725 ;
        RECT 67.785 55.685 68.160 55.845 ;
        RECT 69.080 55.685 69.250 55.855 ;
        RECT 67.785 55.475 68.270 55.685 ;
        RECT 68.460 55.475 68.910 55.685 ;
        RECT 69.080 55.475 69.415 55.685 ;
        RECT 69.585 55.305 69.835 56.275 ;
        RECT 70.005 55.870 70.295 57.035 ;
        RECT 70.470 56.645 70.805 56.865 ;
        RECT 71.810 56.655 72.165 57.035 ;
        RECT 70.470 56.025 70.725 56.645 ;
        RECT 70.975 56.485 71.205 56.525 ;
        RECT 72.335 56.485 72.585 56.865 ;
        RECT 70.975 56.285 72.585 56.485 ;
        RECT 70.975 56.195 71.160 56.285 ;
        RECT 71.750 56.275 72.585 56.285 ;
        RECT 72.835 56.255 73.085 57.035 ;
        RECT 73.255 56.185 73.515 56.865 ;
        RECT 74.235 56.365 74.405 56.865 ;
        RECT 74.575 56.535 74.905 57.035 ;
        RECT 74.235 56.195 74.900 56.365 ;
        RECT 71.315 56.085 71.645 56.115 ;
        RECT 71.315 56.025 73.115 56.085 ;
        RECT 70.470 55.915 73.175 56.025 ;
        RECT 70.470 55.855 71.645 55.915 ;
        RECT 72.975 55.880 73.175 55.915 ;
        RECT 70.465 55.475 70.955 55.675 ;
        RECT 71.145 55.475 71.620 55.685 ;
        RECT 62.655 54.700 62.985 55.210 ;
        RECT 63.155 55.055 65.520 55.225 ;
        RECT 63.155 54.485 63.485 54.885 ;
        RECT 64.535 54.715 64.865 55.055 ;
        RECT 66.025 55.045 66.535 55.225 ;
        RECT 66.940 55.135 68.640 55.305 ;
        RECT 66.940 55.045 67.325 55.135 ;
        RECT 65.035 54.485 65.365 54.885 ;
        RECT 66.025 54.655 66.355 55.045 ;
        RECT 66.525 54.705 67.710 54.875 ;
        RECT 67.970 54.485 68.140 54.955 ;
        RECT 68.310 54.670 68.640 55.135 ;
        RECT 68.810 54.485 68.980 55.305 ;
        RECT 69.150 54.665 69.835 55.305 ;
        RECT 70.005 54.485 70.295 55.210 ;
        RECT 70.470 54.485 70.925 55.250 ;
        RECT 71.400 55.075 71.620 55.475 ;
        RECT 71.865 55.475 72.195 55.685 ;
        RECT 71.865 55.075 72.075 55.475 ;
        RECT 72.365 55.440 72.775 55.745 ;
        RECT 73.005 55.305 73.175 55.880 ;
        RECT 72.905 55.185 73.175 55.305 ;
        RECT 72.330 55.140 73.175 55.185 ;
        RECT 72.330 55.015 73.085 55.140 ;
        RECT 72.330 54.865 72.500 55.015 ;
        RECT 73.345 54.985 73.515 56.185 ;
        RECT 74.150 55.375 74.500 56.025 ;
        RECT 74.670 55.205 74.900 56.195 ;
        RECT 71.200 54.655 72.500 54.865 ;
        RECT 72.755 54.485 73.085 54.845 ;
        RECT 73.255 54.655 73.515 54.985 ;
        RECT 74.235 55.035 74.900 55.205 ;
        RECT 74.235 54.745 74.405 55.035 ;
        RECT 74.575 54.485 74.905 54.865 ;
        RECT 75.075 54.745 75.260 56.865 ;
        RECT 75.500 56.575 75.765 57.035 ;
        RECT 75.935 56.440 76.185 56.865 ;
        RECT 76.395 56.590 77.500 56.760 ;
        RECT 75.880 56.310 76.185 56.440 ;
        RECT 75.430 55.115 75.710 56.065 ;
        RECT 75.880 55.205 76.050 56.310 ;
        RECT 76.220 55.525 76.460 56.120 ;
        RECT 76.630 56.055 77.160 56.420 ;
        RECT 76.630 55.355 76.800 56.055 ;
        RECT 77.330 55.975 77.500 56.590 ;
        RECT 77.670 56.235 77.840 57.035 ;
        RECT 78.010 56.535 78.260 56.865 ;
        RECT 78.485 56.565 79.370 56.735 ;
        RECT 77.330 55.885 77.840 55.975 ;
        RECT 75.880 55.075 76.105 55.205 ;
        RECT 76.275 55.135 76.800 55.355 ;
        RECT 76.970 55.715 77.840 55.885 ;
        RECT 75.515 54.485 75.765 54.945 ;
        RECT 75.935 54.935 76.105 55.075 ;
        RECT 76.970 54.935 77.140 55.715 ;
        RECT 77.670 55.645 77.840 55.715 ;
        RECT 77.350 55.465 77.550 55.495 ;
        RECT 78.010 55.465 78.180 56.535 ;
        RECT 78.350 55.645 78.540 56.365 ;
        RECT 77.350 55.165 78.180 55.465 ;
        RECT 78.710 55.435 79.030 56.395 ;
        RECT 75.935 54.765 76.270 54.935 ;
        RECT 76.465 54.765 77.140 54.935 ;
        RECT 77.460 54.485 77.830 54.985 ;
        RECT 78.010 54.935 78.180 55.165 ;
        RECT 78.565 55.105 79.030 55.435 ;
        RECT 79.200 55.725 79.370 56.565 ;
        RECT 79.550 56.535 79.865 57.035 ;
        RECT 80.095 56.305 80.435 56.865 ;
        RECT 79.540 55.930 80.435 56.305 ;
        RECT 80.605 56.025 80.775 57.035 ;
        RECT 80.245 55.725 80.435 55.930 ;
        RECT 80.945 55.975 81.275 56.820 ;
        RECT 80.945 55.895 81.335 55.975 ;
        RECT 81.120 55.845 81.335 55.895 ;
        RECT 79.200 55.395 80.075 55.725 ;
        RECT 80.245 55.395 80.995 55.725 ;
        RECT 79.200 54.935 79.370 55.395 ;
        RECT 80.245 55.225 80.445 55.395 ;
        RECT 81.165 55.265 81.335 55.845 ;
        RECT 81.110 55.225 81.335 55.265 ;
        RECT 78.010 54.765 78.415 54.935 ;
        RECT 78.585 54.765 79.370 54.935 ;
        RECT 79.645 54.485 79.855 55.015 ;
        RECT 80.115 54.700 80.445 55.225 ;
        RECT 80.955 55.140 81.335 55.225 ;
        RECT 81.505 55.960 81.775 56.865 ;
        RECT 81.945 56.275 82.275 57.035 ;
        RECT 82.455 56.105 82.625 56.865 ;
        RECT 81.505 55.160 81.675 55.960 ;
        RECT 81.960 55.935 82.625 56.105 ;
        RECT 82.885 55.945 84.095 57.035 ;
        RECT 81.960 55.790 82.130 55.935 ;
        RECT 81.845 55.460 82.130 55.790 ;
        RECT 81.960 55.205 82.130 55.460 ;
        RECT 82.365 55.385 82.695 55.755 ;
        RECT 82.885 55.405 83.405 55.945 ;
        RECT 83.575 55.235 84.095 55.775 ;
        RECT 80.615 54.485 80.785 55.095 ;
        RECT 80.955 54.705 81.285 55.140 ;
        RECT 81.505 54.655 81.765 55.160 ;
        RECT 81.960 55.035 82.625 55.205 ;
        RECT 81.945 54.485 82.275 54.865 ;
        RECT 82.455 54.655 82.625 55.035 ;
        RECT 82.885 54.485 84.095 55.235 ;
        RECT 5.520 54.315 84.180 54.485 ;
        RECT 5.605 53.565 6.815 54.315 ;
        RECT 6.985 53.565 8.195 54.315 ;
        RECT 5.605 53.025 6.125 53.565 ;
        RECT 6.295 52.855 6.815 53.395 ;
        RECT 6.985 53.025 7.505 53.565 ;
        RECT 8.365 53.515 8.705 54.145 ;
        RECT 8.875 53.515 9.125 54.315 ;
        RECT 9.315 53.665 9.645 54.145 ;
        RECT 9.815 53.855 10.040 54.315 ;
        RECT 10.210 53.665 10.540 54.145 ;
        RECT 7.675 52.855 8.195 53.395 ;
        RECT 5.605 51.765 6.815 52.855 ;
        RECT 6.985 51.765 8.195 52.855 ;
        RECT 8.365 52.905 8.540 53.515 ;
        RECT 9.315 53.495 10.540 53.665 ;
        RECT 11.170 53.535 11.670 54.145 ;
        RECT 8.710 53.155 9.405 53.325 ;
        RECT 9.235 52.905 9.405 53.155 ;
        RECT 9.580 53.125 10.000 53.325 ;
        RECT 10.170 53.125 10.500 53.325 ;
        RECT 10.670 53.125 11.000 53.325 ;
        RECT 11.170 52.905 11.340 53.535 ;
        RECT 12.045 53.515 12.385 54.145 ;
        RECT 12.555 53.515 12.805 54.315 ;
        RECT 12.995 53.665 13.325 54.145 ;
        RECT 13.495 53.855 13.720 54.315 ;
        RECT 13.890 53.665 14.220 54.145 ;
        RECT 11.525 53.075 11.875 53.325 ;
        RECT 12.045 52.905 12.220 53.515 ;
        RECT 12.995 53.495 14.220 53.665 ;
        RECT 14.850 53.535 15.350 54.145 ;
        RECT 15.775 53.775 16.000 54.135 ;
        RECT 16.180 53.945 16.510 54.315 ;
        RECT 16.690 53.775 16.945 54.135 ;
        RECT 17.510 53.945 18.255 54.315 ;
        RECT 15.775 53.585 18.260 53.775 ;
        RECT 12.390 53.155 13.085 53.325 ;
        RECT 12.915 52.905 13.085 53.155 ;
        RECT 13.260 53.125 13.680 53.325 ;
        RECT 13.850 53.125 14.180 53.325 ;
        RECT 14.350 53.125 14.680 53.325 ;
        RECT 14.850 52.905 15.020 53.535 ;
        RECT 15.205 53.075 15.555 53.325 ;
        RECT 15.735 53.075 16.005 53.405 ;
        RECT 16.185 53.075 16.620 53.405 ;
        RECT 16.800 53.075 17.375 53.405 ;
        RECT 17.555 53.075 17.835 53.405 ;
        RECT 8.365 51.935 8.705 52.905 ;
        RECT 8.875 51.765 9.045 52.905 ;
        RECT 9.235 52.735 11.670 52.905 ;
        RECT 9.315 51.765 9.565 52.565 ;
        RECT 10.210 51.935 10.540 52.735 ;
        RECT 10.840 51.765 11.170 52.565 ;
        RECT 11.340 51.935 11.670 52.735 ;
        RECT 12.045 51.935 12.385 52.905 ;
        RECT 12.555 51.765 12.725 52.905 ;
        RECT 12.915 52.735 15.350 52.905 ;
        RECT 18.035 52.895 18.260 53.585 ;
        RECT 12.995 51.765 13.245 52.565 ;
        RECT 13.890 51.935 14.220 52.735 ;
        RECT 14.520 51.765 14.850 52.565 ;
        RECT 15.020 51.935 15.350 52.735 ;
        RECT 15.765 52.715 18.260 52.895 ;
        RECT 18.435 52.715 18.770 54.135 ;
        RECT 19.150 53.535 19.650 54.145 ;
        RECT 18.945 53.075 19.295 53.325 ;
        RECT 19.480 52.905 19.650 53.535 ;
        RECT 20.280 53.665 20.610 54.145 ;
        RECT 20.780 53.855 21.005 54.315 ;
        RECT 21.175 53.665 21.505 54.145 ;
        RECT 20.280 53.495 21.505 53.665 ;
        RECT 21.695 53.515 21.945 54.315 ;
        RECT 22.115 53.515 22.455 54.145 ;
        RECT 22.715 53.765 22.885 54.055 ;
        RECT 23.055 53.935 23.385 54.315 ;
        RECT 22.715 53.595 23.380 53.765 ;
        RECT 22.225 53.465 22.455 53.515 ;
        RECT 19.820 53.125 20.150 53.325 ;
        RECT 20.320 53.125 20.650 53.325 ;
        RECT 20.820 53.125 21.240 53.325 ;
        RECT 21.415 53.155 22.110 53.325 ;
        RECT 21.415 52.905 21.585 53.155 ;
        RECT 22.280 52.905 22.455 53.465 ;
        RECT 15.765 51.945 16.055 52.715 ;
        RECT 16.625 52.305 17.815 52.535 ;
        RECT 16.625 51.945 16.885 52.305 ;
        RECT 17.055 51.765 17.385 52.135 ;
        RECT 17.555 51.945 17.815 52.305 ;
        RECT 18.005 51.765 18.335 52.485 ;
        RECT 18.505 51.945 18.770 52.715 ;
        RECT 19.150 52.735 21.585 52.905 ;
        RECT 19.150 51.935 19.480 52.735 ;
        RECT 19.650 51.765 19.980 52.565 ;
        RECT 20.280 51.935 20.610 52.735 ;
        RECT 21.255 51.765 21.505 52.565 ;
        RECT 21.775 51.765 21.945 52.905 ;
        RECT 22.115 51.935 22.455 52.905 ;
        RECT 22.630 52.775 22.980 53.425 ;
        RECT 23.150 52.605 23.380 53.595 ;
        RECT 22.715 52.435 23.380 52.605 ;
        RECT 22.715 51.935 22.885 52.435 ;
        RECT 23.055 51.765 23.385 52.265 ;
        RECT 23.555 51.935 23.740 54.055 ;
        RECT 23.995 53.855 24.245 54.315 ;
        RECT 24.415 53.865 24.750 54.035 ;
        RECT 24.945 53.865 25.620 54.035 ;
        RECT 24.415 53.725 24.585 53.865 ;
        RECT 23.910 52.735 24.190 53.685 ;
        RECT 24.360 53.595 24.585 53.725 ;
        RECT 24.360 52.490 24.530 53.595 ;
        RECT 24.755 53.445 25.280 53.665 ;
        RECT 24.700 52.680 24.940 53.275 ;
        RECT 25.110 52.745 25.280 53.445 ;
        RECT 25.450 53.085 25.620 53.865 ;
        RECT 25.940 53.815 26.310 54.315 ;
        RECT 26.490 53.865 26.895 54.035 ;
        RECT 27.065 53.865 27.850 54.035 ;
        RECT 26.490 53.635 26.660 53.865 ;
        RECT 25.830 53.335 26.660 53.635 ;
        RECT 27.045 53.365 27.510 53.695 ;
        RECT 25.830 53.305 26.030 53.335 ;
        RECT 26.150 53.085 26.320 53.155 ;
        RECT 25.450 52.915 26.320 53.085 ;
        RECT 25.810 52.825 26.320 52.915 ;
        RECT 24.360 52.360 24.665 52.490 ;
        RECT 25.110 52.380 25.640 52.745 ;
        RECT 23.980 51.765 24.245 52.225 ;
        RECT 24.415 51.935 24.665 52.360 ;
        RECT 25.810 52.210 25.980 52.825 ;
        RECT 24.875 52.040 25.980 52.210 ;
        RECT 26.150 51.765 26.320 52.565 ;
        RECT 26.490 52.265 26.660 53.335 ;
        RECT 26.830 52.435 27.020 53.155 ;
        RECT 27.190 52.405 27.510 53.365 ;
        RECT 27.680 53.405 27.850 53.865 ;
        RECT 28.125 53.785 28.335 54.315 ;
        RECT 28.595 53.575 28.925 54.100 ;
        RECT 29.095 53.705 29.265 54.315 ;
        RECT 29.435 53.660 29.765 54.095 ;
        RECT 29.435 53.575 29.815 53.660 ;
        RECT 28.725 53.405 28.925 53.575 ;
        RECT 29.590 53.535 29.815 53.575 ;
        RECT 27.680 53.075 28.555 53.405 ;
        RECT 28.725 53.075 29.475 53.405 ;
        RECT 26.490 51.935 26.740 52.265 ;
        RECT 27.680 52.235 27.850 53.075 ;
        RECT 28.725 52.870 28.915 53.075 ;
        RECT 29.645 52.955 29.815 53.535 ;
        RECT 29.985 53.565 31.195 54.315 ;
        RECT 31.365 53.590 31.655 54.315 ;
        RECT 31.830 53.575 32.085 54.145 ;
        RECT 32.255 53.915 32.585 54.315 ;
        RECT 33.010 53.780 33.540 54.145 ;
        RECT 33.010 53.745 33.185 53.780 ;
        RECT 32.255 53.575 33.185 53.745 ;
        RECT 29.985 53.025 30.505 53.565 ;
        RECT 29.600 52.905 29.815 52.955 ;
        RECT 28.020 52.495 28.915 52.870 ;
        RECT 29.425 52.825 29.815 52.905 ;
        RECT 30.675 52.855 31.195 53.395 ;
        RECT 26.965 52.065 27.850 52.235 ;
        RECT 28.030 51.765 28.345 52.265 ;
        RECT 28.575 51.935 28.915 52.495 ;
        RECT 29.085 51.765 29.255 52.775 ;
        RECT 29.425 51.980 29.755 52.825 ;
        RECT 29.985 51.765 31.195 52.855 ;
        RECT 31.365 51.765 31.655 52.930 ;
        RECT 31.830 52.905 32.000 53.575 ;
        RECT 32.255 53.405 32.425 53.575 ;
        RECT 32.170 53.075 32.425 53.405 ;
        RECT 32.650 53.075 32.845 53.405 ;
        RECT 31.830 51.935 32.165 52.905 ;
        RECT 32.335 51.765 32.505 52.905 ;
        RECT 32.675 52.105 32.845 53.075 ;
        RECT 33.015 52.445 33.185 53.575 ;
        RECT 33.355 52.785 33.525 53.585 ;
        RECT 33.730 53.295 34.005 54.145 ;
        RECT 33.725 53.125 34.005 53.295 ;
        RECT 33.730 52.985 34.005 53.125 ;
        RECT 34.175 52.785 34.365 54.145 ;
        RECT 34.545 53.780 35.055 54.315 ;
        RECT 35.275 53.505 35.520 54.110 ;
        RECT 35.965 53.575 36.350 54.145 ;
        RECT 36.520 53.855 36.845 54.315 ;
        RECT 37.365 53.685 37.645 54.145 ;
        RECT 34.565 53.335 35.795 53.505 ;
        RECT 33.355 52.615 34.365 52.785 ;
        RECT 34.535 52.770 35.285 52.960 ;
        RECT 33.015 52.275 34.140 52.445 ;
        RECT 34.535 52.105 34.705 52.770 ;
        RECT 35.455 52.525 35.795 53.335 ;
        RECT 32.675 51.935 34.705 52.105 ;
        RECT 34.875 51.765 35.045 52.525 ;
        RECT 35.280 52.115 35.795 52.525 ;
        RECT 35.965 52.905 36.245 53.575 ;
        RECT 36.520 53.515 37.645 53.685 ;
        RECT 36.520 53.405 36.970 53.515 ;
        RECT 36.415 53.075 36.970 53.405 ;
        RECT 37.835 53.345 38.235 54.145 ;
        RECT 38.635 53.855 38.905 54.315 ;
        RECT 39.075 53.685 39.360 54.145 ;
        RECT 35.965 51.935 36.350 52.905 ;
        RECT 36.520 52.615 36.970 53.075 ;
        RECT 37.140 52.785 38.235 53.345 ;
        RECT 36.520 52.395 37.645 52.615 ;
        RECT 36.520 51.765 36.845 52.225 ;
        RECT 37.365 51.935 37.645 52.395 ;
        RECT 37.835 51.935 38.235 52.785 ;
        RECT 38.405 53.515 39.360 53.685 ;
        RECT 38.405 52.615 38.615 53.515 ;
        RECT 38.785 52.785 39.475 53.345 ;
        RECT 39.650 52.715 39.985 54.135 ;
        RECT 40.165 53.945 40.910 54.315 ;
        RECT 41.475 53.775 41.730 54.135 ;
        RECT 41.910 53.945 42.240 54.315 ;
        RECT 42.420 53.775 42.645 54.135 ;
        RECT 40.160 53.585 42.645 53.775 ;
        RECT 40.160 52.895 40.385 53.585 ;
        RECT 42.865 53.545 44.535 54.315 ;
        RECT 44.710 53.575 44.965 54.145 ;
        RECT 45.135 53.915 45.465 54.315 ;
        RECT 45.890 53.780 46.420 54.145 ;
        RECT 45.890 53.745 46.065 53.780 ;
        RECT 45.135 53.575 46.065 53.745 ;
        RECT 40.585 53.075 40.865 53.405 ;
        RECT 41.045 53.075 41.620 53.405 ;
        RECT 41.800 53.075 42.235 53.405 ;
        RECT 42.415 53.075 42.685 53.405 ;
        RECT 42.865 53.025 43.615 53.545 ;
        RECT 40.160 52.715 42.655 52.895 ;
        RECT 43.785 52.855 44.535 53.375 ;
        RECT 38.405 52.395 39.360 52.615 ;
        RECT 38.635 51.765 38.905 52.225 ;
        RECT 39.075 51.935 39.360 52.395 ;
        RECT 39.650 51.945 39.915 52.715 ;
        RECT 40.085 51.765 40.415 52.485 ;
        RECT 40.605 52.305 41.795 52.535 ;
        RECT 40.605 51.945 40.865 52.305 ;
        RECT 41.035 51.765 41.365 52.135 ;
        RECT 41.535 51.945 41.795 52.305 ;
        RECT 42.365 51.945 42.655 52.715 ;
        RECT 42.865 51.765 44.535 52.855 ;
        RECT 44.710 52.905 44.880 53.575 ;
        RECT 45.135 53.405 45.305 53.575 ;
        RECT 45.050 53.075 45.305 53.405 ;
        RECT 45.530 53.075 45.725 53.405 ;
        RECT 44.710 51.935 45.045 52.905 ;
        RECT 45.215 51.765 45.385 52.905 ;
        RECT 45.555 52.105 45.725 53.075 ;
        RECT 45.895 52.445 46.065 53.575 ;
        RECT 46.235 52.785 46.405 53.585 ;
        RECT 46.610 53.295 46.885 54.145 ;
        RECT 46.605 53.125 46.885 53.295 ;
        RECT 46.610 52.985 46.885 53.125 ;
        RECT 47.055 52.785 47.245 54.145 ;
        RECT 47.425 53.780 47.935 54.315 ;
        RECT 48.155 53.505 48.400 54.110 ;
        RECT 48.845 53.575 49.230 54.145 ;
        RECT 49.400 53.855 49.725 54.315 ;
        RECT 50.245 53.685 50.525 54.145 ;
        RECT 47.445 53.335 48.675 53.505 ;
        RECT 46.235 52.615 47.245 52.785 ;
        RECT 47.415 52.770 48.165 52.960 ;
        RECT 45.895 52.275 47.020 52.445 ;
        RECT 47.415 52.105 47.585 52.770 ;
        RECT 48.335 52.525 48.675 53.335 ;
        RECT 45.555 51.935 47.585 52.105 ;
        RECT 47.755 51.765 47.925 52.525 ;
        RECT 48.160 52.115 48.675 52.525 ;
        RECT 48.845 52.905 49.125 53.575 ;
        RECT 49.400 53.515 50.525 53.685 ;
        RECT 49.400 53.405 49.850 53.515 ;
        RECT 49.295 53.075 49.850 53.405 ;
        RECT 50.715 53.345 51.115 54.145 ;
        RECT 51.515 53.855 51.785 54.315 ;
        RECT 51.955 53.685 52.240 54.145 ;
        RECT 48.845 51.935 49.230 52.905 ;
        RECT 49.400 52.615 49.850 53.075 ;
        RECT 50.020 52.785 51.115 53.345 ;
        RECT 49.400 52.395 50.525 52.615 ;
        RECT 49.400 51.765 49.725 52.225 ;
        RECT 50.245 51.935 50.525 52.395 ;
        RECT 50.715 51.935 51.115 52.785 ;
        RECT 51.285 53.515 52.240 53.685 ;
        RECT 52.985 53.575 53.370 54.145 ;
        RECT 53.540 53.855 53.865 54.315 ;
        RECT 54.385 53.685 54.665 54.145 ;
        RECT 51.285 52.615 51.495 53.515 ;
        RECT 51.665 52.785 52.355 53.345 ;
        RECT 52.985 52.905 53.265 53.575 ;
        RECT 53.540 53.515 54.665 53.685 ;
        RECT 53.540 53.405 53.990 53.515 ;
        RECT 53.435 53.075 53.990 53.405 ;
        RECT 54.855 53.345 55.255 54.145 ;
        RECT 55.655 53.855 55.925 54.315 ;
        RECT 56.095 53.685 56.380 54.145 ;
        RECT 51.285 52.395 52.240 52.615 ;
        RECT 51.515 51.765 51.785 52.225 ;
        RECT 51.955 51.935 52.240 52.395 ;
        RECT 52.985 51.935 53.370 52.905 ;
        RECT 53.540 52.615 53.990 53.075 ;
        RECT 54.160 52.785 55.255 53.345 ;
        RECT 53.540 52.395 54.665 52.615 ;
        RECT 53.540 51.765 53.865 52.225 ;
        RECT 54.385 51.935 54.665 52.395 ;
        RECT 54.855 51.935 55.255 52.785 ;
        RECT 55.425 53.515 56.380 53.685 ;
        RECT 57.125 53.590 57.415 54.315 ;
        RECT 57.700 53.685 57.985 54.145 ;
        RECT 58.155 53.855 58.425 54.315 ;
        RECT 57.700 53.515 58.655 53.685 ;
        RECT 55.425 52.615 55.635 53.515 ;
        RECT 55.805 52.785 56.495 53.345 ;
        RECT 55.425 52.395 56.380 52.615 ;
        RECT 55.655 51.765 55.925 52.225 ;
        RECT 56.095 51.935 56.380 52.395 ;
        RECT 57.125 51.765 57.415 52.930 ;
        RECT 57.585 52.785 58.275 53.345 ;
        RECT 58.445 52.615 58.655 53.515 ;
        RECT 57.700 52.395 58.655 52.615 ;
        RECT 58.825 53.345 59.225 54.145 ;
        RECT 59.415 53.685 59.695 54.145 ;
        RECT 60.215 53.855 60.540 54.315 ;
        RECT 59.415 53.515 60.540 53.685 ;
        RECT 60.710 53.575 61.095 54.145 ;
        RECT 61.275 53.805 62.505 54.145 ;
        RECT 62.675 53.825 62.930 54.315 ;
        RECT 61.275 53.575 61.605 53.805 ;
        RECT 60.090 53.405 60.540 53.515 ;
        RECT 58.825 52.785 59.920 53.345 ;
        RECT 60.090 53.075 60.645 53.405 ;
        RECT 57.700 51.935 57.985 52.395 ;
        RECT 58.155 51.765 58.425 52.225 ;
        RECT 58.825 51.935 59.225 52.785 ;
        RECT 60.090 52.615 60.540 53.075 ;
        RECT 60.815 52.905 61.095 53.575 ;
        RECT 61.265 53.075 61.575 53.405 ;
        RECT 61.780 53.075 62.155 53.635 ;
        RECT 62.325 52.905 62.505 53.805 ;
        RECT 62.690 53.075 62.910 53.655 ;
        RECT 63.195 53.635 63.365 54.010 ;
        RECT 63.165 53.465 63.365 53.635 ;
        RECT 63.555 53.785 63.785 54.090 ;
        RECT 63.955 53.955 64.285 54.315 ;
        RECT 64.480 53.785 64.770 54.135 ;
        RECT 65.905 53.805 66.305 54.315 ;
        RECT 63.555 53.615 64.770 53.785 ;
        RECT 66.880 53.700 67.050 54.145 ;
        RECT 67.220 53.915 67.940 54.315 ;
        RECT 68.110 53.745 68.280 54.145 ;
        RECT 68.515 53.870 68.945 54.315 ;
        RECT 63.195 53.445 63.365 53.465 ;
        RECT 63.195 53.275 63.715 53.445 ;
        RECT 59.415 52.395 60.540 52.615 ;
        RECT 59.415 51.935 59.695 52.395 ;
        RECT 60.215 51.765 60.540 52.225 ;
        RECT 60.710 51.935 61.095 52.905 ;
        RECT 61.275 52.735 62.505 52.905 ;
        RECT 61.275 51.935 61.605 52.735 ;
        RECT 61.775 51.765 62.005 52.565 ;
        RECT 62.175 51.935 62.505 52.735 ;
        RECT 62.675 51.765 62.930 52.905 ;
        RECT 63.110 52.745 63.355 53.105 ;
        RECT 63.545 52.895 63.715 53.275 ;
        RECT 63.885 53.075 64.270 53.405 ;
        RECT 64.450 53.295 64.710 53.405 ;
        RECT 64.450 53.125 64.715 53.295 ;
        RECT 64.450 53.075 64.710 53.125 ;
        RECT 63.545 52.615 63.895 52.895 ;
        RECT 63.110 51.765 63.365 52.565 ;
        RECT 63.565 51.935 63.895 52.615 ;
        RECT 64.075 52.025 64.270 53.075 ;
        RECT 64.450 51.765 64.770 52.905 ;
        RECT 65.920 52.745 66.180 53.635 ;
        RECT 66.380 53.045 66.640 53.635 ;
        RECT 66.880 53.530 67.230 53.700 ;
        RECT 66.380 52.745 66.860 53.045 ;
        RECT 65.945 52.395 66.885 52.565 ;
        RECT 65.945 51.935 66.125 52.395 ;
        RECT 66.295 51.765 66.545 52.225 ;
        RECT 66.715 52.145 66.885 52.395 ;
        RECT 67.060 52.505 67.230 53.530 ;
        RECT 67.400 53.575 68.280 53.745 ;
        RECT 69.115 53.590 69.375 54.145 ;
        RECT 67.400 52.855 67.570 53.575 ;
        RECT 67.760 53.025 68.050 53.405 ;
        RECT 67.400 52.685 67.920 52.855 ;
        RECT 68.220 52.785 68.550 53.405 ;
        RECT 68.775 53.075 69.030 53.405 ;
        RECT 67.060 52.335 67.470 52.505 ;
        RECT 67.750 52.495 67.920 52.685 ;
        RECT 68.775 52.595 68.945 53.075 ;
        RECT 69.200 52.875 69.375 53.590 ;
        RECT 69.565 53.585 69.895 54.315 ;
        RECT 70.065 53.405 70.275 54.025 ;
        RECT 70.455 53.605 70.885 54.135 ;
        RECT 69.580 53.055 69.870 53.405 ;
        RECT 70.065 53.055 70.460 53.405 ;
        RECT 70.640 53.355 70.885 53.605 ;
        RECT 71.065 53.535 71.295 54.315 ;
        RECT 71.475 53.685 71.855 54.135 ;
        RECT 72.855 53.765 73.025 54.055 ;
        RECT 73.195 53.935 73.525 54.315 ;
        RECT 70.640 53.055 71.175 53.355 ;
        RECT 71.475 53.235 71.705 53.685 ;
        RECT 72.855 53.595 73.520 53.765 ;
        RECT 67.215 52.200 67.470 52.335 ;
        RECT 68.185 52.425 68.945 52.595 ;
        RECT 68.185 52.200 68.355 52.425 ;
        RECT 66.715 51.975 67.045 52.145 ;
        RECT 67.215 52.030 68.355 52.200 ;
        RECT 67.215 51.935 67.470 52.030 ;
        RECT 68.615 51.765 68.945 52.165 ;
        RECT 69.115 51.935 69.375 52.875 ;
        RECT 69.635 52.675 70.675 52.875 ;
        RECT 69.635 51.945 69.805 52.675 ;
        RECT 69.985 51.765 70.315 52.495 ;
        RECT 70.485 51.945 70.675 52.675 ;
        RECT 70.845 51.945 71.175 53.055 ;
        RECT 71.365 52.555 71.705 53.235 ;
        RECT 71.885 52.735 72.115 53.425 ;
        RECT 72.770 52.775 73.120 53.425 ;
        RECT 73.290 52.605 73.520 53.595 ;
        RECT 71.365 52.355 72.125 52.555 ;
        RECT 71.365 51.765 71.695 52.175 ;
        RECT 71.865 51.965 72.125 52.355 ;
        RECT 72.855 52.435 73.520 52.605 ;
        RECT 72.855 51.935 73.025 52.435 ;
        RECT 73.195 51.765 73.525 52.265 ;
        RECT 73.695 51.935 73.880 54.055 ;
        RECT 74.135 53.855 74.385 54.315 ;
        RECT 74.555 53.865 74.890 54.035 ;
        RECT 75.085 53.865 75.760 54.035 ;
        RECT 74.555 53.725 74.725 53.865 ;
        RECT 74.050 52.735 74.330 53.685 ;
        RECT 74.500 53.595 74.725 53.725 ;
        RECT 74.500 52.490 74.670 53.595 ;
        RECT 74.895 53.445 75.420 53.665 ;
        RECT 74.840 52.680 75.080 53.275 ;
        RECT 75.250 52.745 75.420 53.445 ;
        RECT 75.590 53.085 75.760 53.865 ;
        RECT 76.080 53.815 76.450 54.315 ;
        RECT 76.630 53.865 77.035 54.035 ;
        RECT 77.205 53.865 77.990 54.035 ;
        RECT 76.630 53.635 76.800 53.865 ;
        RECT 75.970 53.335 76.800 53.635 ;
        RECT 77.185 53.365 77.650 53.695 ;
        RECT 75.970 53.305 76.170 53.335 ;
        RECT 76.290 53.085 76.460 53.155 ;
        RECT 75.590 52.915 76.460 53.085 ;
        RECT 75.950 52.825 76.460 52.915 ;
        RECT 74.500 52.360 74.805 52.490 ;
        RECT 75.250 52.380 75.780 52.745 ;
        RECT 74.120 51.765 74.385 52.225 ;
        RECT 74.555 51.935 74.805 52.360 ;
        RECT 75.950 52.210 76.120 52.825 ;
        RECT 75.015 52.040 76.120 52.210 ;
        RECT 76.290 51.765 76.460 52.565 ;
        RECT 76.630 52.265 76.800 53.335 ;
        RECT 76.970 52.435 77.160 53.155 ;
        RECT 77.330 52.405 77.650 53.365 ;
        RECT 77.820 53.405 77.990 53.865 ;
        RECT 78.265 53.785 78.475 54.315 ;
        RECT 78.735 53.575 79.065 54.100 ;
        RECT 79.235 53.705 79.405 54.315 ;
        RECT 79.575 53.660 79.905 54.095 ;
        RECT 81.135 53.765 81.305 54.145 ;
        RECT 81.520 53.935 81.850 54.315 ;
        RECT 79.575 53.575 79.955 53.660 ;
        RECT 81.135 53.595 81.850 53.765 ;
        RECT 78.865 53.405 79.065 53.575 ;
        RECT 79.730 53.535 79.955 53.575 ;
        RECT 77.820 53.075 78.695 53.405 ;
        RECT 78.865 53.075 79.615 53.405 ;
        RECT 76.630 51.935 76.880 52.265 ;
        RECT 77.820 52.235 77.990 53.075 ;
        RECT 78.865 52.870 79.055 53.075 ;
        RECT 79.785 52.955 79.955 53.535 ;
        RECT 81.045 53.045 81.400 53.415 ;
        RECT 81.680 53.405 81.850 53.595 ;
        RECT 82.020 53.570 82.275 54.145 ;
        RECT 81.680 53.075 81.935 53.405 ;
        RECT 79.740 52.905 79.955 52.955 ;
        RECT 78.160 52.495 79.055 52.870 ;
        RECT 79.565 52.825 79.955 52.905 ;
        RECT 81.680 52.865 81.850 53.075 ;
        RECT 77.105 52.065 77.990 52.235 ;
        RECT 78.170 51.765 78.485 52.265 ;
        RECT 78.715 51.935 79.055 52.495 ;
        RECT 79.225 51.765 79.395 52.775 ;
        RECT 79.565 51.980 79.895 52.825 ;
        RECT 81.135 52.695 81.850 52.865 ;
        RECT 82.105 52.840 82.275 53.570 ;
        RECT 82.450 53.475 82.710 54.315 ;
        RECT 82.885 53.565 84.095 54.315 ;
        RECT 81.135 51.935 81.305 52.695 ;
        RECT 81.520 51.765 81.850 52.525 ;
        RECT 82.020 51.935 82.275 52.840 ;
        RECT 82.450 51.765 82.710 52.915 ;
        RECT 82.885 52.855 83.405 53.395 ;
        RECT 83.575 53.025 84.095 53.565 ;
        RECT 82.885 51.765 84.095 52.855 ;
        RECT 5.520 51.595 84.180 51.765 ;
        RECT 5.605 50.505 6.815 51.595 ;
        RECT 5.605 49.795 6.125 50.335 ;
        RECT 6.295 49.965 6.815 50.505 ;
        RECT 7.170 50.625 7.560 50.800 ;
        RECT 8.045 50.795 8.375 51.595 ;
        RECT 8.545 50.805 9.080 51.425 ;
        RECT 7.170 50.455 8.595 50.625 ;
        RECT 5.605 49.045 6.815 49.795 ;
        RECT 7.045 49.725 7.400 50.285 ;
        RECT 7.570 49.555 7.740 50.455 ;
        RECT 7.910 49.725 8.175 50.285 ;
        RECT 8.425 49.955 8.595 50.455 ;
        RECT 8.765 49.785 9.080 50.805 ;
        RECT 9.375 50.925 9.545 51.425 ;
        RECT 9.715 51.095 10.045 51.595 ;
        RECT 9.375 50.755 10.040 50.925 ;
        RECT 9.290 49.935 9.640 50.585 ;
        RECT 7.150 49.045 7.390 49.555 ;
        RECT 7.570 49.225 7.850 49.555 ;
        RECT 8.080 49.045 8.295 49.555 ;
        RECT 8.465 49.215 9.080 49.785 ;
        RECT 9.810 49.765 10.040 50.755 ;
        RECT 9.375 49.595 10.040 49.765 ;
        RECT 9.375 49.305 9.545 49.595 ;
        RECT 9.715 49.045 10.045 49.425 ;
        RECT 10.215 49.305 10.400 51.425 ;
        RECT 10.640 51.135 10.905 51.595 ;
        RECT 11.075 51.000 11.325 51.425 ;
        RECT 11.535 51.150 12.640 51.320 ;
        RECT 11.020 50.870 11.325 51.000 ;
        RECT 10.570 49.675 10.850 50.625 ;
        RECT 11.020 49.765 11.190 50.870 ;
        RECT 11.360 50.085 11.600 50.680 ;
        RECT 11.770 50.615 12.300 50.980 ;
        RECT 11.770 49.915 11.940 50.615 ;
        RECT 12.470 50.535 12.640 51.150 ;
        RECT 12.810 50.795 12.980 51.595 ;
        RECT 13.150 51.095 13.400 51.425 ;
        RECT 13.625 51.125 14.510 51.295 ;
        RECT 12.470 50.445 12.980 50.535 ;
        RECT 11.020 49.635 11.245 49.765 ;
        RECT 11.415 49.695 11.940 49.915 ;
        RECT 12.110 50.275 12.980 50.445 ;
        RECT 10.655 49.045 10.905 49.505 ;
        RECT 11.075 49.495 11.245 49.635 ;
        RECT 12.110 49.495 12.280 50.275 ;
        RECT 12.810 50.205 12.980 50.275 ;
        RECT 12.490 50.025 12.690 50.055 ;
        RECT 13.150 50.025 13.320 51.095 ;
        RECT 13.490 50.205 13.680 50.925 ;
        RECT 12.490 49.725 13.320 50.025 ;
        RECT 13.850 49.995 14.170 50.955 ;
        RECT 11.075 49.325 11.410 49.495 ;
        RECT 11.605 49.325 12.280 49.495 ;
        RECT 12.600 49.045 12.970 49.545 ;
        RECT 13.150 49.495 13.320 49.725 ;
        RECT 13.705 49.665 14.170 49.995 ;
        RECT 14.340 50.285 14.510 51.125 ;
        RECT 14.690 51.095 15.005 51.595 ;
        RECT 15.235 50.865 15.575 51.425 ;
        RECT 14.680 50.490 15.575 50.865 ;
        RECT 15.745 50.585 15.915 51.595 ;
        RECT 15.385 50.285 15.575 50.490 ;
        RECT 16.085 50.535 16.415 51.380 ;
        RECT 16.085 50.455 16.475 50.535 ;
        RECT 16.645 50.505 18.315 51.595 ;
        RECT 16.260 50.405 16.475 50.455 ;
        RECT 14.340 49.955 15.215 50.285 ;
        RECT 15.385 49.955 16.135 50.285 ;
        RECT 14.340 49.495 14.510 49.955 ;
        RECT 15.385 49.785 15.585 49.955 ;
        RECT 16.305 49.825 16.475 50.405 ;
        RECT 16.250 49.785 16.475 49.825 ;
        RECT 13.150 49.325 13.555 49.495 ;
        RECT 13.725 49.325 14.510 49.495 ;
        RECT 14.785 49.045 14.995 49.575 ;
        RECT 15.255 49.260 15.585 49.785 ;
        RECT 16.095 49.700 16.475 49.785 ;
        RECT 16.645 49.815 17.395 50.335 ;
        RECT 17.565 49.985 18.315 50.505 ;
        RECT 18.485 50.430 18.775 51.595 ;
        RECT 18.955 50.485 19.250 51.595 ;
        RECT 19.430 50.285 19.680 51.420 ;
        RECT 19.850 50.485 20.110 51.595 ;
        RECT 20.280 50.695 20.540 51.420 ;
        RECT 20.710 50.865 20.970 51.595 ;
        RECT 21.140 50.695 21.400 51.420 ;
        RECT 21.570 50.865 21.830 51.595 ;
        RECT 22.000 50.695 22.260 51.420 ;
        RECT 22.430 50.865 22.690 51.595 ;
        RECT 22.860 50.695 23.120 51.420 ;
        RECT 23.290 50.865 23.585 51.595 ;
        RECT 20.280 50.455 23.590 50.695 ;
        RECT 24.045 50.645 24.335 51.415 ;
        RECT 24.905 51.055 25.165 51.415 ;
        RECT 25.335 51.225 25.665 51.595 ;
        RECT 25.835 51.055 26.095 51.415 ;
        RECT 24.905 50.825 26.095 51.055 ;
        RECT 26.285 50.875 26.615 51.595 ;
        RECT 26.785 50.645 27.050 51.415 ;
        RECT 27.225 51.160 32.570 51.595 ;
        RECT 32.745 51.160 38.090 51.595 ;
        RECT 24.045 50.465 26.540 50.645 ;
        RECT 15.755 49.045 15.925 49.655 ;
        RECT 16.095 49.265 16.425 49.700 ;
        RECT 16.645 49.045 18.315 49.815 ;
        RECT 18.485 49.045 18.775 49.770 ;
        RECT 18.945 49.675 19.260 50.285 ;
        RECT 19.430 50.035 22.450 50.285 ;
        RECT 19.005 49.045 19.250 49.505 ;
        RECT 19.430 49.225 19.680 50.035 ;
        RECT 22.620 49.865 23.590 50.455 ;
        RECT 24.015 49.955 24.285 50.285 ;
        RECT 24.465 49.955 24.900 50.285 ;
        RECT 25.080 49.955 25.655 50.285 ;
        RECT 25.835 49.955 26.115 50.285 ;
        RECT 20.280 49.695 23.590 49.865 ;
        RECT 26.315 49.775 26.540 50.465 ;
        RECT 19.850 49.045 20.110 49.570 ;
        RECT 20.280 49.240 20.540 49.695 ;
        RECT 20.710 49.045 20.970 49.525 ;
        RECT 21.140 49.240 21.400 49.695 ;
        RECT 21.570 49.045 21.830 49.525 ;
        RECT 22.000 49.240 22.260 49.695 ;
        RECT 22.430 49.045 22.690 49.525 ;
        RECT 22.860 49.240 23.120 49.695 ;
        RECT 24.055 49.585 26.540 49.775 ;
        RECT 23.290 49.045 23.590 49.525 ;
        RECT 24.055 49.225 24.280 49.585 ;
        RECT 24.460 49.045 24.790 49.415 ;
        RECT 24.970 49.225 25.225 49.585 ;
        RECT 25.790 49.045 26.535 49.415 ;
        RECT 26.715 49.225 27.050 50.645 ;
        RECT 28.810 49.590 29.150 50.420 ;
        RECT 30.630 49.910 30.980 51.160 ;
        RECT 34.330 49.590 34.670 50.420 ;
        RECT 36.150 49.910 36.500 51.160 ;
        RECT 38.265 50.505 40.855 51.595 ;
        RECT 38.265 49.815 39.475 50.335 ;
        RECT 39.645 49.985 40.855 50.505 ;
        RECT 41.030 50.645 41.295 51.415 ;
        RECT 41.465 50.875 41.795 51.595 ;
        RECT 41.985 51.055 42.245 51.415 ;
        RECT 42.415 51.225 42.745 51.595 ;
        RECT 42.915 51.055 43.175 51.415 ;
        RECT 41.985 50.825 43.175 51.055 ;
        RECT 43.745 50.645 44.035 51.415 ;
        RECT 27.225 49.045 32.570 49.590 ;
        RECT 32.745 49.045 38.090 49.590 ;
        RECT 38.265 49.045 40.855 49.815 ;
        RECT 41.030 49.225 41.365 50.645 ;
        RECT 41.540 50.465 44.035 50.645 ;
        RECT 41.540 49.775 41.765 50.465 ;
        RECT 44.245 50.430 44.535 51.595 ;
        RECT 45.715 50.925 45.885 51.425 ;
        RECT 46.055 51.095 46.385 51.595 ;
        RECT 45.715 50.755 46.380 50.925 ;
        RECT 41.965 49.955 42.245 50.285 ;
        RECT 42.425 49.955 43.000 50.285 ;
        RECT 43.180 49.955 43.615 50.285 ;
        RECT 43.795 49.955 44.065 50.285 ;
        RECT 45.630 49.935 45.980 50.585 ;
        RECT 41.540 49.585 44.025 49.775 ;
        RECT 41.545 49.045 42.290 49.415 ;
        RECT 42.855 49.225 43.110 49.585 ;
        RECT 43.290 49.045 43.620 49.415 ;
        RECT 43.800 49.225 44.025 49.585 ;
        RECT 44.245 49.045 44.535 49.770 ;
        RECT 46.150 49.765 46.380 50.755 ;
        RECT 45.715 49.595 46.380 49.765 ;
        RECT 45.715 49.305 45.885 49.595 ;
        RECT 46.055 49.045 46.385 49.425 ;
        RECT 46.555 49.305 46.740 51.425 ;
        RECT 46.980 51.135 47.245 51.595 ;
        RECT 47.415 51.000 47.665 51.425 ;
        RECT 47.875 51.150 48.980 51.320 ;
        RECT 47.360 50.870 47.665 51.000 ;
        RECT 46.910 49.675 47.190 50.625 ;
        RECT 47.360 49.765 47.530 50.870 ;
        RECT 47.700 50.085 47.940 50.680 ;
        RECT 48.110 50.615 48.640 50.980 ;
        RECT 48.110 49.915 48.280 50.615 ;
        RECT 48.810 50.535 48.980 51.150 ;
        RECT 49.150 50.795 49.320 51.595 ;
        RECT 49.490 51.095 49.740 51.425 ;
        RECT 49.965 51.125 50.850 51.295 ;
        RECT 48.810 50.445 49.320 50.535 ;
        RECT 47.360 49.635 47.585 49.765 ;
        RECT 47.755 49.695 48.280 49.915 ;
        RECT 48.450 50.275 49.320 50.445 ;
        RECT 46.995 49.045 47.245 49.505 ;
        RECT 47.415 49.495 47.585 49.635 ;
        RECT 48.450 49.495 48.620 50.275 ;
        RECT 49.150 50.205 49.320 50.275 ;
        RECT 48.830 50.025 49.030 50.055 ;
        RECT 49.490 50.025 49.660 51.095 ;
        RECT 49.830 50.205 50.020 50.925 ;
        RECT 48.830 49.725 49.660 50.025 ;
        RECT 50.190 49.995 50.510 50.955 ;
        RECT 47.415 49.325 47.750 49.495 ;
        RECT 47.945 49.325 48.620 49.495 ;
        RECT 48.940 49.045 49.310 49.545 ;
        RECT 49.490 49.495 49.660 49.725 ;
        RECT 50.045 49.665 50.510 49.995 ;
        RECT 50.680 50.285 50.850 51.125 ;
        RECT 51.030 51.095 51.345 51.595 ;
        RECT 51.575 50.865 51.915 51.425 ;
        RECT 51.020 50.490 51.915 50.865 ;
        RECT 52.085 50.585 52.255 51.595 ;
        RECT 51.725 50.285 51.915 50.490 ;
        RECT 52.425 50.535 52.755 51.380 ;
        RECT 53.045 50.535 53.375 51.380 ;
        RECT 53.545 50.585 53.715 51.595 ;
        RECT 53.885 50.865 54.225 51.425 ;
        RECT 54.455 51.095 54.770 51.595 ;
        RECT 54.950 51.125 55.835 51.295 ;
        RECT 52.425 50.455 52.815 50.535 ;
        RECT 52.600 50.405 52.815 50.455 ;
        RECT 50.680 49.955 51.555 50.285 ;
        RECT 51.725 49.955 52.475 50.285 ;
        RECT 50.680 49.495 50.850 49.955 ;
        RECT 51.725 49.785 51.925 49.955 ;
        RECT 52.645 49.825 52.815 50.405 ;
        RECT 52.590 49.785 52.815 49.825 ;
        RECT 49.490 49.325 49.895 49.495 ;
        RECT 50.065 49.325 50.850 49.495 ;
        RECT 51.125 49.045 51.335 49.575 ;
        RECT 51.595 49.260 51.925 49.785 ;
        RECT 52.435 49.700 52.815 49.785 ;
        RECT 52.985 50.455 53.375 50.535 ;
        RECT 53.885 50.490 54.780 50.865 ;
        RECT 52.985 50.405 53.200 50.455 ;
        RECT 52.985 49.825 53.155 50.405 ;
        RECT 53.885 50.285 54.075 50.490 ;
        RECT 54.950 50.285 55.120 51.125 ;
        RECT 56.060 51.095 56.310 51.425 ;
        RECT 53.325 49.955 54.075 50.285 ;
        RECT 54.245 49.955 55.120 50.285 ;
        RECT 52.985 49.785 53.210 49.825 ;
        RECT 53.875 49.785 54.075 49.955 ;
        RECT 52.985 49.700 53.365 49.785 ;
        RECT 52.095 49.045 52.265 49.655 ;
        RECT 52.435 49.265 52.765 49.700 ;
        RECT 53.035 49.265 53.365 49.700 ;
        RECT 53.535 49.045 53.705 49.655 ;
        RECT 53.875 49.260 54.205 49.785 ;
        RECT 54.465 49.045 54.675 49.575 ;
        RECT 54.950 49.495 55.120 49.955 ;
        RECT 55.290 49.995 55.610 50.955 ;
        RECT 55.780 50.205 55.970 50.925 ;
        RECT 56.140 50.025 56.310 51.095 ;
        RECT 56.480 50.795 56.650 51.595 ;
        RECT 56.820 51.150 57.925 51.320 ;
        RECT 56.820 50.535 56.990 51.150 ;
        RECT 58.135 51.000 58.385 51.425 ;
        RECT 58.555 51.135 58.820 51.595 ;
        RECT 57.160 50.615 57.690 50.980 ;
        RECT 58.135 50.870 58.440 51.000 ;
        RECT 56.480 50.445 56.990 50.535 ;
        RECT 56.480 50.275 57.350 50.445 ;
        RECT 56.480 50.205 56.650 50.275 ;
        RECT 56.770 50.025 56.970 50.055 ;
        RECT 55.290 49.665 55.755 49.995 ;
        RECT 56.140 49.725 56.970 50.025 ;
        RECT 56.140 49.495 56.310 49.725 ;
        RECT 54.950 49.325 55.735 49.495 ;
        RECT 55.905 49.325 56.310 49.495 ;
        RECT 56.490 49.045 56.860 49.545 ;
        RECT 57.180 49.495 57.350 50.275 ;
        RECT 57.520 49.915 57.690 50.615 ;
        RECT 57.860 50.085 58.100 50.680 ;
        RECT 57.520 49.695 58.045 49.915 ;
        RECT 58.270 49.765 58.440 50.870 ;
        RECT 58.215 49.635 58.440 49.765 ;
        RECT 58.610 49.675 58.890 50.625 ;
        RECT 58.215 49.495 58.385 49.635 ;
        RECT 57.180 49.325 57.855 49.495 ;
        RECT 58.050 49.325 58.385 49.495 ;
        RECT 58.555 49.045 58.805 49.505 ;
        RECT 59.060 49.305 59.245 51.425 ;
        RECT 59.415 51.095 59.745 51.595 ;
        RECT 59.915 50.925 60.085 51.425 ;
        RECT 59.420 50.755 60.085 50.925 ;
        RECT 59.420 49.765 59.650 50.755 ;
        RECT 59.820 49.935 60.170 50.585 ;
        RECT 60.405 50.535 60.735 51.380 ;
        RECT 60.905 50.585 61.075 51.595 ;
        RECT 61.245 50.865 61.585 51.425 ;
        RECT 61.815 51.095 62.130 51.595 ;
        RECT 62.310 51.125 63.195 51.295 ;
        RECT 60.345 50.455 60.735 50.535 ;
        RECT 61.245 50.490 62.140 50.865 ;
        RECT 60.345 50.405 60.560 50.455 ;
        RECT 60.345 49.825 60.515 50.405 ;
        RECT 61.245 50.285 61.435 50.490 ;
        RECT 62.310 50.285 62.480 51.125 ;
        RECT 63.420 51.095 63.670 51.425 ;
        RECT 60.685 49.955 61.435 50.285 ;
        RECT 61.605 49.955 62.480 50.285 ;
        RECT 60.345 49.785 60.570 49.825 ;
        RECT 61.235 49.785 61.435 49.955 ;
        RECT 59.420 49.595 60.085 49.765 ;
        RECT 60.345 49.700 60.725 49.785 ;
        RECT 59.415 49.045 59.745 49.425 ;
        RECT 59.915 49.305 60.085 49.595 ;
        RECT 60.395 49.265 60.725 49.700 ;
        RECT 60.895 49.045 61.065 49.655 ;
        RECT 61.235 49.260 61.565 49.785 ;
        RECT 61.825 49.045 62.035 49.575 ;
        RECT 62.310 49.495 62.480 49.955 ;
        RECT 62.650 49.995 62.970 50.955 ;
        RECT 63.140 50.205 63.330 50.925 ;
        RECT 63.500 50.025 63.670 51.095 ;
        RECT 63.840 50.795 64.010 51.595 ;
        RECT 64.180 51.150 65.285 51.320 ;
        RECT 64.180 50.535 64.350 51.150 ;
        RECT 65.495 51.000 65.745 51.425 ;
        RECT 65.915 51.135 66.180 51.595 ;
        RECT 64.520 50.615 65.050 50.980 ;
        RECT 65.495 50.870 65.800 51.000 ;
        RECT 63.840 50.445 64.350 50.535 ;
        RECT 63.840 50.275 64.710 50.445 ;
        RECT 63.840 50.205 64.010 50.275 ;
        RECT 64.130 50.025 64.330 50.055 ;
        RECT 62.650 49.665 63.115 49.995 ;
        RECT 63.500 49.725 64.330 50.025 ;
        RECT 63.500 49.495 63.670 49.725 ;
        RECT 62.310 49.325 63.095 49.495 ;
        RECT 63.265 49.325 63.670 49.495 ;
        RECT 63.850 49.045 64.220 49.545 ;
        RECT 64.540 49.495 64.710 50.275 ;
        RECT 64.880 49.915 65.050 50.615 ;
        RECT 65.220 50.085 65.460 50.680 ;
        RECT 64.880 49.695 65.405 49.915 ;
        RECT 65.630 49.765 65.800 50.870 ;
        RECT 65.575 49.635 65.800 49.765 ;
        RECT 65.970 49.675 66.250 50.625 ;
        RECT 65.575 49.495 65.745 49.635 ;
        RECT 64.540 49.325 65.215 49.495 ;
        RECT 65.410 49.325 65.745 49.495 ;
        RECT 65.915 49.045 66.165 49.505 ;
        RECT 66.420 49.305 66.605 51.425 ;
        RECT 66.775 51.095 67.105 51.595 ;
        RECT 67.275 50.925 67.445 51.425 ;
        RECT 66.780 50.755 67.445 50.925 ;
        RECT 66.780 49.765 67.010 50.755 ;
        RECT 67.180 49.935 67.530 50.585 ;
        RECT 67.705 50.455 67.985 51.595 ;
        RECT 68.155 50.445 68.485 51.425 ;
        RECT 68.655 50.455 68.915 51.595 ;
        RECT 67.715 50.015 68.050 50.285 ;
        RECT 68.220 49.845 68.390 50.445 ;
        RECT 70.005 50.430 70.295 51.595 ;
        RECT 70.465 50.455 70.850 51.425 ;
        RECT 71.020 51.135 71.345 51.595 ;
        RECT 71.865 50.965 72.145 51.425 ;
        RECT 71.020 50.745 72.145 50.965 ;
        RECT 68.560 50.035 68.895 50.285 ;
        RECT 66.780 49.595 67.445 49.765 ;
        RECT 66.775 49.045 67.105 49.425 ;
        RECT 67.275 49.305 67.445 49.595 ;
        RECT 67.705 49.045 68.015 49.845 ;
        RECT 68.220 49.215 68.915 49.845 ;
        RECT 70.465 49.785 70.745 50.455 ;
        RECT 71.020 50.285 71.470 50.745 ;
        RECT 72.335 50.575 72.735 51.425 ;
        RECT 73.135 51.135 73.405 51.595 ;
        RECT 73.575 50.965 73.860 51.425 ;
        RECT 70.915 49.955 71.470 50.285 ;
        RECT 71.640 50.015 72.735 50.575 ;
        RECT 71.020 49.845 71.470 49.955 ;
        RECT 70.005 49.045 70.295 49.770 ;
        RECT 70.465 49.215 70.850 49.785 ;
        RECT 71.020 49.675 72.145 49.845 ;
        RECT 71.020 49.045 71.345 49.505 ;
        RECT 71.865 49.215 72.145 49.675 ;
        RECT 72.335 49.215 72.735 50.015 ;
        RECT 72.905 50.745 73.860 50.965 ;
        RECT 72.905 49.845 73.115 50.745 ;
        RECT 73.285 50.015 73.975 50.575 ;
        RECT 74.610 50.455 74.945 51.425 ;
        RECT 75.115 50.455 75.285 51.595 ;
        RECT 75.455 51.255 77.485 51.425 ;
        RECT 72.905 49.675 73.860 49.845 ;
        RECT 73.135 49.045 73.405 49.505 ;
        RECT 73.575 49.215 73.860 49.675 ;
        RECT 74.610 49.785 74.780 50.455 ;
        RECT 75.455 50.285 75.625 51.255 ;
        RECT 74.950 49.955 75.205 50.285 ;
        RECT 75.430 49.955 75.625 50.285 ;
        RECT 75.795 50.915 76.920 51.085 ;
        RECT 75.035 49.785 75.205 49.955 ;
        RECT 75.795 49.785 75.965 50.915 ;
        RECT 74.610 49.215 74.865 49.785 ;
        RECT 75.035 49.615 75.965 49.785 ;
        RECT 76.135 50.575 77.145 50.745 ;
        RECT 76.135 49.775 76.305 50.575 ;
        RECT 75.790 49.580 75.965 49.615 ;
        RECT 75.035 49.045 75.365 49.445 ;
        RECT 75.790 49.215 76.320 49.580 ;
        RECT 76.510 49.555 76.785 50.375 ;
        RECT 76.505 49.385 76.785 49.555 ;
        RECT 76.510 49.215 76.785 49.385 ;
        RECT 76.955 49.215 77.145 50.575 ;
        RECT 77.315 50.590 77.485 51.255 ;
        RECT 77.655 50.835 77.825 51.595 ;
        RECT 78.060 50.835 78.575 51.245 ;
        RECT 77.315 50.400 78.065 50.590 ;
        RECT 78.235 50.025 78.575 50.835 ;
        RECT 77.345 49.855 78.575 50.025 ;
        RECT 78.745 50.455 79.130 51.425 ;
        RECT 79.300 51.135 79.625 51.595 ;
        RECT 80.145 50.965 80.425 51.425 ;
        RECT 79.300 50.745 80.425 50.965 ;
        RECT 77.325 49.045 77.835 49.580 ;
        RECT 78.055 49.250 78.300 49.855 ;
        RECT 78.745 49.785 79.025 50.455 ;
        RECT 79.300 50.285 79.750 50.745 ;
        RECT 80.615 50.575 81.015 51.425 ;
        RECT 81.415 51.135 81.685 51.595 ;
        RECT 81.855 50.965 82.140 51.425 ;
        RECT 79.195 49.955 79.750 50.285 ;
        RECT 79.920 50.015 81.015 50.575 ;
        RECT 79.300 49.845 79.750 49.955 ;
        RECT 78.745 49.215 79.130 49.785 ;
        RECT 79.300 49.675 80.425 49.845 ;
        RECT 79.300 49.045 79.625 49.505 ;
        RECT 80.145 49.215 80.425 49.675 ;
        RECT 80.615 49.215 81.015 50.015 ;
        RECT 81.185 50.745 82.140 50.965 ;
        RECT 81.185 49.845 81.395 50.745 ;
        RECT 81.565 50.015 82.255 50.575 ;
        RECT 82.885 50.505 84.095 51.595 ;
        RECT 82.885 49.965 83.405 50.505 ;
        RECT 81.185 49.675 82.140 49.845 ;
        RECT 83.575 49.795 84.095 50.335 ;
        RECT 81.415 49.045 81.685 49.505 ;
        RECT 81.855 49.215 82.140 49.675 ;
        RECT 82.885 49.045 84.095 49.795 ;
        RECT 5.520 48.875 84.180 49.045 ;
        RECT 5.605 48.125 6.815 48.875 ;
        RECT 5.605 47.585 6.125 48.125 ;
        RECT 6.990 48.035 7.250 48.875 ;
        RECT 7.425 48.130 7.680 48.705 ;
        RECT 7.850 48.495 8.180 48.875 ;
        RECT 8.395 48.325 8.565 48.705 ;
        RECT 7.850 48.155 8.565 48.325 ;
        RECT 6.295 47.415 6.815 47.955 ;
        RECT 5.605 46.325 6.815 47.415 ;
        RECT 6.990 46.325 7.250 47.475 ;
        RECT 7.425 47.400 7.595 48.130 ;
        RECT 7.850 47.965 8.020 48.155 ;
        RECT 8.830 48.035 9.090 48.875 ;
        RECT 9.265 48.130 9.520 48.705 ;
        RECT 9.690 48.495 10.020 48.875 ;
        RECT 10.235 48.325 10.405 48.705 ;
        RECT 10.665 48.330 16.010 48.875 ;
        RECT 16.810 48.365 17.050 48.875 ;
        RECT 17.230 48.365 17.510 48.695 ;
        RECT 17.740 48.365 17.955 48.875 ;
        RECT 9.690 48.155 10.405 48.325 ;
        RECT 7.765 47.635 8.020 47.965 ;
        RECT 7.850 47.425 8.020 47.635 ;
        RECT 8.300 47.605 8.655 47.975 ;
        RECT 7.425 46.495 7.680 47.400 ;
        RECT 7.850 47.255 8.565 47.425 ;
        RECT 7.850 46.325 8.180 47.085 ;
        RECT 8.395 46.495 8.565 47.255 ;
        RECT 8.830 46.325 9.090 47.475 ;
        RECT 9.265 47.400 9.435 48.130 ;
        RECT 9.690 47.965 9.860 48.155 ;
        RECT 9.605 47.635 9.860 47.965 ;
        RECT 9.690 47.425 9.860 47.635 ;
        RECT 10.140 47.605 10.495 47.975 ;
        RECT 12.250 47.500 12.590 48.330 ;
        RECT 9.265 46.495 9.520 47.400 ;
        RECT 9.690 47.255 10.405 47.425 ;
        RECT 9.690 46.325 10.020 47.085 ;
        RECT 10.235 46.495 10.405 47.255 ;
        RECT 14.070 46.760 14.420 48.010 ;
        RECT 16.705 47.635 17.060 48.195 ;
        RECT 17.230 47.465 17.400 48.365 ;
        RECT 17.570 47.635 17.835 48.195 ;
        RECT 18.125 48.135 18.740 48.705 ;
        RECT 19.190 48.395 19.490 48.875 ;
        RECT 19.660 48.225 19.920 48.680 ;
        RECT 20.090 48.395 20.350 48.875 ;
        RECT 20.520 48.225 20.780 48.680 ;
        RECT 20.950 48.395 21.210 48.875 ;
        RECT 21.380 48.225 21.640 48.680 ;
        RECT 21.810 48.395 22.070 48.875 ;
        RECT 22.240 48.225 22.500 48.680 ;
        RECT 22.670 48.350 22.930 48.875 ;
        RECT 18.085 47.465 18.255 47.965 ;
        RECT 16.830 47.295 18.255 47.465 ;
        RECT 16.830 47.120 17.220 47.295 ;
        RECT 10.665 46.325 16.010 46.760 ;
        RECT 17.705 46.325 18.035 47.125 ;
        RECT 18.425 47.115 18.740 48.135 ;
        RECT 19.190 48.055 22.500 48.225 ;
        RECT 19.190 47.465 20.160 48.055 ;
        RECT 23.100 47.885 23.350 48.695 ;
        RECT 23.530 48.415 23.775 48.875 ;
        RECT 24.170 48.365 24.410 48.875 ;
        RECT 24.590 48.365 24.870 48.695 ;
        RECT 25.100 48.365 25.315 48.875 ;
        RECT 20.330 47.635 23.350 47.885 ;
        RECT 23.520 47.635 23.835 48.245 ;
        RECT 24.065 47.635 24.420 48.195 ;
        RECT 19.190 47.225 22.500 47.465 ;
        RECT 18.205 46.495 18.740 47.115 ;
        RECT 19.195 46.325 19.490 47.055 ;
        RECT 19.660 46.500 19.920 47.225 ;
        RECT 20.090 46.325 20.350 47.055 ;
        RECT 20.520 46.500 20.780 47.225 ;
        RECT 20.950 46.325 21.210 47.055 ;
        RECT 21.380 46.500 21.640 47.225 ;
        RECT 21.810 46.325 22.070 47.055 ;
        RECT 22.240 46.500 22.500 47.225 ;
        RECT 22.670 46.325 22.930 47.435 ;
        RECT 23.100 46.500 23.350 47.635 ;
        RECT 24.590 47.465 24.760 48.365 ;
        RECT 24.930 47.635 25.195 48.195 ;
        RECT 25.485 48.135 26.100 48.705 ;
        RECT 25.445 47.465 25.615 47.965 ;
        RECT 23.530 46.325 23.825 47.435 ;
        RECT 24.190 47.295 25.615 47.465 ;
        RECT 24.190 47.120 24.580 47.295 ;
        RECT 25.065 46.325 25.395 47.125 ;
        RECT 25.785 47.115 26.100 48.135 ;
        RECT 26.305 48.105 27.975 48.875 ;
        RECT 28.665 48.405 28.965 48.875 ;
        RECT 29.135 48.235 29.390 48.680 ;
        RECT 29.560 48.405 29.820 48.875 ;
        RECT 29.990 48.235 30.250 48.680 ;
        RECT 30.420 48.405 30.715 48.875 ;
        RECT 26.305 47.585 27.055 48.105 ;
        RECT 28.145 48.065 31.175 48.235 ;
        RECT 31.365 48.150 31.655 48.875 ;
        RECT 27.225 47.415 27.975 47.935 ;
        RECT 25.565 46.495 26.100 47.115 ;
        RECT 26.305 46.325 27.975 47.415 ;
        RECT 28.145 47.500 28.445 48.065 ;
        RECT 28.620 47.670 30.835 47.895 ;
        RECT 31.005 47.500 31.175 48.065 ;
        RECT 28.145 47.330 31.175 47.500 ;
        RECT 28.145 46.325 28.530 47.160 ;
        RECT 28.700 46.525 28.960 47.330 ;
        RECT 29.130 46.325 29.390 47.160 ;
        RECT 29.560 46.525 29.815 47.330 ;
        RECT 29.990 46.325 30.250 47.160 ;
        RECT 30.420 46.525 30.675 47.330 ;
        RECT 30.850 46.325 31.195 47.160 ;
        RECT 31.365 46.325 31.655 47.490 ;
        RECT 32.290 47.275 32.625 48.695 ;
        RECT 32.805 48.505 33.550 48.875 ;
        RECT 34.115 48.335 34.370 48.695 ;
        RECT 34.550 48.505 34.880 48.875 ;
        RECT 35.060 48.335 35.285 48.695 ;
        RECT 32.800 48.145 35.285 48.335 ;
        RECT 36.055 48.325 36.225 48.615 ;
        RECT 36.395 48.495 36.725 48.875 ;
        RECT 36.055 48.155 36.720 48.325 ;
        RECT 32.800 47.455 33.025 48.145 ;
        RECT 33.225 47.635 33.505 47.965 ;
        RECT 33.685 47.635 34.260 47.965 ;
        RECT 34.440 47.635 34.875 47.965 ;
        RECT 35.055 47.635 35.325 47.965 ;
        RECT 32.800 47.275 35.295 47.455 ;
        RECT 35.970 47.335 36.320 47.985 ;
        RECT 32.290 46.505 32.555 47.275 ;
        RECT 32.725 46.325 33.055 47.045 ;
        RECT 33.245 46.865 34.435 47.095 ;
        RECT 33.245 46.505 33.505 46.865 ;
        RECT 33.675 46.325 34.005 46.695 ;
        RECT 34.175 46.505 34.435 46.865 ;
        RECT 35.005 46.505 35.295 47.275 ;
        RECT 36.490 47.165 36.720 48.155 ;
        RECT 36.055 46.995 36.720 47.165 ;
        RECT 36.055 46.495 36.225 46.995 ;
        RECT 36.395 46.325 36.725 46.825 ;
        RECT 36.895 46.495 37.080 48.615 ;
        RECT 37.335 48.415 37.585 48.875 ;
        RECT 37.755 48.425 38.090 48.595 ;
        RECT 38.285 48.425 38.960 48.595 ;
        RECT 37.755 48.285 37.925 48.425 ;
        RECT 37.250 47.295 37.530 48.245 ;
        RECT 37.700 48.155 37.925 48.285 ;
        RECT 37.700 47.050 37.870 48.155 ;
        RECT 38.095 48.005 38.620 48.225 ;
        RECT 38.040 47.240 38.280 47.835 ;
        RECT 38.450 47.305 38.620 48.005 ;
        RECT 38.790 47.645 38.960 48.425 ;
        RECT 39.280 48.375 39.650 48.875 ;
        RECT 39.830 48.425 40.235 48.595 ;
        RECT 40.405 48.425 41.190 48.595 ;
        RECT 39.830 48.195 40.000 48.425 ;
        RECT 39.170 47.895 40.000 48.195 ;
        RECT 40.385 47.925 40.850 48.255 ;
        RECT 39.170 47.865 39.370 47.895 ;
        RECT 39.490 47.645 39.660 47.715 ;
        RECT 38.790 47.475 39.660 47.645 ;
        RECT 39.150 47.385 39.660 47.475 ;
        RECT 37.700 46.920 38.005 47.050 ;
        RECT 38.450 46.940 38.980 47.305 ;
        RECT 37.320 46.325 37.585 46.785 ;
        RECT 37.755 46.495 38.005 46.920 ;
        RECT 39.150 46.770 39.320 47.385 ;
        RECT 38.215 46.600 39.320 46.770 ;
        RECT 39.490 46.325 39.660 47.125 ;
        RECT 39.830 46.825 40.000 47.895 ;
        RECT 40.170 46.995 40.360 47.715 ;
        RECT 40.530 46.965 40.850 47.925 ;
        RECT 41.020 47.965 41.190 48.425 ;
        RECT 41.465 48.345 41.675 48.875 ;
        RECT 41.935 48.135 42.265 48.660 ;
        RECT 42.435 48.265 42.605 48.875 ;
        RECT 42.775 48.220 43.105 48.655 ;
        RECT 43.415 48.325 43.585 48.615 ;
        RECT 43.755 48.495 44.085 48.875 ;
        RECT 42.775 48.135 43.155 48.220 ;
        RECT 43.415 48.155 44.080 48.325 ;
        RECT 42.065 47.965 42.265 48.135 ;
        RECT 42.930 48.095 43.155 48.135 ;
        RECT 41.020 47.635 41.895 47.965 ;
        RECT 42.065 47.635 42.815 47.965 ;
        RECT 39.830 46.495 40.080 46.825 ;
        RECT 41.020 46.795 41.190 47.635 ;
        RECT 42.065 47.430 42.255 47.635 ;
        RECT 42.985 47.515 43.155 48.095 ;
        RECT 42.940 47.465 43.155 47.515 ;
        RECT 41.360 47.055 42.255 47.430 ;
        RECT 42.765 47.385 43.155 47.465 ;
        RECT 40.305 46.625 41.190 46.795 ;
        RECT 41.370 46.325 41.685 46.825 ;
        RECT 41.915 46.495 42.255 47.055 ;
        RECT 42.425 46.325 42.595 47.335 ;
        RECT 42.765 46.540 43.095 47.385 ;
        RECT 43.330 47.335 43.680 47.985 ;
        RECT 43.850 47.165 44.080 48.155 ;
        RECT 43.415 46.995 44.080 47.165 ;
        RECT 43.415 46.495 43.585 46.995 ;
        RECT 43.755 46.325 44.085 46.825 ;
        RECT 44.255 46.495 44.440 48.615 ;
        RECT 44.695 48.415 44.945 48.875 ;
        RECT 45.115 48.425 45.450 48.595 ;
        RECT 45.645 48.425 46.320 48.595 ;
        RECT 45.115 48.285 45.285 48.425 ;
        RECT 44.610 47.295 44.890 48.245 ;
        RECT 45.060 48.155 45.285 48.285 ;
        RECT 45.060 47.050 45.230 48.155 ;
        RECT 45.455 48.005 45.980 48.225 ;
        RECT 45.400 47.240 45.640 47.835 ;
        RECT 45.810 47.305 45.980 48.005 ;
        RECT 46.150 47.645 46.320 48.425 ;
        RECT 46.640 48.375 47.010 48.875 ;
        RECT 47.190 48.425 47.595 48.595 ;
        RECT 47.765 48.425 48.550 48.595 ;
        RECT 47.190 48.195 47.360 48.425 ;
        RECT 46.530 47.895 47.360 48.195 ;
        RECT 47.745 47.925 48.210 48.255 ;
        RECT 46.530 47.865 46.730 47.895 ;
        RECT 46.850 47.645 47.020 47.715 ;
        RECT 46.150 47.475 47.020 47.645 ;
        RECT 46.510 47.385 47.020 47.475 ;
        RECT 45.060 46.920 45.365 47.050 ;
        RECT 45.810 46.940 46.340 47.305 ;
        RECT 44.680 46.325 44.945 46.785 ;
        RECT 45.115 46.495 45.365 46.920 ;
        RECT 46.510 46.770 46.680 47.385 ;
        RECT 45.575 46.600 46.680 46.770 ;
        RECT 46.850 46.325 47.020 47.125 ;
        RECT 47.190 46.825 47.360 47.895 ;
        RECT 47.530 46.995 47.720 47.715 ;
        RECT 47.890 46.965 48.210 47.925 ;
        RECT 48.380 47.965 48.550 48.425 ;
        RECT 48.825 48.345 49.035 48.875 ;
        RECT 49.295 48.135 49.625 48.660 ;
        RECT 49.795 48.265 49.965 48.875 ;
        RECT 50.135 48.220 50.465 48.655 ;
        RECT 50.135 48.135 50.515 48.220 ;
        RECT 49.425 47.965 49.625 48.135 ;
        RECT 50.290 48.095 50.515 48.135 ;
        RECT 48.380 47.635 49.255 47.965 ;
        RECT 49.425 47.635 50.175 47.965 ;
        RECT 47.190 46.495 47.440 46.825 ;
        RECT 48.380 46.795 48.550 47.635 ;
        RECT 49.425 47.430 49.615 47.635 ;
        RECT 50.345 47.515 50.515 48.095 ;
        RECT 50.300 47.465 50.515 47.515 ;
        RECT 48.720 47.055 49.615 47.430 ;
        RECT 50.125 47.385 50.515 47.465 ;
        RECT 50.690 48.135 50.945 48.705 ;
        RECT 51.115 48.475 51.445 48.875 ;
        RECT 51.870 48.340 52.400 48.705 ;
        RECT 52.590 48.535 52.865 48.705 ;
        RECT 52.585 48.365 52.865 48.535 ;
        RECT 51.870 48.305 52.045 48.340 ;
        RECT 51.115 48.135 52.045 48.305 ;
        RECT 50.690 47.465 50.860 48.135 ;
        RECT 51.115 47.965 51.285 48.135 ;
        RECT 51.030 47.635 51.285 47.965 ;
        RECT 51.510 47.635 51.705 47.965 ;
        RECT 47.665 46.625 48.550 46.795 ;
        RECT 48.730 46.325 49.045 46.825 ;
        RECT 49.275 46.495 49.615 47.055 ;
        RECT 49.785 46.325 49.955 47.335 ;
        RECT 50.125 46.540 50.455 47.385 ;
        RECT 50.690 46.495 51.025 47.465 ;
        RECT 51.195 46.325 51.365 47.465 ;
        RECT 51.535 46.665 51.705 47.635 ;
        RECT 51.875 47.005 52.045 48.135 ;
        RECT 52.215 47.345 52.385 48.145 ;
        RECT 52.590 47.545 52.865 48.365 ;
        RECT 53.035 47.345 53.225 48.705 ;
        RECT 53.405 48.340 53.915 48.875 ;
        RECT 54.135 48.065 54.380 48.670 ;
        RECT 54.825 48.105 56.495 48.875 ;
        RECT 57.125 48.150 57.415 48.875 ;
        RECT 57.585 48.330 62.930 48.875 ;
        RECT 63.105 48.330 68.450 48.875 ;
        RECT 53.425 47.895 54.655 48.065 ;
        RECT 52.215 47.175 53.225 47.345 ;
        RECT 53.395 47.330 54.145 47.520 ;
        RECT 51.875 46.835 53.000 47.005 ;
        RECT 53.395 46.665 53.565 47.330 ;
        RECT 54.315 47.085 54.655 47.895 ;
        RECT 54.825 47.585 55.575 48.105 ;
        RECT 55.745 47.415 56.495 47.935 ;
        RECT 59.170 47.500 59.510 48.330 ;
        RECT 51.535 46.495 53.565 46.665 ;
        RECT 53.735 46.325 53.905 47.085 ;
        RECT 54.140 46.675 54.655 47.085 ;
        RECT 54.825 46.325 56.495 47.415 ;
        RECT 57.125 46.325 57.415 47.490 ;
        RECT 60.990 46.760 61.340 48.010 ;
        RECT 64.690 47.500 65.030 48.330 ;
        RECT 68.625 48.105 70.295 48.875 ;
        RECT 66.510 46.760 66.860 48.010 ;
        RECT 68.625 47.585 69.375 48.105 ;
        RECT 70.505 48.055 70.735 48.875 ;
        RECT 70.905 48.075 71.235 48.705 ;
        RECT 69.545 47.415 70.295 47.935 ;
        RECT 70.485 47.635 70.815 47.885 ;
        RECT 70.985 47.475 71.235 48.075 ;
        RECT 71.405 48.055 71.615 48.875 ;
        RECT 71.845 48.330 77.190 48.875 ;
        RECT 73.430 47.500 73.770 48.330 ;
        RECT 77.365 48.105 80.875 48.875 ;
        RECT 81.505 48.200 81.765 48.705 ;
        RECT 81.945 48.495 82.275 48.875 ;
        RECT 82.455 48.325 82.625 48.705 ;
        RECT 57.585 46.325 62.930 46.760 ;
        RECT 63.105 46.325 68.450 46.760 ;
        RECT 68.625 46.325 70.295 47.415 ;
        RECT 70.505 46.325 70.735 47.465 ;
        RECT 70.905 46.495 71.235 47.475 ;
        RECT 71.405 46.325 71.615 47.465 ;
        RECT 75.250 46.760 75.600 48.010 ;
        RECT 77.365 47.585 79.015 48.105 ;
        RECT 79.185 47.415 80.875 47.935 ;
        RECT 71.845 46.325 77.190 46.760 ;
        RECT 77.365 46.325 80.875 47.415 ;
        RECT 81.505 47.400 81.675 48.200 ;
        RECT 81.960 48.155 82.625 48.325 ;
        RECT 81.960 47.900 82.130 48.155 ;
        RECT 82.885 48.125 84.095 48.875 ;
        RECT 81.845 47.570 82.130 47.900 ;
        RECT 82.365 47.605 82.695 47.975 ;
        RECT 81.960 47.425 82.130 47.570 ;
        RECT 81.505 46.495 81.775 47.400 ;
        RECT 81.960 47.255 82.625 47.425 ;
        RECT 81.945 46.325 82.275 47.085 ;
        RECT 82.455 46.495 82.625 47.255 ;
        RECT 82.885 47.415 83.405 47.955 ;
        RECT 83.575 47.585 84.095 48.125 ;
        RECT 82.885 46.325 84.095 47.415 ;
        RECT 5.520 46.155 84.180 46.325 ;
        RECT 5.605 45.065 6.815 46.155 ;
        RECT 5.605 44.355 6.125 44.895 ;
        RECT 6.295 44.525 6.815 45.065 ;
        RECT 6.990 45.005 7.250 46.155 ;
        RECT 7.425 45.080 7.680 45.985 ;
        RECT 7.850 45.395 8.180 46.155 ;
        RECT 8.395 45.225 8.565 45.985 ;
        RECT 5.605 43.605 6.815 44.355 ;
        RECT 6.990 43.605 7.250 44.445 ;
        RECT 7.425 44.350 7.595 45.080 ;
        RECT 7.850 45.055 8.565 45.225 ;
        RECT 9.950 45.185 10.280 45.985 ;
        RECT 10.450 45.355 10.780 46.155 ;
        RECT 11.080 45.185 11.410 45.985 ;
        RECT 12.055 45.355 12.305 46.155 ;
        RECT 7.850 44.845 8.020 45.055 ;
        RECT 9.950 45.015 12.385 45.185 ;
        RECT 12.575 45.015 12.745 46.155 ;
        RECT 12.915 45.015 13.255 45.985 ;
        RECT 7.765 44.515 8.020 44.845 ;
        RECT 7.425 43.775 7.680 44.350 ;
        RECT 7.850 44.325 8.020 44.515 ;
        RECT 8.300 44.505 8.655 44.875 ;
        RECT 9.745 44.595 10.095 44.845 ;
        RECT 10.280 44.385 10.450 45.015 ;
        RECT 10.620 44.595 10.950 44.795 ;
        RECT 11.120 44.595 11.450 44.795 ;
        RECT 11.620 44.595 12.040 44.795 ;
        RECT 12.215 44.765 12.385 45.015 ;
        RECT 12.215 44.595 12.910 44.765 ;
        RECT 7.850 44.155 8.565 44.325 ;
        RECT 7.850 43.605 8.180 43.985 ;
        RECT 8.395 43.775 8.565 44.155 ;
        RECT 9.950 43.775 10.450 44.385 ;
        RECT 11.080 44.255 12.305 44.425 ;
        RECT 13.080 44.405 13.255 45.015 ;
        RECT 13.430 45.005 13.690 46.155 ;
        RECT 13.865 45.080 14.120 45.985 ;
        RECT 14.290 45.395 14.620 46.155 ;
        RECT 14.835 45.225 15.005 45.985 ;
        RECT 11.080 43.775 11.410 44.255 ;
        RECT 11.580 43.605 11.805 44.065 ;
        RECT 11.975 43.775 12.305 44.255 ;
        RECT 12.495 43.605 12.745 44.405 ;
        RECT 12.915 43.775 13.255 44.405 ;
        RECT 13.430 43.605 13.690 44.445 ;
        RECT 13.865 44.350 14.035 45.080 ;
        RECT 14.290 45.055 15.005 45.225 ;
        RECT 15.265 45.065 17.855 46.155 ;
        RECT 14.290 44.845 14.460 45.055 ;
        RECT 14.205 44.515 14.460 44.845 ;
        RECT 13.865 43.775 14.120 44.350 ;
        RECT 14.290 44.325 14.460 44.515 ;
        RECT 14.740 44.505 15.095 44.875 ;
        RECT 15.265 44.375 16.475 44.895 ;
        RECT 16.645 44.545 17.855 45.065 ;
        RECT 18.485 44.990 18.775 46.155 ;
        RECT 19.610 45.185 19.940 45.985 ;
        RECT 20.110 45.355 20.440 46.155 ;
        RECT 20.740 45.185 21.070 45.985 ;
        RECT 21.715 45.355 21.965 46.155 ;
        RECT 19.610 45.015 22.045 45.185 ;
        RECT 22.235 45.015 22.405 46.155 ;
        RECT 22.575 45.015 22.915 45.985 ;
        RECT 23.175 45.485 23.345 45.985 ;
        RECT 23.515 45.655 23.845 46.155 ;
        RECT 23.175 45.315 23.840 45.485 ;
        RECT 19.405 44.595 19.755 44.845 ;
        RECT 19.940 44.385 20.110 45.015 ;
        RECT 20.280 44.595 20.610 44.795 ;
        RECT 20.780 44.595 21.110 44.795 ;
        RECT 21.280 44.595 21.700 44.795 ;
        RECT 21.875 44.765 22.045 45.015 ;
        RECT 21.875 44.595 22.570 44.765 ;
        RECT 22.740 44.455 22.915 45.015 ;
        RECT 23.090 44.495 23.440 45.145 ;
        RECT 14.290 44.155 15.005 44.325 ;
        RECT 14.290 43.605 14.620 43.985 ;
        RECT 14.835 43.775 15.005 44.155 ;
        RECT 15.265 43.605 17.855 44.375 ;
        RECT 18.485 43.605 18.775 44.330 ;
        RECT 19.610 43.775 20.110 44.385 ;
        RECT 20.740 44.255 21.965 44.425 ;
        RECT 22.685 44.405 22.915 44.455 ;
        RECT 20.740 43.775 21.070 44.255 ;
        RECT 21.240 43.605 21.465 44.065 ;
        RECT 21.635 43.775 21.965 44.255 ;
        RECT 22.155 43.605 22.405 44.405 ;
        RECT 22.575 43.775 22.915 44.405 ;
        RECT 23.610 44.325 23.840 45.315 ;
        RECT 23.175 44.155 23.840 44.325 ;
        RECT 23.175 43.865 23.345 44.155 ;
        RECT 23.515 43.605 23.845 43.985 ;
        RECT 24.015 43.865 24.200 45.985 ;
        RECT 24.440 45.695 24.705 46.155 ;
        RECT 24.875 45.560 25.125 45.985 ;
        RECT 25.335 45.710 26.440 45.880 ;
        RECT 24.820 45.430 25.125 45.560 ;
        RECT 24.370 44.235 24.650 45.185 ;
        RECT 24.820 44.325 24.990 45.430 ;
        RECT 25.160 44.645 25.400 45.240 ;
        RECT 25.570 45.175 26.100 45.540 ;
        RECT 25.570 44.475 25.740 45.175 ;
        RECT 26.270 45.095 26.440 45.710 ;
        RECT 26.610 45.355 26.780 46.155 ;
        RECT 26.950 45.655 27.200 45.985 ;
        RECT 27.425 45.685 28.310 45.855 ;
        RECT 26.270 45.005 26.780 45.095 ;
        RECT 24.820 44.195 25.045 44.325 ;
        RECT 25.215 44.255 25.740 44.475 ;
        RECT 25.910 44.835 26.780 45.005 ;
        RECT 24.455 43.605 24.705 44.065 ;
        RECT 24.875 44.055 25.045 44.195 ;
        RECT 25.910 44.055 26.080 44.835 ;
        RECT 26.610 44.765 26.780 44.835 ;
        RECT 26.290 44.585 26.490 44.615 ;
        RECT 26.950 44.585 27.120 45.655 ;
        RECT 27.290 44.765 27.480 45.485 ;
        RECT 26.290 44.285 27.120 44.585 ;
        RECT 27.650 44.555 27.970 45.515 ;
        RECT 24.875 43.885 25.210 44.055 ;
        RECT 25.405 43.885 26.080 44.055 ;
        RECT 26.400 43.605 26.770 44.105 ;
        RECT 26.950 44.055 27.120 44.285 ;
        RECT 27.505 44.225 27.970 44.555 ;
        RECT 28.140 44.845 28.310 45.685 ;
        RECT 28.490 45.655 28.805 46.155 ;
        RECT 29.035 45.425 29.375 45.985 ;
        RECT 28.480 45.050 29.375 45.425 ;
        RECT 29.545 45.145 29.715 46.155 ;
        RECT 29.185 44.845 29.375 45.050 ;
        RECT 29.885 45.095 30.215 45.940 ;
        RECT 30.535 45.485 30.705 45.985 ;
        RECT 30.875 45.655 31.205 46.155 ;
        RECT 30.535 45.315 31.200 45.485 ;
        RECT 29.885 45.015 30.275 45.095 ;
        RECT 30.060 44.965 30.275 45.015 ;
        RECT 28.140 44.515 29.015 44.845 ;
        RECT 29.185 44.515 29.935 44.845 ;
        RECT 28.140 44.055 28.310 44.515 ;
        RECT 29.185 44.345 29.385 44.515 ;
        RECT 30.105 44.385 30.275 44.965 ;
        RECT 30.450 44.495 30.800 45.145 ;
        RECT 30.050 44.345 30.275 44.385 ;
        RECT 26.950 43.885 27.355 44.055 ;
        RECT 27.525 43.885 28.310 44.055 ;
        RECT 28.585 43.605 28.795 44.135 ;
        RECT 29.055 43.820 29.385 44.345 ;
        RECT 29.895 44.260 30.275 44.345 ;
        RECT 30.970 44.325 31.200 45.315 ;
        RECT 29.555 43.605 29.725 44.215 ;
        RECT 29.895 43.825 30.225 44.260 ;
        RECT 30.535 44.155 31.200 44.325 ;
        RECT 30.535 43.865 30.705 44.155 ;
        RECT 30.875 43.605 31.205 43.985 ;
        RECT 31.375 43.865 31.560 45.985 ;
        RECT 31.800 45.695 32.065 46.155 ;
        RECT 32.235 45.560 32.485 45.985 ;
        RECT 32.695 45.710 33.800 45.880 ;
        RECT 32.180 45.430 32.485 45.560 ;
        RECT 31.730 44.235 32.010 45.185 ;
        RECT 32.180 44.325 32.350 45.430 ;
        RECT 32.520 44.645 32.760 45.240 ;
        RECT 32.930 45.175 33.460 45.540 ;
        RECT 32.930 44.475 33.100 45.175 ;
        RECT 33.630 45.095 33.800 45.710 ;
        RECT 33.970 45.355 34.140 46.155 ;
        RECT 34.310 45.655 34.560 45.985 ;
        RECT 34.785 45.685 35.670 45.855 ;
        RECT 33.630 45.005 34.140 45.095 ;
        RECT 32.180 44.195 32.405 44.325 ;
        RECT 32.575 44.255 33.100 44.475 ;
        RECT 33.270 44.835 34.140 45.005 ;
        RECT 31.815 43.605 32.065 44.065 ;
        RECT 32.235 44.055 32.405 44.195 ;
        RECT 33.270 44.055 33.440 44.835 ;
        RECT 33.970 44.765 34.140 44.835 ;
        RECT 33.650 44.585 33.850 44.615 ;
        RECT 34.310 44.585 34.480 45.655 ;
        RECT 34.650 44.765 34.840 45.485 ;
        RECT 33.650 44.285 34.480 44.585 ;
        RECT 35.010 44.555 35.330 45.515 ;
        RECT 32.235 43.885 32.570 44.055 ;
        RECT 32.765 43.885 33.440 44.055 ;
        RECT 33.760 43.605 34.130 44.105 ;
        RECT 34.310 44.055 34.480 44.285 ;
        RECT 34.865 44.225 35.330 44.555 ;
        RECT 35.500 44.845 35.670 45.685 ;
        RECT 35.850 45.655 36.165 46.155 ;
        RECT 36.395 45.425 36.735 45.985 ;
        RECT 35.840 45.050 36.735 45.425 ;
        RECT 36.905 45.145 37.075 46.155 ;
        RECT 36.545 44.845 36.735 45.050 ;
        RECT 37.245 45.095 37.575 45.940 ;
        RECT 37.245 45.015 37.635 45.095 ;
        RECT 37.420 44.965 37.635 45.015 ;
        RECT 35.500 44.515 36.375 44.845 ;
        RECT 36.545 44.515 37.295 44.845 ;
        RECT 35.500 44.055 35.670 44.515 ;
        RECT 36.545 44.345 36.745 44.515 ;
        RECT 37.465 44.385 37.635 44.965 ;
        RECT 37.410 44.345 37.635 44.385 ;
        RECT 34.310 43.885 34.715 44.055 ;
        RECT 34.885 43.885 35.670 44.055 ;
        RECT 35.945 43.605 36.155 44.135 ;
        RECT 36.415 43.820 36.745 44.345 ;
        RECT 37.255 44.260 37.635 44.345 ;
        RECT 37.810 45.015 38.145 45.985 ;
        RECT 38.315 45.015 38.485 46.155 ;
        RECT 38.655 45.815 40.685 45.985 ;
        RECT 37.810 44.345 37.980 45.015 ;
        RECT 38.655 44.845 38.825 45.815 ;
        RECT 38.150 44.515 38.405 44.845 ;
        RECT 38.630 44.515 38.825 44.845 ;
        RECT 38.995 45.475 40.120 45.645 ;
        RECT 38.235 44.345 38.405 44.515 ;
        RECT 38.995 44.345 39.165 45.475 ;
        RECT 36.915 43.605 37.085 44.215 ;
        RECT 37.255 43.825 37.585 44.260 ;
        RECT 37.810 43.775 38.065 44.345 ;
        RECT 38.235 44.175 39.165 44.345 ;
        RECT 39.335 45.135 40.345 45.305 ;
        RECT 39.335 44.335 39.505 45.135 ;
        RECT 39.710 44.455 39.985 44.935 ;
        RECT 39.705 44.285 39.985 44.455 ;
        RECT 38.990 44.140 39.165 44.175 ;
        RECT 38.235 43.605 38.565 44.005 ;
        RECT 38.990 43.775 39.520 44.140 ;
        RECT 39.710 43.775 39.985 44.285 ;
        RECT 40.155 43.775 40.345 45.135 ;
        RECT 40.515 45.150 40.685 45.815 ;
        RECT 40.855 45.395 41.025 46.155 ;
        RECT 41.260 45.395 41.775 45.805 ;
        RECT 40.515 44.960 41.265 45.150 ;
        RECT 41.435 44.585 41.775 45.395 ;
        RECT 41.945 45.065 43.615 46.155 ;
        RECT 40.545 44.415 41.775 44.585 ;
        RECT 40.525 43.605 41.035 44.140 ;
        RECT 41.255 43.810 41.500 44.415 ;
        RECT 41.945 44.375 42.695 44.895 ;
        RECT 42.865 44.545 43.615 45.065 ;
        RECT 44.245 44.990 44.535 46.155 ;
        RECT 44.705 45.015 45.090 45.985 ;
        RECT 45.260 45.695 45.585 46.155 ;
        RECT 46.105 45.525 46.385 45.985 ;
        RECT 45.260 45.305 46.385 45.525 ;
        RECT 41.945 43.605 43.615 44.375 ;
        RECT 44.705 44.345 44.985 45.015 ;
        RECT 45.260 44.845 45.710 45.305 ;
        RECT 46.575 45.135 46.975 45.985 ;
        RECT 47.375 45.695 47.645 46.155 ;
        RECT 47.815 45.525 48.100 45.985 ;
        RECT 48.385 45.650 49.015 46.155 ;
        RECT 45.155 44.515 45.710 44.845 ;
        RECT 45.880 44.575 46.975 45.135 ;
        RECT 45.260 44.405 45.710 44.515 ;
        RECT 44.245 43.605 44.535 44.330 ;
        RECT 44.705 43.775 45.090 44.345 ;
        RECT 45.260 44.235 46.385 44.405 ;
        RECT 45.260 43.605 45.585 44.065 ;
        RECT 46.105 43.775 46.385 44.235 ;
        RECT 46.575 43.775 46.975 44.575 ;
        RECT 47.145 45.305 48.100 45.525 ;
        RECT 47.145 44.405 47.355 45.305 ;
        RECT 47.525 44.575 48.215 45.135 ;
        RECT 48.400 45.115 48.655 45.480 ;
        RECT 48.825 45.475 49.015 45.650 ;
        RECT 49.195 45.645 49.670 45.985 ;
        RECT 48.825 45.285 49.155 45.475 ;
        RECT 49.380 45.115 49.630 45.410 ;
        RECT 49.855 45.310 50.070 46.155 ;
        RECT 50.270 45.315 50.545 45.985 ;
        RECT 48.400 44.945 50.190 45.115 ;
        RECT 50.375 44.965 50.545 45.315 ;
        RECT 50.715 45.145 50.975 46.155 ;
        RECT 51.145 45.185 51.415 45.955 ;
        RECT 51.585 45.375 51.915 46.155 ;
        RECT 52.120 45.550 52.305 45.955 ;
        RECT 52.475 45.730 52.810 46.155 ;
        RECT 52.120 45.375 52.785 45.550 ;
        RECT 51.145 45.015 52.275 45.185 ;
        RECT 47.145 44.235 48.100 44.405 ;
        RECT 48.385 44.285 48.770 44.765 ;
        RECT 47.375 43.605 47.645 44.065 ;
        RECT 47.815 43.775 48.100 44.235 ;
        RECT 48.940 44.090 49.195 44.945 ;
        RECT 48.405 43.825 49.195 44.090 ;
        RECT 49.365 44.270 49.775 44.765 ;
        RECT 49.960 44.515 50.190 44.945 ;
        RECT 50.360 44.445 50.975 44.965 ;
        RECT 49.365 43.825 49.595 44.270 ;
        RECT 50.360 44.235 50.530 44.445 ;
        RECT 49.775 43.605 50.105 44.100 ;
        RECT 50.280 43.775 50.530 44.235 ;
        RECT 50.700 43.605 50.975 44.265 ;
        RECT 51.145 44.105 51.315 45.015 ;
        RECT 51.485 44.265 51.845 44.845 ;
        RECT 52.025 44.515 52.275 45.015 ;
        RECT 52.445 44.345 52.785 45.375 ;
        RECT 52.985 45.065 54.195 46.155 ;
        RECT 52.100 44.175 52.785 44.345 ;
        RECT 52.985 44.355 53.505 44.895 ;
        RECT 53.675 44.525 54.195 45.065 ;
        RECT 54.365 45.305 54.625 45.985 ;
        RECT 54.795 45.375 55.045 46.155 ;
        RECT 55.295 45.605 55.545 45.985 ;
        RECT 55.715 45.775 56.070 46.155 ;
        RECT 57.075 45.765 57.410 45.985 ;
        RECT 56.675 45.605 56.905 45.645 ;
        RECT 55.295 45.405 56.905 45.605 ;
        RECT 55.295 45.395 56.130 45.405 ;
        RECT 56.720 45.315 56.905 45.405 ;
        RECT 51.145 43.775 51.405 44.105 ;
        RECT 51.615 43.605 51.890 44.085 ;
        RECT 52.100 43.775 52.305 44.175 ;
        RECT 52.475 43.605 52.810 44.005 ;
        RECT 52.985 43.605 54.195 44.355 ;
        RECT 54.365 44.105 54.535 45.305 ;
        RECT 56.235 45.205 56.565 45.235 ;
        RECT 54.765 45.145 56.565 45.205 ;
        RECT 57.155 45.145 57.410 45.765 ;
        RECT 57.585 45.560 58.020 45.985 ;
        RECT 58.190 45.730 58.575 46.155 ;
        RECT 57.585 45.390 58.575 45.560 ;
        RECT 54.705 45.035 57.410 45.145 ;
        RECT 54.705 45.000 54.905 45.035 ;
        RECT 54.705 44.425 54.875 45.000 ;
        RECT 56.235 44.975 57.410 45.035 ;
        RECT 55.105 44.560 55.515 44.865 ;
        RECT 55.685 44.595 56.015 44.805 ;
        RECT 54.705 44.305 54.975 44.425 ;
        RECT 54.705 44.260 55.550 44.305 ;
        RECT 54.795 44.135 55.550 44.260 ;
        RECT 55.805 44.195 56.015 44.595 ;
        RECT 56.260 44.595 56.735 44.805 ;
        RECT 56.925 44.595 57.415 44.795 ;
        RECT 56.260 44.195 56.480 44.595 ;
        RECT 57.585 44.515 58.070 45.220 ;
        RECT 58.240 44.845 58.575 45.390 ;
        RECT 58.745 45.195 59.170 45.985 ;
        RECT 59.340 45.560 59.615 45.985 ;
        RECT 59.785 45.730 60.170 46.155 ;
        RECT 59.340 45.365 60.170 45.560 ;
        RECT 58.745 45.015 59.650 45.195 ;
        RECT 58.240 44.515 58.650 44.845 ;
        RECT 58.820 44.515 59.650 45.015 ;
        RECT 59.820 44.845 60.170 45.365 ;
        RECT 60.340 45.195 60.585 45.985 ;
        RECT 60.775 45.560 61.030 45.985 ;
        RECT 61.200 45.730 61.585 46.155 ;
        RECT 60.775 45.365 61.585 45.560 ;
        RECT 60.340 45.015 61.065 45.195 ;
        RECT 59.820 44.515 60.245 44.845 ;
        RECT 60.415 44.515 61.065 45.015 ;
        RECT 61.235 44.845 61.585 45.365 ;
        RECT 61.755 45.015 62.015 45.985 ;
        RECT 61.235 44.515 61.660 44.845 ;
        RECT 54.365 43.775 54.625 44.105 ;
        RECT 55.380 43.985 55.550 44.135 ;
        RECT 54.795 43.605 55.125 43.965 ;
        RECT 55.380 43.775 56.680 43.985 ;
        RECT 56.955 43.605 57.410 44.370 ;
        RECT 58.240 44.345 58.575 44.515 ;
        RECT 58.820 44.345 59.170 44.515 ;
        RECT 59.820 44.345 60.170 44.515 ;
        RECT 60.415 44.345 60.585 44.515 ;
        RECT 61.235 44.345 61.585 44.515 ;
        RECT 61.830 44.345 62.015 45.015 ;
        RECT 62.190 45.765 62.525 45.985 ;
        RECT 63.530 45.775 63.885 46.155 ;
        RECT 62.190 45.145 62.445 45.765 ;
        RECT 62.695 45.605 62.925 45.645 ;
        RECT 64.055 45.605 64.305 45.985 ;
        RECT 62.695 45.405 64.305 45.605 ;
        RECT 62.695 45.315 62.880 45.405 ;
        RECT 63.470 45.395 64.305 45.405 ;
        RECT 64.555 45.375 64.805 46.155 ;
        RECT 64.975 45.305 65.235 45.985 ;
        RECT 63.035 45.205 63.365 45.235 ;
        RECT 63.035 45.145 64.835 45.205 ;
        RECT 62.190 45.035 64.895 45.145 ;
        RECT 62.190 44.975 63.365 45.035 ;
        RECT 64.695 45.000 64.895 45.035 ;
        RECT 62.185 44.595 62.675 44.795 ;
        RECT 62.865 44.595 63.340 44.805 ;
        RECT 57.585 44.175 58.575 44.345 ;
        RECT 57.585 43.775 58.020 44.175 ;
        RECT 58.190 43.605 58.575 44.005 ;
        RECT 58.745 43.775 59.170 44.345 ;
        RECT 59.360 44.175 60.170 44.345 ;
        RECT 59.360 43.775 59.615 44.175 ;
        RECT 59.785 43.605 60.170 44.005 ;
        RECT 60.340 43.775 60.585 44.345 ;
        RECT 60.775 44.175 61.585 44.345 ;
        RECT 60.775 43.775 61.030 44.175 ;
        RECT 61.200 43.605 61.585 44.005 ;
        RECT 61.755 43.775 62.015 44.345 ;
        RECT 62.190 43.605 62.645 44.370 ;
        RECT 63.120 44.195 63.340 44.595 ;
        RECT 63.585 44.595 63.915 44.805 ;
        RECT 63.585 44.195 63.795 44.595 ;
        RECT 64.085 44.560 64.495 44.865 ;
        RECT 64.725 44.425 64.895 45.000 ;
        RECT 64.625 44.305 64.895 44.425 ;
        RECT 64.050 44.260 64.895 44.305 ;
        RECT 64.050 44.135 64.805 44.260 ;
        RECT 64.050 43.985 64.220 44.135 ;
        RECT 65.065 44.105 65.235 45.305 ;
        RECT 62.920 43.775 64.220 43.985 ;
        RECT 64.475 43.605 64.805 43.965 ;
        RECT 64.975 43.775 65.235 44.105 ;
        RECT 65.440 45.365 65.975 45.985 ;
        RECT 65.440 44.345 65.755 45.365 ;
        RECT 66.145 45.355 66.475 46.155 ;
        RECT 66.960 45.185 67.350 45.360 ;
        RECT 65.925 45.015 67.350 45.185 ;
        RECT 67.705 45.065 69.375 46.155 ;
        RECT 65.925 44.515 66.095 45.015 ;
        RECT 65.440 43.775 66.055 44.345 ;
        RECT 66.345 44.285 66.610 44.845 ;
        RECT 66.780 44.115 66.950 45.015 ;
        RECT 67.120 44.285 67.475 44.845 ;
        RECT 67.705 44.375 68.455 44.895 ;
        RECT 68.625 44.545 69.375 45.065 ;
        RECT 70.005 44.990 70.295 46.155 ;
        RECT 70.670 45.185 71.000 45.985 ;
        RECT 71.170 45.355 71.500 46.155 ;
        RECT 71.800 45.185 72.130 45.985 ;
        RECT 72.775 45.355 73.025 46.155 ;
        RECT 70.670 45.015 73.105 45.185 ;
        RECT 73.295 45.015 73.465 46.155 ;
        RECT 73.635 45.015 73.975 45.985 ;
        RECT 74.145 45.720 79.490 46.155 ;
        RECT 70.465 44.595 70.815 44.845 ;
        RECT 71.000 44.385 71.170 45.015 ;
        RECT 71.340 44.595 71.670 44.795 ;
        RECT 71.840 44.595 72.170 44.795 ;
        RECT 72.340 44.595 72.760 44.795 ;
        RECT 72.935 44.765 73.105 45.015 ;
        RECT 72.935 44.595 73.630 44.765 ;
        RECT 66.225 43.605 66.440 44.115 ;
        RECT 66.670 43.785 66.950 44.115 ;
        RECT 67.130 43.605 67.370 44.115 ;
        RECT 67.705 43.605 69.375 44.375 ;
        RECT 70.005 43.605 70.295 44.330 ;
        RECT 70.670 43.775 71.170 44.385 ;
        RECT 71.800 44.255 73.025 44.425 ;
        RECT 73.800 44.405 73.975 45.015 ;
        RECT 71.800 43.775 72.130 44.255 ;
        RECT 72.300 43.605 72.525 44.065 ;
        RECT 72.695 43.775 73.025 44.255 ;
        RECT 73.215 43.605 73.465 44.405 ;
        RECT 73.635 43.775 73.975 44.405 ;
        RECT 75.730 44.150 76.070 44.980 ;
        RECT 77.550 44.470 77.900 45.720 ;
        RECT 79.665 45.065 82.255 46.155 ;
        RECT 79.665 44.375 80.875 44.895 ;
        RECT 81.045 44.545 82.255 45.065 ;
        RECT 82.885 45.065 84.095 46.155 ;
        RECT 82.885 44.525 83.405 45.065 ;
        RECT 74.145 43.605 79.490 44.150 ;
        RECT 79.665 43.605 82.255 44.375 ;
        RECT 83.575 44.355 84.095 44.895 ;
        RECT 82.885 43.605 84.095 44.355 ;
        RECT 5.520 43.435 84.180 43.605 ;
        RECT 5.605 42.685 6.815 43.435 ;
        RECT 6.985 42.685 8.195 43.435 ;
        RECT 8.530 42.925 8.770 43.435 ;
        RECT 8.950 42.925 9.230 43.255 ;
        RECT 9.460 42.925 9.675 43.435 ;
        RECT 5.605 42.145 6.125 42.685 ;
        RECT 6.295 41.975 6.815 42.515 ;
        RECT 6.985 42.145 7.505 42.685 ;
        RECT 7.675 41.975 8.195 42.515 ;
        RECT 8.425 42.195 8.780 42.755 ;
        RECT 8.950 42.025 9.120 42.925 ;
        RECT 9.290 42.195 9.555 42.755 ;
        RECT 9.845 42.695 10.460 43.265 ;
        RECT 10.755 42.885 10.925 43.175 ;
        RECT 11.095 43.055 11.425 43.435 ;
        RECT 10.755 42.715 11.420 42.885 ;
        RECT 9.805 42.025 9.975 42.525 ;
        RECT 5.605 40.885 6.815 41.975 ;
        RECT 6.985 40.885 8.195 41.975 ;
        RECT 8.550 41.855 9.975 42.025 ;
        RECT 8.550 41.680 8.940 41.855 ;
        RECT 9.425 40.885 9.755 41.685 ;
        RECT 10.145 41.675 10.460 42.695 ;
        RECT 10.670 41.895 11.020 42.545 ;
        RECT 11.190 41.725 11.420 42.715 ;
        RECT 9.925 41.055 10.460 41.675 ;
        RECT 10.755 41.555 11.420 41.725 ;
        RECT 10.755 41.055 10.925 41.555 ;
        RECT 11.095 40.885 11.425 41.385 ;
        RECT 11.595 41.055 11.780 43.175 ;
        RECT 12.035 42.975 12.285 43.435 ;
        RECT 12.455 42.985 12.790 43.155 ;
        RECT 12.985 42.985 13.660 43.155 ;
        RECT 12.455 42.845 12.625 42.985 ;
        RECT 11.950 41.855 12.230 42.805 ;
        RECT 12.400 42.715 12.625 42.845 ;
        RECT 12.400 41.610 12.570 42.715 ;
        RECT 12.795 42.565 13.320 42.785 ;
        RECT 12.740 41.800 12.980 42.395 ;
        RECT 13.150 41.865 13.320 42.565 ;
        RECT 13.490 42.205 13.660 42.985 ;
        RECT 13.980 42.935 14.350 43.435 ;
        RECT 14.530 42.985 14.935 43.155 ;
        RECT 15.105 42.985 15.890 43.155 ;
        RECT 14.530 42.755 14.700 42.985 ;
        RECT 13.870 42.455 14.700 42.755 ;
        RECT 15.085 42.485 15.550 42.815 ;
        RECT 13.870 42.425 14.070 42.455 ;
        RECT 14.190 42.205 14.360 42.275 ;
        RECT 13.490 42.035 14.360 42.205 ;
        RECT 13.850 41.945 14.360 42.035 ;
        RECT 12.400 41.480 12.705 41.610 ;
        RECT 13.150 41.500 13.680 41.865 ;
        RECT 12.020 40.885 12.285 41.345 ;
        RECT 12.455 41.055 12.705 41.480 ;
        RECT 13.850 41.330 14.020 41.945 ;
        RECT 12.915 41.160 14.020 41.330 ;
        RECT 14.190 40.885 14.360 41.685 ;
        RECT 14.530 41.385 14.700 42.455 ;
        RECT 14.870 41.555 15.060 42.275 ;
        RECT 15.230 41.525 15.550 42.485 ;
        RECT 15.720 42.525 15.890 42.985 ;
        RECT 16.165 42.905 16.375 43.435 ;
        RECT 16.635 42.695 16.965 43.220 ;
        RECT 17.135 42.825 17.305 43.435 ;
        RECT 17.475 42.780 17.805 43.215 ;
        RECT 18.190 42.925 18.430 43.435 ;
        RECT 18.610 42.925 18.890 43.255 ;
        RECT 19.120 42.925 19.335 43.435 ;
        RECT 17.475 42.695 17.855 42.780 ;
        RECT 16.765 42.525 16.965 42.695 ;
        RECT 17.630 42.655 17.855 42.695 ;
        RECT 15.720 42.195 16.595 42.525 ;
        RECT 16.765 42.195 17.515 42.525 ;
        RECT 14.530 41.055 14.780 41.385 ;
        RECT 15.720 41.355 15.890 42.195 ;
        RECT 16.765 41.990 16.955 42.195 ;
        RECT 17.685 42.075 17.855 42.655 ;
        RECT 18.085 42.195 18.440 42.755 ;
        RECT 17.640 42.025 17.855 42.075 ;
        RECT 18.610 42.025 18.780 42.925 ;
        RECT 18.950 42.195 19.215 42.755 ;
        RECT 19.505 42.695 20.120 43.265 ;
        RECT 19.465 42.025 19.635 42.525 ;
        RECT 16.060 41.615 16.955 41.990 ;
        RECT 17.465 41.945 17.855 42.025 ;
        RECT 15.005 41.185 15.890 41.355 ;
        RECT 16.070 40.885 16.385 41.385 ;
        RECT 16.615 41.055 16.955 41.615 ;
        RECT 17.125 40.885 17.295 41.895 ;
        RECT 17.465 41.100 17.795 41.945 ;
        RECT 18.210 41.855 19.635 42.025 ;
        RECT 18.210 41.680 18.600 41.855 ;
        RECT 19.085 40.885 19.415 41.685 ;
        RECT 19.805 41.675 20.120 42.695 ;
        RECT 20.530 42.655 21.030 43.265 ;
        RECT 20.325 42.195 20.675 42.445 ;
        RECT 20.860 42.025 21.030 42.655 ;
        RECT 21.660 42.785 21.990 43.265 ;
        RECT 22.160 42.975 22.385 43.435 ;
        RECT 22.555 42.785 22.885 43.265 ;
        RECT 21.660 42.615 22.885 42.785 ;
        RECT 23.075 42.635 23.325 43.435 ;
        RECT 23.495 42.635 23.835 43.265 ;
        RECT 24.095 42.885 24.265 43.175 ;
        RECT 24.435 43.055 24.765 43.435 ;
        RECT 24.095 42.715 24.760 42.885 ;
        RECT 21.200 42.245 21.530 42.445 ;
        RECT 21.700 42.245 22.030 42.445 ;
        RECT 22.200 42.245 22.620 42.445 ;
        RECT 22.795 42.275 23.490 42.445 ;
        RECT 22.795 42.025 22.965 42.275 ;
        RECT 23.660 42.075 23.835 42.635 ;
        RECT 23.605 42.025 23.835 42.075 ;
        RECT 19.585 41.055 20.120 41.675 ;
        RECT 20.530 41.855 22.965 42.025 ;
        RECT 20.530 41.055 20.860 41.855 ;
        RECT 21.030 40.885 21.360 41.685 ;
        RECT 21.660 41.055 21.990 41.855 ;
        RECT 22.635 40.885 22.885 41.685 ;
        RECT 23.155 40.885 23.325 42.025 ;
        RECT 23.495 41.055 23.835 42.025 ;
        RECT 24.010 41.895 24.360 42.545 ;
        RECT 24.530 41.725 24.760 42.715 ;
        RECT 24.095 41.555 24.760 41.725 ;
        RECT 24.095 41.055 24.265 41.555 ;
        RECT 24.435 40.885 24.765 41.385 ;
        RECT 24.935 41.055 25.120 43.175 ;
        RECT 25.375 42.975 25.625 43.435 ;
        RECT 25.795 42.985 26.130 43.155 ;
        RECT 26.325 42.985 27.000 43.155 ;
        RECT 25.795 42.845 25.965 42.985 ;
        RECT 25.290 41.855 25.570 42.805 ;
        RECT 25.740 42.715 25.965 42.845 ;
        RECT 25.740 41.610 25.910 42.715 ;
        RECT 26.135 42.565 26.660 42.785 ;
        RECT 26.080 41.800 26.320 42.395 ;
        RECT 26.490 41.865 26.660 42.565 ;
        RECT 26.830 42.205 27.000 42.985 ;
        RECT 27.320 42.935 27.690 43.435 ;
        RECT 27.870 42.985 28.275 43.155 ;
        RECT 28.445 42.985 29.230 43.155 ;
        RECT 27.870 42.755 28.040 42.985 ;
        RECT 27.210 42.455 28.040 42.755 ;
        RECT 28.425 42.485 28.890 42.815 ;
        RECT 27.210 42.425 27.410 42.455 ;
        RECT 27.530 42.205 27.700 42.275 ;
        RECT 26.830 42.035 27.700 42.205 ;
        RECT 27.190 41.945 27.700 42.035 ;
        RECT 25.740 41.480 26.045 41.610 ;
        RECT 26.490 41.500 27.020 41.865 ;
        RECT 25.360 40.885 25.625 41.345 ;
        RECT 25.795 41.055 26.045 41.480 ;
        RECT 27.190 41.330 27.360 41.945 ;
        RECT 26.255 41.160 27.360 41.330 ;
        RECT 27.530 40.885 27.700 41.685 ;
        RECT 27.870 41.385 28.040 42.455 ;
        RECT 28.210 41.555 28.400 42.275 ;
        RECT 28.570 41.525 28.890 42.485 ;
        RECT 29.060 42.525 29.230 42.985 ;
        RECT 29.505 42.905 29.715 43.435 ;
        RECT 29.975 42.695 30.305 43.220 ;
        RECT 30.475 42.825 30.645 43.435 ;
        RECT 30.815 42.780 31.145 43.215 ;
        RECT 30.815 42.695 31.195 42.780 ;
        RECT 31.365 42.710 31.655 43.435 ;
        RECT 31.885 42.975 32.130 43.435 ;
        RECT 30.105 42.525 30.305 42.695 ;
        RECT 30.970 42.655 31.195 42.695 ;
        RECT 29.060 42.195 29.935 42.525 ;
        RECT 30.105 42.195 30.855 42.525 ;
        RECT 27.870 41.055 28.120 41.385 ;
        RECT 29.060 41.355 29.230 42.195 ;
        RECT 30.105 41.990 30.295 42.195 ;
        RECT 31.025 42.075 31.195 42.655 ;
        RECT 31.825 42.195 32.140 42.805 ;
        RECT 32.310 42.445 32.560 43.255 ;
        RECT 32.730 42.910 32.990 43.435 ;
        RECT 33.160 42.785 33.420 43.240 ;
        RECT 33.590 42.955 33.850 43.435 ;
        RECT 34.020 42.785 34.280 43.240 ;
        RECT 34.450 42.955 34.710 43.435 ;
        RECT 34.880 42.785 35.140 43.240 ;
        RECT 35.310 42.955 35.570 43.435 ;
        RECT 35.740 42.785 36.000 43.240 ;
        RECT 36.170 42.955 36.470 43.435 ;
        RECT 33.160 42.615 36.470 42.785 ;
        RECT 32.310 42.195 35.330 42.445 ;
        RECT 30.980 42.025 31.195 42.075 ;
        RECT 29.400 41.615 30.295 41.990 ;
        RECT 30.805 41.945 31.195 42.025 ;
        RECT 28.345 41.185 29.230 41.355 ;
        RECT 29.410 40.885 29.725 41.385 ;
        RECT 29.955 41.055 30.295 41.615 ;
        RECT 30.465 40.885 30.635 41.895 ;
        RECT 30.805 41.100 31.135 41.945 ;
        RECT 31.365 40.885 31.655 42.050 ;
        RECT 31.835 40.885 32.130 41.995 ;
        RECT 32.310 41.060 32.560 42.195 ;
        RECT 35.500 42.025 36.470 42.615 ;
        RECT 32.730 40.885 32.990 41.995 ;
        RECT 33.160 41.785 36.470 42.025 ;
        RECT 36.885 42.695 37.270 43.265 ;
        RECT 37.440 42.975 37.765 43.435 ;
        RECT 38.285 42.805 38.565 43.265 ;
        RECT 36.885 42.025 37.165 42.695 ;
        RECT 37.440 42.635 38.565 42.805 ;
        RECT 37.440 42.525 37.890 42.635 ;
        RECT 37.335 42.195 37.890 42.525 ;
        RECT 38.755 42.465 39.155 43.265 ;
        RECT 39.555 42.975 39.825 43.435 ;
        RECT 39.995 42.805 40.280 43.265 ;
        RECT 33.160 41.060 33.420 41.785 ;
        RECT 33.590 40.885 33.850 41.615 ;
        RECT 34.020 41.060 34.280 41.785 ;
        RECT 34.450 40.885 34.710 41.615 ;
        RECT 34.880 41.060 35.140 41.785 ;
        RECT 35.310 40.885 35.570 41.615 ;
        RECT 35.740 41.060 36.000 41.785 ;
        RECT 36.170 40.885 36.465 41.615 ;
        RECT 36.885 41.055 37.270 42.025 ;
        RECT 37.440 41.735 37.890 42.195 ;
        RECT 38.060 41.905 39.155 42.465 ;
        RECT 37.440 41.515 38.565 41.735 ;
        RECT 37.440 40.885 37.765 41.345 ;
        RECT 38.285 41.055 38.565 41.515 ;
        RECT 38.755 41.055 39.155 41.905 ;
        RECT 39.325 42.635 40.280 42.805 ;
        RECT 40.565 42.935 40.865 43.265 ;
        RECT 41.035 42.955 41.310 43.435 ;
        RECT 39.325 41.735 39.535 42.635 ;
        RECT 39.705 41.905 40.395 42.465 ;
        RECT 40.565 42.025 40.735 42.935 ;
        RECT 41.490 42.785 41.785 43.175 ;
        RECT 41.955 42.955 42.210 43.435 ;
        RECT 42.385 42.785 42.645 43.175 ;
        RECT 42.815 42.955 43.095 43.435 ;
        RECT 40.905 42.195 41.255 42.765 ;
        RECT 41.490 42.615 43.140 42.785 ;
        RECT 43.330 42.615 43.605 43.435 ;
        RECT 43.775 42.795 44.105 43.265 ;
        RECT 44.275 42.965 44.445 43.435 ;
        RECT 44.615 42.795 44.945 43.265 ;
        RECT 45.115 42.965 45.825 43.435 ;
        RECT 45.995 42.795 46.325 43.265 ;
        RECT 46.495 42.965 46.785 43.435 ;
        RECT 43.775 42.615 46.835 42.795 ;
        RECT 41.425 42.275 42.565 42.445 ;
        RECT 41.425 42.025 41.595 42.275 ;
        RECT 42.735 42.105 43.140 42.615 ;
        RECT 43.375 42.235 44.205 42.445 ;
        RECT 44.375 42.235 45.425 42.445 ;
        RECT 45.615 42.235 46.205 42.445 ;
        RECT 40.565 41.855 41.595 42.025 ;
        RECT 42.385 41.935 43.140 42.105 ;
        RECT 39.325 41.515 40.280 41.735 ;
        RECT 39.555 40.885 39.825 41.345 ;
        RECT 39.995 41.055 40.280 41.515 ;
        RECT 40.565 41.055 40.875 41.855 ;
        RECT 42.385 41.685 42.645 41.935 ;
        RECT 43.390 41.895 45.325 42.065 ;
        RECT 45.615 41.895 45.880 42.235 ;
        RECT 46.375 42.065 46.835 42.615 ;
        RECT 47.005 42.665 48.675 43.435 ;
        RECT 48.855 42.945 49.185 43.435 ;
        RECT 49.355 42.840 49.975 43.265 ;
        RECT 47.005 42.145 47.755 42.665 ;
        RECT 46.075 41.895 46.835 42.065 ;
        RECT 47.925 41.975 48.675 42.495 ;
        RECT 48.845 42.195 49.185 42.775 ;
        RECT 49.355 42.505 49.715 42.840 ;
        RECT 50.435 42.745 50.765 43.435 ;
        RECT 52.635 43.055 53.805 43.265 ;
        RECT 52.635 43.035 52.965 43.055 ;
        RECT 52.525 42.615 53.385 42.865 ;
        RECT 53.555 42.805 53.805 43.055 ;
        RECT 53.975 42.975 54.145 43.435 ;
        RECT 54.315 42.805 54.655 43.265 ;
        RECT 53.555 42.635 54.655 42.805 ;
        RECT 54.825 42.665 56.495 43.435 ;
        RECT 57.125 42.710 57.415 43.435 ;
        RECT 57.585 42.665 59.255 43.435 ;
        RECT 59.430 42.965 59.760 43.435 ;
        RECT 59.930 42.795 60.155 43.240 ;
        RECT 60.325 42.910 60.620 43.435 ;
        RECT 61.325 42.975 61.570 43.435 ;
        RECT 49.355 42.225 50.775 42.505 ;
        RECT 41.045 40.885 41.355 41.685 ;
        RECT 41.525 41.515 42.645 41.685 ;
        RECT 41.525 41.055 41.785 41.515 ;
        RECT 41.955 40.885 42.210 41.345 ;
        RECT 42.385 41.055 42.645 41.515 ;
        RECT 42.815 40.885 43.100 41.755 ;
        RECT 43.390 41.055 43.645 41.895 ;
        RECT 43.815 40.885 44.065 41.725 ;
        RECT 44.235 41.055 44.485 41.895 ;
        RECT 44.655 41.225 44.905 41.725 ;
        RECT 45.075 41.395 45.325 41.895 ;
        RECT 45.655 41.225 45.865 41.725 ;
        RECT 46.075 41.395 46.285 41.895 ;
        RECT 46.455 41.225 46.705 41.725 ;
        RECT 44.655 41.055 46.705 41.225 ;
        RECT 47.005 40.885 48.675 41.975 ;
        RECT 48.855 40.885 49.185 42.025 ;
        RECT 49.355 41.055 49.715 42.225 ;
        RECT 49.915 40.885 50.245 42.055 ;
        RECT 50.445 41.055 50.775 42.225 ;
        RECT 50.975 40.885 51.305 42.055 ;
        RECT 52.525 42.025 52.805 42.615 ;
        RECT 52.975 42.195 53.725 42.445 ;
        RECT 53.895 42.195 54.655 42.445 ;
        RECT 54.825 42.145 55.575 42.665 ;
        RECT 52.525 41.855 54.225 42.025 ;
        RECT 52.630 40.885 52.885 41.685 ;
        RECT 53.055 41.055 53.385 41.855 ;
        RECT 53.555 40.885 53.725 41.685 ;
        RECT 53.895 41.055 54.225 41.855 ;
        RECT 54.395 40.885 54.655 42.025 ;
        RECT 55.745 41.975 56.495 42.495 ;
        RECT 57.585 42.145 58.335 42.665 ;
        RECT 59.425 42.625 60.155 42.795 ;
        RECT 54.825 40.885 56.495 41.975 ;
        RECT 57.125 40.885 57.415 42.050 ;
        RECT 58.505 41.975 59.255 42.495 ;
        RECT 57.585 40.885 59.255 41.975 ;
        RECT 59.425 42.060 59.705 42.625 ;
        RECT 59.875 42.230 61.095 42.455 ;
        RECT 61.265 42.195 61.580 42.805 ;
        RECT 61.750 42.445 62.000 43.255 ;
        RECT 62.170 42.910 62.430 43.435 ;
        RECT 62.600 42.785 62.860 43.240 ;
        RECT 63.030 42.955 63.290 43.435 ;
        RECT 63.460 42.785 63.720 43.240 ;
        RECT 63.890 42.955 64.150 43.435 ;
        RECT 64.320 42.785 64.580 43.240 ;
        RECT 64.750 42.955 65.010 43.435 ;
        RECT 65.180 42.785 65.440 43.240 ;
        RECT 65.610 42.955 65.910 43.435 ;
        RECT 66.415 42.885 66.585 43.175 ;
        RECT 66.755 43.055 67.085 43.435 ;
        RECT 62.600 42.615 65.910 42.785 ;
        RECT 66.415 42.715 67.080 42.885 ;
        RECT 61.750 42.195 64.770 42.445 ;
        RECT 59.425 41.890 61.025 42.060 ;
        RECT 59.485 40.885 59.740 41.720 ;
        RECT 59.910 41.085 60.170 41.890 ;
        RECT 60.340 40.885 60.600 41.720 ;
        RECT 60.770 41.085 61.025 41.890 ;
        RECT 61.275 40.885 61.570 41.995 ;
        RECT 61.750 41.060 62.000 42.195 ;
        RECT 64.940 42.025 65.910 42.615 ;
        RECT 62.170 40.885 62.430 41.995 ;
        RECT 62.600 41.785 65.910 42.025 ;
        RECT 66.330 41.895 66.680 42.545 ;
        RECT 62.600 41.060 62.860 41.785 ;
        RECT 63.030 40.885 63.290 41.615 ;
        RECT 63.460 41.060 63.720 41.785 ;
        RECT 63.890 40.885 64.150 41.615 ;
        RECT 64.320 41.060 64.580 41.785 ;
        RECT 64.750 40.885 65.010 41.615 ;
        RECT 65.180 41.060 65.440 41.785 ;
        RECT 66.850 41.725 67.080 42.715 ;
        RECT 65.610 40.885 65.905 41.615 ;
        RECT 66.415 41.555 67.080 41.725 ;
        RECT 66.415 41.055 66.585 41.555 ;
        RECT 66.755 40.885 67.085 41.385 ;
        RECT 67.255 41.055 67.440 43.175 ;
        RECT 67.695 42.975 67.945 43.435 ;
        RECT 68.115 42.985 68.450 43.155 ;
        RECT 68.645 42.985 69.320 43.155 ;
        RECT 68.115 42.845 68.285 42.985 ;
        RECT 67.610 41.855 67.890 42.805 ;
        RECT 68.060 42.715 68.285 42.845 ;
        RECT 68.060 41.610 68.230 42.715 ;
        RECT 68.455 42.565 68.980 42.785 ;
        RECT 68.400 41.800 68.640 42.395 ;
        RECT 68.810 41.865 68.980 42.565 ;
        RECT 69.150 42.205 69.320 42.985 ;
        RECT 69.640 42.935 70.010 43.435 ;
        RECT 70.190 42.985 70.595 43.155 ;
        RECT 70.765 42.985 71.550 43.155 ;
        RECT 70.190 42.755 70.360 42.985 ;
        RECT 69.530 42.455 70.360 42.755 ;
        RECT 70.745 42.485 71.210 42.815 ;
        RECT 69.530 42.425 69.730 42.455 ;
        RECT 69.850 42.205 70.020 42.275 ;
        RECT 69.150 42.035 70.020 42.205 ;
        RECT 69.510 41.945 70.020 42.035 ;
        RECT 68.060 41.480 68.365 41.610 ;
        RECT 68.810 41.500 69.340 41.865 ;
        RECT 67.680 40.885 67.945 41.345 ;
        RECT 68.115 41.055 68.365 41.480 ;
        RECT 69.510 41.330 69.680 41.945 ;
        RECT 68.575 41.160 69.680 41.330 ;
        RECT 69.850 40.885 70.020 41.685 ;
        RECT 70.190 41.385 70.360 42.455 ;
        RECT 70.530 41.555 70.720 42.275 ;
        RECT 70.890 41.525 71.210 42.485 ;
        RECT 71.380 42.525 71.550 42.985 ;
        RECT 71.825 42.905 72.035 43.435 ;
        RECT 72.295 42.695 72.625 43.220 ;
        RECT 72.795 42.825 72.965 43.435 ;
        RECT 73.135 42.780 73.465 43.215 ;
        RECT 73.685 42.890 79.030 43.435 ;
        RECT 73.135 42.695 73.515 42.780 ;
        RECT 72.425 42.525 72.625 42.695 ;
        RECT 73.290 42.655 73.515 42.695 ;
        RECT 71.380 42.195 72.255 42.525 ;
        RECT 72.425 42.195 73.175 42.525 ;
        RECT 70.190 41.055 70.440 41.385 ;
        RECT 71.380 41.355 71.550 42.195 ;
        RECT 72.425 41.990 72.615 42.195 ;
        RECT 73.345 42.075 73.515 42.655 ;
        RECT 73.300 42.025 73.515 42.075 ;
        RECT 75.270 42.060 75.610 42.890 ;
        RECT 79.205 42.665 80.875 43.435 ;
        RECT 81.135 42.885 81.305 43.265 ;
        RECT 81.520 43.055 81.850 43.435 ;
        RECT 81.135 42.715 81.850 42.885 ;
        RECT 71.720 41.615 72.615 41.990 ;
        RECT 73.125 41.945 73.515 42.025 ;
        RECT 70.665 41.185 71.550 41.355 ;
        RECT 71.730 40.885 72.045 41.385 ;
        RECT 72.275 41.055 72.615 41.615 ;
        RECT 72.785 40.885 72.955 41.895 ;
        RECT 73.125 41.100 73.455 41.945 ;
        RECT 77.090 41.320 77.440 42.570 ;
        RECT 79.205 42.145 79.955 42.665 ;
        RECT 80.125 41.975 80.875 42.495 ;
        RECT 81.045 42.165 81.400 42.535 ;
        RECT 81.680 42.525 81.850 42.715 ;
        RECT 82.020 42.690 82.275 43.265 ;
        RECT 81.680 42.195 81.935 42.525 ;
        RECT 81.680 41.985 81.850 42.195 ;
        RECT 73.685 40.885 79.030 41.320 ;
        RECT 79.205 40.885 80.875 41.975 ;
        RECT 81.135 41.815 81.850 41.985 ;
        RECT 82.105 41.960 82.275 42.690 ;
        RECT 82.450 42.595 82.710 43.435 ;
        RECT 82.885 42.685 84.095 43.435 ;
        RECT 81.135 41.055 81.305 41.815 ;
        RECT 81.520 40.885 81.850 41.645 ;
        RECT 82.020 41.055 82.275 41.960 ;
        RECT 82.450 40.885 82.710 42.035 ;
        RECT 82.885 41.975 83.405 42.515 ;
        RECT 83.575 42.145 84.095 42.685 ;
        RECT 82.885 40.885 84.095 41.975 ;
        RECT 5.520 40.715 84.180 40.885 ;
        RECT 5.605 39.625 6.815 40.715 ;
        RECT 7.075 40.045 7.245 40.545 ;
        RECT 7.415 40.215 7.745 40.715 ;
        RECT 7.075 39.875 7.740 40.045 ;
        RECT 5.605 38.915 6.125 39.455 ;
        RECT 6.295 39.085 6.815 39.625 ;
        RECT 6.990 39.055 7.340 39.705 ;
        RECT 5.605 38.165 6.815 38.915 ;
        RECT 7.510 38.885 7.740 39.875 ;
        RECT 7.075 38.715 7.740 38.885 ;
        RECT 7.075 38.425 7.245 38.715 ;
        RECT 7.415 38.165 7.745 38.545 ;
        RECT 7.915 38.425 8.100 40.545 ;
        RECT 8.340 40.255 8.605 40.715 ;
        RECT 8.775 40.120 9.025 40.545 ;
        RECT 9.235 40.270 10.340 40.440 ;
        RECT 8.720 39.990 9.025 40.120 ;
        RECT 8.270 38.795 8.550 39.745 ;
        RECT 8.720 38.885 8.890 39.990 ;
        RECT 9.060 39.205 9.300 39.800 ;
        RECT 9.470 39.735 10.000 40.100 ;
        RECT 9.470 39.035 9.640 39.735 ;
        RECT 10.170 39.655 10.340 40.270 ;
        RECT 10.510 39.915 10.680 40.715 ;
        RECT 10.850 40.215 11.100 40.545 ;
        RECT 11.325 40.245 12.210 40.415 ;
        RECT 10.170 39.565 10.680 39.655 ;
        RECT 8.720 38.755 8.945 38.885 ;
        RECT 9.115 38.815 9.640 39.035 ;
        RECT 9.810 39.395 10.680 39.565 ;
        RECT 8.355 38.165 8.605 38.625 ;
        RECT 8.775 38.615 8.945 38.755 ;
        RECT 9.810 38.615 9.980 39.395 ;
        RECT 10.510 39.325 10.680 39.395 ;
        RECT 10.190 39.145 10.390 39.175 ;
        RECT 10.850 39.145 11.020 40.215 ;
        RECT 11.190 39.325 11.380 40.045 ;
        RECT 10.190 38.845 11.020 39.145 ;
        RECT 11.550 39.115 11.870 40.075 ;
        RECT 8.775 38.445 9.110 38.615 ;
        RECT 9.305 38.445 9.980 38.615 ;
        RECT 10.300 38.165 10.670 38.665 ;
        RECT 10.850 38.615 11.020 38.845 ;
        RECT 11.405 38.785 11.870 39.115 ;
        RECT 12.040 39.405 12.210 40.245 ;
        RECT 12.390 40.215 12.705 40.715 ;
        RECT 12.935 39.985 13.275 40.545 ;
        RECT 12.380 39.610 13.275 39.985 ;
        RECT 13.445 39.705 13.615 40.715 ;
        RECT 13.085 39.405 13.275 39.610 ;
        RECT 13.785 39.655 14.115 40.500 ;
        RECT 13.785 39.575 14.175 39.655 ;
        RECT 13.960 39.525 14.175 39.575 ;
        RECT 14.350 39.565 14.610 40.715 ;
        RECT 14.785 39.640 15.040 40.545 ;
        RECT 15.210 39.955 15.540 40.715 ;
        RECT 15.755 39.785 15.925 40.545 ;
        RECT 12.040 39.075 12.915 39.405 ;
        RECT 13.085 39.075 13.835 39.405 ;
        RECT 12.040 38.615 12.210 39.075 ;
        RECT 13.085 38.905 13.285 39.075 ;
        RECT 14.005 38.945 14.175 39.525 ;
        RECT 13.950 38.905 14.175 38.945 ;
        RECT 10.850 38.445 11.255 38.615 ;
        RECT 11.425 38.445 12.210 38.615 ;
        RECT 12.485 38.165 12.695 38.695 ;
        RECT 12.955 38.380 13.285 38.905 ;
        RECT 13.795 38.820 14.175 38.905 ;
        RECT 13.455 38.165 13.625 38.775 ;
        RECT 13.795 38.385 14.125 38.820 ;
        RECT 14.350 38.165 14.610 39.005 ;
        RECT 14.785 38.910 14.955 39.640 ;
        RECT 15.210 39.615 15.925 39.785 ;
        RECT 16.185 39.625 17.855 40.715 ;
        RECT 15.210 39.405 15.380 39.615 ;
        RECT 15.125 39.075 15.380 39.405 ;
        RECT 14.785 38.335 15.040 38.910 ;
        RECT 15.210 38.885 15.380 39.075 ;
        RECT 15.660 39.065 16.015 39.435 ;
        RECT 16.185 38.935 16.935 39.455 ;
        RECT 17.105 39.105 17.855 39.625 ;
        RECT 18.485 39.550 18.775 40.715 ;
        RECT 18.985 39.765 19.275 40.535 ;
        RECT 19.845 40.175 20.105 40.535 ;
        RECT 20.275 40.345 20.605 40.715 ;
        RECT 20.775 40.175 21.035 40.535 ;
        RECT 19.845 39.945 21.035 40.175 ;
        RECT 21.225 39.995 21.555 40.715 ;
        RECT 21.725 39.765 21.990 40.535 ;
        RECT 22.270 40.255 22.440 40.715 ;
        RECT 22.610 40.085 22.940 40.545 ;
        RECT 18.985 39.585 21.480 39.765 ;
        RECT 18.955 39.075 19.225 39.405 ;
        RECT 19.405 39.075 19.840 39.405 ;
        RECT 20.020 39.075 20.595 39.405 ;
        RECT 20.775 39.075 21.055 39.405 ;
        RECT 15.210 38.715 15.925 38.885 ;
        RECT 15.210 38.165 15.540 38.545 ;
        RECT 15.755 38.335 15.925 38.715 ;
        RECT 16.185 38.165 17.855 38.935 ;
        RECT 21.255 38.895 21.480 39.585 ;
        RECT 18.485 38.165 18.775 38.890 ;
        RECT 18.995 38.705 21.480 38.895 ;
        RECT 18.995 38.345 19.220 38.705 ;
        RECT 19.400 38.165 19.730 38.535 ;
        RECT 19.910 38.345 20.165 38.705 ;
        RECT 20.730 38.165 21.475 38.535 ;
        RECT 21.655 38.345 21.990 39.765 ;
        RECT 22.165 39.915 22.940 40.085 ;
        RECT 23.110 39.915 23.280 40.715 ;
        RECT 22.165 38.905 22.595 39.915 ;
        RECT 23.865 39.745 24.225 39.920 ;
        RECT 22.765 39.575 24.225 39.745 ;
        RECT 24.505 39.575 24.735 40.715 ;
        RECT 22.765 39.075 22.935 39.575 ;
        RECT 22.165 38.735 22.860 38.905 ;
        RECT 23.105 38.845 23.515 39.405 ;
        RECT 22.190 38.165 22.520 38.565 ;
        RECT 22.690 38.465 22.860 38.735 ;
        RECT 23.685 38.675 23.865 39.575 ;
        RECT 24.905 39.565 25.235 40.545 ;
        RECT 25.405 39.575 25.615 40.715 ;
        RECT 25.845 40.280 31.190 40.715 ;
        RECT 24.035 39.355 24.230 39.405 ;
        RECT 24.035 39.185 24.235 39.355 ;
        RECT 24.035 38.845 24.230 39.185 ;
        RECT 24.485 39.155 24.815 39.405 ;
        RECT 23.030 38.165 23.345 38.675 ;
        RECT 23.575 38.335 23.865 38.675 ;
        RECT 24.035 38.165 24.275 38.675 ;
        RECT 24.505 38.165 24.735 38.985 ;
        RECT 24.985 38.965 25.235 39.565 ;
        RECT 24.905 38.335 25.235 38.965 ;
        RECT 25.405 38.165 25.615 38.985 ;
        RECT 27.430 38.710 27.770 39.540 ;
        RECT 29.250 39.030 29.600 40.280 ;
        RECT 31.830 39.575 32.165 40.545 ;
        RECT 32.335 39.575 32.505 40.715 ;
        RECT 32.675 40.375 34.705 40.545 ;
        RECT 31.830 38.905 32.000 39.575 ;
        RECT 32.675 39.405 32.845 40.375 ;
        RECT 32.170 39.075 32.425 39.405 ;
        RECT 32.650 39.075 32.845 39.405 ;
        RECT 33.015 40.035 34.140 40.205 ;
        RECT 32.255 38.905 32.425 39.075 ;
        RECT 33.015 38.905 33.185 40.035 ;
        RECT 25.845 38.165 31.190 38.710 ;
        RECT 31.830 38.335 32.085 38.905 ;
        RECT 32.255 38.735 33.185 38.905 ;
        RECT 33.355 39.695 34.365 39.865 ;
        RECT 33.355 38.895 33.525 39.695 ;
        RECT 33.730 39.355 34.005 39.495 ;
        RECT 33.725 39.185 34.005 39.355 ;
        RECT 33.010 38.700 33.185 38.735 ;
        RECT 32.255 38.165 32.585 38.565 ;
        RECT 33.010 38.335 33.540 38.700 ;
        RECT 33.730 38.335 34.005 39.185 ;
        RECT 34.175 38.335 34.365 39.695 ;
        RECT 34.535 39.710 34.705 40.375 ;
        RECT 34.875 39.955 35.045 40.715 ;
        RECT 35.280 39.955 35.795 40.365 ;
        RECT 34.535 39.520 35.285 39.710 ;
        RECT 35.455 39.145 35.795 39.955 ;
        RECT 36.975 40.045 37.145 40.545 ;
        RECT 37.315 40.215 37.645 40.715 ;
        RECT 36.975 39.875 37.640 40.045 ;
        RECT 34.565 38.975 35.795 39.145 ;
        RECT 36.890 39.055 37.240 39.705 ;
        RECT 34.545 38.165 35.055 38.700 ;
        RECT 35.275 38.370 35.520 38.975 ;
        RECT 37.410 38.885 37.640 39.875 ;
        RECT 36.975 38.715 37.640 38.885 ;
        RECT 36.975 38.425 37.145 38.715 ;
        RECT 37.315 38.165 37.645 38.545 ;
        RECT 37.815 38.425 38.000 40.545 ;
        RECT 38.240 40.255 38.505 40.715 ;
        RECT 38.675 40.120 38.925 40.545 ;
        RECT 39.135 40.270 40.240 40.440 ;
        RECT 38.620 39.990 38.925 40.120 ;
        RECT 38.170 38.795 38.450 39.745 ;
        RECT 38.620 38.885 38.790 39.990 ;
        RECT 38.960 39.205 39.200 39.800 ;
        RECT 39.370 39.735 39.900 40.100 ;
        RECT 39.370 39.035 39.540 39.735 ;
        RECT 40.070 39.655 40.240 40.270 ;
        RECT 40.410 39.915 40.580 40.715 ;
        RECT 40.750 40.215 41.000 40.545 ;
        RECT 41.225 40.245 42.110 40.415 ;
        RECT 40.070 39.565 40.580 39.655 ;
        RECT 38.620 38.755 38.845 38.885 ;
        RECT 39.015 38.815 39.540 39.035 ;
        RECT 39.710 39.395 40.580 39.565 ;
        RECT 38.255 38.165 38.505 38.625 ;
        RECT 38.675 38.615 38.845 38.755 ;
        RECT 39.710 38.615 39.880 39.395 ;
        RECT 40.410 39.325 40.580 39.395 ;
        RECT 40.090 39.145 40.290 39.175 ;
        RECT 40.750 39.145 40.920 40.215 ;
        RECT 41.090 39.325 41.280 40.045 ;
        RECT 40.090 38.845 40.920 39.145 ;
        RECT 41.450 39.115 41.770 40.075 ;
        RECT 38.675 38.445 39.010 38.615 ;
        RECT 39.205 38.445 39.880 38.615 ;
        RECT 40.200 38.165 40.570 38.665 ;
        RECT 40.750 38.615 40.920 38.845 ;
        RECT 41.305 38.785 41.770 39.115 ;
        RECT 41.940 39.405 42.110 40.245 ;
        RECT 42.290 40.215 42.605 40.715 ;
        RECT 42.835 39.985 43.175 40.545 ;
        RECT 42.280 39.610 43.175 39.985 ;
        RECT 43.345 39.705 43.515 40.715 ;
        RECT 42.985 39.405 43.175 39.610 ;
        RECT 43.685 39.655 44.015 40.500 ;
        RECT 43.685 39.575 44.075 39.655 ;
        RECT 43.860 39.525 44.075 39.575 ;
        RECT 44.245 39.550 44.535 40.715 ;
        RECT 44.745 39.575 44.975 40.715 ;
        RECT 45.145 39.565 45.475 40.545 ;
        RECT 45.645 39.575 45.855 40.715 ;
        RECT 46.175 40.045 46.345 40.545 ;
        RECT 46.515 40.215 46.845 40.715 ;
        RECT 46.175 39.875 46.840 40.045 ;
        RECT 41.940 39.075 42.815 39.405 ;
        RECT 42.985 39.075 43.735 39.405 ;
        RECT 41.940 38.615 42.110 39.075 ;
        RECT 42.985 38.905 43.185 39.075 ;
        RECT 43.905 38.945 44.075 39.525 ;
        RECT 44.725 39.155 45.055 39.405 ;
        RECT 43.850 38.905 44.075 38.945 ;
        RECT 40.750 38.445 41.155 38.615 ;
        RECT 41.325 38.445 42.110 38.615 ;
        RECT 42.385 38.165 42.595 38.695 ;
        RECT 42.855 38.380 43.185 38.905 ;
        RECT 43.695 38.820 44.075 38.905 ;
        RECT 43.355 38.165 43.525 38.775 ;
        RECT 43.695 38.385 44.025 38.820 ;
        RECT 44.245 38.165 44.535 38.890 ;
        RECT 44.745 38.165 44.975 38.985 ;
        RECT 45.225 38.965 45.475 39.565 ;
        RECT 46.090 39.055 46.440 39.705 ;
        RECT 45.145 38.335 45.475 38.965 ;
        RECT 45.645 38.165 45.855 38.985 ;
        RECT 46.610 38.885 46.840 39.875 ;
        RECT 46.175 38.715 46.840 38.885 ;
        RECT 46.175 38.425 46.345 38.715 ;
        RECT 46.515 38.165 46.845 38.545 ;
        RECT 47.015 38.425 47.200 40.545 ;
        RECT 47.440 40.255 47.705 40.715 ;
        RECT 47.875 40.120 48.125 40.545 ;
        RECT 48.335 40.270 49.440 40.440 ;
        RECT 47.820 39.990 48.125 40.120 ;
        RECT 47.370 38.795 47.650 39.745 ;
        RECT 47.820 38.885 47.990 39.990 ;
        RECT 48.160 39.205 48.400 39.800 ;
        RECT 48.570 39.735 49.100 40.100 ;
        RECT 48.570 39.035 48.740 39.735 ;
        RECT 49.270 39.655 49.440 40.270 ;
        RECT 49.610 39.915 49.780 40.715 ;
        RECT 49.950 40.215 50.200 40.545 ;
        RECT 50.425 40.245 51.310 40.415 ;
        RECT 49.270 39.565 49.780 39.655 ;
        RECT 47.820 38.755 48.045 38.885 ;
        RECT 48.215 38.815 48.740 39.035 ;
        RECT 48.910 39.395 49.780 39.565 ;
        RECT 47.455 38.165 47.705 38.625 ;
        RECT 47.875 38.615 48.045 38.755 ;
        RECT 48.910 38.615 49.080 39.395 ;
        RECT 49.610 39.325 49.780 39.395 ;
        RECT 49.290 39.145 49.490 39.175 ;
        RECT 49.950 39.145 50.120 40.215 ;
        RECT 50.290 39.325 50.480 40.045 ;
        RECT 49.290 38.845 50.120 39.145 ;
        RECT 50.650 39.115 50.970 40.075 ;
        RECT 47.875 38.445 48.210 38.615 ;
        RECT 48.405 38.445 49.080 38.615 ;
        RECT 49.400 38.165 49.770 38.665 ;
        RECT 49.950 38.615 50.120 38.845 ;
        RECT 50.505 38.785 50.970 39.115 ;
        RECT 51.140 39.405 51.310 40.245 ;
        RECT 51.490 40.215 51.805 40.715 ;
        RECT 52.035 39.985 52.375 40.545 ;
        RECT 51.480 39.610 52.375 39.985 ;
        RECT 52.545 39.705 52.715 40.715 ;
        RECT 52.185 39.405 52.375 39.610 ;
        RECT 52.885 39.655 53.215 40.500 ;
        RECT 54.455 40.045 54.625 40.545 ;
        RECT 54.795 40.215 55.125 40.715 ;
        RECT 54.455 39.875 55.120 40.045 ;
        RECT 52.885 39.575 53.275 39.655 ;
        RECT 53.060 39.525 53.275 39.575 ;
        RECT 51.140 39.075 52.015 39.405 ;
        RECT 52.185 39.075 52.935 39.405 ;
        RECT 51.140 38.615 51.310 39.075 ;
        RECT 52.185 38.905 52.385 39.075 ;
        RECT 53.105 38.945 53.275 39.525 ;
        RECT 54.370 39.055 54.720 39.705 ;
        RECT 53.050 38.905 53.275 38.945 ;
        RECT 49.950 38.445 50.355 38.615 ;
        RECT 50.525 38.445 51.310 38.615 ;
        RECT 51.585 38.165 51.795 38.695 ;
        RECT 52.055 38.380 52.385 38.905 ;
        RECT 52.895 38.820 53.275 38.905 ;
        RECT 54.890 38.885 55.120 39.875 ;
        RECT 52.555 38.165 52.725 38.775 ;
        RECT 52.895 38.385 53.225 38.820 ;
        RECT 54.455 38.715 55.120 38.885 ;
        RECT 54.455 38.425 54.625 38.715 ;
        RECT 54.795 38.165 55.125 38.545 ;
        RECT 55.295 38.425 55.480 40.545 ;
        RECT 55.720 40.255 55.985 40.715 ;
        RECT 56.155 40.120 56.405 40.545 ;
        RECT 56.615 40.270 57.720 40.440 ;
        RECT 56.100 39.990 56.405 40.120 ;
        RECT 55.650 38.795 55.930 39.745 ;
        RECT 56.100 38.885 56.270 39.990 ;
        RECT 56.440 39.205 56.680 39.800 ;
        RECT 56.850 39.735 57.380 40.100 ;
        RECT 56.850 39.035 57.020 39.735 ;
        RECT 57.550 39.655 57.720 40.270 ;
        RECT 57.890 39.915 58.060 40.715 ;
        RECT 58.230 40.215 58.480 40.545 ;
        RECT 58.705 40.245 59.590 40.415 ;
        RECT 57.550 39.565 58.060 39.655 ;
        RECT 56.100 38.755 56.325 38.885 ;
        RECT 56.495 38.815 57.020 39.035 ;
        RECT 57.190 39.395 58.060 39.565 ;
        RECT 55.735 38.165 55.985 38.625 ;
        RECT 56.155 38.615 56.325 38.755 ;
        RECT 57.190 38.615 57.360 39.395 ;
        RECT 57.890 39.325 58.060 39.395 ;
        RECT 57.570 39.145 57.770 39.175 ;
        RECT 58.230 39.145 58.400 40.215 ;
        RECT 58.570 39.325 58.760 40.045 ;
        RECT 57.570 38.845 58.400 39.145 ;
        RECT 58.930 39.115 59.250 40.075 ;
        RECT 56.155 38.445 56.490 38.615 ;
        RECT 56.685 38.445 57.360 38.615 ;
        RECT 57.680 38.165 58.050 38.665 ;
        RECT 58.230 38.615 58.400 38.845 ;
        RECT 58.785 38.785 59.250 39.115 ;
        RECT 59.420 39.405 59.590 40.245 ;
        RECT 59.770 40.215 60.085 40.715 ;
        RECT 60.315 39.985 60.655 40.545 ;
        RECT 59.760 39.610 60.655 39.985 ;
        RECT 60.825 39.705 60.995 40.715 ;
        RECT 60.465 39.405 60.655 39.610 ;
        RECT 61.165 39.655 61.495 40.500 ;
        RECT 62.850 39.745 63.180 40.545 ;
        RECT 63.350 39.915 63.680 40.715 ;
        RECT 63.980 39.745 64.310 40.545 ;
        RECT 64.955 39.915 65.205 40.715 ;
        RECT 61.165 39.575 61.555 39.655 ;
        RECT 62.850 39.575 65.285 39.745 ;
        RECT 65.475 39.575 65.645 40.715 ;
        RECT 65.815 39.575 66.155 40.545 ;
        RECT 66.510 39.745 66.900 39.920 ;
        RECT 67.385 39.915 67.715 40.715 ;
        RECT 67.885 39.925 68.420 40.545 ;
        RECT 66.510 39.575 67.935 39.745 ;
        RECT 61.340 39.525 61.555 39.575 ;
        RECT 59.420 39.075 60.295 39.405 ;
        RECT 60.465 39.075 61.215 39.405 ;
        RECT 59.420 38.615 59.590 39.075 ;
        RECT 60.465 38.905 60.665 39.075 ;
        RECT 61.385 38.945 61.555 39.525 ;
        RECT 62.645 39.155 62.995 39.405 ;
        RECT 63.180 38.945 63.350 39.575 ;
        RECT 63.520 39.155 63.850 39.355 ;
        RECT 64.020 39.155 64.350 39.355 ;
        RECT 64.520 39.155 64.940 39.355 ;
        RECT 65.115 39.325 65.285 39.575 ;
        RECT 65.115 39.155 65.810 39.325 ;
        RECT 61.330 38.905 61.555 38.945 ;
        RECT 58.230 38.445 58.635 38.615 ;
        RECT 58.805 38.445 59.590 38.615 ;
        RECT 59.865 38.165 60.075 38.695 ;
        RECT 60.335 38.380 60.665 38.905 ;
        RECT 61.175 38.820 61.555 38.905 ;
        RECT 60.835 38.165 61.005 38.775 ;
        RECT 61.175 38.385 61.505 38.820 ;
        RECT 62.850 38.335 63.350 38.945 ;
        RECT 63.980 38.815 65.205 38.985 ;
        RECT 65.980 38.965 66.155 39.575 ;
        RECT 63.980 38.335 64.310 38.815 ;
        RECT 64.480 38.165 64.705 38.625 ;
        RECT 64.875 38.335 65.205 38.815 ;
        RECT 65.395 38.165 65.645 38.965 ;
        RECT 65.815 38.335 66.155 38.965 ;
        RECT 66.385 38.845 66.740 39.405 ;
        RECT 66.910 38.675 67.080 39.575 ;
        RECT 67.250 38.845 67.515 39.405 ;
        RECT 67.765 39.075 67.935 39.575 ;
        RECT 68.105 38.905 68.420 39.925 ;
        RECT 68.625 39.625 69.835 40.715 ;
        RECT 66.490 38.165 66.730 38.675 ;
        RECT 66.910 38.345 67.190 38.675 ;
        RECT 67.420 38.165 67.635 38.675 ;
        RECT 67.805 38.335 68.420 38.905 ;
        RECT 68.625 38.915 69.145 39.455 ;
        RECT 69.315 39.085 69.835 39.625 ;
        RECT 70.005 39.550 70.295 40.715 ;
        RECT 70.555 40.045 70.725 40.545 ;
        RECT 70.895 40.215 71.225 40.715 ;
        RECT 70.555 39.875 71.220 40.045 ;
        RECT 70.470 39.055 70.820 39.705 ;
        RECT 68.625 38.165 69.835 38.915 ;
        RECT 70.005 38.165 70.295 38.890 ;
        RECT 70.990 38.885 71.220 39.875 ;
        RECT 70.555 38.715 71.220 38.885 ;
        RECT 70.555 38.425 70.725 38.715 ;
        RECT 70.895 38.165 71.225 38.545 ;
        RECT 71.395 38.425 71.580 40.545 ;
        RECT 71.820 40.255 72.085 40.715 ;
        RECT 72.255 40.120 72.505 40.545 ;
        RECT 72.715 40.270 73.820 40.440 ;
        RECT 72.200 39.990 72.505 40.120 ;
        RECT 71.750 38.795 72.030 39.745 ;
        RECT 72.200 38.885 72.370 39.990 ;
        RECT 72.540 39.205 72.780 39.800 ;
        RECT 72.950 39.735 73.480 40.100 ;
        RECT 72.950 39.035 73.120 39.735 ;
        RECT 73.650 39.655 73.820 40.270 ;
        RECT 73.990 39.915 74.160 40.715 ;
        RECT 74.330 40.215 74.580 40.545 ;
        RECT 74.805 40.245 75.690 40.415 ;
        RECT 73.650 39.565 74.160 39.655 ;
        RECT 72.200 38.755 72.425 38.885 ;
        RECT 72.595 38.815 73.120 39.035 ;
        RECT 73.290 39.395 74.160 39.565 ;
        RECT 71.835 38.165 72.085 38.625 ;
        RECT 72.255 38.615 72.425 38.755 ;
        RECT 73.290 38.615 73.460 39.395 ;
        RECT 73.990 39.325 74.160 39.395 ;
        RECT 73.670 39.145 73.870 39.175 ;
        RECT 74.330 39.145 74.500 40.215 ;
        RECT 74.670 39.325 74.860 40.045 ;
        RECT 73.670 38.845 74.500 39.145 ;
        RECT 75.030 39.115 75.350 40.075 ;
        RECT 72.255 38.445 72.590 38.615 ;
        RECT 72.785 38.445 73.460 38.615 ;
        RECT 73.780 38.165 74.150 38.665 ;
        RECT 74.330 38.615 74.500 38.845 ;
        RECT 74.885 38.785 75.350 39.115 ;
        RECT 75.520 39.405 75.690 40.245 ;
        RECT 75.870 40.215 76.185 40.715 ;
        RECT 76.415 39.985 76.755 40.545 ;
        RECT 75.860 39.610 76.755 39.985 ;
        RECT 76.925 39.705 77.095 40.715 ;
        RECT 76.565 39.405 76.755 39.610 ;
        RECT 77.265 39.655 77.595 40.500 ;
        RECT 77.265 39.575 77.655 39.655 ;
        RECT 77.825 39.625 81.335 40.715 ;
        RECT 81.505 39.625 82.715 40.715 ;
        RECT 77.440 39.525 77.655 39.575 ;
        RECT 75.520 39.075 76.395 39.405 ;
        RECT 76.565 39.075 77.315 39.405 ;
        RECT 75.520 38.615 75.690 39.075 ;
        RECT 76.565 38.905 76.765 39.075 ;
        RECT 77.485 38.945 77.655 39.525 ;
        RECT 77.430 38.905 77.655 38.945 ;
        RECT 74.330 38.445 74.735 38.615 ;
        RECT 74.905 38.445 75.690 38.615 ;
        RECT 75.965 38.165 76.175 38.695 ;
        RECT 76.435 38.380 76.765 38.905 ;
        RECT 77.275 38.820 77.655 38.905 ;
        RECT 77.825 38.935 79.475 39.455 ;
        RECT 79.645 39.105 81.335 39.625 ;
        RECT 76.935 38.165 77.105 38.775 ;
        RECT 77.275 38.385 77.605 38.820 ;
        RECT 77.825 38.165 81.335 38.935 ;
        RECT 81.505 38.915 82.025 39.455 ;
        RECT 82.195 39.085 82.715 39.625 ;
        RECT 82.885 39.625 84.095 40.715 ;
        RECT 82.885 39.085 83.405 39.625 ;
        RECT 83.575 38.915 84.095 39.455 ;
        RECT 81.505 38.165 82.715 38.915 ;
        RECT 82.885 38.165 84.095 38.915 ;
        RECT 5.520 37.995 84.180 38.165 ;
        RECT 5.605 37.245 6.815 37.995 ;
        RECT 5.605 36.705 6.125 37.245 ;
        RECT 7.905 37.195 8.245 37.825 ;
        RECT 8.415 37.195 8.665 37.995 ;
        RECT 8.855 37.345 9.185 37.825 ;
        RECT 9.355 37.535 9.580 37.995 ;
        RECT 9.750 37.345 10.080 37.825 ;
        RECT 6.295 36.535 6.815 37.075 ;
        RECT 5.605 35.445 6.815 36.535 ;
        RECT 7.905 36.585 8.080 37.195 ;
        RECT 8.855 37.175 10.080 37.345 ;
        RECT 10.710 37.215 11.210 37.825 ;
        RECT 11.620 37.255 12.235 37.825 ;
        RECT 12.405 37.485 12.620 37.995 ;
        RECT 12.850 37.485 13.130 37.815 ;
        RECT 13.310 37.485 13.550 37.995 ;
        RECT 8.250 36.835 8.945 37.005 ;
        RECT 8.775 36.585 8.945 36.835 ;
        RECT 9.120 36.805 9.540 37.005 ;
        RECT 9.710 36.805 10.040 37.005 ;
        RECT 10.210 36.805 10.540 37.005 ;
        RECT 10.710 36.585 10.880 37.215 ;
        RECT 11.065 36.755 11.415 37.005 ;
        RECT 7.905 35.615 8.245 36.585 ;
        RECT 8.415 35.445 8.585 36.585 ;
        RECT 8.775 36.415 11.210 36.585 ;
        RECT 8.855 35.445 9.105 36.245 ;
        RECT 9.750 35.615 10.080 36.415 ;
        RECT 10.380 35.445 10.710 36.245 ;
        RECT 10.880 35.615 11.210 36.415 ;
        RECT 11.620 36.235 11.935 37.255 ;
        RECT 12.105 36.585 12.275 37.085 ;
        RECT 12.525 36.755 12.790 37.315 ;
        RECT 12.960 36.585 13.130 37.485 ;
        RECT 13.300 36.755 13.655 37.315 ;
        RECT 13.890 37.230 14.345 37.995 ;
        RECT 14.620 37.615 15.920 37.825 ;
        RECT 16.175 37.635 16.505 37.995 ;
        RECT 15.750 37.465 15.920 37.615 ;
        RECT 16.675 37.495 16.935 37.825 ;
        RECT 16.705 37.485 16.935 37.495 ;
        RECT 14.820 37.005 15.040 37.405 ;
        RECT 13.885 36.805 14.375 37.005 ;
        RECT 14.565 36.795 15.040 37.005 ;
        RECT 15.285 37.005 15.495 37.405 ;
        RECT 15.750 37.340 16.505 37.465 ;
        RECT 15.750 37.295 16.595 37.340 ;
        RECT 16.325 37.175 16.595 37.295 ;
        RECT 15.285 36.795 15.615 37.005 ;
        RECT 15.785 36.735 16.195 37.040 ;
        RECT 12.105 36.415 13.530 36.585 ;
        RECT 11.620 35.615 12.155 36.235 ;
        RECT 12.325 35.445 12.655 36.245 ;
        RECT 13.140 36.240 13.530 36.415 ;
        RECT 13.890 36.565 15.065 36.625 ;
        RECT 16.425 36.600 16.595 37.175 ;
        RECT 16.395 36.565 16.595 36.600 ;
        RECT 13.890 36.455 16.595 36.565 ;
        RECT 13.890 35.835 14.145 36.455 ;
        RECT 14.735 36.395 16.535 36.455 ;
        RECT 14.735 36.365 15.065 36.395 ;
        RECT 16.765 36.295 16.935 37.485 ;
        RECT 17.105 37.225 20.615 37.995 ;
        RECT 17.105 36.705 18.755 37.225 ;
        RECT 21.265 37.185 21.505 37.995 ;
        RECT 21.675 37.185 22.005 37.825 ;
        RECT 22.175 37.185 22.445 37.995 ;
        RECT 22.625 37.245 23.835 37.995 ;
        RECT 24.005 37.535 24.565 37.825 ;
        RECT 24.735 37.535 24.985 37.995 ;
        RECT 18.925 36.535 20.615 37.055 ;
        RECT 21.245 36.755 21.595 37.005 ;
        RECT 21.765 36.585 21.935 37.185 ;
        RECT 22.105 36.755 22.455 37.005 ;
        RECT 22.625 36.705 23.145 37.245 ;
        RECT 14.395 36.195 14.580 36.285 ;
        RECT 15.170 36.195 16.005 36.205 ;
        RECT 14.395 35.995 16.005 36.195 ;
        RECT 14.395 35.955 14.625 35.995 ;
        RECT 13.890 35.615 14.225 35.835 ;
        RECT 15.230 35.445 15.585 35.825 ;
        RECT 15.755 35.615 16.005 35.995 ;
        RECT 16.255 35.445 16.505 36.225 ;
        RECT 16.675 35.615 16.935 36.295 ;
        RECT 17.105 35.445 20.615 36.535 ;
        RECT 21.255 36.415 21.935 36.585 ;
        RECT 21.255 35.630 21.585 36.415 ;
        RECT 22.115 35.445 22.445 36.585 ;
        RECT 23.315 36.535 23.835 37.075 ;
        RECT 22.625 35.445 23.835 36.535 ;
        RECT 24.005 36.165 24.255 37.535 ;
        RECT 25.605 37.365 25.935 37.725 ;
        RECT 24.545 37.175 25.935 37.365 ;
        RECT 26.305 37.225 29.815 37.995 ;
        RECT 29.985 37.245 31.195 37.995 ;
        RECT 31.365 37.270 31.655 37.995 ;
        RECT 24.545 37.085 24.715 37.175 ;
        RECT 24.425 36.755 24.715 37.085 ;
        RECT 24.885 36.755 25.225 37.005 ;
        RECT 25.445 36.755 26.120 37.005 ;
        RECT 24.545 36.505 24.715 36.755 ;
        RECT 24.545 36.335 25.485 36.505 ;
        RECT 25.855 36.395 26.120 36.755 ;
        RECT 26.305 36.705 27.955 37.225 ;
        RECT 28.125 36.535 29.815 37.055 ;
        RECT 29.985 36.705 30.505 37.245 ;
        RECT 31.825 37.225 33.495 37.995 ;
        RECT 30.675 36.535 31.195 37.075 ;
        RECT 31.825 36.705 32.575 37.225 ;
        RECT 24.005 35.615 24.465 36.165 ;
        RECT 24.655 35.445 24.985 36.165 ;
        RECT 25.185 35.785 25.485 36.335 ;
        RECT 25.655 35.445 25.935 36.115 ;
        RECT 26.305 35.445 29.815 36.535 ;
        RECT 29.985 35.445 31.195 36.535 ;
        RECT 31.365 35.445 31.655 36.610 ;
        RECT 32.745 36.535 33.495 37.055 ;
        RECT 31.825 35.445 33.495 36.535 ;
        RECT 33.670 36.395 34.005 37.815 ;
        RECT 34.185 37.625 34.930 37.995 ;
        RECT 35.495 37.455 35.750 37.815 ;
        RECT 35.930 37.625 36.260 37.995 ;
        RECT 36.440 37.455 36.665 37.815 ;
        RECT 34.180 37.265 36.665 37.455 ;
        RECT 34.180 36.575 34.405 37.265 ;
        RECT 36.885 37.225 39.475 37.995 ;
        RECT 40.110 37.255 40.365 37.825 ;
        RECT 40.535 37.595 40.865 37.995 ;
        RECT 41.290 37.460 41.820 37.825 ;
        RECT 42.010 37.655 42.285 37.825 ;
        RECT 42.005 37.485 42.285 37.655 ;
        RECT 41.290 37.425 41.465 37.460 ;
        RECT 40.535 37.255 41.465 37.425 ;
        RECT 34.605 36.755 34.885 37.085 ;
        RECT 35.065 36.755 35.640 37.085 ;
        RECT 35.820 36.755 36.255 37.085 ;
        RECT 36.435 36.755 36.705 37.085 ;
        RECT 36.885 36.705 38.095 37.225 ;
        RECT 34.180 36.395 36.675 36.575 ;
        RECT 38.265 36.535 39.475 37.055 ;
        RECT 33.670 35.625 33.935 36.395 ;
        RECT 34.105 35.445 34.435 36.165 ;
        RECT 34.625 35.985 35.815 36.215 ;
        RECT 34.625 35.625 34.885 35.985 ;
        RECT 35.055 35.445 35.385 35.815 ;
        RECT 35.555 35.625 35.815 35.985 ;
        RECT 36.385 35.625 36.675 36.395 ;
        RECT 36.885 35.445 39.475 36.535 ;
        RECT 40.110 36.585 40.280 37.255 ;
        RECT 40.535 37.085 40.705 37.255 ;
        RECT 40.450 36.755 40.705 37.085 ;
        RECT 40.930 36.755 41.125 37.085 ;
        RECT 40.110 35.615 40.445 36.585 ;
        RECT 40.615 35.445 40.785 36.585 ;
        RECT 40.955 35.785 41.125 36.755 ;
        RECT 41.295 36.125 41.465 37.255 ;
        RECT 41.635 36.465 41.805 37.265 ;
        RECT 42.010 36.665 42.285 37.485 ;
        RECT 42.455 36.465 42.645 37.825 ;
        RECT 42.825 37.460 43.335 37.995 ;
        RECT 43.555 37.185 43.800 37.790 ;
        RECT 44.245 37.335 44.520 37.995 ;
        RECT 44.690 37.365 44.940 37.825 ;
        RECT 45.115 37.500 45.445 37.995 ;
        RECT 42.845 37.015 44.075 37.185 ;
        RECT 44.690 37.155 44.860 37.365 ;
        RECT 45.625 37.330 45.855 37.775 ;
        RECT 41.635 36.295 42.645 36.465 ;
        RECT 42.815 36.450 43.565 36.640 ;
        RECT 41.295 35.955 42.420 36.125 ;
        RECT 42.815 35.785 42.985 36.450 ;
        RECT 43.735 36.205 44.075 37.015 ;
        RECT 44.245 36.635 44.860 37.155 ;
        RECT 45.030 36.655 45.260 37.085 ;
        RECT 45.445 36.835 45.855 37.330 ;
        RECT 46.025 37.510 46.815 37.775 ;
        RECT 46.025 36.655 46.280 37.510 ;
        RECT 46.450 36.835 46.835 37.315 ;
        RECT 47.525 37.175 47.735 37.995 ;
        RECT 47.905 37.195 48.235 37.825 ;
        RECT 40.955 35.615 42.985 35.785 ;
        RECT 43.155 35.445 43.325 36.205 ;
        RECT 43.560 35.795 44.075 36.205 ;
        RECT 44.245 35.445 44.505 36.455 ;
        RECT 44.675 36.285 44.845 36.635 ;
        RECT 45.030 36.485 46.820 36.655 ;
        RECT 47.905 36.595 48.155 37.195 ;
        RECT 48.405 37.175 48.635 37.995 ;
        RECT 49.090 37.515 49.390 37.995 ;
        RECT 49.560 37.345 49.820 37.800 ;
        RECT 49.990 37.515 50.250 37.995 ;
        RECT 50.420 37.345 50.680 37.800 ;
        RECT 50.850 37.515 51.110 37.995 ;
        RECT 51.280 37.345 51.540 37.800 ;
        RECT 51.710 37.515 51.970 37.995 ;
        RECT 52.140 37.345 52.400 37.800 ;
        RECT 52.570 37.470 52.830 37.995 ;
        RECT 49.090 37.175 52.400 37.345 ;
        RECT 48.325 36.755 48.655 37.005 ;
        RECT 44.675 35.615 44.950 36.285 ;
        RECT 45.150 35.445 45.365 36.290 ;
        RECT 45.590 36.190 45.840 36.485 ;
        RECT 46.065 36.125 46.395 36.315 ;
        RECT 45.550 35.615 46.025 35.955 ;
        RECT 46.205 35.950 46.395 36.125 ;
        RECT 46.565 36.120 46.820 36.485 ;
        RECT 46.205 35.445 46.835 35.950 ;
        RECT 47.525 35.445 47.735 36.585 ;
        RECT 47.905 35.615 48.235 36.595 ;
        RECT 49.090 36.585 50.060 37.175 ;
        RECT 53.000 37.005 53.250 37.815 ;
        RECT 53.430 37.535 53.675 37.995 ;
        RECT 54.105 37.365 54.435 37.725 ;
        RECT 55.065 37.535 55.315 37.995 ;
        RECT 55.485 37.535 56.035 37.825 ;
        RECT 50.230 36.755 53.250 37.005 ;
        RECT 53.420 36.755 53.735 37.365 ;
        RECT 54.105 37.175 55.495 37.365 ;
        RECT 55.325 37.085 55.495 37.175 ;
        RECT 53.905 36.755 54.595 37.005 ;
        RECT 54.825 36.755 55.155 37.005 ;
        RECT 55.325 36.755 55.615 37.085 ;
        RECT 48.405 35.445 48.635 36.585 ;
        RECT 49.090 36.345 52.400 36.585 ;
        RECT 49.095 35.445 49.390 36.175 ;
        RECT 49.560 35.620 49.820 36.345 ;
        RECT 49.990 35.445 50.250 36.175 ;
        RECT 50.420 35.620 50.680 36.345 ;
        RECT 50.850 35.445 51.110 36.175 ;
        RECT 51.280 35.620 51.540 36.345 ;
        RECT 51.710 35.445 51.970 36.175 ;
        RECT 52.140 35.620 52.400 36.345 ;
        RECT 52.570 35.445 52.830 36.555 ;
        RECT 53.000 35.620 53.250 36.755 ;
        RECT 53.430 35.445 53.725 36.555 ;
        RECT 53.905 36.315 54.220 36.755 ;
        RECT 55.325 36.505 55.495 36.755 ;
        RECT 54.555 36.335 55.495 36.505 ;
        RECT 54.105 35.445 54.385 36.115 ;
        RECT 54.555 35.785 54.855 36.335 ;
        RECT 55.785 36.165 56.035 37.535 ;
        RECT 56.205 37.195 56.495 37.995 ;
        RECT 57.125 37.270 57.415 37.995 ;
        RECT 57.585 37.195 57.925 37.825 ;
        RECT 58.095 37.195 58.345 37.995 ;
        RECT 58.535 37.345 58.865 37.825 ;
        RECT 59.035 37.535 59.260 37.995 ;
        RECT 59.430 37.345 59.760 37.825 ;
        RECT 55.065 35.445 55.395 36.165 ;
        RECT 55.585 35.615 56.035 36.165 ;
        RECT 56.205 35.445 56.495 36.585 ;
        RECT 57.125 35.445 57.415 36.610 ;
        RECT 57.585 36.585 57.760 37.195 ;
        RECT 58.535 37.175 59.760 37.345 ;
        RECT 60.390 37.215 60.890 37.825 ;
        RECT 61.890 37.485 62.130 37.995 ;
        RECT 62.310 37.485 62.590 37.815 ;
        RECT 62.820 37.485 63.035 37.995 ;
        RECT 57.930 36.835 58.625 37.005 ;
        RECT 58.455 36.585 58.625 36.835 ;
        RECT 58.800 36.805 59.220 37.005 ;
        RECT 59.390 36.805 59.720 37.005 ;
        RECT 59.890 36.805 60.220 37.005 ;
        RECT 60.390 36.585 60.560 37.215 ;
        RECT 60.745 36.755 61.095 37.005 ;
        RECT 61.785 36.755 62.140 37.315 ;
        RECT 62.310 36.585 62.480 37.485 ;
        RECT 62.650 36.755 62.915 37.315 ;
        RECT 63.205 37.255 63.820 37.825 ;
        RECT 63.165 36.585 63.335 37.085 ;
        RECT 57.585 35.615 57.925 36.585 ;
        RECT 58.095 35.445 58.265 36.585 ;
        RECT 58.455 36.415 60.890 36.585 ;
        RECT 58.535 35.445 58.785 36.245 ;
        RECT 59.430 35.615 59.760 36.415 ;
        RECT 60.060 35.445 60.390 36.245 ;
        RECT 60.560 35.615 60.890 36.415 ;
        RECT 61.910 36.415 63.335 36.585 ;
        RECT 61.910 36.240 62.300 36.415 ;
        RECT 62.785 35.445 63.115 36.245 ;
        RECT 63.505 36.235 63.820 37.255 ;
        RECT 64.025 37.365 64.365 37.825 ;
        RECT 64.535 37.535 64.705 37.995 ;
        RECT 64.875 37.615 66.045 37.825 ;
        RECT 64.875 37.365 65.125 37.615 ;
        RECT 65.715 37.595 66.045 37.615 ;
        RECT 64.025 37.195 65.125 37.365 ;
        RECT 65.295 37.175 66.155 37.425 ;
        RECT 66.525 37.365 66.855 37.725 ;
        RECT 67.475 37.535 67.725 37.995 ;
        RECT 67.895 37.535 68.455 37.825 ;
        RECT 66.525 37.175 67.915 37.365 ;
        RECT 64.025 36.755 64.785 37.005 ;
        RECT 64.955 36.755 65.705 37.005 ;
        RECT 65.875 36.585 66.155 37.175 ;
        RECT 67.745 37.085 67.915 37.175 ;
        RECT 63.285 35.615 63.820 36.235 ;
        RECT 64.025 35.445 64.285 36.585 ;
        RECT 64.455 36.415 66.155 36.585 ;
        RECT 66.340 36.755 67.015 37.005 ;
        RECT 67.235 36.755 67.575 37.005 ;
        RECT 67.745 36.755 68.035 37.085 ;
        RECT 64.455 35.615 64.785 36.415 ;
        RECT 64.955 35.445 65.125 36.245 ;
        RECT 65.295 35.615 65.625 36.415 ;
        RECT 66.340 36.395 66.605 36.755 ;
        RECT 67.745 36.505 67.915 36.755 ;
        RECT 66.975 36.335 67.915 36.505 ;
        RECT 65.795 35.445 66.050 36.245 ;
        RECT 66.525 35.445 66.805 36.115 ;
        RECT 66.975 35.785 67.275 36.335 ;
        RECT 68.205 36.165 68.455 37.535 ;
        RECT 68.625 37.225 72.135 37.995 ;
        RECT 68.625 36.705 70.275 37.225 ;
        RECT 72.510 37.215 73.010 37.825 ;
        RECT 70.445 36.535 72.135 37.055 ;
        RECT 72.305 36.755 72.655 37.005 ;
        RECT 72.840 36.585 73.010 37.215 ;
        RECT 73.640 37.345 73.970 37.825 ;
        RECT 74.140 37.535 74.365 37.995 ;
        RECT 74.535 37.345 74.865 37.825 ;
        RECT 73.640 37.175 74.865 37.345 ;
        RECT 75.055 37.195 75.305 37.995 ;
        RECT 75.475 37.195 75.815 37.825 ;
        RECT 73.180 36.805 73.510 37.005 ;
        RECT 73.680 36.805 74.010 37.005 ;
        RECT 74.180 36.805 74.600 37.005 ;
        RECT 74.775 36.835 75.470 37.005 ;
        RECT 74.775 36.585 74.945 36.835 ;
        RECT 75.640 36.585 75.815 37.195 ;
        RECT 67.475 35.445 67.805 36.165 ;
        RECT 67.995 35.615 68.455 36.165 ;
        RECT 68.625 35.445 72.135 36.535 ;
        RECT 72.510 36.415 74.945 36.585 ;
        RECT 72.510 35.615 72.840 36.415 ;
        RECT 73.010 35.445 73.340 36.245 ;
        RECT 73.640 35.615 73.970 36.415 ;
        RECT 74.615 35.445 74.865 36.245 ;
        RECT 75.135 35.445 75.305 36.585 ;
        RECT 75.475 35.615 75.815 36.585 ;
        RECT 75.985 37.320 76.245 37.825 ;
        RECT 76.425 37.615 76.755 37.995 ;
        RECT 76.935 37.445 77.105 37.825 ;
        RECT 77.365 37.450 82.710 37.995 ;
        RECT 75.985 36.520 76.165 37.320 ;
        RECT 76.440 37.275 77.105 37.445 ;
        RECT 76.440 37.020 76.610 37.275 ;
        RECT 76.335 36.690 76.610 37.020 ;
        RECT 76.835 36.725 77.175 37.095 ;
        RECT 76.440 36.545 76.610 36.690 ;
        RECT 78.950 36.620 79.290 37.450 ;
        RECT 82.885 37.245 84.095 37.995 ;
        RECT 75.985 35.615 76.255 36.520 ;
        RECT 76.440 36.375 77.115 36.545 ;
        RECT 76.425 35.445 76.755 36.205 ;
        RECT 76.935 35.615 77.115 36.375 ;
        RECT 80.770 35.880 81.120 37.130 ;
        RECT 82.885 36.535 83.405 37.075 ;
        RECT 83.575 36.705 84.095 37.245 ;
        RECT 77.365 35.445 82.710 35.880 ;
        RECT 82.885 35.445 84.095 36.535 ;
        RECT 5.520 35.275 84.180 35.445 ;
        RECT 5.605 34.185 6.815 35.275 ;
        RECT 6.985 34.185 9.575 35.275 ;
        RECT 10.295 34.605 10.465 35.105 ;
        RECT 10.635 34.775 10.965 35.275 ;
        RECT 10.295 34.435 10.960 34.605 ;
        RECT 5.605 33.475 6.125 34.015 ;
        RECT 6.295 33.645 6.815 34.185 ;
        RECT 6.985 33.495 8.195 34.015 ;
        RECT 8.365 33.665 9.575 34.185 ;
        RECT 10.210 33.615 10.560 34.265 ;
        RECT 5.605 32.725 6.815 33.475 ;
        RECT 6.985 32.725 9.575 33.495 ;
        RECT 10.730 33.445 10.960 34.435 ;
        RECT 10.295 33.275 10.960 33.445 ;
        RECT 10.295 32.985 10.465 33.275 ;
        RECT 10.635 32.725 10.965 33.105 ;
        RECT 11.135 32.985 11.320 35.105 ;
        RECT 11.560 34.815 11.825 35.275 ;
        RECT 11.995 34.680 12.245 35.105 ;
        RECT 12.455 34.830 13.560 35.000 ;
        RECT 11.940 34.550 12.245 34.680 ;
        RECT 11.490 33.355 11.770 34.305 ;
        RECT 11.940 33.445 12.110 34.550 ;
        RECT 12.280 33.765 12.520 34.360 ;
        RECT 12.690 34.295 13.220 34.660 ;
        RECT 12.690 33.595 12.860 34.295 ;
        RECT 13.390 34.215 13.560 34.830 ;
        RECT 13.730 34.475 13.900 35.275 ;
        RECT 14.070 34.775 14.320 35.105 ;
        RECT 14.545 34.805 15.430 34.975 ;
        RECT 13.390 34.125 13.900 34.215 ;
        RECT 11.940 33.315 12.165 33.445 ;
        RECT 12.335 33.375 12.860 33.595 ;
        RECT 13.030 33.955 13.900 34.125 ;
        RECT 11.575 32.725 11.825 33.185 ;
        RECT 11.995 33.175 12.165 33.315 ;
        RECT 13.030 33.175 13.200 33.955 ;
        RECT 13.730 33.885 13.900 33.955 ;
        RECT 13.410 33.705 13.610 33.735 ;
        RECT 14.070 33.705 14.240 34.775 ;
        RECT 14.410 33.885 14.600 34.605 ;
        RECT 13.410 33.405 14.240 33.705 ;
        RECT 14.770 33.675 15.090 34.635 ;
        RECT 11.995 33.005 12.330 33.175 ;
        RECT 12.525 33.005 13.200 33.175 ;
        RECT 13.520 32.725 13.890 33.225 ;
        RECT 14.070 33.175 14.240 33.405 ;
        RECT 14.625 33.345 15.090 33.675 ;
        RECT 15.260 33.965 15.430 34.805 ;
        RECT 15.610 34.775 15.925 35.275 ;
        RECT 16.155 34.545 16.495 35.105 ;
        RECT 15.600 34.170 16.495 34.545 ;
        RECT 16.665 34.265 16.835 35.275 ;
        RECT 16.305 33.965 16.495 34.170 ;
        RECT 17.005 34.215 17.335 35.060 ;
        RECT 17.005 34.135 17.395 34.215 ;
        RECT 17.180 34.085 17.395 34.135 ;
        RECT 18.485 34.110 18.775 35.275 ;
        RECT 18.980 34.485 19.515 35.105 ;
        RECT 15.260 33.635 16.135 33.965 ;
        RECT 16.305 33.635 17.055 33.965 ;
        RECT 15.260 33.175 15.430 33.635 ;
        RECT 16.305 33.465 16.505 33.635 ;
        RECT 17.225 33.505 17.395 34.085 ;
        RECT 17.170 33.465 17.395 33.505 ;
        RECT 14.070 33.005 14.475 33.175 ;
        RECT 14.645 33.005 15.430 33.175 ;
        RECT 15.705 32.725 15.915 33.255 ;
        RECT 16.175 32.940 16.505 33.465 ;
        RECT 17.015 33.380 17.395 33.465 ;
        RECT 18.980 33.465 19.295 34.485 ;
        RECT 19.685 34.475 20.015 35.275 ;
        RECT 20.500 34.305 20.890 34.480 ;
        RECT 19.465 34.135 20.890 34.305 ;
        RECT 22.370 34.305 22.700 35.105 ;
        RECT 22.870 34.475 23.200 35.275 ;
        RECT 23.500 34.305 23.830 35.105 ;
        RECT 24.475 34.475 24.725 35.275 ;
        RECT 22.370 34.135 24.805 34.305 ;
        RECT 24.995 34.135 25.165 35.275 ;
        RECT 25.335 34.135 25.675 35.105 ;
        RECT 25.950 34.475 26.205 35.275 ;
        RECT 26.375 34.305 26.705 35.105 ;
        RECT 26.875 34.475 27.045 35.275 ;
        RECT 27.215 34.305 27.545 35.105 ;
        RECT 19.465 33.635 19.635 34.135 ;
        RECT 16.675 32.725 16.845 33.335 ;
        RECT 17.015 32.945 17.345 33.380 ;
        RECT 18.485 32.725 18.775 33.450 ;
        RECT 18.980 32.895 19.595 33.465 ;
        RECT 19.885 33.405 20.150 33.965 ;
        RECT 20.320 33.235 20.490 34.135 ;
        RECT 20.660 33.405 21.015 33.965 ;
        RECT 22.165 33.715 22.515 33.965 ;
        RECT 22.700 33.505 22.870 34.135 ;
        RECT 23.040 33.715 23.370 33.915 ;
        RECT 23.540 33.715 23.870 33.915 ;
        RECT 24.040 33.715 24.460 33.915 ;
        RECT 24.635 33.885 24.805 34.135 ;
        RECT 24.635 33.715 25.330 33.885 ;
        RECT 19.765 32.725 19.980 33.235 ;
        RECT 20.210 32.905 20.490 33.235 ;
        RECT 20.670 32.725 20.910 33.235 ;
        RECT 22.370 32.895 22.870 33.505 ;
        RECT 23.500 33.375 24.725 33.545 ;
        RECT 25.500 33.525 25.675 34.135 ;
        RECT 23.500 32.895 23.830 33.375 ;
        RECT 24.000 32.725 24.225 33.185 ;
        RECT 24.395 32.895 24.725 33.375 ;
        RECT 24.915 32.725 25.165 33.525 ;
        RECT 25.335 32.895 25.675 33.525 ;
        RECT 25.845 34.135 27.545 34.305 ;
        RECT 27.715 34.135 27.975 35.275 ;
        RECT 28.145 34.185 29.815 35.275 ;
        RECT 30.045 34.215 30.375 35.060 ;
        RECT 30.545 34.265 30.715 35.275 ;
        RECT 30.885 34.545 31.225 35.105 ;
        RECT 31.455 34.775 31.770 35.275 ;
        RECT 31.950 34.805 32.835 34.975 ;
        RECT 25.845 33.545 26.125 34.135 ;
        RECT 26.295 33.715 27.045 33.965 ;
        RECT 27.215 33.715 27.975 33.965 ;
        RECT 25.845 33.295 26.705 33.545 ;
        RECT 26.875 33.355 27.975 33.525 ;
        RECT 25.955 33.105 26.285 33.125 ;
        RECT 26.875 33.105 27.125 33.355 ;
        RECT 25.955 32.895 27.125 33.105 ;
        RECT 27.295 32.725 27.465 33.185 ;
        RECT 27.635 32.895 27.975 33.355 ;
        RECT 28.145 33.495 28.895 34.015 ;
        RECT 29.065 33.665 29.815 34.185 ;
        RECT 29.985 34.135 30.375 34.215 ;
        RECT 30.885 34.170 31.780 34.545 ;
        RECT 29.985 34.085 30.200 34.135 ;
        RECT 29.985 33.505 30.155 34.085 ;
        RECT 30.885 33.965 31.075 34.170 ;
        RECT 31.950 33.965 32.120 34.805 ;
        RECT 33.060 34.775 33.310 35.105 ;
        RECT 30.325 33.635 31.075 33.965 ;
        RECT 31.245 33.635 32.120 33.965 ;
        RECT 28.145 32.725 29.815 33.495 ;
        RECT 29.985 33.465 30.210 33.505 ;
        RECT 30.875 33.465 31.075 33.635 ;
        RECT 29.985 33.380 30.365 33.465 ;
        RECT 30.035 32.945 30.365 33.380 ;
        RECT 30.535 32.725 30.705 33.335 ;
        RECT 30.875 32.940 31.205 33.465 ;
        RECT 31.465 32.725 31.675 33.255 ;
        RECT 31.950 33.175 32.120 33.635 ;
        RECT 32.290 33.675 32.610 34.635 ;
        RECT 32.780 33.885 32.970 34.605 ;
        RECT 33.140 33.705 33.310 34.775 ;
        RECT 33.480 34.475 33.650 35.275 ;
        RECT 33.820 34.830 34.925 35.000 ;
        RECT 33.820 34.215 33.990 34.830 ;
        RECT 35.135 34.680 35.385 35.105 ;
        RECT 35.555 34.815 35.820 35.275 ;
        RECT 34.160 34.295 34.690 34.660 ;
        RECT 35.135 34.550 35.440 34.680 ;
        RECT 33.480 34.125 33.990 34.215 ;
        RECT 33.480 33.955 34.350 34.125 ;
        RECT 33.480 33.885 33.650 33.955 ;
        RECT 33.770 33.705 33.970 33.735 ;
        RECT 32.290 33.345 32.755 33.675 ;
        RECT 33.140 33.405 33.970 33.705 ;
        RECT 33.140 33.175 33.310 33.405 ;
        RECT 31.950 33.005 32.735 33.175 ;
        RECT 32.905 33.005 33.310 33.175 ;
        RECT 33.490 32.725 33.860 33.225 ;
        RECT 34.180 33.175 34.350 33.955 ;
        RECT 34.520 33.595 34.690 34.295 ;
        RECT 34.860 33.765 35.100 34.360 ;
        RECT 34.520 33.375 35.045 33.595 ;
        RECT 35.270 33.445 35.440 34.550 ;
        RECT 35.215 33.315 35.440 33.445 ;
        RECT 35.610 33.355 35.890 34.305 ;
        RECT 35.215 33.175 35.385 33.315 ;
        RECT 34.180 33.005 34.855 33.175 ;
        RECT 35.050 33.005 35.385 33.175 ;
        RECT 35.555 32.725 35.805 33.185 ;
        RECT 36.060 32.985 36.245 35.105 ;
        RECT 36.415 34.775 36.745 35.275 ;
        RECT 36.915 34.605 37.085 35.105 ;
        RECT 36.420 34.435 37.085 34.605 ;
        RECT 36.420 33.445 36.650 34.435 ;
        RECT 36.820 33.615 37.170 34.265 ;
        RECT 37.345 34.135 37.685 35.105 ;
        RECT 37.855 34.135 38.025 35.275 ;
        RECT 38.295 34.475 38.545 35.275 ;
        RECT 39.190 34.305 39.520 35.105 ;
        RECT 39.820 34.475 40.150 35.275 ;
        RECT 40.320 34.305 40.650 35.105 ;
        RECT 38.215 34.135 40.650 34.305 ;
        RECT 41.025 34.185 43.615 35.275 ;
        RECT 37.345 33.575 37.520 34.135 ;
        RECT 38.215 33.885 38.385 34.135 ;
        RECT 37.690 33.715 38.385 33.885 ;
        RECT 38.560 33.715 38.980 33.915 ;
        RECT 39.150 33.715 39.480 33.915 ;
        RECT 39.650 33.715 39.980 33.915 ;
        RECT 37.345 33.525 37.575 33.575 ;
        RECT 36.420 33.275 37.085 33.445 ;
        RECT 36.415 32.725 36.745 33.105 ;
        RECT 36.915 32.985 37.085 33.275 ;
        RECT 37.345 32.895 37.685 33.525 ;
        RECT 37.855 32.725 38.105 33.525 ;
        RECT 38.295 33.375 39.520 33.545 ;
        RECT 38.295 32.895 38.625 33.375 ;
        RECT 38.795 32.725 39.020 33.185 ;
        RECT 39.190 32.895 39.520 33.375 ;
        RECT 40.150 33.505 40.320 34.135 ;
        RECT 40.505 33.715 40.855 33.965 ;
        RECT 40.150 32.895 40.650 33.505 ;
        RECT 41.025 33.495 42.235 34.015 ;
        RECT 42.405 33.665 43.615 34.185 ;
        RECT 44.245 34.110 44.535 35.275 ;
        RECT 44.705 34.185 47.295 35.275 ;
        RECT 44.705 33.495 45.915 34.015 ;
        RECT 46.085 33.665 47.295 34.185 ;
        RECT 47.470 34.135 47.805 35.105 ;
        RECT 47.975 34.135 48.145 35.275 ;
        RECT 48.315 34.935 50.345 35.105 ;
        RECT 41.025 32.725 43.615 33.495 ;
        RECT 44.245 32.725 44.535 33.450 ;
        RECT 44.705 32.725 47.295 33.495 ;
        RECT 47.470 33.465 47.640 34.135 ;
        RECT 48.315 33.965 48.485 34.935 ;
        RECT 47.810 33.635 48.065 33.965 ;
        RECT 48.290 33.635 48.485 33.965 ;
        RECT 48.655 34.595 49.780 34.765 ;
        RECT 47.895 33.465 48.065 33.635 ;
        RECT 48.655 33.465 48.825 34.595 ;
        RECT 47.470 32.895 47.725 33.465 ;
        RECT 47.895 33.295 48.825 33.465 ;
        RECT 48.995 34.255 50.005 34.425 ;
        RECT 48.995 33.455 49.165 34.255 ;
        RECT 49.370 33.575 49.645 34.055 ;
        RECT 49.365 33.405 49.645 33.575 ;
        RECT 48.650 33.260 48.825 33.295 ;
        RECT 47.895 32.725 48.225 33.125 ;
        RECT 48.650 32.895 49.180 33.260 ;
        RECT 49.370 32.895 49.645 33.405 ;
        RECT 49.815 32.895 50.005 34.255 ;
        RECT 50.175 34.270 50.345 34.935 ;
        RECT 50.515 34.515 50.685 35.275 ;
        RECT 50.920 34.515 51.435 34.925 ;
        RECT 50.175 34.080 50.925 34.270 ;
        RECT 51.095 33.705 51.435 34.515 ;
        RECT 50.205 33.535 51.435 33.705 ;
        RECT 51.605 34.135 51.990 35.105 ;
        RECT 52.160 34.815 52.485 35.275 ;
        RECT 53.005 34.645 53.285 35.105 ;
        RECT 52.160 34.425 53.285 34.645 ;
        RECT 50.185 32.725 50.695 33.260 ;
        RECT 50.915 32.930 51.160 33.535 ;
        RECT 51.605 33.465 51.885 34.135 ;
        RECT 52.160 33.965 52.610 34.425 ;
        RECT 53.475 34.255 53.875 35.105 ;
        RECT 54.275 34.815 54.545 35.275 ;
        RECT 54.715 34.645 55.000 35.105 ;
        RECT 52.055 33.635 52.610 33.965 ;
        RECT 52.780 33.695 53.875 34.255 ;
        RECT 52.160 33.525 52.610 33.635 ;
        RECT 51.605 32.895 51.990 33.465 ;
        RECT 52.160 33.355 53.285 33.525 ;
        RECT 52.160 32.725 52.485 33.185 ;
        RECT 53.005 32.895 53.285 33.355 ;
        RECT 53.475 32.895 53.875 33.695 ;
        RECT 54.045 34.425 55.000 34.645 ;
        RECT 54.045 33.525 54.255 34.425 ;
        RECT 55.285 34.305 55.555 35.075 ;
        RECT 55.725 34.495 56.055 35.275 ;
        RECT 56.260 34.670 56.445 35.075 ;
        RECT 56.615 34.850 56.950 35.275 ;
        RECT 57.125 34.840 62.470 35.275 ;
        RECT 56.260 34.495 56.925 34.670 ;
        RECT 54.425 33.695 55.115 34.255 ;
        RECT 55.285 34.135 56.415 34.305 ;
        RECT 54.045 33.355 55.000 33.525 ;
        RECT 54.275 32.725 54.545 33.185 ;
        RECT 54.715 32.895 55.000 33.355 ;
        RECT 55.285 33.225 55.455 34.135 ;
        RECT 55.625 33.385 55.985 33.965 ;
        RECT 56.165 33.635 56.415 34.135 ;
        RECT 56.585 33.465 56.925 34.495 ;
        RECT 56.240 33.295 56.925 33.465 ;
        RECT 55.285 32.895 55.545 33.225 ;
        RECT 55.755 32.725 56.030 33.205 ;
        RECT 56.240 32.895 56.445 33.295 ;
        RECT 58.710 33.270 59.050 34.100 ;
        RECT 60.530 33.590 60.880 34.840 ;
        RECT 62.645 34.185 66.155 35.275 ;
        RECT 66.325 34.185 67.535 35.275 ;
        RECT 62.645 33.495 64.295 34.015 ;
        RECT 64.465 33.665 66.155 34.185 ;
        RECT 56.615 32.725 56.950 33.125 ;
        RECT 57.125 32.725 62.470 33.270 ;
        RECT 62.645 32.725 66.155 33.495 ;
        RECT 66.325 33.475 66.845 34.015 ;
        RECT 67.015 33.645 67.535 34.185 ;
        RECT 67.890 34.305 68.280 34.480 ;
        RECT 68.765 34.475 69.095 35.275 ;
        RECT 69.265 34.485 69.800 35.105 ;
        RECT 67.890 34.135 69.315 34.305 ;
        RECT 66.325 32.725 67.535 33.475 ;
        RECT 67.765 33.405 68.120 33.965 ;
        RECT 68.290 33.235 68.460 34.135 ;
        RECT 68.630 33.405 68.895 33.965 ;
        RECT 69.145 33.635 69.315 34.135 ;
        RECT 69.485 33.465 69.800 34.485 ;
        RECT 70.005 34.110 70.295 35.275 ;
        RECT 71.590 34.305 71.920 35.105 ;
        RECT 72.090 34.475 72.420 35.275 ;
        RECT 72.720 34.305 73.050 35.105 ;
        RECT 73.695 34.475 73.945 35.275 ;
        RECT 71.590 34.135 74.025 34.305 ;
        RECT 74.215 34.135 74.385 35.275 ;
        RECT 74.555 34.135 74.895 35.105 ;
        RECT 75.155 34.605 75.325 35.105 ;
        RECT 75.495 34.775 75.825 35.275 ;
        RECT 75.155 34.435 75.820 34.605 ;
        RECT 71.385 33.715 71.735 33.965 ;
        RECT 71.920 33.505 72.090 34.135 ;
        RECT 72.260 33.715 72.590 33.915 ;
        RECT 72.760 33.715 73.090 33.915 ;
        RECT 73.260 33.715 73.680 33.915 ;
        RECT 73.855 33.885 74.025 34.135 ;
        RECT 73.855 33.715 74.550 33.885 ;
        RECT 74.720 33.575 74.895 34.135 ;
        RECT 75.070 33.615 75.420 34.265 ;
        RECT 67.870 32.725 68.110 33.235 ;
        RECT 68.290 32.905 68.570 33.235 ;
        RECT 68.800 32.725 69.015 33.235 ;
        RECT 69.185 32.895 69.800 33.465 ;
        RECT 70.005 32.725 70.295 33.450 ;
        RECT 71.590 32.895 72.090 33.505 ;
        RECT 72.720 33.375 73.945 33.545 ;
        RECT 74.665 33.525 74.895 33.575 ;
        RECT 72.720 32.895 73.050 33.375 ;
        RECT 73.220 32.725 73.445 33.185 ;
        RECT 73.615 32.895 73.945 33.375 ;
        RECT 74.135 32.725 74.385 33.525 ;
        RECT 74.555 32.895 74.895 33.525 ;
        RECT 75.590 33.445 75.820 34.435 ;
        RECT 75.155 33.275 75.820 33.445 ;
        RECT 75.155 32.985 75.325 33.275 ;
        RECT 75.495 32.725 75.825 33.105 ;
        RECT 75.995 32.985 76.180 35.105 ;
        RECT 76.420 34.815 76.685 35.275 ;
        RECT 76.855 34.680 77.105 35.105 ;
        RECT 77.315 34.830 78.420 35.000 ;
        RECT 76.800 34.550 77.105 34.680 ;
        RECT 76.350 33.355 76.630 34.305 ;
        RECT 76.800 33.445 76.970 34.550 ;
        RECT 77.140 33.765 77.380 34.360 ;
        RECT 77.550 34.295 78.080 34.660 ;
        RECT 77.550 33.595 77.720 34.295 ;
        RECT 78.250 34.215 78.420 34.830 ;
        RECT 78.590 34.475 78.760 35.275 ;
        RECT 78.930 34.775 79.180 35.105 ;
        RECT 79.405 34.805 80.290 34.975 ;
        RECT 78.250 34.125 78.760 34.215 ;
        RECT 76.800 33.315 77.025 33.445 ;
        RECT 77.195 33.375 77.720 33.595 ;
        RECT 77.890 33.955 78.760 34.125 ;
        RECT 76.435 32.725 76.685 33.185 ;
        RECT 76.855 33.175 77.025 33.315 ;
        RECT 77.890 33.175 78.060 33.955 ;
        RECT 78.590 33.885 78.760 33.955 ;
        RECT 78.270 33.705 78.470 33.735 ;
        RECT 78.930 33.705 79.100 34.775 ;
        RECT 79.270 33.885 79.460 34.605 ;
        RECT 78.270 33.405 79.100 33.705 ;
        RECT 79.630 33.675 79.950 34.635 ;
        RECT 76.855 33.005 77.190 33.175 ;
        RECT 77.385 33.005 78.060 33.175 ;
        RECT 78.380 32.725 78.750 33.225 ;
        RECT 78.930 33.175 79.100 33.405 ;
        RECT 79.485 33.345 79.950 33.675 ;
        RECT 80.120 33.965 80.290 34.805 ;
        RECT 80.470 34.775 80.785 35.275 ;
        RECT 81.015 34.545 81.355 35.105 ;
        RECT 80.460 34.170 81.355 34.545 ;
        RECT 81.525 34.265 81.695 35.275 ;
        RECT 81.165 33.965 81.355 34.170 ;
        RECT 81.865 34.215 82.195 35.060 ;
        RECT 81.865 34.135 82.255 34.215 ;
        RECT 82.040 34.085 82.255 34.135 ;
        RECT 80.120 33.635 80.995 33.965 ;
        RECT 81.165 33.635 81.915 33.965 ;
        RECT 80.120 33.175 80.290 33.635 ;
        RECT 81.165 33.465 81.365 33.635 ;
        RECT 82.085 33.505 82.255 34.085 ;
        RECT 82.885 34.185 84.095 35.275 ;
        RECT 82.885 33.645 83.405 34.185 ;
        RECT 82.030 33.465 82.255 33.505 ;
        RECT 83.575 33.475 84.095 34.015 ;
        RECT 78.930 33.005 79.335 33.175 ;
        RECT 79.505 33.005 80.290 33.175 ;
        RECT 80.565 32.725 80.775 33.255 ;
        RECT 81.035 32.940 81.365 33.465 ;
        RECT 81.875 33.380 82.255 33.465 ;
        RECT 81.535 32.725 81.705 33.335 ;
        RECT 81.875 32.945 82.205 33.380 ;
        RECT 82.885 32.725 84.095 33.475 ;
        RECT 5.520 32.555 84.180 32.725 ;
        RECT 5.605 31.805 6.815 32.555 ;
        RECT 6.985 32.010 12.330 32.555 ;
        RECT 5.605 31.265 6.125 31.805 ;
        RECT 6.295 31.095 6.815 31.635 ;
        RECT 8.570 31.180 8.910 32.010 ;
        RECT 13.425 31.755 13.765 32.385 ;
        RECT 13.935 31.755 14.185 32.555 ;
        RECT 14.375 31.905 14.705 32.385 ;
        RECT 14.875 32.095 15.100 32.555 ;
        RECT 15.270 31.905 15.600 32.385 ;
        RECT 5.605 30.005 6.815 31.095 ;
        RECT 10.390 30.440 10.740 31.690 ;
        RECT 13.425 31.145 13.600 31.755 ;
        RECT 14.375 31.735 15.600 31.905 ;
        RECT 16.230 31.775 16.730 32.385 ;
        RECT 17.195 32.005 17.365 32.385 ;
        RECT 17.580 32.175 17.910 32.555 ;
        RECT 17.195 31.835 17.910 32.005 ;
        RECT 13.770 31.395 14.465 31.565 ;
        RECT 14.295 31.145 14.465 31.395 ;
        RECT 14.640 31.365 15.060 31.565 ;
        RECT 15.230 31.365 15.560 31.565 ;
        RECT 15.730 31.365 16.060 31.565 ;
        RECT 16.230 31.145 16.400 31.775 ;
        RECT 16.585 31.315 16.935 31.565 ;
        RECT 17.105 31.285 17.460 31.655 ;
        RECT 17.740 31.645 17.910 31.835 ;
        RECT 18.080 31.810 18.335 32.385 ;
        RECT 17.740 31.315 17.995 31.645 ;
        RECT 6.985 30.005 12.330 30.440 ;
        RECT 13.425 30.175 13.765 31.145 ;
        RECT 13.935 30.005 14.105 31.145 ;
        RECT 14.295 30.975 16.730 31.145 ;
        RECT 17.740 31.105 17.910 31.315 ;
        RECT 14.375 30.005 14.625 30.805 ;
        RECT 15.270 30.175 15.600 30.975 ;
        RECT 15.900 30.005 16.230 30.805 ;
        RECT 16.400 30.175 16.730 30.975 ;
        RECT 17.195 30.935 17.910 31.105 ;
        RECT 18.165 31.080 18.335 31.810 ;
        RECT 18.510 31.715 18.770 32.555 ;
        RECT 18.945 31.785 20.615 32.555 ;
        RECT 20.950 32.045 21.190 32.555 ;
        RECT 21.370 32.045 21.650 32.375 ;
        RECT 21.880 32.045 22.095 32.555 ;
        RECT 18.945 31.265 19.695 31.785 ;
        RECT 17.195 30.175 17.365 30.935 ;
        RECT 17.580 30.005 17.910 30.765 ;
        RECT 18.080 30.175 18.335 31.080 ;
        RECT 18.510 30.005 18.770 31.155 ;
        RECT 19.865 31.095 20.615 31.615 ;
        RECT 20.845 31.315 21.200 31.875 ;
        RECT 21.370 31.145 21.540 32.045 ;
        RECT 21.710 31.315 21.975 31.875 ;
        RECT 22.265 31.815 22.880 32.385 ;
        RECT 23.175 32.005 23.345 32.295 ;
        RECT 23.515 32.175 23.845 32.555 ;
        RECT 23.175 31.835 23.840 32.005 ;
        RECT 22.225 31.145 22.395 31.645 ;
        RECT 18.945 30.005 20.615 31.095 ;
        RECT 20.970 30.975 22.395 31.145 ;
        RECT 20.970 30.800 21.360 30.975 ;
        RECT 21.845 30.005 22.175 30.805 ;
        RECT 22.565 30.795 22.880 31.815 ;
        RECT 23.090 31.015 23.440 31.665 ;
        RECT 23.610 30.845 23.840 31.835 ;
        RECT 22.345 30.175 22.880 30.795 ;
        RECT 23.175 30.675 23.840 30.845 ;
        RECT 23.175 30.175 23.345 30.675 ;
        RECT 23.515 30.005 23.845 30.505 ;
        RECT 24.015 30.175 24.200 32.295 ;
        RECT 24.455 32.095 24.705 32.555 ;
        RECT 24.875 32.105 25.210 32.275 ;
        RECT 25.405 32.105 26.080 32.275 ;
        RECT 24.875 31.965 25.045 32.105 ;
        RECT 24.370 30.975 24.650 31.925 ;
        RECT 24.820 31.835 25.045 31.965 ;
        RECT 24.820 30.730 24.990 31.835 ;
        RECT 25.215 31.685 25.740 31.905 ;
        RECT 25.160 30.920 25.400 31.515 ;
        RECT 25.570 30.985 25.740 31.685 ;
        RECT 25.910 31.325 26.080 32.105 ;
        RECT 26.400 32.055 26.770 32.555 ;
        RECT 26.950 32.105 27.355 32.275 ;
        RECT 27.525 32.105 28.310 32.275 ;
        RECT 26.950 31.875 27.120 32.105 ;
        RECT 26.290 31.575 27.120 31.875 ;
        RECT 27.505 31.605 27.970 31.935 ;
        RECT 26.290 31.545 26.490 31.575 ;
        RECT 26.610 31.325 26.780 31.395 ;
        RECT 25.910 31.155 26.780 31.325 ;
        RECT 26.270 31.065 26.780 31.155 ;
        RECT 24.820 30.600 25.125 30.730 ;
        RECT 25.570 30.620 26.100 30.985 ;
        RECT 24.440 30.005 24.705 30.465 ;
        RECT 24.875 30.175 25.125 30.600 ;
        RECT 26.270 30.450 26.440 31.065 ;
        RECT 25.335 30.280 26.440 30.450 ;
        RECT 26.610 30.005 26.780 30.805 ;
        RECT 26.950 30.505 27.120 31.575 ;
        RECT 27.290 30.675 27.480 31.395 ;
        RECT 27.650 30.645 27.970 31.605 ;
        RECT 28.140 31.645 28.310 32.105 ;
        RECT 28.585 32.025 28.795 32.555 ;
        RECT 29.055 31.815 29.385 32.340 ;
        RECT 29.555 31.945 29.725 32.555 ;
        RECT 29.895 31.900 30.225 32.335 ;
        RECT 29.895 31.815 30.275 31.900 ;
        RECT 31.365 31.830 31.655 32.555 ;
        RECT 29.185 31.645 29.385 31.815 ;
        RECT 30.050 31.775 30.275 31.815 ;
        RECT 31.830 31.790 32.285 32.555 ;
        RECT 32.560 32.175 33.860 32.385 ;
        RECT 34.115 32.195 34.445 32.555 ;
        RECT 33.690 32.025 33.860 32.175 ;
        RECT 34.615 32.055 34.875 32.385 ;
        RECT 34.645 32.045 34.875 32.055 ;
        RECT 35.210 32.045 35.450 32.555 ;
        RECT 35.630 32.045 35.910 32.375 ;
        RECT 36.140 32.045 36.355 32.555 ;
        RECT 28.140 31.315 29.015 31.645 ;
        RECT 29.185 31.315 29.935 31.645 ;
        RECT 26.950 30.175 27.200 30.505 ;
        RECT 28.140 30.475 28.310 31.315 ;
        RECT 29.185 31.110 29.375 31.315 ;
        RECT 30.105 31.195 30.275 31.775 ;
        RECT 32.760 31.565 32.980 31.965 ;
        RECT 31.825 31.365 32.315 31.565 ;
        RECT 32.505 31.355 32.980 31.565 ;
        RECT 33.225 31.565 33.435 31.965 ;
        RECT 33.690 31.900 34.445 32.025 ;
        RECT 33.690 31.855 34.535 31.900 ;
        RECT 34.265 31.735 34.535 31.855 ;
        RECT 33.225 31.355 33.555 31.565 ;
        RECT 33.725 31.295 34.135 31.600 ;
        RECT 30.060 31.145 30.275 31.195 ;
        RECT 28.480 30.735 29.375 31.110 ;
        RECT 29.885 31.065 30.275 31.145 ;
        RECT 27.425 30.305 28.310 30.475 ;
        RECT 28.490 30.005 28.805 30.505 ;
        RECT 29.035 30.175 29.375 30.735 ;
        RECT 29.545 30.005 29.715 31.015 ;
        RECT 29.885 30.220 30.215 31.065 ;
        RECT 31.365 30.005 31.655 31.170 ;
        RECT 31.830 31.125 33.005 31.185 ;
        RECT 34.365 31.160 34.535 31.735 ;
        RECT 34.335 31.125 34.535 31.160 ;
        RECT 31.830 31.015 34.535 31.125 ;
        RECT 31.830 30.395 32.085 31.015 ;
        RECT 32.675 30.955 34.475 31.015 ;
        RECT 32.675 30.925 33.005 30.955 ;
        RECT 34.705 30.855 34.875 32.045 ;
        RECT 35.105 31.315 35.460 31.875 ;
        RECT 35.630 31.145 35.800 32.045 ;
        RECT 35.970 31.315 36.235 31.875 ;
        RECT 36.525 31.815 37.140 32.385 ;
        RECT 37.345 32.010 42.690 32.555 ;
        RECT 36.485 31.145 36.655 31.645 ;
        RECT 32.335 30.755 32.520 30.845 ;
        RECT 33.110 30.755 33.945 30.765 ;
        RECT 32.335 30.555 33.945 30.755 ;
        RECT 32.335 30.515 32.565 30.555 ;
        RECT 31.830 30.175 32.165 30.395 ;
        RECT 33.170 30.005 33.525 30.385 ;
        RECT 33.695 30.175 33.945 30.555 ;
        RECT 34.195 30.005 34.445 30.785 ;
        RECT 34.615 30.175 34.875 30.855 ;
        RECT 35.230 30.975 36.655 31.145 ;
        RECT 35.230 30.800 35.620 30.975 ;
        RECT 36.105 30.005 36.435 30.805 ;
        RECT 36.825 30.795 37.140 31.815 ;
        RECT 38.930 31.180 39.270 32.010 ;
        RECT 42.865 31.785 44.535 32.555 ;
        RECT 36.605 30.175 37.140 30.795 ;
        RECT 40.750 30.440 41.100 31.690 ;
        RECT 42.865 31.265 43.615 31.785 ;
        RECT 44.710 31.735 44.985 32.555 ;
        RECT 45.155 31.915 45.485 32.385 ;
        RECT 45.655 32.085 45.825 32.555 ;
        RECT 45.995 31.915 46.325 32.385 ;
        RECT 46.495 32.085 47.205 32.555 ;
        RECT 47.375 31.915 47.705 32.385 ;
        RECT 47.875 32.085 48.165 32.555 ;
        RECT 45.155 31.735 48.215 31.915 ;
        RECT 43.785 31.095 44.535 31.615 ;
        RECT 44.755 31.355 45.585 31.565 ;
        RECT 45.755 31.355 46.805 31.565 ;
        RECT 46.995 31.355 47.585 31.565 ;
        RECT 37.345 30.005 42.690 30.440 ;
        RECT 42.865 30.005 44.535 31.095 ;
        RECT 44.770 31.015 46.705 31.185 ;
        RECT 46.995 31.015 47.260 31.355 ;
        RECT 47.755 31.185 48.215 31.735 ;
        RECT 48.385 31.805 49.595 32.555 ;
        RECT 49.855 32.005 50.025 32.295 ;
        RECT 50.195 32.175 50.525 32.555 ;
        RECT 49.855 31.835 50.520 32.005 ;
        RECT 48.385 31.265 48.905 31.805 ;
        RECT 47.455 31.015 48.215 31.185 ;
        RECT 49.075 31.095 49.595 31.635 ;
        RECT 44.770 30.175 45.025 31.015 ;
        RECT 45.195 30.005 45.445 30.845 ;
        RECT 45.615 30.175 45.865 31.015 ;
        RECT 46.035 30.345 46.285 30.845 ;
        RECT 46.455 30.515 46.705 31.015 ;
        RECT 47.035 30.345 47.245 30.845 ;
        RECT 47.455 30.515 47.665 31.015 ;
        RECT 47.835 30.345 48.085 30.845 ;
        RECT 46.035 30.175 48.085 30.345 ;
        RECT 48.385 30.005 49.595 31.095 ;
        RECT 49.770 31.015 50.120 31.665 ;
        RECT 50.290 30.845 50.520 31.835 ;
        RECT 49.855 30.675 50.520 30.845 ;
        RECT 49.855 30.175 50.025 30.675 ;
        RECT 50.195 30.005 50.525 30.505 ;
        RECT 50.695 30.175 50.880 32.295 ;
        RECT 51.135 32.095 51.385 32.555 ;
        RECT 51.555 32.105 51.890 32.275 ;
        RECT 52.085 32.105 52.760 32.275 ;
        RECT 51.555 31.965 51.725 32.105 ;
        RECT 51.050 30.975 51.330 31.925 ;
        RECT 51.500 31.835 51.725 31.965 ;
        RECT 51.500 30.730 51.670 31.835 ;
        RECT 51.895 31.685 52.420 31.905 ;
        RECT 51.840 30.920 52.080 31.515 ;
        RECT 52.250 30.985 52.420 31.685 ;
        RECT 52.590 31.325 52.760 32.105 ;
        RECT 53.080 32.055 53.450 32.555 ;
        RECT 53.630 32.105 54.035 32.275 ;
        RECT 54.205 32.105 54.990 32.275 ;
        RECT 53.630 31.875 53.800 32.105 ;
        RECT 52.970 31.575 53.800 31.875 ;
        RECT 54.185 31.605 54.650 31.935 ;
        RECT 52.970 31.545 53.170 31.575 ;
        RECT 53.290 31.325 53.460 31.395 ;
        RECT 52.590 31.155 53.460 31.325 ;
        RECT 52.950 31.065 53.460 31.155 ;
        RECT 51.500 30.600 51.805 30.730 ;
        RECT 52.250 30.620 52.780 30.985 ;
        RECT 51.120 30.005 51.385 30.465 ;
        RECT 51.555 30.175 51.805 30.600 ;
        RECT 52.950 30.450 53.120 31.065 ;
        RECT 52.015 30.280 53.120 30.450 ;
        RECT 53.290 30.005 53.460 30.805 ;
        RECT 53.630 30.505 53.800 31.575 ;
        RECT 53.970 30.675 54.160 31.395 ;
        RECT 54.330 30.645 54.650 31.605 ;
        RECT 54.820 31.645 54.990 32.105 ;
        RECT 55.265 32.025 55.475 32.555 ;
        RECT 55.735 31.815 56.065 32.340 ;
        RECT 56.235 31.945 56.405 32.555 ;
        RECT 56.575 31.900 56.905 32.335 ;
        RECT 56.575 31.815 56.955 31.900 ;
        RECT 57.125 31.830 57.415 32.555 ;
        RECT 55.865 31.645 56.065 31.815 ;
        RECT 56.730 31.775 56.955 31.815 ;
        RECT 54.820 31.315 55.695 31.645 ;
        RECT 55.865 31.315 56.615 31.645 ;
        RECT 53.630 30.175 53.880 30.505 ;
        RECT 54.820 30.475 54.990 31.315 ;
        RECT 55.865 31.110 56.055 31.315 ;
        RECT 56.785 31.195 56.955 31.775 ;
        RECT 57.585 31.785 61.095 32.555 ;
        RECT 57.585 31.265 59.235 31.785 ;
        RECT 61.725 31.755 62.015 32.555 ;
        RECT 62.185 32.095 62.735 32.385 ;
        RECT 62.905 32.095 63.155 32.555 ;
        RECT 56.740 31.145 56.955 31.195 ;
        RECT 55.160 30.735 56.055 31.110 ;
        RECT 56.565 31.065 56.955 31.145 ;
        RECT 54.105 30.305 54.990 30.475 ;
        RECT 55.170 30.005 55.485 30.505 ;
        RECT 55.715 30.175 56.055 30.735 ;
        RECT 56.225 30.005 56.395 31.015 ;
        RECT 56.565 30.220 56.895 31.065 ;
        RECT 57.125 30.005 57.415 31.170 ;
        RECT 59.405 31.095 61.095 31.615 ;
        RECT 57.585 30.005 61.095 31.095 ;
        RECT 61.725 30.005 62.015 31.145 ;
        RECT 62.185 30.725 62.435 32.095 ;
        RECT 63.785 31.925 64.115 32.285 ;
        RECT 62.725 31.735 64.115 31.925 ;
        RECT 64.485 31.925 64.825 32.385 ;
        RECT 64.995 32.095 65.165 32.555 ;
        RECT 65.335 32.175 66.505 32.385 ;
        RECT 65.335 31.925 65.585 32.175 ;
        RECT 66.175 32.155 66.505 32.175 ;
        RECT 64.485 31.755 65.585 31.925 ;
        RECT 65.755 31.735 66.615 31.985 ;
        RECT 62.725 31.645 62.895 31.735 ;
        RECT 62.605 31.315 62.895 31.645 ;
        RECT 63.065 31.315 63.395 31.565 ;
        RECT 63.625 31.315 64.315 31.565 ;
        RECT 64.485 31.315 65.245 31.565 ;
        RECT 65.415 31.315 66.165 31.565 ;
        RECT 62.725 31.065 62.895 31.315 ;
        RECT 62.725 30.895 63.665 31.065 ;
        RECT 62.185 30.175 62.635 30.725 ;
        RECT 62.825 30.005 63.155 30.725 ;
        RECT 63.365 30.345 63.665 30.895 ;
        RECT 64.000 30.875 64.315 31.315 ;
        RECT 66.335 31.145 66.615 31.735 ;
        RECT 66.785 31.785 68.455 32.555 ;
        RECT 69.250 32.045 69.490 32.555 ;
        RECT 69.670 32.045 69.950 32.375 ;
        RECT 70.180 32.045 70.395 32.555 ;
        RECT 66.785 31.265 67.535 31.785 ;
        RECT 63.835 30.005 64.115 30.675 ;
        RECT 64.485 30.005 64.745 31.145 ;
        RECT 64.915 30.975 66.615 31.145 ;
        RECT 67.705 31.095 68.455 31.615 ;
        RECT 69.145 31.315 69.500 31.875 ;
        RECT 69.670 31.145 69.840 32.045 ;
        RECT 70.010 31.315 70.275 31.875 ;
        RECT 70.565 31.815 71.180 32.385 ;
        RECT 70.525 31.145 70.695 31.645 ;
        RECT 64.915 30.175 65.245 30.975 ;
        RECT 65.415 30.005 65.585 30.805 ;
        RECT 65.755 30.175 66.085 30.975 ;
        RECT 66.255 30.005 66.510 30.805 ;
        RECT 66.785 30.005 68.455 31.095 ;
        RECT 69.270 30.975 70.695 31.145 ;
        RECT 69.270 30.800 69.660 30.975 ;
        RECT 70.145 30.005 70.475 30.805 ;
        RECT 70.865 30.795 71.180 31.815 ;
        RECT 70.645 30.175 71.180 30.795 ;
        RECT 71.385 32.055 71.645 32.385 ;
        RECT 71.815 32.195 72.145 32.555 ;
        RECT 72.400 32.175 73.700 32.385 ;
        RECT 71.385 30.855 71.555 32.055 ;
        RECT 72.400 32.025 72.570 32.175 ;
        RECT 71.815 31.900 72.570 32.025 ;
        RECT 71.725 31.855 72.570 31.900 ;
        RECT 71.725 31.735 71.995 31.855 ;
        RECT 71.725 31.160 71.895 31.735 ;
        RECT 72.125 31.295 72.535 31.600 ;
        RECT 72.825 31.565 73.035 31.965 ;
        RECT 72.705 31.355 73.035 31.565 ;
        RECT 73.280 31.565 73.500 31.965 ;
        RECT 73.975 31.790 74.430 32.555 ;
        RECT 75.615 32.005 75.785 32.295 ;
        RECT 75.955 32.175 76.285 32.555 ;
        RECT 75.615 31.835 76.280 32.005 ;
        RECT 73.280 31.355 73.755 31.565 ;
        RECT 73.945 31.365 74.435 31.565 ;
        RECT 71.725 31.125 71.925 31.160 ;
        RECT 73.255 31.125 74.430 31.185 ;
        RECT 71.725 31.015 74.430 31.125 ;
        RECT 75.530 31.015 75.880 31.665 ;
        RECT 71.785 30.955 73.585 31.015 ;
        RECT 73.255 30.925 73.585 30.955 ;
        RECT 71.385 30.175 71.645 30.855 ;
        RECT 71.815 30.005 72.065 30.785 ;
        RECT 72.315 30.755 73.150 30.765 ;
        RECT 73.740 30.755 73.925 30.845 ;
        RECT 72.315 30.555 73.925 30.755 ;
        RECT 72.315 30.175 72.565 30.555 ;
        RECT 73.695 30.515 73.925 30.555 ;
        RECT 74.175 30.395 74.430 31.015 ;
        RECT 76.050 30.845 76.280 31.835 ;
        RECT 72.735 30.005 73.090 30.385 ;
        RECT 74.095 30.175 74.430 30.395 ;
        RECT 75.615 30.675 76.280 30.845 ;
        RECT 75.615 30.175 75.785 30.675 ;
        RECT 75.955 30.005 76.285 30.505 ;
        RECT 76.455 30.175 76.640 32.295 ;
        RECT 76.895 32.095 77.145 32.555 ;
        RECT 77.315 32.105 77.650 32.275 ;
        RECT 77.845 32.105 78.520 32.275 ;
        RECT 77.315 31.965 77.485 32.105 ;
        RECT 76.810 30.975 77.090 31.925 ;
        RECT 77.260 31.835 77.485 31.965 ;
        RECT 77.260 30.730 77.430 31.835 ;
        RECT 77.655 31.685 78.180 31.905 ;
        RECT 77.600 30.920 77.840 31.515 ;
        RECT 78.010 30.985 78.180 31.685 ;
        RECT 78.350 31.325 78.520 32.105 ;
        RECT 78.840 32.055 79.210 32.555 ;
        RECT 79.390 32.105 79.795 32.275 ;
        RECT 79.965 32.105 80.750 32.275 ;
        RECT 79.390 31.875 79.560 32.105 ;
        RECT 78.730 31.575 79.560 31.875 ;
        RECT 79.945 31.605 80.410 31.935 ;
        RECT 78.730 31.545 78.930 31.575 ;
        RECT 79.050 31.325 79.220 31.395 ;
        RECT 78.350 31.155 79.220 31.325 ;
        RECT 78.710 31.065 79.220 31.155 ;
        RECT 77.260 30.600 77.565 30.730 ;
        RECT 78.010 30.620 78.540 30.985 ;
        RECT 76.880 30.005 77.145 30.465 ;
        RECT 77.315 30.175 77.565 30.600 ;
        RECT 78.710 30.450 78.880 31.065 ;
        RECT 77.775 30.280 78.880 30.450 ;
        RECT 79.050 30.005 79.220 30.805 ;
        RECT 79.390 30.505 79.560 31.575 ;
        RECT 79.730 30.675 79.920 31.395 ;
        RECT 80.090 30.645 80.410 31.605 ;
        RECT 80.580 31.645 80.750 32.105 ;
        RECT 81.025 32.025 81.235 32.555 ;
        RECT 81.495 31.815 81.825 32.340 ;
        RECT 81.995 31.945 82.165 32.555 ;
        RECT 82.335 31.900 82.665 32.335 ;
        RECT 82.335 31.815 82.715 31.900 ;
        RECT 81.625 31.645 81.825 31.815 ;
        RECT 82.490 31.775 82.715 31.815 ;
        RECT 82.885 31.805 84.095 32.555 ;
        RECT 80.580 31.315 81.455 31.645 ;
        RECT 81.625 31.315 82.375 31.645 ;
        RECT 79.390 30.175 79.640 30.505 ;
        RECT 80.580 30.475 80.750 31.315 ;
        RECT 81.625 31.110 81.815 31.315 ;
        RECT 82.545 31.195 82.715 31.775 ;
        RECT 82.500 31.145 82.715 31.195 ;
        RECT 80.920 30.735 81.815 31.110 ;
        RECT 82.325 31.065 82.715 31.145 ;
        RECT 82.885 31.095 83.405 31.635 ;
        RECT 83.575 31.265 84.095 31.805 ;
        RECT 79.865 30.305 80.750 30.475 ;
        RECT 80.930 30.005 81.245 30.505 ;
        RECT 81.475 30.175 81.815 30.735 ;
        RECT 81.985 30.005 82.155 31.015 ;
        RECT 82.325 30.220 82.655 31.065 ;
        RECT 82.885 30.005 84.095 31.095 ;
        RECT 5.520 29.835 84.180 30.005 ;
        RECT 5.605 28.745 6.815 29.835 ;
        RECT 5.605 28.035 6.125 28.575 ;
        RECT 6.295 28.205 6.815 28.745 ;
        RECT 6.990 28.685 7.250 29.835 ;
        RECT 7.425 28.760 7.680 29.665 ;
        RECT 7.850 29.075 8.180 29.835 ;
        RECT 8.395 28.905 8.565 29.665 ;
        RECT 5.605 27.285 6.815 28.035 ;
        RECT 6.990 27.285 7.250 28.125 ;
        RECT 7.425 28.030 7.595 28.760 ;
        RECT 7.850 28.735 8.565 28.905 ;
        RECT 9.320 29.045 9.855 29.665 ;
        RECT 7.850 28.525 8.020 28.735 ;
        RECT 7.765 28.195 8.020 28.525 ;
        RECT 7.425 27.455 7.680 28.030 ;
        RECT 7.850 28.005 8.020 28.195 ;
        RECT 8.300 28.185 8.655 28.555 ;
        RECT 9.320 28.025 9.635 29.045 ;
        RECT 10.025 29.035 10.355 29.835 ;
        RECT 10.840 28.865 11.230 29.040 ;
        RECT 9.805 28.695 11.230 28.865 ;
        RECT 11.585 28.745 13.255 29.835 ;
        RECT 9.805 28.195 9.975 28.695 ;
        RECT 7.850 27.835 8.565 28.005 ;
        RECT 7.850 27.285 8.180 27.665 ;
        RECT 8.395 27.455 8.565 27.835 ;
        RECT 9.320 27.455 9.935 28.025 ;
        RECT 10.225 27.965 10.490 28.525 ;
        RECT 10.660 27.795 10.830 28.695 ;
        RECT 11.000 27.965 11.355 28.525 ;
        RECT 11.585 28.055 12.335 28.575 ;
        RECT 12.505 28.225 13.255 28.745 ;
        RECT 13.885 28.695 14.225 29.665 ;
        RECT 14.395 28.695 14.565 29.835 ;
        RECT 14.835 29.035 15.085 29.835 ;
        RECT 15.730 28.865 16.060 29.665 ;
        RECT 16.360 29.035 16.690 29.835 ;
        RECT 16.860 28.865 17.190 29.665 ;
        RECT 14.755 28.695 17.190 28.865 ;
        RECT 13.885 28.085 14.060 28.695 ;
        RECT 14.755 28.445 14.925 28.695 ;
        RECT 14.230 28.275 14.925 28.445 ;
        RECT 15.100 28.275 15.520 28.475 ;
        RECT 15.690 28.275 16.020 28.475 ;
        RECT 16.190 28.275 16.520 28.475 ;
        RECT 10.105 27.285 10.320 27.795 ;
        RECT 10.550 27.465 10.830 27.795 ;
        RECT 11.010 27.285 11.250 27.795 ;
        RECT 11.585 27.285 13.255 28.055 ;
        RECT 13.885 27.455 14.225 28.085 ;
        RECT 14.395 27.285 14.645 28.085 ;
        RECT 14.835 27.935 16.060 28.105 ;
        RECT 14.835 27.455 15.165 27.935 ;
        RECT 15.335 27.285 15.560 27.745 ;
        RECT 15.730 27.455 16.060 27.935 ;
        RECT 16.690 28.065 16.860 28.695 ;
        RECT 18.485 28.670 18.775 29.835 ;
        RECT 18.945 29.400 24.290 29.835 ;
        RECT 24.465 29.400 29.810 29.835 ;
        RECT 29.985 29.400 35.330 29.835 ;
        RECT 17.045 28.275 17.395 28.525 ;
        RECT 16.690 27.455 17.190 28.065 ;
        RECT 18.485 27.285 18.775 28.010 ;
        RECT 20.530 27.830 20.870 28.660 ;
        RECT 22.350 28.150 22.700 29.400 ;
        RECT 26.050 27.830 26.390 28.660 ;
        RECT 27.870 28.150 28.220 29.400 ;
        RECT 31.570 27.830 31.910 28.660 ;
        RECT 33.390 28.150 33.740 29.400 ;
        RECT 36.610 28.865 37.000 29.040 ;
        RECT 37.485 29.035 37.815 29.835 ;
        RECT 37.985 29.045 38.520 29.665 ;
        RECT 36.610 28.695 38.035 28.865 ;
        RECT 36.485 27.965 36.840 28.525 ;
        RECT 18.945 27.285 24.290 27.830 ;
        RECT 24.465 27.285 29.810 27.830 ;
        RECT 29.985 27.285 35.330 27.830 ;
        RECT 37.010 27.795 37.180 28.695 ;
        RECT 37.350 27.965 37.615 28.525 ;
        RECT 37.865 28.195 38.035 28.695 ;
        RECT 38.205 28.025 38.520 29.045 ;
        RECT 38.725 28.745 40.395 29.835 ;
        RECT 36.590 27.285 36.830 27.795 ;
        RECT 37.010 27.465 37.290 27.795 ;
        RECT 37.520 27.285 37.735 27.795 ;
        RECT 37.905 27.455 38.520 28.025 ;
        RECT 38.725 28.055 39.475 28.575 ;
        RECT 39.645 28.225 40.395 28.745 ;
        RECT 41.030 29.445 41.365 29.665 ;
        RECT 42.370 29.455 42.725 29.835 ;
        RECT 41.030 28.825 41.285 29.445 ;
        RECT 41.535 29.285 41.765 29.325 ;
        RECT 42.895 29.285 43.145 29.665 ;
        RECT 41.535 29.085 43.145 29.285 ;
        RECT 41.535 28.995 41.720 29.085 ;
        RECT 42.310 29.075 43.145 29.085 ;
        RECT 43.395 29.055 43.645 29.835 ;
        RECT 43.815 28.985 44.075 29.665 ;
        RECT 41.875 28.885 42.205 28.915 ;
        RECT 41.875 28.825 43.675 28.885 ;
        RECT 41.030 28.715 43.735 28.825 ;
        RECT 41.030 28.655 42.205 28.715 ;
        RECT 43.535 28.680 43.735 28.715 ;
        RECT 41.025 28.275 41.515 28.475 ;
        RECT 41.705 28.275 42.180 28.485 ;
        RECT 38.725 27.285 40.395 28.055 ;
        RECT 41.030 27.285 41.485 28.050 ;
        RECT 41.960 27.875 42.180 28.275 ;
        RECT 42.425 28.275 42.755 28.485 ;
        RECT 42.425 27.875 42.635 28.275 ;
        RECT 42.925 28.240 43.335 28.545 ;
        RECT 43.565 28.105 43.735 28.680 ;
        RECT 43.465 27.985 43.735 28.105 ;
        RECT 42.890 27.940 43.735 27.985 ;
        RECT 42.890 27.815 43.645 27.940 ;
        RECT 42.890 27.665 43.060 27.815 ;
        RECT 43.905 27.785 44.075 28.985 ;
        RECT 44.245 28.670 44.535 29.835 ;
        RECT 44.705 28.745 45.915 29.835 ;
        RECT 44.705 28.035 45.225 28.575 ;
        RECT 45.395 28.205 45.915 28.745 ;
        RECT 46.290 28.865 46.620 29.665 ;
        RECT 46.790 29.035 47.120 29.835 ;
        RECT 47.420 28.865 47.750 29.665 ;
        RECT 48.395 29.035 48.645 29.835 ;
        RECT 46.290 28.695 48.725 28.865 ;
        RECT 48.915 28.695 49.085 29.835 ;
        RECT 49.255 28.695 49.595 29.665 ;
        RECT 46.085 28.275 46.435 28.525 ;
        RECT 46.620 28.065 46.790 28.695 ;
        RECT 46.960 28.275 47.290 28.475 ;
        RECT 47.460 28.275 47.790 28.475 ;
        RECT 47.960 28.275 48.380 28.475 ;
        RECT 48.555 28.445 48.725 28.695 ;
        RECT 48.555 28.275 49.250 28.445 ;
        RECT 41.760 27.455 43.060 27.665 ;
        RECT 43.315 27.285 43.645 27.645 ;
        RECT 43.815 27.455 44.075 27.785 ;
        RECT 44.245 27.285 44.535 28.010 ;
        RECT 44.705 27.285 45.915 28.035 ;
        RECT 46.290 27.455 46.790 28.065 ;
        RECT 47.420 27.935 48.645 28.105 ;
        RECT 49.420 28.085 49.595 28.695 ;
        RECT 47.420 27.455 47.750 27.935 ;
        RECT 47.920 27.285 48.145 27.745 ;
        RECT 48.315 27.455 48.645 27.935 ;
        RECT 48.835 27.285 49.085 28.085 ;
        RECT 49.255 27.455 49.595 28.085 ;
        RECT 49.800 29.045 50.335 29.665 ;
        RECT 49.800 28.025 50.115 29.045 ;
        RECT 50.505 29.035 50.835 29.835 ;
        RECT 52.155 29.165 52.325 29.665 ;
        RECT 52.495 29.335 52.825 29.835 ;
        RECT 51.320 28.865 51.710 29.040 ;
        RECT 52.155 28.995 52.820 29.165 ;
        RECT 50.285 28.695 51.710 28.865 ;
        RECT 50.285 28.195 50.455 28.695 ;
        RECT 49.800 27.455 50.415 28.025 ;
        RECT 50.705 27.965 50.970 28.525 ;
        RECT 51.140 27.795 51.310 28.695 ;
        RECT 51.480 27.965 51.835 28.525 ;
        RECT 52.070 28.175 52.420 28.825 ;
        RECT 52.590 28.005 52.820 28.995 ;
        RECT 52.155 27.835 52.820 28.005 ;
        RECT 50.585 27.285 50.800 27.795 ;
        RECT 51.030 27.465 51.310 27.795 ;
        RECT 51.490 27.285 51.730 27.795 ;
        RECT 52.155 27.545 52.325 27.835 ;
        RECT 52.495 27.285 52.825 27.665 ;
        RECT 52.995 27.545 53.180 29.665 ;
        RECT 53.420 29.375 53.685 29.835 ;
        RECT 53.855 29.240 54.105 29.665 ;
        RECT 54.315 29.390 55.420 29.560 ;
        RECT 53.800 29.110 54.105 29.240 ;
        RECT 53.350 27.915 53.630 28.865 ;
        RECT 53.800 28.005 53.970 29.110 ;
        RECT 54.140 28.325 54.380 28.920 ;
        RECT 54.550 28.855 55.080 29.220 ;
        RECT 54.550 28.155 54.720 28.855 ;
        RECT 55.250 28.775 55.420 29.390 ;
        RECT 55.590 29.035 55.760 29.835 ;
        RECT 55.930 29.335 56.180 29.665 ;
        RECT 56.405 29.365 57.290 29.535 ;
        RECT 55.250 28.685 55.760 28.775 ;
        RECT 53.800 27.875 54.025 28.005 ;
        RECT 54.195 27.935 54.720 28.155 ;
        RECT 54.890 28.515 55.760 28.685 ;
        RECT 53.435 27.285 53.685 27.745 ;
        RECT 53.855 27.735 54.025 27.875 ;
        RECT 54.890 27.735 55.060 28.515 ;
        RECT 55.590 28.445 55.760 28.515 ;
        RECT 55.270 28.265 55.470 28.295 ;
        RECT 55.930 28.265 56.100 29.335 ;
        RECT 56.270 28.445 56.460 29.165 ;
        RECT 55.270 27.965 56.100 28.265 ;
        RECT 56.630 28.235 56.950 29.195 ;
        RECT 53.855 27.565 54.190 27.735 ;
        RECT 54.385 27.565 55.060 27.735 ;
        RECT 55.380 27.285 55.750 27.785 ;
        RECT 55.930 27.735 56.100 27.965 ;
        RECT 56.485 27.905 56.950 28.235 ;
        RECT 57.120 28.525 57.290 29.365 ;
        RECT 57.470 29.335 57.785 29.835 ;
        RECT 58.015 29.105 58.355 29.665 ;
        RECT 57.460 28.730 58.355 29.105 ;
        RECT 58.525 28.825 58.695 29.835 ;
        RECT 58.165 28.525 58.355 28.730 ;
        RECT 58.865 28.775 59.195 29.620 ;
        RECT 59.460 29.045 59.995 29.665 ;
        RECT 58.865 28.695 59.255 28.775 ;
        RECT 59.040 28.645 59.255 28.695 ;
        RECT 57.120 28.195 57.995 28.525 ;
        RECT 58.165 28.195 58.915 28.525 ;
        RECT 57.120 27.735 57.290 28.195 ;
        RECT 58.165 28.025 58.365 28.195 ;
        RECT 59.085 28.065 59.255 28.645 ;
        RECT 59.030 28.025 59.255 28.065 ;
        RECT 55.930 27.565 56.335 27.735 ;
        RECT 56.505 27.565 57.290 27.735 ;
        RECT 57.565 27.285 57.775 27.815 ;
        RECT 58.035 27.500 58.365 28.025 ;
        RECT 58.875 27.940 59.255 28.025 ;
        RECT 59.460 28.025 59.775 29.045 ;
        RECT 60.165 29.035 60.495 29.835 ;
        RECT 61.815 29.165 61.985 29.665 ;
        RECT 62.155 29.335 62.485 29.835 ;
        RECT 60.980 28.865 61.370 29.040 ;
        RECT 61.815 28.995 62.480 29.165 ;
        RECT 59.945 28.695 61.370 28.865 ;
        RECT 59.945 28.195 60.115 28.695 ;
        RECT 58.535 27.285 58.705 27.895 ;
        RECT 58.875 27.505 59.205 27.940 ;
        RECT 59.460 27.455 60.075 28.025 ;
        RECT 60.365 27.965 60.630 28.525 ;
        RECT 60.800 27.795 60.970 28.695 ;
        RECT 61.140 27.965 61.495 28.525 ;
        RECT 61.730 28.175 62.080 28.825 ;
        RECT 62.250 28.005 62.480 28.995 ;
        RECT 61.815 27.835 62.480 28.005 ;
        RECT 60.245 27.285 60.460 27.795 ;
        RECT 60.690 27.465 60.970 27.795 ;
        RECT 61.150 27.285 61.390 27.795 ;
        RECT 61.815 27.545 61.985 27.835 ;
        RECT 62.155 27.285 62.485 27.665 ;
        RECT 62.655 27.545 62.840 29.665 ;
        RECT 63.080 29.375 63.345 29.835 ;
        RECT 63.515 29.240 63.765 29.665 ;
        RECT 63.975 29.390 65.080 29.560 ;
        RECT 63.460 29.110 63.765 29.240 ;
        RECT 63.010 27.915 63.290 28.865 ;
        RECT 63.460 28.005 63.630 29.110 ;
        RECT 63.800 28.325 64.040 28.920 ;
        RECT 64.210 28.855 64.740 29.220 ;
        RECT 64.210 28.155 64.380 28.855 ;
        RECT 64.910 28.775 65.080 29.390 ;
        RECT 65.250 29.035 65.420 29.835 ;
        RECT 65.590 29.335 65.840 29.665 ;
        RECT 66.065 29.365 66.950 29.535 ;
        RECT 64.910 28.685 65.420 28.775 ;
        RECT 63.460 27.875 63.685 28.005 ;
        RECT 63.855 27.935 64.380 28.155 ;
        RECT 64.550 28.515 65.420 28.685 ;
        RECT 63.095 27.285 63.345 27.745 ;
        RECT 63.515 27.735 63.685 27.875 ;
        RECT 64.550 27.735 64.720 28.515 ;
        RECT 65.250 28.445 65.420 28.515 ;
        RECT 64.930 28.265 65.130 28.295 ;
        RECT 65.590 28.265 65.760 29.335 ;
        RECT 65.930 28.445 66.120 29.165 ;
        RECT 64.930 27.965 65.760 28.265 ;
        RECT 66.290 28.235 66.610 29.195 ;
        RECT 63.515 27.565 63.850 27.735 ;
        RECT 64.045 27.565 64.720 27.735 ;
        RECT 65.040 27.285 65.410 27.785 ;
        RECT 65.590 27.735 65.760 27.965 ;
        RECT 66.145 27.905 66.610 28.235 ;
        RECT 66.780 28.525 66.950 29.365 ;
        RECT 67.130 29.335 67.445 29.835 ;
        RECT 67.675 29.105 68.015 29.665 ;
        RECT 67.120 28.730 68.015 29.105 ;
        RECT 68.185 28.825 68.355 29.835 ;
        RECT 67.825 28.525 68.015 28.730 ;
        RECT 68.525 28.775 68.855 29.620 ;
        RECT 68.525 28.695 68.915 28.775 ;
        RECT 68.700 28.645 68.915 28.695 ;
        RECT 70.005 28.670 70.295 29.835 ;
        RECT 71.110 28.865 71.500 29.040 ;
        RECT 71.985 29.035 72.315 29.835 ;
        RECT 72.485 29.045 73.020 29.665 ;
        RECT 73.225 29.400 78.570 29.835 ;
        RECT 71.110 28.695 72.535 28.865 ;
        RECT 66.780 28.195 67.655 28.525 ;
        RECT 67.825 28.195 68.575 28.525 ;
        RECT 66.780 27.735 66.950 28.195 ;
        RECT 67.825 28.025 68.025 28.195 ;
        RECT 68.745 28.065 68.915 28.645 ;
        RECT 68.690 28.025 68.915 28.065 ;
        RECT 65.590 27.565 65.995 27.735 ;
        RECT 66.165 27.565 66.950 27.735 ;
        RECT 67.225 27.285 67.435 27.815 ;
        RECT 67.695 27.500 68.025 28.025 ;
        RECT 68.535 27.940 68.915 28.025 ;
        RECT 68.195 27.285 68.365 27.895 ;
        RECT 68.535 27.505 68.865 27.940 ;
        RECT 70.005 27.285 70.295 28.010 ;
        RECT 70.985 27.965 71.340 28.525 ;
        RECT 71.510 27.795 71.680 28.695 ;
        RECT 71.850 27.965 72.115 28.525 ;
        RECT 72.365 28.195 72.535 28.695 ;
        RECT 72.705 28.025 73.020 29.045 ;
        RECT 71.090 27.285 71.330 27.795 ;
        RECT 71.510 27.465 71.790 27.795 ;
        RECT 72.020 27.285 72.235 27.795 ;
        RECT 72.405 27.455 73.020 28.025 ;
        RECT 74.810 27.830 75.150 28.660 ;
        RECT 76.630 28.150 76.980 29.400 ;
        RECT 78.745 28.745 80.415 29.835 ;
        RECT 78.745 28.055 79.495 28.575 ;
        RECT 79.665 28.225 80.415 28.745 ;
        RECT 81.135 28.905 81.305 29.665 ;
        RECT 81.520 29.075 81.850 29.835 ;
        RECT 81.135 28.735 81.850 28.905 ;
        RECT 82.020 28.760 82.275 29.665 ;
        RECT 81.045 28.185 81.400 28.555 ;
        RECT 81.680 28.525 81.850 28.735 ;
        RECT 81.680 28.195 81.935 28.525 ;
        RECT 73.225 27.285 78.570 27.830 ;
        RECT 78.745 27.285 80.415 28.055 ;
        RECT 81.680 28.005 81.850 28.195 ;
        RECT 82.105 28.030 82.275 28.760 ;
        RECT 82.450 28.685 82.710 29.835 ;
        RECT 82.885 28.745 84.095 29.835 ;
        RECT 82.885 28.205 83.405 28.745 ;
        RECT 81.135 27.835 81.850 28.005 ;
        RECT 81.135 27.455 81.305 27.835 ;
        RECT 81.520 27.285 81.850 27.665 ;
        RECT 82.020 27.455 82.275 28.030 ;
        RECT 82.450 27.285 82.710 28.125 ;
        RECT 83.575 28.035 84.095 28.575 ;
        RECT 82.885 27.285 84.095 28.035 ;
        RECT 5.520 27.115 84.180 27.285 ;
        RECT 5.605 26.365 6.815 27.115 ;
        RECT 5.605 25.825 6.125 26.365 ;
        RECT 7.445 26.315 7.785 26.945 ;
        RECT 7.955 26.315 8.205 27.115 ;
        RECT 8.395 26.465 8.725 26.945 ;
        RECT 8.895 26.655 9.120 27.115 ;
        RECT 9.290 26.465 9.620 26.945 ;
        RECT 6.295 25.655 6.815 26.195 ;
        RECT 5.605 24.565 6.815 25.655 ;
        RECT 7.445 25.705 7.620 26.315 ;
        RECT 8.395 26.295 9.620 26.465 ;
        RECT 10.250 26.335 10.750 26.945 ;
        RECT 11.215 26.565 11.385 26.855 ;
        RECT 11.555 26.735 11.885 27.115 ;
        RECT 11.215 26.395 11.880 26.565 ;
        RECT 7.790 25.955 8.485 26.125 ;
        RECT 8.315 25.705 8.485 25.955 ;
        RECT 8.660 25.925 9.080 26.125 ;
        RECT 9.250 25.925 9.580 26.125 ;
        RECT 9.750 25.925 10.080 26.125 ;
        RECT 10.250 25.705 10.420 26.335 ;
        RECT 10.605 25.875 10.955 26.125 ;
        RECT 7.445 24.735 7.785 25.705 ;
        RECT 7.955 24.565 8.125 25.705 ;
        RECT 8.315 25.535 10.750 25.705 ;
        RECT 11.130 25.575 11.480 26.225 ;
        RECT 8.395 24.565 8.645 25.365 ;
        RECT 9.290 24.735 9.620 25.535 ;
        RECT 9.920 24.565 10.250 25.365 ;
        RECT 10.420 24.735 10.750 25.535 ;
        RECT 11.650 25.405 11.880 26.395 ;
        RECT 11.215 25.235 11.880 25.405 ;
        RECT 11.215 24.735 11.385 25.235 ;
        RECT 11.555 24.565 11.885 25.065 ;
        RECT 12.055 24.735 12.240 26.855 ;
        RECT 12.495 26.655 12.745 27.115 ;
        RECT 12.915 26.665 13.250 26.835 ;
        RECT 13.445 26.665 14.120 26.835 ;
        RECT 12.915 26.525 13.085 26.665 ;
        RECT 12.410 25.535 12.690 26.485 ;
        RECT 12.860 26.395 13.085 26.525 ;
        RECT 12.860 25.290 13.030 26.395 ;
        RECT 13.255 26.245 13.780 26.465 ;
        RECT 13.200 25.480 13.440 26.075 ;
        RECT 13.610 25.545 13.780 26.245 ;
        RECT 13.950 25.885 14.120 26.665 ;
        RECT 14.440 26.615 14.810 27.115 ;
        RECT 14.990 26.665 15.395 26.835 ;
        RECT 15.565 26.665 16.350 26.835 ;
        RECT 14.990 26.435 15.160 26.665 ;
        RECT 14.330 26.135 15.160 26.435 ;
        RECT 15.545 26.165 16.010 26.495 ;
        RECT 14.330 26.105 14.530 26.135 ;
        RECT 14.650 25.885 14.820 25.955 ;
        RECT 13.950 25.715 14.820 25.885 ;
        RECT 14.310 25.625 14.820 25.715 ;
        RECT 12.860 25.160 13.165 25.290 ;
        RECT 13.610 25.180 14.140 25.545 ;
        RECT 12.480 24.565 12.745 25.025 ;
        RECT 12.915 24.735 13.165 25.160 ;
        RECT 14.310 25.010 14.480 25.625 ;
        RECT 13.375 24.840 14.480 25.010 ;
        RECT 14.650 24.565 14.820 25.365 ;
        RECT 14.990 25.065 15.160 26.135 ;
        RECT 15.330 25.235 15.520 25.955 ;
        RECT 15.690 25.205 16.010 26.165 ;
        RECT 16.180 26.205 16.350 26.665 ;
        RECT 16.625 26.585 16.835 27.115 ;
        RECT 17.095 26.375 17.425 26.900 ;
        RECT 17.595 26.505 17.765 27.115 ;
        RECT 17.935 26.460 18.265 26.895 ;
        RECT 17.935 26.375 18.315 26.460 ;
        RECT 17.225 26.205 17.425 26.375 ;
        RECT 18.090 26.335 18.315 26.375 ;
        RECT 16.180 25.875 17.055 26.205 ;
        RECT 17.225 25.875 17.975 26.205 ;
        RECT 14.990 24.735 15.240 25.065 ;
        RECT 16.180 25.035 16.350 25.875 ;
        RECT 17.225 25.670 17.415 25.875 ;
        RECT 18.145 25.755 18.315 26.335 ;
        RECT 18.100 25.705 18.315 25.755 ;
        RECT 16.520 25.295 17.415 25.670 ;
        RECT 17.925 25.625 18.315 25.705 ;
        RECT 18.520 26.375 19.135 26.945 ;
        RECT 19.305 26.605 19.520 27.115 ;
        RECT 19.750 26.605 20.030 26.935 ;
        RECT 20.210 26.605 20.450 27.115 ;
        RECT 15.465 24.865 16.350 25.035 ;
        RECT 16.530 24.565 16.845 25.065 ;
        RECT 17.075 24.735 17.415 25.295 ;
        RECT 17.585 24.565 17.755 25.575 ;
        RECT 17.925 24.780 18.255 25.625 ;
        RECT 18.520 25.355 18.835 26.375 ;
        RECT 19.005 25.705 19.175 26.205 ;
        RECT 19.425 25.875 19.690 26.435 ;
        RECT 19.860 25.705 20.030 26.605 ;
        RECT 20.200 25.875 20.555 26.435 ;
        RECT 21.245 26.315 21.585 26.945 ;
        RECT 21.755 26.315 22.005 27.115 ;
        RECT 22.195 26.465 22.525 26.945 ;
        RECT 22.695 26.655 22.920 27.115 ;
        RECT 23.090 26.465 23.420 26.945 ;
        RECT 21.245 25.705 21.420 26.315 ;
        RECT 22.195 26.295 23.420 26.465 ;
        RECT 24.050 26.335 24.550 26.945 ;
        RECT 25.590 26.335 26.090 26.945 ;
        RECT 21.590 25.955 22.285 26.125 ;
        RECT 22.115 25.705 22.285 25.955 ;
        RECT 22.460 25.925 22.880 26.125 ;
        RECT 23.050 25.925 23.380 26.125 ;
        RECT 23.550 25.925 23.880 26.125 ;
        RECT 24.050 25.705 24.220 26.335 ;
        RECT 24.405 25.875 24.755 26.125 ;
        RECT 25.385 25.875 25.735 26.125 ;
        RECT 25.920 25.705 26.090 26.335 ;
        RECT 26.720 26.465 27.050 26.945 ;
        RECT 27.220 26.655 27.445 27.115 ;
        RECT 27.615 26.465 27.945 26.945 ;
        RECT 26.720 26.295 27.945 26.465 ;
        RECT 28.135 26.315 28.385 27.115 ;
        RECT 28.555 26.315 28.895 26.945 ;
        RECT 29.230 26.605 29.470 27.115 ;
        RECT 29.650 26.605 29.930 26.935 ;
        RECT 30.160 26.605 30.375 27.115 ;
        RECT 26.260 25.925 26.590 26.125 ;
        RECT 26.760 25.925 27.090 26.125 ;
        RECT 27.260 25.925 27.680 26.125 ;
        RECT 27.855 25.955 28.550 26.125 ;
        RECT 27.855 25.705 28.025 25.955 ;
        RECT 28.720 25.705 28.895 26.315 ;
        RECT 29.125 25.875 29.480 26.435 ;
        RECT 29.650 25.705 29.820 26.605 ;
        RECT 29.990 25.875 30.255 26.435 ;
        RECT 30.545 26.375 31.160 26.945 ;
        RECT 31.365 26.390 31.655 27.115 ;
        RECT 30.505 25.705 30.675 26.205 ;
        RECT 19.005 25.535 20.430 25.705 ;
        RECT 18.520 24.735 19.055 25.355 ;
        RECT 19.225 24.565 19.555 25.365 ;
        RECT 20.040 25.360 20.430 25.535 ;
        RECT 21.245 24.735 21.585 25.705 ;
        RECT 21.755 24.565 21.925 25.705 ;
        RECT 22.115 25.535 24.550 25.705 ;
        RECT 22.195 24.565 22.445 25.365 ;
        RECT 23.090 24.735 23.420 25.535 ;
        RECT 23.720 24.565 24.050 25.365 ;
        RECT 24.220 24.735 24.550 25.535 ;
        RECT 25.590 25.535 28.025 25.705 ;
        RECT 25.590 24.735 25.920 25.535 ;
        RECT 26.090 24.565 26.420 25.365 ;
        RECT 26.720 24.735 27.050 25.535 ;
        RECT 27.695 24.565 27.945 25.365 ;
        RECT 28.215 24.565 28.385 25.705 ;
        RECT 28.555 24.735 28.895 25.705 ;
        RECT 29.250 25.535 30.675 25.705 ;
        RECT 29.250 25.360 29.640 25.535 ;
        RECT 30.125 24.565 30.455 25.365 ;
        RECT 30.845 25.355 31.160 26.375 ;
        RECT 31.825 26.345 34.415 27.115 ;
        RECT 34.675 26.565 34.845 26.855 ;
        RECT 35.015 26.735 35.345 27.115 ;
        RECT 34.675 26.395 35.340 26.565 ;
        RECT 31.825 25.825 33.035 26.345 ;
        RECT 30.625 24.735 31.160 25.355 ;
        RECT 31.365 24.565 31.655 25.730 ;
        RECT 33.205 25.655 34.415 26.175 ;
        RECT 31.825 24.565 34.415 25.655 ;
        RECT 34.590 25.575 34.940 26.225 ;
        RECT 35.110 25.405 35.340 26.395 ;
        RECT 34.675 25.235 35.340 25.405 ;
        RECT 34.675 24.735 34.845 25.235 ;
        RECT 35.015 24.565 35.345 25.065 ;
        RECT 35.515 24.735 35.700 26.855 ;
        RECT 35.955 26.655 36.205 27.115 ;
        RECT 36.375 26.665 36.710 26.835 ;
        RECT 36.905 26.665 37.580 26.835 ;
        RECT 36.375 26.525 36.545 26.665 ;
        RECT 35.870 25.535 36.150 26.485 ;
        RECT 36.320 26.395 36.545 26.525 ;
        RECT 36.320 25.290 36.490 26.395 ;
        RECT 36.715 26.245 37.240 26.465 ;
        RECT 36.660 25.480 36.900 26.075 ;
        RECT 37.070 25.545 37.240 26.245 ;
        RECT 37.410 25.885 37.580 26.665 ;
        RECT 37.900 26.615 38.270 27.115 ;
        RECT 38.450 26.665 38.855 26.835 ;
        RECT 39.025 26.665 39.810 26.835 ;
        RECT 38.450 26.435 38.620 26.665 ;
        RECT 37.790 26.135 38.620 26.435 ;
        RECT 39.005 26.165 39.470 26.495 ;
        RECT 37.790 26.105 37.990 26.135 ;
        RECT 38.110 25.885 38.280 25.955 ;
        RECT 37.410 25.715 38.280 25.885 ;
        RECT 37.770 25.625 38.280 25.715 ;
        RECT 36.320 25.160 36.625 25.290 ;
        RECT 37.070 25.180 37.600 25.545 ;
        RECT 35.940 24.565 36.205 25.025 ;
        RECT 36.375 24.735 36.625 25.160 ;
        RECT 37.770 25.010 37.940 25.625 ;
        RECT 36.835 24.840 37.940 25.010 ;
        RECT 38.110 24.565 38.280 25.365 ;
        RECT 38.450 25.065 38.620 26.135 ;
        RECT 38.790 25.235 38.980 25.955 ;
        RECT 39.150 25.205 39.470 26.165 ;
        RECT 39.640 26.205 39.810 26.665 ;
        RECT 40.085 26.585 40.295 27.115 ;
        RECT 40.555 26.375 40.885 26.900 ;
        RECT 41.055 26.505 41.225 27.115 ;
        RECT 41.395 26.460 41.725 26.895 ;
        RECT 41.395 26.375 41.775 26.460 ;
        RECT 40.685 26.205 40.885 26.375 ;
        RECT 41.550 26.335 41.775 26.375 ;
        RECT 39.640 25.875 40.515 26.205 ;
        RECT 40.685 25.875 41.435 26.205 ;
        RECT 38.450 24.735 38.700 25.065 ;
        RECT 39.640 25.035 39.810 25.875 ;
        RECT 40.685 25.670 40.875 25.875 ;
        RECT 41.605 25.755 41.775 26.335 ;
        RECT 41.945 26.365 43.155 27.115 ;
        RECT 43.415 26.565 43.585 26.855 ;
        RECT 43.755 26.735 44.085 27.115 ;
        RECT 43.415 26.395 44.080 26.565 ;
        RECT 41.945 25.825 42.465 26.365 ;
        RECT 41.560 25.705 41.775 25.755 ;
        RECT 39.980 25.295 40.875 25.670 ;
        RECT 41.385 25.625 41.775 25.705 ;
        RECT 42.635 25.655 43.155 26.195 ;
        RECT 38.925 24.865 39.810 25.035 ;
        RECT 39.990 24.565 40.305 25.065 ;
        RECT 40.535 24.735 40.875 25.295 ;
        RECT 41.045 24.565 41.215 25.575 ;
        RECT 41.385 24.780 41.715 25.625 ;
        RECT 41.945 24.565 43.155 25.655 ;
        RECT 43.330 25.575 43.680 26.225 ;
        RECT 43.850 25.405 44.080 26.395 ;
        RECT 43.415 25.235 44.080 25.405 ;
        RECT 43.415 24.735 43.585 25.235 ;
        RECT 43.755 24.565 44.085 25.065 ;
        RECT 44.255 24.735 44.440 26.855 ;
        RECT 44.695 26.655 44.945 27.115 ;
        RECT 45.115 26.665 45.450 26.835 ;
        RECT 45.645 26.665 46.320 26.835 ;
        RECT 45.115 26.525 45.285 26.665 ;
        RECT 44.610 25.535 44.890 26.485 ;
        RECT 45.060 26.395 45.285 26.525 ;
        RECT 45.060 25.290 45.230 26.395 ;
        RECT 45.455 26.245 45.980 26.465 ;
        RECT 45.400 25.480 45.640 26.075 ;
        RECT 45.810 25.545 45.980 26.245 ;
        RECT 46.150 25.885 46.320 26.665 ;
        RECT 46.640 26.615 47.010 27.115 ;
        RECT 47.190 26.665 47.595 26.835 ;
        RECT 47.765 26.665 48.550 26.835 ;
        RECT 47.190 26.435 47.360 26.665 ;
        RECT 46.530 26.135 47.360 26.435 ;
        RECT 47.745 26.165 48.210 26.495 ;
        RECT 46.530 26.105 46.730 26.135 ;
        RECT 46.850 25.885 47.020 25.955 ;
        RECT 46.150 25.715 47.020 25.885 ;
        RECT 46.510 25.625 47.020 25.715 ;
        RECT 45.060 25.160 45.365 25.290 ;
        RECT 45.810 25.180 46.340 25.545 ;
        RECT 44.680 24.565 44.945 25.025 ;
        RECT 45.115 24.735 45.365 25.160 ;
        RECT 46.510 25.010 46.680 25.625 ;
        RECT 45.575 24.840 46.680 25.010 ;
        RECT 46.850 24.565 47.020 25.365 ;
        RECT 47.190 25.065 47.360 26.135 ;
        RECT 47.530 25.235 47.720 25.955 ;
        RECT 47.890 25.205 48.210 26.165 ;
        RECT 48.380 26.205 48.550 26.665 ;
        RECT 48.825 26.585 49.035 27.115 ;
        RECT 49.295 26.375 49.625 26.900 ;
        RECT 49.795 26.505 49.965 27.115 ;
        RECT 50.135 26.460 50.465 26.895 ;
        RECT 50.135 26.375 50.515 26.460 ;
        RECT 49.425 26.205 49.625 26.375 ;
        RECT 50.290 26.335 50.515 26.375 ;
        RECT 48.380 25.875 49.255 26.205 ;
        RECT 49.425 25.875 50.175 26.205 ;
        RECT 47.190 24.735 47.440 25.065 ;
        RECT 48.380 25.035 48.550 25.875 ;
        RECT 49.425 25.670 49.615 25.875 ;
        RECT 50.345 25.755 50.515 26.335 ;
        RECT 50.300 25.705 50.515 25.755 ;
        RECT 48.720 25.295 49.615 25.670 ;
        RECT 50.125 25.625 50.515 25.705 ;
        RECT 51.145 26.315 51.485 26.945 ;
        RECT 51.655 26.315 51.905 27.115 ;
        RECT 52.095 26.465 52.425 26.945 ;
        RECT 52.595 26.655 52.820 27.115 ;
        RECT 52.990 26.465 53.320 26.945 ;
        RECT 51.145 25.705 51.320 26.315 ;
        RECT 52.095 26.295 53.320 26.465 ;
        RECT 53.950 26.335 54.450 26.945 ;
        RECT 54.860 26.375 55.475 26.945 ;
        RECT 55.645 26.605 55.860 27.115 ;
        RECT 56.090 26.605 56.370 26.935 ;
        RECT 56.550 26.605 56.790 27.115 ;
        RECT 51.490 25.955 52.185 26.125 ;
        RECT 52.015 25.705 52.185 25.955 ;
        RECT 52.360 25.925 52.780 26.125 ;
        RECT 52.950 25.925 53.280 26.125 ;
        RECT 53.450 25.925 53.780 26.125 ;
        RECT 53.950 25.705 54.120 26.335 ;
        RECT 54.305 25.875 54.655 26.125 ;
        RECT 47.665 24.865 48.550 25.035 ;
        RECT 48.730 24.565 49.045 25.065 ;
        RECT 49.275 24.735 49.615 25.295 ;
        RECT 49.785 24.565 49.955 25.575 ;
        RECT 50.125 24.780 50.455 25.625 ;
        RECT 51.145 24.735 51.485 25.705 ;
        RECT 51.655 24.565 51.825 25.705 ;
        RECT 52.015 25.535 54.450 25.705 ;
        RECT 52.095 24.565 52.345 25.365 ;
        RECT 52.990 24.735 53.320 25.535 ;
        RECT 53.620 24.565 53.950 25.365 ;
        RECT 54.120 24.735 54.450 25.535 ;
        RECT 54.860 25.355 55.175 26.375 ;
        RECT 55.345 25.705 55.515 26.205 ;
        RECT 55.765 25.875 56.030 26.435 ;
        RECT 56.200 25.705 56.370 26.605 ;
        RECT 56.540 25.875 56.895 26.435 ;
        RECT 57.125 26.390 57.415 27.115 ;
        RECT 58.505 26.615 58.765 26.945 ;
        RECT 58.935 26.755 59.265 27.115 ;
        RECT 59.520 26.735 60.820 26.945 ;
        RECT 58.505 26.605 58.735 26.615 ;
        RECT 55.345 25.535 56.770 25.705 ;
        RECT 54.860 24.735 55.395 25.355 ;
        RECT 55.565 24.565 55.895 25.365 ;
        RECT 56.380 25.360 56.770 25.535 ;
        RECT 57.125 24.565 57.415 25.730 ;
        RECT 58.505 25.415 58.675 26.605 ;
        RECT 59.520 26.585 59.690 26.735 ;
        RECT 58.935 26.460 59.690 26.585 ;
        RECT 58.845 26.415 59.690 26.460 ;
        RECT 58.845 26.295 59.115 26.415 ;
        RECT 58.845 25.720 59.015 26.295 ;
        RECT 59.245 25.855 59.655 26.160 ;
        RECT 59.945 26.125 60.155 26.525 ;
        RECT 59.825 25.915 60.155 26.125 ;
        RECT 60.400 26.125 60.620 26.525 ;
        RECT 61.095 26.350 61.550 27.115 ;
        RECT 61.930 26.335 62.430 26.945 ;
        RECT 60.400 25.915 60.875 26.125 ;
        RECT 61.065 25.925 61.555 26.125 ;
        RECT 61.725 25.875 62.075 26.125 ;
        RECT 58.845 25.685 59.045 25.720 ;
        RECT 60.375 25.685 61.550 25.745 ;
        RECT 62.260 25.705 62.430 26.335 ;
        RECT 63.060 26.465 63.390 26.945 ;
        RECT 63.560 26.655 63.785 27.115 ;
        RECT 63.955 26.465 64.285 26.945 ;
        RECT 63.060 26.295 64.285 26.465 ;
        RECT 64.475 26.315 64.725 27.115 ;
        RECT 64.895 26.315 65.235 26.945 ;
        RECT 62.600 25.925 62.930 26.125 ;
        RECT 63.100 25.925 63.430 26.125 ;
        RECT 63.600 25.925 64.020 26.125 ;
        RECT 64.195 25.955 64.890 26.125 ;
        RECT 64.195 25.705 64.365 25.955 ;
        RECT 65.060 25.705 65.235 26.315 ;
        RECT 65.405 26.345 67.075 27.115 ;
        RECT 67.795 26.565 67.965 26.855 ;
        RECT 68.135 26.735 68.465 27.115 ;
        RECT 67.795 26.395 68.460 26.565 ;
        RECT 65.405 25.825 66.155 26.345 ;
        RECT 58.845 25.575 61.550 25.685 ;
        RECT 58.905 25.515 60.705 25.575 ;
        RECT 60.375 25.485 60.705 25.515 ;
        RECT 58.505 24.735 58.765 25.415 ;
        RECT 58.935 24.565 59.185 25.345 ;
        RECT 59.435 25.315 60.270 25.325 ;
        RECT 60.860 25.315 61.045 25.405 ;
        RECT 59.435 25.115 61.045 25.315 ;
        RECT 59.435 24.735 59.685 25.115 ;
        RECT 60.815 25.075 61.045 25.115 ;
        RECT 61.295 24.955 61.550 25.575 ;
        RECT 59.855 24.565 60.210 24.945 ;
        RECT 61.215 24.735 61.550 24.955 ;
        RECT 61.930 25.535 64.365 25.705 ;
        RECT 61.930 24.735 62.260 25.535 ;
        RECT 62.430 24.565 62.760 25.365 ;
        RECT 63.060 24.735 63.390 25.535 ;
        RECT 64.035 24.565 64.285 25.365 ;
        RECT 64.555 24.565 64.725 25.705 ;
        RECT 64.895 24.735 65.235 25.705 ;
        RECT 66.325 25.655 67.075 26.175 ;
        RECT 65.405 24.565 67.075 25.655 ;
        RECT 67.710 25.575 68.060 26.225 ;
        RECT 68.230 25.405 68.460 26.395 ;
        RECT 67.795 25.235 68.460 25.405 ;
        RECT 67.795 24.735 67.965 25.235 ;
        RECT 68.135 24.565 68.465 25.065 ;
        RECT 68.635 24.735 68.820 26.855 ;
        RECT 69.075 26.655 69.325 27.115 ;
        RECT 69.495 26.665 69.830 26.835 ;
        RECT 70.025 26.665 70.700 26.835 ;
        RECT 69.495 26.525 69.665 26.665 ;
        RECT 68.990 25.535 69.270 26.485 ;
        RECT 69.440 26.395 69.665 26.525 ;
        RECT 69.440 25.290 69.610 26.395 ;
        RECT 69.835 26.245 70.360 26.465 ;
        RECT 69.780 25.480 70.020 26.075 ;
        RECT 70.190 25.545 70.360 26.245 ;
        RECT 70.530 25.885 70.700 26.665 ;
        RECT 71.020 26.615 71.390 27.115 ;
        RECT 71.570 26.665 71.975 26.835 ;
        RECT 72.145 26.665 72.930 26.835 ;
        RECT 71.570 26.435 71.740 26.665 ;
        RECT 70.910 26.135 71.740 26.435 ;
        RECT 72.125 26.165 72.590 26.495 ;
        RECT 70.910 26.105 71.110 26.135 ;
        RECT 71.230 25.885 71.400 25.955 ;
        RECT 70.530 25.715 71.400 25.885 ;
        RECT 70.890 25.625 71.400 25.715 ;
        RECT 69.440 25.160 69.745 25.290 ;
        RECT 70.190 25.180 70.720 25.545 ;
        RECT 69.060 24.565 69.325 25.025 ;
        RECT 69.495 24.735 69.745 25.160 ;
        RECT 70.890 25.010 71.060 25.625 ;
        RECT 69.955 24.840 71.060 25.010 ;
        RECT 71.230 24.565 71.400 25.365 ;
        RECT 71.570 25.065 71.740 26.135 ;
        RECT 71.910 25.235 72.100 25.955 ;
        RECT 72.270 25.205 72.590 26.165 ;
        RECT 72.760 26.205 72.930 26.665 ;
        RECT 73.205 26.585 73.415 27.115 ;
        RECT 73.675 26.375 74.005 26.900 ;
        RECT 74.175 26.505 74.345 27.115 ;
        RECT 74.515 26.460 74.845 26.895 ;
        RECT 75.065 26.615 75.325 26.945 ;
        RECT 75.495 26.755 75.825 27.115 ;
        RECT 76.080 26.735 77.380 26.945 ;
        RECT 74.515 26.375 74.895 26.460 ;
        RECT 73.805 26.205 74.005 26.375 ;
        RECT 74.670 26.335 74.895 26.375 ;
        RECT 72.760 25.875 73.635 26.205 ;
        RECT 73.805 25.875 74.555 26.205 ;
        RECT 71.570 24.735 71.820 25.065 ;
        RECT 72.760 25.035 72.930 25.875 ;
        RECT 73.805 25.670 73.995 25.875 ;
        RECT 74.725 25.755 74.895 26.335 ;
        RECT 74.680 25.705 74.895 25.755 ;
        RECT 73.100 25.295 73.995 25.670 ;
        RECT 74.505 25.625 74.895 25.705 ;
        RECT 72.045 24.865 72.930 25.035 ;
        RECT 73.110 24.565 73.425 25.065 ;
        RECT 73.655 24.735 73.995 25.295 ;
        RECT 74.165 24.565 74.335 25.575 ;
        RECT 74.505 24.780 74.835 25.625 ;
        RECT 75.065 25.415 75.235 26.615 ;
        RECT 76.080 26.585 76.250 26.735 ;
        RECT 75.495 26.460 76.250 26.585 ;
        RECT 75.405 26.415 76.250 26.460 ;
        RECT 75.405 26.295 75.675 26.415 ;
        RECT 75.405 25.720 75.575 26.295 ;
        RECT 75.805 25.855 76.215 26.160 ;
        RECT 76.505 26.125 76.715 26.525 ;
        RECT 76.385 25.915 76.715 26.125 ;
        RECT 76.960 26.125 77.180 26.525 ;
        RECT 77.655 26.350 78.110 27.115 ;
        RECT 78.285 26.345 81.795 27.115 ;
        RECT 82.885 26.365 84.095 27.115 ;
        RECT 76.960 25.915 77.435 26.125 ;
        RECT 77.625 25.925 78.115 26.125 ;
        RECT 78.285 25.825 79.935 26.345 ;
        RECT 75.405 25.685 75.605 25.720 ;
        RECT 76.935 25.685 78.110 25.745 ;
        RECT 75.405 25.575 78.110 25.685 ;
        RECT 80.105 25.655 81.795 26.175 ;
        RECT 75.465 25.515 77.265 25.575 ;
        RECT 76.935 25.485 77.265 25.515 ;
        RECT 75.065 24.735 75.325 25.415 ;
        RECT 75.495 24.565 75.745 25.345 ;
        RECT 75.995 25.315 76.830 25.325 ;
        RECT 77.420 25.315 77.605 25.405 ;
        RECT 75.995 25.115 77.605 25.315 ;
        RECT 75.995 24.735 76.245 25.115 ;
        RECT 77.375 25.075 77.605 25.115 ;
        RECT 77.855 24.955 78.110 25.575 ;
        RECT 76.415 24.565 76.770 24.945 ;
        RECT 77.775 24.735 78.110 24.955 ;
        RECT 78.285 24.565 81.795 25.655 ;
        RECT 82.885 25.655 83.405 26.195 ;
        RECT 83.575 25.825 84.095 26.365 ;
        RECT 82.885 24.565 84.095 25.655 ;
        RECT 5.520 24.395 84.180 24.565 ;
        RECT 5.605 23.305 6.815 24.395 ;
        RECT 7.075 23.725 7.245 24.225 ;
        RECT 7.415 23.895 7.745 24.395 ;
        RECT 7.075 23.555 7.740 23.725 ;
        RECT 5.605 22.595 6.125 23.135 ;
        RECT 6.295 22.765 6.815 23.305 ;
        RECT 6.990 22.735 7.340 23.385 ;
        RECT 5.605 21.845 6.815 22.595 ;
        RECT 7.510 22.565 7.740 23.555 ;
        RECT 7.075 22.395 7.740 22.565 ;
        RECT 7.075 22.105 7.245 22.395 ;
        RECT 7.415 21.845 7.745 22.225 ;
        RECT 7.915 22.105 8.100 24.225 ;
        RECT 8.340 23.935 8.605 24.395 ;
        RECT 8.775 23.800 9.025 24.225 ;
        RECT 9.235 23.950 10.340 24.120 ;
        RECT 8.720 23.670 9.025 23.800 ;
        RECT 8.270 22.475 8.550 23.425 ;
        RECT 8.720 22.565 8.890 23.670 ;
        RECT 9.060 22.885 9.300 23.480 ;
        RECT 9.470 23.415 10.000 23.780 ;
        RECT 9.470 22.715 9.640 23.415 ;
        RECT 10.170 23.335 10.340 23.950 ;
        RECT 10.510 23.595 10.680 24.395 ;
        RECT 10.850 23.895 11.100 24.225 ;
        RECT 11.325 23.925 12.210 24.095 ;
        RECT 10.170 23.245 10.680 23.335 ;
        RECT 8.720 22.435 8.945 22.565 ;
        RECT 9.115 22.495 9.640 22.715 ;
        RECT 9.810 23.075 10.680 23.245 ;
        RECT 8.355 21.845 8.605 22.305 ;
        RECT 8.775 22.295 8.945 22.435 ;
        RECT 9.810 22.295 9.980 23.075 ;
        RECT 10.510 23.005 10.680 23.075 ;
        RECT 10.190 22.825 10.390 22.855 ;
        RECT 10.850 22.825 11.020 23.895 ;
        RECT 11.190 23.005 11.380 23.725 ;
        RECT 10.190 22.525 11.020 22.825 ;
        RECT 11.550 22.795 11.870 23.755 ;
        RECT 8.775 22.125 9.110 22.295 ;
        RECT 9.305 22.125 9.980 22.295 ;
        RECT 10.300 21.845 10.670 22.345 ;
        RECT 10.850 22.295 11.020 22.525 ;
        RECT 11.405 22.465 11.870 22.795 ;
        RECT 12.040 23.085 12.210 23.925 ;
        RECT 12.390 23.895 12.705 24.395 ;
        RECT 12.935 23.665 13.275 24.225 ;
        RECT 12.380 23.290 13.275 23.665 ;
        RECT 13.445 23.385 13.615 24.395 ;
        RECT 13.085 23.085 13.275 23.290 ;
        RECT 13.785 23.335 14.115 24.180 ;
        RECT 14.350 24.005 14.685 24.225 ;
        RECT 15.690 24.015 16.045 24.395 ;
        RECT 14.350 23.385 14.605 24.005 ;
        RECT 14.855 23.845 15.085 23.885 ;
        RECT 16.215 23.845 16.465 24.225 ;
        RECT 14.855 23.645 16.465 23.845 ;
        RECT 14.855 23.555 15.040 23.645 ;
        RECT 15.630 23.635 16.465 23.645 ;
        RECT 16.715 23.615 16.965 24.395 ;
        RECT 17.135 23.545 17.395 24.225 ;
        RECT 15.195 23.445 15.525 23.475 ;
        RECT 15.195 23.385 16.995 23.445 ;
        RECT 13.785 23.255 14.175 23.335 ;
        RECT 13.960 23.205 14.175 23.255 ;
        RECT 14.350 23.275 17.055 23.385 ;
        RECT 14.350 23.215 15.525 23.275 ;
        RECT 16.855 23.240 17.055 23.275 ;
        RECT 12.040 22.755 12.915 23.085 ;
        RECT 13.085 22.755 13.835 23.085 ;
        RECT 12.040 22.295 12.210 22.755 ;
        RECT 13.085 22.585 13.285 22.755 ;
        RECT 14.005 22.625 14.175 23.205 ;
        RECT 14.345 22.835 14.835 23.035 ;
        RECT 15.025 22.835 15.500 23.045 ;
        RECT 13.950 22.585 14.175 22.625 ;
        RECT 10.850 22.125 11.255 22.295 ;
        RECT 11.425 22.125 12.210 22.295 ;
        RECT 12.485 21.845 12.695 22.375 ;
        RECT 12.955 22.060 13.285 22.585 ;
        RECT 13.795 22.500 14.175 22.585 ;
        RECT 13.455 21.845 13.625 22.455 ;
        RECT 13.795 22.065 14.125 22.500 ;
        RECT 14.350 21.845 14.805 22.610 ;
        RECT 15.280 22.435 15.500 22.835 ;
        RECT 15.745 22.835 16.075 23.045 ;
        RECT 15.745 22.435 15.955 22.835 ;
        RECT 16.245 22.800 16.655 23.105 ;
        RECT 16.885 22.665 17.055 23.240 ;
        RECT 16.785 22.545 17.055 22.665 ;
        RECT 16.210 22.500 17.055 22.545 ;
        RECT 16.210 22.375 16.965 22.500 ;
        RECT 16.210 22.225 16.380 22.375 ;
        RECT 17.225 22.345 17.395 23.545 ;
        RECT 18.485 23.230 18.775 24.395 ;
        RECT 18.945 23.305 20.155 24.395 ;
        RECT 20.415 23.725 20.585 24.225 ;
        RECT 20.755 23.895 21.085 24.395 ;
        RECT 20.415 23.555 21.080 23.725 ;
        RECT 18.945 22.595 19.465 23.135 ;
        RECT 19.635 22.765 20.155 23.305 ;
        RECT 20.330 22.735 20.680 23.385 ;
        RECT 15.080 22.015 16.380 22.225 ;
        RECT 16.635 21.845 16.965 22.205 ;
        RECT 17.135 22.015 17.395 22.345 ;
        RECT 18.485 21.845 18.775 22.570 ;
        RECT 18.945 21.845 20.155 22.595 ;
        RECT 20.850 22.565 21.080 23.555 ;
        RECT 20.415 22.395 21.080 22.565 ;
        RECT 20.415 22.105 20.585 22.395 ;
        RECT 20.755 21.845 21.085 22.225 ;
        RECT 21.255 22.105 21.440 24.225 ;
        RECT 21.680 23.935 21.945 24.395 ;
        RECT 22.115 23.800 22.365 24.225 ;
        RECT 22.575 23.950 23.680 24.120 ;
        RECT 22.060 23.670 22.365 23.800 ;
        RECT 21.610 22.475 21.890 23.425 ;
        RECT 22.060 22.565 22.230 23.670 ;
        RECT 22.400 22.885 22.640 23.480 ;
        RECT 22.810 23.415 23.340 23.780 ;
        RECT 22.810 22.715 22.980 23.415 ;
        RECT 23.510 23.335 23.680 23.950 ;
        RECT 23.850 23.595 24.020 24.395 ;
        RECT 24.190 23.895 24.440 24.225 ;
        RECT 24.665 23.925 25.550 24.095 ;
        RECT 23.510 23.245 24.020 23.335 ;
        RECT 22.060 22.435 22.285 22.565 ;
        RECT 22.455 22.495 22.980 22.715 ;
        RECT 23.150 23.075 24.020 23.245 ;
        RECT 21.695 21.845 21.945 22.305 ;
        RECT 22.115 22.295 22.285 22.435 ;
        RECT 23.150 22.295 23.320 23.075 ;
        RECT 23.850 23.005 24.020 23.075 ;
        RECT 23.530 22.825 23.730 22.855 ;
        RECT 24.190 22.825 24.360 23.895 ;
        RECT 24.530 23.005 24.720 23.725 ;
        RECT 23.530 22.525 24.360 22.825 ;
        RECT 24.890 22.795 25.210 23.755 ;
        RECT 22.115 22.125 22.450 22.295 ;
        RECT 22.645 22.125 23.320 22.295 ;
        RECT 23.640 21.845 24.010 22.345 ;
        RECT 24.190 22.295 24.360 22.525 ;
        RECT 24.745 22.465 25.210 22.795 ;
        RECT 25.380 23.085 25.550 23.925 ;
        RECT 25.730 23.895 26.045 24.395 ;
        RECT 26.275 23.665 26.615 24.225 ;
        RECT 25.720 23.290 26.615 23.665 ;
        RECT 26.785 23.385 26.955 24.395 ;
        RECT 26.425 23.085 26.615 23.290 ;
        RECT 27.125 23.335 27.455 24.180 ;
        RECT 27.775 23.725 27.945 24.225 ;
        RECT 28.115 23.895 28.445 24.395 ;
        RECT 27.775 23.555 28.440 23.725 ;
        RECT 27.125 23.255 27.515 23.335 ;
        RECT 27.300 23.205 27.515 23.255 ;
        RECT 25.380 22.755 26.255 23.085 ;
        RECT 26.425 22.755 27.175 23.085 ;
        RECT 25.380 22.295 25.550 22.755 ;
        RECT 26.425 22.585 26.625 22.755 ;
        RECT 27.345 22.625 27.515 23.205 ;
        RECT 27.690 22.735 28.040 23.385 ;
        RECT 27.290 22.585 27.515 22.625 ;
        RECT 24.190 22.125 24.595 22.295 ;
        RECT 24.765 22.125 25.550 22.295 ;
        RECT 25.825 21.845 26.035 22.375 ;
        RECT 26.295 22.060 26.625 22.585 ;
        RECT 27.135 22.500 27.515 22.585 ;
        RECT 28.210 22.565 28.440 23.555 ;
        RECT 26.795 21.845 26.965 22.455 ;
        RECT 27.135 22.065 27.465 22.500 ;
        RECT 27.775 22.395 28.440 22.565 ;
        RECT 27.775 22.105 27.945 22.395 ;
        RECT 28.115 21.845 28.445 22.225 ;
        RECT 28.615 22.105 28.800 24.225 ;
        RECT 29.040 23.935 29.305 24.395 ;
        RECT 29.475 23.800 29.725 24.225 ;
        RECT 29.935 23.950 31.040 24.120 ;
        RECT 29.420 23.670 29.725 23.800 ;
        RECT 28.970 22.475 29.250 23.425 ;
        RECT 29.420 22.565 29.590 23.670 ;
        RECT 29.760 22.885 30.000 23.480 ;
        RECT 30.170 23.415 30.700 23.780 ;
        RECT 30.170 22.715 30.340 23.415 ;
        RECT 30.870 23.335 31.040 23.950 ;
        RECT 31.210 23.595 31.380 24.395 ;
        RECT 31.550 23.895 31.800 24.225 ;
        RECT 32.025 23.925 32.910 24.095 ;
        RECT 30.870 23.245 31.380 23.335 ;
        RECT 29.420 22.435 29.645 22.565 ;
        RECT 29.815 22.495 30.340 22.715 ;
        RECT 30.510 23.075 31.380 23.245 ;
        RECT 29.055 21.845 29.305 22.305 ;
        RECT 29.475 22.295 29.645 22.435 ;
        RECT 30.510 22.295 30.680 23.075 ;
        RECT 31.210 23.005 31.380 23.075 ;
        RECT 30.890 22.825 31.090 22.855 ;
        RECT 31.550 22.825 31.720 23.895 ;
        RECT 31.890 23.005 32.080 23.725 ;
        RECT 30.890 22.525 31.720 22.825 ;
        RECT 32.250 22.795 32.570 23.755 ;
        RECT 29.475 22.125 29.810 22.295 ;
        RECT 30.005 22.125 30.680 22.295 ;
        RECT 31.000 21.845 31.370 22.345 ;
        RECT 31.550 22.295 31.720 22.525 ;
        RECT 32.105 22.465 32.570 22.795 ;
        RECT 32.740 23.085 32.910 23.925 ;
        RECT 33.090 23.895 33.405 24.395 ;
        RECT 33.635 23.665 33.975 24.225 ;
        RECT 33.080 23.290 33.975 23.665 ;
        RECT 34.145 23.385 34.315 24.395 ;
        RECT 33.785 23.085 33.975 23.290 ;
        RECT 34.485 23.335 34.815 24.180 ;
        RECT 34.485 23.255 34.875 23.335 ;
        RECT 34.660 23.205 34.875 23.255 ;
        RECT 32.740 22.755 33.615 23.085 ;
        RECT 33.785 22.755 34.535 23.085 ;
        RECT 32.740 22.295 32.910 22.755 ;
        RECT 33.785 22.585 33.985 22.755 ;
        RECT 34.705 22.625 34.875 23.205 ;
        RECT 34.650 22.585 34.875 22.625 ;
        RECT 31.550 22.125 31.955 22.295 ;
        RECT 32.125 22.125 32.910 22.295 ;
        RECT 33.185 21.845 33.395 22.375 ;
        RECT 33.655 22.060 33.985 22.585 ;
        RECT 34.495 22.500 34.875 22.585 ;
        RECT 35.965 23.255 36.305 24.225 ;
        RECT 36.475 23.255 36.645 24.395 ;
        RECT 36.915 23.595 37.165 24.395 ;
        RECT 37.810 23.425 38.140 24.225 ;
        RECT 38.440 23.595 38.770 24.395 ;
        RECT 38.940 23.425 39.270 24.225 ;
        RECT 36.835 23.255 39.270 23.425 ;
        RECT 39.645 23.305 41.315 24.395 ;
        RECT 35.965 22.645 36.140 23.255 ;
        RECT 36.835 23.005 37.005 23.255 ;
        RECT 36.310 22.835 37.005 23.005 ;
        RECT 37.180 22.835 37.600 23.035 ;
        RECT 37.770 22.835 38.100 23.035 ;
        RECT 38.270 22.835 38.600 23.035 ;
        RECT 34.155 21.845 34.325 22.455 ;
        RECT 34.495 22.065 34.825 22.500 ;
        RECT 35.965 22.015 36.305 22.645 ;
        RECT 36.475 21.845 36.725 22.645 ;
        RECT 36.915 22.495 38.140 22.665 ;
        RECT 36.915 22.015 37.245 22.495 ;
        RECT 37.415 21.845 37.640 22.305 ;
        RECT 37.810 22.015 38.140 22.495 ;
        RECT 38.770 22.625 38.940 23.255 ;
        RECT 39.125 22.835 39.475 23.085 ;
        RECT 38.770 22.015 39.270 22.625 ;
        RECT 39.645 22.615 40.395 23.135 ;
        RECT 40.565 22.785 41.315 23.305 ;
        RECT 42.130 23.425 42.520 23.600 ;
        RECT 43.005 23.595 43.335 24.395 ;
        RECT 43.505 23.605 44.040 24.225 ;
        RECT 42.130 23.255 43.555 23.425 ;
        RECT 39.645 21.845 41.315 22.615 ;
        RECT 42.005 22.525 42.360 23.085 ;
        RECT 42.530 22.355 42.700 23.255 ;
        RECT 42.870 22.525 43.135 23.085 ;
        RECT 43.385 22.755 43.555 23.255 ;
        RECT 43.725 22.585 44.040 23.605 ;
        RECT 44.245 23.230 44.535 24.395 ;
        RECT 44.705 23.255 45.045 24.225 ;
        RECT 45.215 23.255 45.385 24.395 ;
        RECT 45.655 23.595 45.905 24.395 ;
        RECT 46.550 23.425 46.880 24.225 ;
        RECT 47.180 23.595 47.510 24.395 ;
        RECT 47.680 23.425 48.010 24.225 ;
        RECT 45.575 23.255 48.010 23.425 ;
        RECT 48.385 23.305 50.055 24.395 ;
        RECT 42.110 21.845 42.350 22.355 ;
        RECT 42.530 22.025 42.810 22.355 ;
        RECT 43.040 21.845 43.255 22.355 ;
        RECT 43.425 22.015 44.040 22.585 ;
        RECT 44.705 22.645 44.880 23.255 ;
        RECT 45.575 23.005 45.745 23.255 ;
        RECT 45.050 22.835 45.745 23.005 ;
        RECT 45.920 22.835 46.340 23.035 ;
        RECT 46.510 22.835 46.840 23.035 ;
        RECT 47.010 22.835 47.340 23.035 ;
        RECT 44.245 21.845 44.535 22.570 ;
        RECT 44.705 22.015 45.045 22.645 ;
        RECT 45.215 21.845 45.465 22.645 ;
        RECT 45.655 22.495 46.880 22.665 ;
        RECT 45.655 22.015 45.985 22.495 ;
        RECT 46.155 21.845 46.380 22.305 ;
        RECT 46.550 22.015 46.880 22.495 ;
        RECT 47.510 22.625 47.680 23.255 ;
        RECT 47.865 22.835 48.215 23.085 ;
        RECT 47.510 22.015 48.010 22.625 ;
        RECT 48.385 22.615 49.135 23.135 ;
        RECT 49.305 22.785 50.055 23.305 ;
        RECT 50.230 23.245 50.490 24.395 ;
        RECT 50.665 23.320 50.920 24.225 ;
        RECT 51.090 23.635 51.420 24.395 ;
        RECT 51.635 23.465 51.805 24.225 ;
        RECT 52.065 23.960 57.410 24.395 ;
        RECT 57.585 23.960 62.930 24.395 ;
        RECT 48.385 21.845 50.055 22.615 ;
        RECT 50.230 21.845 50.490 22.685 ;
        RECT 50.665 22.590 50.835 23.320 ;
        RECT 51.090 23.295 51.805 23.465 ;
        RECT 51.090 23.085 51.260 23.295 ;
        RECT 51.005 22.755 51.260 23.085 ;
        RECT 50.665 22.015 50.920 22.590 ;
        RECT 51.090 22.565 51.260 22.755 ;
        RECT 51.540 22.745 51.895 23.115 ;
        RECT 51.090 22.395 51.805 22.565 ;
        RECT 51.090 21.845 51.420 22.225 ;
        RECT 51.635 22.015 51.805 22.395 ;
        RECT 53.650 22.390 53.990 23.220 ;
        RECT 55.470 22.710 55.820 23.960 ;
        RECT 59.170 22.390 59.510 23.220 ;
        RECT 60.990 22.710 61.340 23.960 ;
        RECT 63.105 23.305 66.615 24.395 ;
        RECT 63.105 22.615 64.755 23.135 ;
        RECT 64.925 22.785 66.615 23.305 ;
        RECT 67.890 23.425 68.280 23.600 ;
        RECT 68.765 23.595 69.095 24.395 ;
        RECT 69.265 23.605 69.800 24.225 ;
        RECT 67.890 23.255 69.315 23.425 ;
        RECT 52.065 21.845 57.410 22.390 ;
        RECT 57.585 21.845 62.930 22.390 ;
        RECT 63.105 21.845 66.615 22.615 ;
        RECT 67.765 22.525 68.120 23.085 ;
        RECT 68.290 22.355 68.460 23.255 ;
        RECT 68.630 22.525 68.895 23.085 ;
        RECT 69.145 22.755 69.315 23.255 ;
        RECT 69.485 22.585 69.800 23.605 ;
        RECT 70.005 23.230 70.295 24.395 ;
        RECT 70.465 23.255 70.805 24.225 ;
        RECT 70.975 23.255 71.145 24.395 ;
        RECT 71.415 23.595 71.665 24.395 ;
        RECT 72.310 23.425 72.640 24.225 ;
        RECT 72.940 23.595 73.270 24.395 ;
        RECT 73.440 23.425 73.770 24.225 ;
        RECT 71.335 23.255 73.770 23.425 ;
        RECT 74.145 23.305 75.355 24.395 ;
        RECT 75.615 23.725 75.785 24.225 ;
        RECT 75.955 23.895 76.285 24.395 ;
        RECT 75.615 23.555 76.280 23.725 ;
        RECT 67.870 21.845 68.110 22.355 ;
        RECT 68.290 22.025 68.570 22.355 ;
        RECT 68.800 21.845 69.015 22.355 ;
        RECT 69.185 22.015 69.800 22.585 ;
        RECT 70.465 22.645 70.640 23.255 ;
        RECT 71.335 23.005 71.505 23.255 ;
        RECT 70.810 22.835 71.505 23.005 ;
        RECT 71.680 22.835 72.100 23.035 ;
        RECT 72.270 22.835 72.600 23.035 ;
        RECT 72.770 22.835 73.100 23.035 ;
        RECT 70.005 21.845 70.295 22.570 ;
        RECT 70.465 22.015 70.805 22.645 ;
        RECT 70.975 21.845 71.225 22.645 ;
        RECT 71.415 22.495 72.640 22.665 ;
        RECT 71.415 22.015 71.745 22.495 ;
        RECT 71.915 21.845 72.140 22.305 ;
        RECT 72.310 22.015 72.640 22.495 ;
        RECT 73.270 22.625 73.440 23.255 ;
        RECT 73.625 22.835 73.975 23.085 ;
        RECT 73.270 22.015 73.770 22.625 ;
        RECT 74.145 22.595 74.665 23.135 ;
        RECT 74.835 22.765 75.355 23.305 ;
        RECT 75.530 22.735 75.880 23.385 ;
        RECT 74.145 21.845 75.355 22.595 ;
        RECT 76.050 22.565 76.280 23.555 ;
        RECT 75.615 22.395 76.280 22.565 ;
        RECT 75.615 22.105 75.785 22.395 ;
        RECT 75.955 21.845 76.285 22.225 ;
        RECT 76.455 22.105 76.640 24.225 ;
        RECT 76.880 23.935 77.145 24.395 ;
        RECT 77.315 23.800 77.565 24.225 ;
        RECT 77.775 23.950 78.880 24.120 ;
        RECT 77.260 23.670 77.565 23.800 ;
        RECT 76.810 22.475 77.090 23.425 ;
        RECT 77.260 22.565 77.430 23.670 ;
        RECT 77.600 22.885 77.840 23.480 ;
        RECT 78.010 23.415 78.540 23.780 ;
        RECT 78.010 22.715 78.180 23.415 ;
        RECT 78.710 23.335 78.880 23.950 ;
        RECT 79.050 23.595 79.220 24.395 ;
        RECT 79.390 23.895 79.640 24.225 ;
        RECT 79.865 23.925 80.750 24.095 ;
        RECT 78.710 23.245 79.220 23.335 ;
        RECT 77.260 22.435 77.485 22.565 ;
        RECT 77.655 22.495 78.180 22.715 ;
        RECT 78.350 23.075 79.220 23.245 ;
        RECT 76.895 21.845 77.145 22.305 ;
        RECT 77.315 22.295 77.485 22.435 ;
        RECT 78.350 22.295 78.520 23.075 ;
        RECT 79.050 23.005 79.220 23.075 ;
        RECT 78.730 22.825 78.930 22.855 ;
        RECT 79.390 22.825 79.560 23.895 ;
        RECT 79.730 23.005 79.920 23.725 ;
        RECT 78.730 22.525 79.560 22.825 ;
        RECT 80.090 22.795 80.410 23.755 ;
        RECT 77.315 22.125 77.650 22.295 ;
        RECT 77.845 22.125 78.520 22.295 ;
        RECT 78.840 21.845 79.210 22.345 ;
        RECT 79.390 22.295 79.560 22.525 ;
        RECT 79.945 22.465 80.410 22.795 ;
        RECT 80.580 23.085 80.750 23.925 ;
        RECT 80.930 23.895 81.245 24.395 ;
        RECT 81.475 23.665 81.815 24.225 ;
        RECT 80.920 23.290 81.815 23.665 ;
        RECT 81.985 23.385 82.155 24.395 ;
        RECT 81.625 23.085 81.815 23.290 ;
        RECT 82.325 23.335 82.655 24.180 ;
        RECT 82.325 23.255 82.715 23.335 ;
        RECT 82.500 23.205 82.715 23.255 ;
        RECT 80.580 22.755 81.455 23.085 ;
        RECT 81.625 22.755 82.375 23.085 ;
        RECT 80.580 22.295 80.750 22.755 ;
        RECT 81.625 22.585 81.825 22.755 ;
        RECT 82.545 22.625 82.715 23.205 ;
        RECT 82.885 23.305 84.095 24.395 ;
        RECT 82.885 22.765 83.405 23.305 ;
        RECT 82.490 22.585 82.715 22.625 ;
        RECT 83.575 22.595 84.095 23.135 ;
        RECT 79.390 22.125 79.795 22.295 ;
        RECT 79.965 22.125 80.750 22.295 ;
        RECT 81.025 21.845 81.235 22.375 ;
        RECT 81.495 22.060 81.825 22.585 ;
        RECT 82.335 22.500 82.715 22.585 ;
        RECT 81.995 21.845 82.165 22.455 ;
        RECT 82.335 22.065 82.665 22.500 ;
        RECT 82.885 21.845 84.095 22.595 ;
        RECT 5.520 21.675 84.180 21.845 ;
        RECT 5.605 20.925 6.815 21.675 ;
        RECT 5.605 20.385 6.125 20.925 ;
        RECT 6.990 20.835 7.250 21.675 ;
        RECT 7.425 20.930 7.680 21.505 ;
        RECT 7.850 21.295 8.180 21.675 ;
        RECT 8.395 21.125 8.565 21.505 ;
        RECT 7.850 20.955 8.565 21.125 ;
        RECT 6.295 20.215 6.815 20.755 ;
        RECT 5.605 19.125 6.815 20.215 ;
        RECT 6.990 19.125 7.250 20.275 ;
        RECT 7.425 20.200 7.595 20.930 ;
        RECT 7.850 20.765 8.020 20.955 ;
        RECT 8.825 20.925 10.035 21.675 ;
        RECT 7.765 20.435 8.020 20.765 ;
        RECT 7.850 20.225 8.020 20.435 ;
        RECT 8.300 20.405 8.655 20.775 ;
        RECT 8.825 20.385 9.345 20.925 ;
        RECT 10.210 20.835 10.470 21.675 ;
        RECT 10.645 20.930 10.900 21.505 ;
        RECT 11.070 21.295 11.400 21.675 ;
        RECT 11.615 21.125 11.785 21.505 ;
        RECT 11.070 20.955 11.785 21.125 ;
        RECT 7.425 19.295 7.680 20.200 ;
        RECT 7.850 20.055 8.565 20.225 ;
        RECT 9.515 20.215 10.035 20.755 ;
        RECT 7.850 19.125 8.180 19.885 ;
        RECT 8.395 19.295 8.565 20.055 ;
        RECT 8.825 19.125 10.035 20.215 ;
        RECT 10.210 19.125 10.470 20.275 ;
        RECT 10.645 20.200 10.815 20.930 ;
        RECT 11.070 20.765 11.240 20.955 ;
        RECT 12.050 20.835 12.310 21.675 ;
        RECT 12.485 20.930 12.740 21.505 ;
        RECT 12.910 21.295 13.240 21.675 ;
        RECT 13.455 21.125 13.625 21.505 ;
        RECT 12.910 20.955 13.625 21.125 ;
        RECT 10.985 20.435 11.240 20.765 ;
        RECT 11.070 20.225 11.240 20.435 ;
        RECT 11.520 20.405 11.875 20.775 ;
        RECT 10.645 19.295 10.900 20.200 ;
        RECT 11.070 20.055 11.785 20.225 ;
        RECT 11.070 19.125 11.400 19.885 ;
        RECT 11.615 19.295 11.785 20.055 ;
        RECT 12.050 19.125 12.310 20.275 ;
        RECT 12.485 20.200 12.655 20.930 ;
        RECT 12.910 20.765 13.080 20.955 ;
        RECT 14.810 20.910 15.265 21.675 ;
        RECT 15.540 21.295 16.840 21.505 ;
        RECT 17.095 21.315 17.425 21.675 ;
        RECT 16.670 21.145 16.840 21.295 ;
        RECT 17.595 21.175 17.855 21.505 ;
        RECT 12.825 20.435 13.080 20.765 ;
        RECT 12.910 20.225 13.080 20.435 ;
        RECT 13.360 20.405 13.715 20.775 ;
        RECT 15.740 20.685 15.960 21.085 ;
        RECT 14.805 20.485 15.295 20.685 ;
        RECT 15.485 20.475 15.960 20.685 ;
        RECT 16.205 20.685 16.415 21.085 ;
        RECT 16.670 21.020 17.425 21.145 ;
        RECT 16.670 20.975 17.515 21.020 ;
        RECT 17.245 20.855 17.515 20.975 ;
        RECT 16.205 20.475 16.535 20.685 ;
        RECT 16.705 20.415 17.115 20.720 ;
        RECT 14.810 20.245 15.985 20.305 ;
        RECT 17.345 20.280 17.515 20.855 ;
        RECT 17.315 20.245 17.515 20.280 ;
        RECT 12.485 19.295 12.740 20.200 ;
        RECT 12.910 20.055 13.625 20.225 ;
        RECT 12.910 19.125 13.240 19.885 ;
        RECT 13.455 19.295 13.625 20.055 ;
        RECT 14.810 20.135 17.515 20.245 ;
        RECT 14.810 19.515 15.065 20.135 ;
        RECT 15.655 20.075 17.455 20.135 ;
        RECT 15.655 20.045 15.985 20.075 ;
        RECT 17.685 19.975 17.855 21.175 ;
        RECT 18.115 21.125 18.285 21.505 ;
        RECT 18.500 21.295 18.830 21.675 ;
        RECT 18.115 20.955 18.830 21.125 ;
        RECT 18.025 20.405 18.380 20.775 ;
        RECT 18.660 20.765 18.830 20.955 ;
        RECT 19.000 20.930 19.255 21.505 ;
        RECT 18.660 20.435 18.915 20.765 ;
        RECT 18.660 20.225 18.830 20.435 ;
        RECT 15.315 19.875 15.500 19.965 ;
        RECT 16.090 19.875 16.925 19.885 ;
        RECT 15.315 19.675 16.925 19.875 ;
        RECT 15.315 19.635 15.545 19.675 ;
        RECT 14.810 19.295 15.145 19.515 ;
        RECT 16.150 19.125 16.505 19.505 ;
        RECT 16.675 19.295 16.925 19.675 ;
        RECT 17.175 19.125 17.425 19.905 ;
        RECT 17.595 19.295 17.855 19.975 ;
        RECT 18.115 20.055 18.830 20.225 ;
        RECT 19.085 20.200 19.255 20.930 ;
        RECT 19.430 20.835 19.690 21.675 ;
        RECT 20.950 21.165 21.190 21.675 ;
        RECT 21.370 21.165 21.650 21.495 ;
        RECT 21.880 21.165 22.095 21.675 ;
        RECT 20.845 20.435 21.200 20.995 ;
        RECT 18.115 19.295 18.285 20.055 ;
        RECT 18.500 19.125 18.830 19.885 ;
        RECT 19.000 19.295 19.255 20.200 ;
        RECT 19.430 19.125 19.690 20.275 ;
        RECT 21.370 20.265 21.540 21.165 ;
        RECT 21.710 20.435 21.975 20.995 ;
        RECT 22.265 20.935 22.880 21.505 ;
        RECT 23.085 21.130 28.430 21.675 ;
        RECT 22.225 20.265 22.395 20.765 ;
        RECT 20.970 20.095 22.395 20.265 ;
        RECT 20.970 19.920 21.360 20.095 ;
        RECT 21.845 19.125 22.175 19.925 ;
        RECT 22.565 19.915 22.880 20.935 ;
        RECT 24.670 20.300 25.010 21.130 ;
        RECT 28.605 20.905 31.195 21.675 ;
        RECT 31.365 20.950 31.655 21.675 ;
        RECT 31.825 20.905 33.495 21.675 ;
        RECT 33.670 20.910 34.125 21.675 ;
        RECT 34.400 21.295 35.700 21.505 ;
        RECT 35.955 21.315 36.285 21.675 ;
        RECT 35.530 21.145 35.700 21.295 ;
        RECT 36.455 21.175 36.715 21.505 ;
        RECT 22.345 19.295 22.880 19.915 ;
        RECT 26.490 19.560 26.840 20.810 ;
        RECT 28.605 20.385 29.815 20.905 ;
        RECT 29.985 20.215 31.195 20.735 ;
        RECT 31.825 20.385 32.575 20.905 ;
        RECT 23.085 19.125 28.430 19.560 ;
        RECT 28.605 19.125 31.195 20.215 ;
        RECT 31.365 19.125 31.655 20.290 ;
        RECT 32.745 20.215 33.495 20.735 ;
        RECT 34.600 20.685 34.820 21.085 ;
        RECT 33.665 20.485 34.155 20.685 ;
        RECT 34.345 20.475 34.820 20.685 ;
        RECT 35.065 20.685 35.275 21.085 ;
        RECT 35.530 21.020 36.285 21.145 ;
        RECT 35.530 20.975 36.375 21.020 ;
        RECT 36.105 20.855 36.375 20.975 ;
        RECT 35.065 20.475 35.395 20.685 ;
        RECT 35.565 20.415 35.975 20.720 ;
        RECT 31.825 19.125 33.495 20.215 ;
        RECT 33.670 20.245 34.845 20.305 ;
        RECT 36.205 20.280 36.375 20.855 ;
        RECT 36.175 20.245 36.375 20.280 ;
        RECT 33.670 20.135 36.375 20.245 ;
        RECT 33.670 19.515 33.925 20.135 ;
        RECT 34.515 20.075 36.315 20.135 ;
        RECT 34.515 20.045 34.845 20.075 ;
        RECT 36.545 19.975 36.715 21.175 ;
        RECT 36.885 20.925 38.095 21.675 ;
        RECT 36.885 20.385 37.405 20.925 ;
        RECT 38.270 20.910 38.725 21.675 ;
        RECT 39.000 21.295 40.300 21.505 ;
        RECT 40.555 21.315 40.885 21.675 ;
        RECT 40.130 21.145 40.300 21.295 ;
        RECT 41.055 21.175 41.315 21.505 ;
        RECT 37.575 20.215 38.095 20.755 ;
        RECT 39.200 20.685 39.420 21.085 ;
        RECT 38.265 20.485 38.755 20.685 ;
        RECT 38.945 20.475 39.420 20.685 ;
        RECT 39.665 20.685 39.875 21.085 ;
        RECT 40.130 21.020 40.885 21.145 ;
        RECT 40.130 20.975 40.975 21.020 ;
        RECT 40.705 20.855 40.975 20.975 ;
        RECT 39.665 20.475 39.995 20.685 ;
        RECT 40.165 20.415 40.575 20.720 ;
        RECT 34.175 19.875 34.360 19.965 ;
        RECT 34.950 19.875 35.785 19.885 ;
        RECT 34.175 19.675 35.785 19.875 ;
        RECT 34.175 19.635 34.405 19.675 ;
        RECT 33.670 19.295 34.005 19.515 ;
        RECT 35.010 19.125 35.365 19.505 ;
        RECT 35.535 19.295 35.785 19.675 ;
        RECT 36.035 19.125 36.285 19.905 ;
        RECT 36.455 19.295 36.715 19.975 ;
        RECT 36.885 19.125 38.095 20.215 ;
        RECT 38.270 20.245 39.445 20.305 ;
        RECT 40.805 20.280 40.975 20.855 ;
        RECT 40.775 20.245 40.975 20.280 ;
        RECT 38.270 20.135 40.975 20.245 ;
        RECT 38.270 19.515 38.525 20.135 ;
        RECT 39.115 20.075 40.915 20.135 ;
        RECT 39.115 20.045 39.445 20.075 ;
        RECT 41.145 19.975 41.315 21.175 ;
        RECT 41.485 21.130 46.830 21.675 ;
        RECT 43.070 20.300 43.410 21.130 ;
        RECT 47.005 20.905 50.515 21.675 ;
        RECT 38.775 19.875 38.960 19.965 ;
        RECT 39.550 19.875 40.385 19.885 ;
        RECT 38.775 19.675 40.385 19.875 ;
        RECT 38.775 19.635 39.005 19.675 ;
        RECT 38.270 19.295 38.605 19.515 ;
        RECT 39.610 19.125 39.965 19.505 ;
        RECT 40.135 19.295 40.385 19.675 ;
        RECT 40.635 19.125 40.885 19.905 ;
        RECT 41.055 19.295 41.315 19.975 ;
        RECT 44.890 19.560 45.240 20.810 ;
        RECT 47.005 20.385 48.655 20.905 ;
        RECT 51.145 20.875 51.485 21.505 ;
        RECT 51.655 20.875 51.905 21.675 ;
        RECT 52.095 21.025 52.425 21.505 ;
        RECT 52.595 21.215 52.820 21.675 ;
        RECT 52.990 21.025 53.320 21.505 ;
        RECT 48.825 20.215 50.515 20.735 ;
        RECT 41.485 19.125 46.830 19.560 ;
        RECT 47.005 19.125 50.515 20.215 ;
        RECT 51.145 20.265 51.320 20.875 ;
        RECT 52.095 20.855 53.320 21.025 ;
        RECT 53.950 20.895 54.450 21.505 ;
        RECT 54.860 20.935 55.475 21.505 ;
        RECT 55.645 21.165 55.860 21.675 ;
        RECT 56.090 21.165 56.370 21.495 ;
        RECT 56.550 21.165 56.790 21.675 ;
        RECT 51.490 20.515 52.185 20.685 ;
        RECT 52.015 20.265 52.185 20.515 ;
        RECT 52.360 20.485 52.780 20.685 ;
        RECT 52.950 20.485 53.280 20.685 ;
        RECT 53.450 20.485 53.780 20.685 ;
        RECT 53.950 20.265 54.120 20.895 ;
        RECT 54.305 20.435 54.655 20.685 ;
        RECT 51.145 19.295 51.485 20.265 ;
        RECT 51.655 19.125 51.825 20.265 ;
        RECT 52.015 20.095 54.450 20.265 ;
        RECT 52.095 19.125 52.345 19.925 ;
        RECT 52.990 19.295 53.320 20.095 ;
        RECT 53.620 19.125 53.950 19.925 ;
        RECT 54.120 19.295 54.450 20.095 ;
        RECT 54.860 19.915 55.175 20.935 ;
        RECT 55.345 20.265 55.515 20.765 ;
        RECT 55.765 20.435 56.030 20.995 ;
        RECT 56.200 20.265 56.370 21.165 ;
        RECT 56.540 20.435 56.895 20.995 ;
        RECT 57.125 20.950 57.415 21.675 ;
        RECT 57.585 21.175 57.845 21.505 ;
        RECT 58.015 21.315 58.345 21.675 ;
        RECT 58.600 21.295 59.900 21.505 ;
        RECT 55.345 20.095 56.770 20.265 ;
        RECT 54.860 19.295 55.395 19.915 ;
        RECT 55.565 19.125 55.895 19.925 ;
        RECT 56.380 19.920 56.770 20.095 ;
        RECT 57.125 19.125 57.415 20.290 ;
        RECT 57.585 19.975 57.755 21.175 ;
        RECT 58.600 21.145 58.770 21.295 ;
        RECT 58.015 21.020 58.770 21.145 ;
        RECT 57.925 20.975 58.770 21.020 ;
        RECT 57.925 20.855 58.195 20.975 ;
        RECT 57.925 20.280 58.095 20.855 ;
        RECT 58.325 20.415 58.735 20.720 ;
        RECT 59.025 20.685 59.235 21.085 ;
        RECT 58.905 20.475 59.235 20.685 ;
        RECT 59.480 20.685 59.700 21.085 ;
        RECT 60.175 20.910 60.630 21.675 ;
        RECT 60.805 20.875 61.145 21.505 ;
        RECT 61.315 20.875 61.565 21.675 ;
        RECT 61.755 21.025 62.085 21.505 ;
        RECT 62.255 21.215 62.480 21.675 ;
        RECT 62.650 21.025 62.980 21.505 ;
        RECT 59.480 20.475 59.955 20.685 ;
        RECT 60.145 20.485 60.635 20.685 ;
        RECT 57.925 20.245 58.125 20.280 ;
        RECT 59.455 20.245 60.630 20.305 ;
        RECT 57.925 20.135 60.630 20.245 ;
        RECT 57.985 20.075 59.785 20.135 ;
        RECT 59.455 20.045 59.785 20.075 ;
        RECT 57.585 19.295 57.845 19.975 ;
        RECT 58.015 19.125 58.265 19.905 ;
        RECT 58.515 19.875 59.350 19.885 ;
        RECT 59.940 19.875 60.125 19.965 ;
        RECT 58.515 19.675 60.125 19.875 ;
        RECT 58.515 19.295 58.765 19.675 ;
        RECT 59.895 19.635 60.125 19.675 ;
        RECT 60.375 19.515 60.630 20.135 ;
        RECT 58.935 19.125 59.290 19.505 ;
        RECT 60.295 19.295 60.630 19.515 ;
        RECT 60.805 20.265 60.980 20.875 ;
        RECT 61.755 20.855 62.980 21.025 ;
        RECT 63.610 20.895 64.110 21.505 ;
        RECT 64.520 20.935 65.135 21.505 ;
        RECT 65.305 21.165 65.520 21.675 ;
        RECT 65.750 21.165 66.030 21.495 ;
        RECT 66.210 21.165 66.450 21.675 ;
        RECT 61.150 20.515 61.845 20.685 ;
        RECT 61.675 20.265 61.845 20.515 ;
        RECT 62.020 20.485 62.440 20.685 ;
        RECT 62.610 20.485 62.940 20.685 ;
        RECT 63.110 20.485 63.440 20.685 ;
        RECT 63.610 20.265 63.780 20.895 ;
        RECT 63.965 20.435 64.315 20.685 ;
        RECT 60.805 19.295 61.145 20.265 ;
        RECT 61.315 19.125 61.485 20.265 ;
        RECT 61.675 20.095 64.110 20.265 ;
        RECT 61.755 19.125 62.005 19.925 ;
        RECT 62.650 19.295 62.980 20.095 ;
        RECT 63.280 19.125 63.610 19.925 ;
        RECT 63.780 19.295 64.110 20.095 ;
        RECT 64.520 19.915 64.835 20.935 ;
        RECT 65.005 20.265 65.175 20.765 ;
        RECT 65.425 20.435 65.690 20.995 ;
        RECT 65.860 20.265 66.030 21.165 ;
        RECT 66.200 20.435 66.555 20.995 ;
        RECT 66.785 20.905 68.455 21.675 ;
        RECT 69.085 21.175 69.345 21.505 ;
        RECT 69.515 21.315 69.845 21.675 ;
        RECT 70.100 21.295 71.400 21.505 ;
        RECT 66.785 20.385 67.535 20.905 ;
        RECT 65.005 20.095 66.430 20.265 ;
        RECT 67.705 20.215 68.455 20.735 ;
        RECT 64.520 19.295 65.055 19.915 ;
        RECT 65.225 19.125 65.555 19.925 ;
        RECT 66.040 19.920 66.430 20.095 ;
        RECT 66.785 19.125 68.455 20.215 ;
        RECT 69.085 19.975 69.255 21.175 ;
        RECT 70.100 21.145 70.270 21.295 ;
        RECT 69.515 21.020 70.270 21.145 ;
        RECT 69.425 20.975 70.270 21.020 ;
        RECT 69.425 20.855 69.695 20.975 ;
        RECT 69.425 20.280 69.595 20.855 ;
        RECT 69.825 20.415 70.235 20.720 ;
        RECT 70.525 20.685 70.735 21.085 ;
        RECT 70.405 20.475 70.735 20.685 ;
        RECT 70.980 20.685 71.200 21.085 ;
        RECT 71.675 20.910 72.130 21.675 ;
        RECT 72.510 20.895 73.010 21.505 ;
        RECT 70.980 20.475 71.455 20.685 ;
        RECT 71.645 20.485 72.135 20.685 ;
        RECT 72.305 20.435 72.655 20.685 ;
        RECT 69.425 20.245 69.625 20.280 ;
        RECT 70.955 20.245 72.130 20.305 ;
        RECT 72.840 20.265 73.010 20.895 ;
        RECT 73.640 21.025 73.970 21.505 ;
        RECT 74.140 21.215 74.365 21.675 ;
        RECT 74.535 21.025 74.865 21.505 ;
        RECT 73.640 20.855 74.865 21.025 ;
        RECT 75.055 20.875 75.305 21.675 ;
        RECT 75.475 20.875 75.815 21.505 ;
        RECT 73.180 20.485 73.510 20.685 ;
        RECT 73.680 20.485 74.010 20.685 ;
        RECT 74.180 20.485 74.600 20.685 ;
        RECT 74.775 20.515 75.470 20.685 ;
        RECT 74.775 20.265 74.945 20.515 ;
        RECT 75.640 20.315 75.815 20.875 ;
        RECT 75.985 20.925 77.195 21.675 ;
        RECT 77.455 21.125 77.625 21.505 ;
        RECT 77.840 21.295 78.170 21.675 ;
        RECT 77.455 20.955 78.170 21.125 ;
        RECT 75.985 20.385 76.505 20.925 ;
        RECT 75.585 20.265 75.815 20.315 ;
        RECT 69.425 20.135 72.130 20.245 ;
        RECT 69.485 20.075 71.285 20.135 ;
        RECT 70.955 20.045 71.285 20.075 ;
        RECT 69.085 19.295 69.345 19.975 ;
        RECT 69.515 19.125 69.765 19.905 ;
        RECT 70.015 19.875 70.850 19.885 ;
        RECT 71.440 19.875 71.625 19.965 ;
        RECT 70.015 19.675 71.625 19.875 ;
        RECT 70.015 19.295 70.265 19.675 ;
        RECT 71.395 19.635 71.625 19.675 ;
        RECT 71.875 19.515 72.130 20.135 ;
        RECT 70.435 19.125 70.790 19.505 ;
        RECT 71.795 19.295 72.130 19.515 ;
        RECT 72.510 20.095 74.945 20.265 ;
        RECT 72.510 19.295 72.840 20.095 ;
        RECT 73.010 19.125 73.340 19.925 ;
        RECT 73.640 19.295 73.970 20.095 ;
        RECT 74.615 19.125 74.865 19.925 ;
        RECT 75.135 19.125 75.305 20.265 ;
        RECT 75.475 19.295 75.815 20.265 ;
        RECT 76.675 20.215 77.195 20.755 ;
        RECT 77.365 20.405 77.720 20.775 ;
        RECT 78.000 20.765 78.170 20.955 ;
        RECT 78.340 20.930 78.595 21.505 ;
        RECT 78.000 20.435 78.255 20.765 ;
        RECT 78.000 20.225 78.170 20.435 ;
        RECT 75.985 19.125 77.195 20.215 ;
        RECT 77.455 20.055 78.170 20.225 ;
        RECT 78.425 20.200 78.595 20.930 ;
        RECT 78.770 20.835 79.030 21.675 ;
        RECT 79.295 21.125 79.465 21.505 ;
        RECT 79.680 21.295 80.010 21.675 ;
        RECT 79.295 20.955 80.010 21.125 ;
        RECT 79.205 20.405 79.560 20.775 ;
        RECT 79.840 20.765 80.010 20.955 ;
        RECT 80.180 20.930 80.435 21.505 ;
        RECT 79.840 20.435 80.095 20.765 ;
        RECT 77.455 19.295 77.625 20.055 ;
        RECT 77.840 19.125 78.170 19.885 ;
        RECT 78.340 19.295 78.595 20.200 ;
        RECT 78.770 19.125 79.030 20.275 ;
        RECT 79.840 20.225 80.010 20.435 ;
        RECT 79.295 20.055 80.010 20.225 ;
        RECT 80.265 20.200 80.435 20.930 ;
        RECT 80.610 20.835 80.870 21.675 ;
        RECT 81.050 20.835 81.310 21.675 ;
        RECT 81.485 20.930 81.740 21.505 ;
        RECT 81.910 21.295 82.240 21.675 ;
        RECT 82.455 21.125 82.625 21.505 ;
        RECT 81.910 20.955 82.625 21.125 ;
        RECT 79.295 19.295 79.465 20.055 ;
        RECT 79.680 19.125 80.010 19.885 ;
        RECT 80.180 19.295 80.435 20.200 ;
        RECT 80.610 19.125 80.870 20.275 ;
        RECT 81.050 19.125 81.310 20.275 ;
        RECT 81.485 20.200 81.655 20.930 ;
        RECT 81.910 20.765 82.080 20.955 ;
        RECT 82.885 20.925 84.095 21.675 ;
        RECT 81.825 20.435 82.080 20.765 ;
        RECT 81.910 20.225 82.080 20.435 ;
        RECT 82.360 20.405 82.715 20.775 ;
        RECT 81.485 19.295 81.740 20.200 ;
        RECT 81.910 20.055 82.625 20.225 ;
        RECT 81.910 19.125 82.240 19.885 ;
        RECT 82.455 19.295 82.625 20.055 ;
        RECT 82.885 20.215 83.405 20.755 ;
        RECT 83.575 20.385 84.095 20.925 ;
        RECT 82.885 19.125 84.095 20.215 ;
        RECT 5.520 18.955 84.180 19.125 ;
        RECT 5.605 17.865 6.815 18.955 ;
        RECT 5.605 17.155 6.125 17.695 ;
        RECT 6.295 17.325 6.815 17.865 ;
        RECT 7.445 17.815 7.785 18.785 ;
        RECT 7.955 17.815 8.125 18.955 ;
        RECT 8.395 18.155 8.645 18.955 ;
        RECT 9.290 17.985 9.620 18.785 ;
        RECT 9.920 18.155 10.250 18.955 ;
        RECT 10.420 17.985 10.750 18.785 ;
        RECT 8.315 17.815 10.750 17.985 ;
        RECT 7.445 17.205 7.620 17.815 ;
        RECT 8.315 17.565 8.485 17.815 ;
        RECT 7.790 17.395 8.485 17.565 ;
        RECT 8.660 17.395 9.080 17.595 ;
        RECT 9.250 17.395 9.580 17.595 ;
        RECT 9.750 17.395 10.080 17.595 ;
        RECT 5.605 16.405 6.815 17.155 ;
        RECT 7.445 16.575 7.785 17.205 ;
        RECT 7.955 16.405 8.205 17.205 ;
        RECT 8.395 17.055 9.620 17.225 ;
        RECT 8.395 16.575 8.725 17.055 ;
        RECT 8.895 16.405 9.120 16.865 ;
        RECT 9.290 16.575 9.620 17.055 ;
        RECT 10.250 17.185 10.420 17.815 ;
        RECT 12.050 17.805 12.310 18.955 ;
        RECT 12.485 17.880 12.740 18.785 ;
        RECT 12.910 18.195 13.240 18.955 ;
        RECT 13.455 18.025 13.625 18.785 ;
        RECT 10.605 17.395 10.955 17.645 ;
        RECT 10.250 16.575 10.750 17.185 ;
        RECT 12.050 16.405 12.310 17.245 ;
        RECT 12.485 17.150 12.655 17.880 ;
        RECT 12.910 17.855 13.625 18.025 ;
        RECT 12.910 17.645 13.080 17.855 ;
        RECT 13.885 17.815 14.225 18.785 ;
        RECT 14.395 17.815 14.565 18.955 ;
        RECT 14.835 18.155 15.085 18.955 ;
        RECT 15.730 17.985 16.060 18.785 ;
        RECT 16.360 18.155 16.690 18.955 ;
        RECT 16.860 17.985 17.190 18.785 ;
        RECT 14.755 17.815 17.190 17.985 ;
        RECT 12.825 17.315 13.080 17.645 ;
        RECT 12.485 16.575 12.740 17.150 ;
        RECT 12.910 17.125 13.080 17.315 ;
        RECT 13.360 17.305 13.715 17.675 ;
        RECT 13.885 17.205 14.060 17.815 ;
        RECT 14.755 17.565 14.925 17.815 ;
        RECT 14.230 17.395 14.925 17.565 ;
        RECT 15.100 17.395 15.520 17.595 ;
        RECT 15.690 17.395 16.020 17.595 ;
        RECT 16.190 17.395 16.520 17.595 ;
        RECT 12.910 16.955 13.625 17.125 ;
        RECT 12.910 16.405 13.240 16.785 ;
        RECT 13.455 16.575 13.625 16.955 ;
        RECT 13.885 16.575 14.225 17.205 ;
        RECT 14.395 16.405 14.645 17.205 ;
        RECT 14.835 17.055 16.060 17.225 ;
        RECT 14.835 16.575 15.165 17.055 ;
        RECT 15.335 16.405 15.560 16.865 ;
        RECT 15.730 16.575 16.060 17.055 ;
        RECT 16.690 17.185 16.860 17.815 ;
        RECT 18.485 17.790 18.775 18.955 ;
        RECT 19.610 17.985 19.940 18.785 ;
        RECT 20.110 18.155 20.440 18.955 ;
        RECT 20.740 17.985 21.070 18.785 ;
        RECT 21.715 18.155 21.965 18.955 ;
        RECT 19.610 17.815 22.045 17.985 ;
        RECT 22.235 17.815 22.405 18.955 ;
        RECT 22.575 17.815 22.915 18.785 ;
        RECT 23.290 17.985 23.620 18.785 ;
        RECT 23.790 18.155 24.120 18.955 ;
        RECT 24.420 17.985 24.750 18.785 ;
        RECT 25.395 18.155 25.645 18.955 ;
        RECT 23.290 17.815 25.725 17.985 ;
        RECT 25.915 17.815 26.085 18.955 ;
        RECT 26.255 17.815 26.595 18.785 ;
        RECT 26.855 18.285 27.025 18.785 ;
        RECT 27.195 18.455 27.525 18.955 ;
        RECT 26.855 18.115 27.520 18.285 ;
        RECT 17.045 17.395 17.395 17.645 ;
        RECT 19.405 17.395 19.755 17.645 ;
        RECT 19.940 17.185 20.110 17.815 ;
        RECT 20.280 17.395 20.610 17.595 ;
        RECT 20.780 17.395 21.110 17.595 ;
        RECT 21.280 17.395 21.700 17.595 ;
        RECT 21.875 17.565 22.045 17.815 ;
        RECT 21.875 17.395 22.570 17.565 ;
        RECT 16.690 16.575 17.190 17.185 ;
        RECT 18.485 16.405 18.775 17.130 ;
        RECT 19.610 16.575 20.110 17.185 ;
        RECT 20.740 17.055 21.965 17.225 ;
        RECT 22.740 17.205 22.915 17.815 ;
        RECT 23.085 17.395 23.435 17.645 ;
        RECT 20.740 16.575 21.070 17.055 ;
        RECT 21.240 16.405 21.465 16.865 ;
        RECT 21.635 16.575 21.965 17.055 ;
        RECT 22.155 16.405 22.405 17.205 ;
        RECT 22.575 16.575 22.915 17.205 ;
        RECT 23.620 17.185 23.790 17.815 ;
        RECT 23.960 17.395 24.290 17.595 ;
        RECT 24.460 17.395 24.790 17.595 ;
        RECT 24.960 17.395 25.380 17.595 ;
        RECT 25.555 17.565 25.725 17.815 ;
        RECT 25.555 17.395 26.250 17.565 ;
        RECT 26.420 17.255 26.595 17.815 ;
        RECT 26.770 17.295 27.120 17.945 ;
        RECT 23.290 16.575 23.790 17.185 ;
        RECT 24.420 17.055 25.645 17.225 ;
        RECT 26.365 17.205 26.595 17.255 ;
        RECT 24.420 16.575 24.750 17.055 ;
        RECT 24.920 16.405 25.145 16.865 ;
        RECT 25.315 16.575 25.645 17.055 ;
        RECT 25.835 16.405 26.085 17.205 ;
        RECT 26.255 16.575 26.595 17.205 ;
        RECT 27.290 17.125 27.520 18.115 ;
        RECT 26.855 16.955 27.520 17.125 ;
        RECT 26.855 16.665 27.025 16.955 ;
        RECT 27.195 16.405 27.525 16.785 ;
        RECT 27.695 16.665 27.880 18.785 ;
        RECT 28.120 18.495 28.385 18.955 ;
        RECT 28.555 18.360 28.805 18.785 ;
        RECT 29.015 18.510 30.120 18.680 ;
        RECT 28.500 18.230 28.805 18.360 ;
        RECT 28.050 17.035 28.330 17.985 ;
        RECT 28.500 17.125 28.670 18.230 ;
        RECT 28.840 17.445 29.080 18.040 ;
        RECT 29.250 17.975 29.780 18.340 ;
        RECT 29.250 17.275 29.420 17.975 ;
        RECT 29.950 17.895 30.120 18.510 ;
        RECT 30.290 18.155 30.460 18.955 ;
        RECT 30.630 18.455 30.880 18.785 ;
        RECT 31.105 18.485 31.990 18.655 ;
        RECT 29.950 17.805 30.460 17.895 ;
        RECT 28.500 16.995 28.725 17.125 ;
        RECT 28.895 17.055 29.420 17.275 ;
        RECT 29.590 17.635 30.460 17.805 ;
        RECT 28.135 16.405 28.385 16.865 ;
        RECT 28.555 16.855 28.725 16.995 ;
        RECT 29.590 16.855 29.760 17.635 ;
        RECT 30.290 17.565 30.460 17.635 ;
        RECT 29.970 17.385 30.170 17.415 ;
        RECT 30.630 17.385 30.800 18.455 ;
        RECT 30.970 17.565 31.160 18.285 ;
        RECT 29.970 17.085 30.800 17.385 ;
        RECT 31.330 17.355 31.650 18.315 ;
        RECT 28.555 16.685 28.890 16.855 ;
        RECT 29.085 16.685 29.760 16.855 ;
        RECT 30.080 16.405 30.450 16.905 ;
        RECT 30.630 16.855 30.800 17.085 ;
        RECT 31.185 17.025 31.650 17.355 ;
        RECT 31.820 17.645 31.990 18.485 ;
        RECT 32.170 18.455 32.485 18.955 ;
        RECT 32.715 18.225 33.055 18.785 ;
        RECT 32.160 17.850 33.055 18.225 ;
        RECT 33.225 17.945 33.395 18.955 ;
        RECT 32.865 17.645 33.055 17.850 ;
        RECT 33.565 17.895 33.895 18.740 ;
        RECT 33.565 17.815 33.955 17.895 ;
        RECT 33.740 17.765 33.955 17.815 ;
        RECT 31.820 17.315 32.695 17.645 ;
        RECT 32.865 17.315 33.615 17.645 ;
        RECT 31.820 16.855 31.990 17.315 ;
        RECT 32.865 17.145 33.065 17.315 ;
        RECT 33.785 17.185 33.955 17.765 ;
        RECT 33.730 17.145 33.955 17.185 ;
        RECT 30.630 16.685 31.035 16.855 ;
        RECT 31.205 16.685 31.990 16.855 ;
        RECT 32.265 16.405 32.475 16.935 ;
        RECT 32.735 16.620 33.065 17.145 ;
        RECT 33.575 17.060 33.955 17.145 ;
        RECT 35.045 17.815 35.385 18.785 ;
        RECT 35.555 17.815 35.725 18.955 ;
        RECT 35.995 18.155 36.245 18.955 ;
        RECT 36.890 17.985 37.220 18.785 ;
        RECT 37.520 18.155 37.850 18.955 ;
        RECT 38.020 17.985 38.350 18.785 ;
        RECT 35.915 17.815 38.350 17.985 ;
        RECT 38.725 17.865 40.395 18.955 ;
        RECT 35.045 17.205 35.220 17.815 ;
        RECT 35.915 17.565 36.085 17.815 ;
        RECT 35.390 17.395 36.085 17.565 ;
        RECT 36.260 17.395 36.680 17.595 ;
        RECT 36.850 17.395 37.180 17.595 ;
        RECT 37.350 17.395 37.680 17.595 ;
        RECT 33.235 16.405 33.405 17.015 ;
        RECT 33.575 16.625 33.905 17.060 ;
        RECT 35.045 16.575 35.385 17.205 ;
        RECT 35.555 16.405 35.805 17.205 ;
        RECT 35.995 17.055 37.220 17.225 ;
        RECT 35.995 16.575 36.325 17.055 ;
        RECT 36.495 16.405 36.720 16.865 ;
        RECT 36.890 16.575 37.220 17.055 ;
        RECT 37.850 17.185 38.020 17.815 ;
        RECT 38.205 17.395 38.555 17.645 ;
        RECT 37.850 16.575 38.350 17.185 ;
        RECT 38.725 17.175 39.475 17.695 ;
        RECT 39.645 17.345 40.395 17.865 ;
        RECT 40.565 17.815 40.905 18.785 ;
        RECT 41.075 17.815 41.245 18.955 ;
        RECT 41.515 18.155 41.765 18.955 ;
        RECT 42.410 17.985 42.740 18.785 ;
        RECT 43.040 18.155 43.370 18.955 ;
        RECT 43.540 17.985 43.870 18.785 ;
        RECT 41.435 17.815 43.870 17.985 ;
        RECT 40.565 17.205 40.740 17.815 ;
        RECT 41.435 17.565 41.605 17.815 ;
        RECT 40.910 17.395 41.605 17.565 ;
        RECT 41.780 17.395 42.200 17.595 ;
        RECT 42.370 17.395 42.700 17.595 ;
        RECT 42.870 17.395 43.200 17.595 ;
        RECT 38.725 16.405 40.395 17.175 ;
        RECT 40.565 16.575 40.905 17.205 ;
        RECT 41.075 16.405 41.325 17.205 ;
        RECT 41.515 17.055 42.740 17.225 ;
        RECT 41.515 16.575 41.845 17.055 ;
        RECT 42.015 16.405 42.240 16.865 ;
        RECT 42.410 16.575 42.740 17.055 ;
        RECT 43.370 17.185 43.540 17.815 ;
        RECT 44.245 17.790 44.535 18.955 ;
        RECT 44.705 17.865 46.375 18.955 ;
        RECT 43.725 17.395 44.075 17.645 ;
        RECT 43.370 16.575 43.870 17.185 ;
        RECT 44.705 17.175 45.455 17.695 ;
        RECT 45.625 17.345 46.375 17.865 ;
        RECT 47.005 17.815 47.345 18.785 ;
        RECT 47.515 17.815 47.685 18.955 ;
        RECT 47.955 18.155 48.205 18.955 ;
        RECT 48.850 17.985 49.180 18.785 ;
        RECT 49.480 18.155 49.810 18.955 ;
        RECT 49.980 17.985 50.310 18.785 ;
        RECT 50.775 18.285 50.945 18.785 ;
        RECT 51.115 18.455 51.445 18.955 ;
        RECT 50.775 18.115 51.440 18.285 ;
        RECT 47.875 17.815 50.310 17.985 ;
        RECT 47.005 17.205 47.180 17.815 ;
        RECT 47.875 17.565 48.045 17.815 ;
        RECT 47.350 17.395 48.045 17.565 ;
        RECT 48.220 17.395 48.640 17.595 ;
        RECT 48.810 17.395 49.140 17.595 ;
        RECT 49.310 17.395 49.640 17.595 ;
        RECT 44.245 16.405 44.535 17.130 ;
        RECT 44.705 16.405 46.375 17.175 ;
        RECT 47.005 16.575 47.345 17.205 ;
        RECT 47.515 16.405 47.765 17.205 ;
        RECT 47.955 17.055 49.180 17.225 ;
        RECT 47.955 16.575 48.285 17.055 ;
        RECT 48.455 16.405 48.680 16.865 ;
        RECT 48.850 16.575 49.180 17.055 ;
        RECT 49.810 17.185 49.980 17.815 ;
        RECT 50.165 17.395 50.515 17.645 ;
        RECT 50.690 17.295 51.040 17.945 ;
        RECT 49.810 16.575 50.310 17.185 ;
        RECT 51.210 17.125 51.440 18.115 ;
        RECT 50.775 16.955 51.440 17.125 ;
        RECT 50.775 16.665 50.945 16.955 ;
        RECT 51.115 16.405 51.445 16.785 ;
        RECT 51.615 16.665 51.800 18.785 ;
        RECT 52.040 18.495 52.305 18.955 ;
        RECT 52.475 18.360 52.725 18.785 ;
        RECT 52.935 18.510 54.040 18.680 ;
        RECT 52.420 18.230 52.725 18.360 ;
        RECT 51.970 17.035 52.250 17.985 ;
        RECT 52.420 17.125 52.590 18.230 ;
        RECT 52.760 17.445 53.000 18.040 ;
        RECT 53.170 17.975 53.700 18.340 ;
        RECT 53.170 17.275 53.340 17.975 ;
        RECT 53.870 17.895 54.040 18.510 ;
        RECT 54.210 18.155 54.380 18.955 ;
        RECT 54.550 18.455 54.800 18.785 ;
        RECT 55.025 18.485 55.910 18.655 ;
        RECT 53.870 17.805 54.380 17.895 ;
        RECT 52.420 16.995 52.645 17.125 ;
        RECT 52.815 17.055 53.340 17.275 ;
        RECT 53.510 17.635 54.380 17.805 ;
        RECT 52.055 16.405 52.305 16.865 ;
        RECT 52.475 16.855 52.645 16.995 ;
        RECT 53.510 16.855 53.680 17.635 ;
        RECT 54.210 17.565 54.380 17.635 ;
        RECT 53.890 17.385 54.090 17.415 ;
        RECT 54.550 17.385 54.720 18.455 ;
        RECT 54.890 17.565 55.080 18.285 ;
        RECT 53.890 17.085 54.720 17.385 ;
        RECT 55.250 17.355 55.570 18.315 ;
        RECT 52.475 16.685 52.810 16.855 ;
        RECT 53.005 16.685 53.680 16.855 ;
        RECT 54.000 16.405 54.370 16.905 ;
        RECT 54.550 16.855 54.720 17.085 ;
        RECT 55.105 17.025 55.570 17.355 ;
        RECT 55.740 17.645 55.910 18.485 ;
        RECT 56.090 18.455 56.405 18.955 ;
        RECT 56.635 18.225 56.975 18.785 ;
        RECT 56.080 17.850 56.975 18.225 ;
        RECT 57.145 17.945 57.315 18.955 ;
        RECT 56.785 17.645 56.975 17.850 ;
        RECT 57.485 17.895 57.815 18.740 ;
        RECT 58.135 18.285 58.305 18.785 ;
        RECT 58.475 18.455 58.805 18.955 ;
        RECT 58.135 18.115 58.800 18.285 ;
        RECT 57.485 17.815 57.875 17.895 ;
        RECT 57.660 17.765 57.875 17.815 ;
        RECT 55.740 17.315 56.615 17.645 ;
        RECT 56.785 17.315 57.535 17.645 ;
        RECT 55.740 16.855 55.910 17.315 ;
        RECT 56.785 17.145 56.985 17.315 ;
        RECT 57.705 17.185 57.875 17.765 ;
        RECT 58.050 17.295 58.400 17.945 ;
        RECT 57.650 17.145 57.875 17.185 ;
        RECT 54.550 16.685 54.955 16.855 ;
        RECT 55.125 16.685 55.910 16.855 ;
        RECT 56.185 16.405 56.395 16.935 ;
        RECT 56.655 16.620 56.985 17.145 ;
        RECT 57.495 17.060 57.875 17.145 ;
        RECT 58.570 17.125 58.800 18.115 ;
        RECT 57.155 16.405 57.325 17.015 ;
        RECT 57.495 16.625 57.825 17.060 ;
        RECT 58.135 16.955 58.800 17.125 ;
        RECT 58.135 16.665 58.305 16.955 ;
        RECT 58.475 16.405 58.805 16.785 ;
        RECT 58.975 16.665 59.160 18.785 ;
        RECT 59.400 18.495 59.665 18.955 ;
        RECT 59.835 18.360 60.085 18.785 ;
        RECT 60.295 18.510 61.400 18.680 ;
        RECT 59.780 18.230 60.085 18.360 ;
        RECT 59.330 17.035 59.610 17.985 ;
        RECT 59.780 17.125 59.950 18.230 ;
        RECT 60.120 17.445 60.360 18.040 ;
        RECT 60.530 17.975 61.060 18.340 ;
        RECT 60.530 17.275 60.700 17.975 ;
        RECT 61.230 17.895 61.400 18.510 ;
        RECT 61.570 18.155 61.740 18.955 ;
        RECT 61.910 18.455 62.160 18.785 ;
        RECT 62.385 18.485 63.270 18.655 ;
        RECT 61.230 17.805 61.740 17.895 ;
        RECT 59.780 16.995 60.005 17.125 ;
        RECT 60.175 17.055 60.700 17.275 ;
        RECT 60.870 17.635 61.740 17.805 ;
        RECT 59.415 16.405 59.665 16.865 ;
        RECT 59.835 16.855 60.005 16.995 ;
        RECT 60.870 16.855 61.040 17.635 ;
        RECT 61.570 17.565 61.740 17.635 ;
        RECT 61.250 17.385 61.450 17.415 ;
        RECT 61.910 17.385 62.080 18.455 ;
        RECT 62.250 17.565 62.440 18.285 ;
        RECT 61.250 17.085 62.080 17.385 ;
        RECT 62.610 17.355 62.930 18.315 ;
        RECT 59.835 16.685 60.170 16.855 ;
        RECT 60.365 16.685 61.040 16.855 ;
        RECT 61.360 16.405 61.730 16.905 ;
        RECT 61.910 16.855 62.080 17.085 ;
        RECT 62.465 17.025 62.930 17.355 ;
        RECT 63.100 17.645 63.270 18.485 ;
        RECT 63.450 18.455 63.765 18.955 ;
        RECT 63.995 18.225 64.335 18.785 ;
        RECT 63.440 17.850 64.335 18.225 ;
        RECT 64.505 17.945 64.675 18.955 ;
        RECT 64.145 17.645 64.335 17.850 ;
        RECT 64.845 17.895 65.175 18.740 ;
        RECT 64.845 17.815 65.235 17.895 ;
        RECT 65.020 17.765 65.235 17.815 ;
        RECT 63.100 17.315 63.975 17.645 ;
        RECT 64.145 17.315 64.895 17.645 ;
        RECT 63.100 16.855 63.270 17.315 ;
        RECT 64.145 17.145 64.345 17.315 ;
        RECT 65.065 17.185 65.235 17.765 ;
        RECT 65.010 17.145 65.235 17.185 ;
        RECT 61.910 16.685 62.315 16.855 ;
        RECT 62.485 16.685 63.270 16.855 ;
        RECT 63.545 16.405 63.755 16.935 ;
        RECT 64.015 16.620 64.345 17.145 ;
        RECT 64.855 17.060 65.235 17.145 ;
        RECT 65.405 17.815 65.745 18.785 ;
        RECT 65.915 17.815 66.085 18.955 ;
        RECT 66.355 18.155 66.605 18.955 ;
        RECT 67.250 17.985 67.580 18.785 ;
        RECT 67.880 18.155 68.210 18.955 ;
        RECT 68.380 17.985 68.710 18.785 ;
        RECT 66.275 17.815 68.710 17.985 ;
        RECT 65.405 17.205 65.580 17.815 ;
        RECT 66.275 17.565 66.445 17.815 ;
        RECT 65.750 17.395 66.445 17.565 ;
        RECT 66.620 17.395 67.040 17.595 ;
        RECT 67.210 17.395 67.540 17.595 ;
        RECT 67.710 17.395 68.040 17.595 ;
        RECT 64.515 16.405 64.685 17.015 ;
        RECT 64.855 16.625 65.185 17.060 ;
        RECT 65.405 16.575 65.745 17.205 ;
        RECT 65.915 16.405 66.165 17.205 ;
        RECT 66.355 17.055 67.580 17.225 ;
        RECT 66.355 16.575 66.685 17.055 ;
        RECT 66.855 16.405 67.080 16.865 ;
        RECT 67.250 16.575 67.580 17.055 ;
        RECT 68.210 17.185 68.380 17.815 ;
        RECT 70.005 17.790 70.295 18.955 ;
        RECT 71.130 17.985 71.460 18.785 ;
        RECT 71.630 18.155 71.960 18.955 ;
        RECT 72.260 17.985 72.590 18.785 ;
        RECT 73.235 18.155 73.485 18.955 ;
        RECT 71.130 17.815 73.565 17.985 ;
        RECT 73.755 17.815 73.925 18.955 ;
        RECT 74.095 17.815 74.435 18.785 ;
        RECT 74.810 17.985 75.140 18.785 ;
        RECT 75.310 18.155 75.640 18.955 ;
        RECT 75.940 17.985 76.270 18.785 ;
        RECT 76.915 18.155 77.165 18.955 ;
        RECT 74.810 17.815 77.245 17.985 ;
        RECT 77.435 17.815 77.605 18.955 ;
        RECT 77.775 17.815 78.115 18.785 ;
        RECT 78.375 18.025 78.545 18.785 ;
        RECT 78.760 18.195 79.090 18.955 ;
        RECT 78.375 17.855 79.090 18.025 ;
        RECT 79.260 17.880 79.515 18.785 ;
        RECT 68.565 17.395 68.915 17.645 ;
        RECT 70.925 17.395 71.275 17.645 ;
        RECT 71.460 17.185 71.630 17.815 ;
        RECT 71.800 17.395 72.130 17.595 ;
        RECT 72.300 17.395 72.630 17.595 ;
        RECT 72.800 17.395 73.220 17.595 ;
        RECT 73.395 17.565 73.565 17.815 ;
        RECT 73.395 17.395 74.090 17.565 ;
        RECT 68.210 16.575 68.710 17.185 ;
        RECT 70.005 16.405 70.295 17.130 ;
        RECT 71.130 16.575 71.630 17.185 ;
        RECT 72.260 17.055 73.485 17.225 ;
        RECT 74.260 17.205 74.435 17.815 ;
        RECT 74.605 17.395 74.955 17.645 ;
        RECT 72.260 16.575 72.590 17.055 ;
        RECT 72.760 16.405 72.985 16.865 ;
        RECT 73.155 16.575 73.485 17.055 ;
        RECT 73.675 16.405 73.925 17.205 ;
        RECT 74.095 16.575 74.435 17.205 ;
        RECT 75.140 17.185 75.310 17.815 ;
        RECT 75.480 17.395 75.810 17.595 ;
        RECT 75.980 17.395 76.310 17.595 ;
        RECT 76.480 17.395 76.900 17.595 ;
        RECT 77.075 17.565 77.245 17.815 ;
        RECT 77.075 17.395 77.770 17.565 ;
        RECT 74.810 16.575 75.310 17.185 ;
        RECT 75.940 17.055 77.165 17.225 ;
        RECT 77.940 17.205 78.115 17.815 ;
        RECT 78.285 17.305 78.640 17.675 ;
        RECT 78.920 17.645 79.090 17.855 ;
        RECT 78.920 17.315 79.175 17.645 ;
        RECT 75.940 16.575 76.270 17.055 ;
        RECT 76.440 16.405 76.665 16.865 ;
        RECT 76.835 16.575 77.165 17.055 ;
        RECT 77.355 16.405 77.605 17.205 ;
        RECT 77.775 16.575 78.115 17.205 ;
        RECT 78.920 17.125 79.090 17.315 ;
        RECT 79.345 17.150 79.515 17.880 ;
        RECT 79.690 17.805 79.950 18.955 ;
        RECT 80.215 18.025 80.385 18.785 ;
        RECT 80.600 18.195 80.930 18.955 ;
        RECT 80.215 17.855 80.930 18.025 ;
        RECT 81.100 17.880 81.355 18.785 ;
        RECT 80.125 17.305 80.480 17.675 ;
        RECT 80.760 17.645 80.930 17.855 ;
        RECT 80.760 17.315 81.015 17.645 ;
        RECT 78.375 16.955 79.090 17.125 ;
        RECT 78.375 16.575 78.545 16.955 ;
        RECT 78.760 16.405 79.090 16.785 ;
        RECT 79.260 16.575 79.515 17.150 ;
        RECT 79.690 16.405 79.950 17.245 ;
        RECT 80.760 17.125 80.930 17.315 ;
        RECT 81.185 17.150 81.355 17.880 ;
        RECT 81.530 17.805 81.790 18.955 ;
        RECT 82.885 17.865 84.095 18.955 ;
        RECT 82.885 17.325 83.405 17.865 ;
        RECT 80.215 16.955 80.930 17.125 ;
        RECT 80.215 16.575 80.385 16.955 ;
        RECT 80.600 16.405 80.930 16.785 ;
        RECT 81.100 16.575 81.355 17.150 ;
        RECT 81.530 16.405 81.790 17.245 ;
        RECT 83.575 17.155 84.095 17.695 ;
        RECT 82.885 16.405 84.095 17.155 ;
        RECT 5.520 16.235 84.180 16.405 ;
        RECT 5.605 15.485 6.815 16.235 ;
        RECT 8.070 15.725 8.310 16.235 ;
        RECT 8.490 15.725 8.770 16.055 ;
        RECT 9.000 15.725 9.215 16.235 ;
        RECT 5.605 14.945 6.125 15.485 ;
        RECT 6.295 14.775 6.815 15.315 ;
        RECT 7.965 14.995 8.320 15.555 ;
        RECT 8.490 14.825 8.660 15.725 ;
        RECT 8.830 14.995 9.095 15.555 ;
        RECT 9.385 15.495 10.000 16.065 ;
        RECT 9.345 14.825 9.515 15.325 ;
        RECT 5.605 13.685 6.815 14.775 ;
        RECT 8.090 14.655 9.515 14.825 ;
        RECT 8.090 14.480 8.480 14.655 ;
        RECT 8.965 13.685 9.295 14.485 ;
        RECT 9.685 14.475 10.000 15.495 ;
        RECT 10.205 15.485 11.415 16.235 ;
        RECT 11.675 15.685 11.845 15.975 ;
        RECT 12.015 15.855 12.345 16.235 ;
        RECT 11.675 15.515 12.340 15.685 ;
        RECT 10.205 14.945 10.725 15.485 ;
        RECT 10.895 14.775 11.415 15.315 ;
        RECT 9.465 13.855 10.000 14.475 ;
        RECT 10.205 13.685 11.415 14.775 ;
        RECT 11.590 14.695 11.940 15.345 ;
        RECT 12.110 14.525 12.340 15.515 ;
        RECT 11.675 14.355 12.340 14.525 ;
        RECT 11.675 13.855 11.845 14.355 ;
        RECT 12.015 13.685 12.345 14.185 ;
        RECT 12.515 13.855 12.700 15.975 ;
        RECT 12.955 15.775 13.205 16.235 ;
        RECT 13.375 15.785 13.710 15.955 ;
        RECT 13.905 15.785 14.580 15.955 ;
        RECT 13.375 15.645 13.545 15.785 ;
        RECT 12.870 14.655 13.150 15.605 ;
        RECT 13.320 15.515 13.545 15.645 ;
        RECT 13.320 14.410 13.490 15.515 ;
        RECT 13.715 15.365 14.240 15.585 ;
        RECT 13.660 14.600 13.900 15.195 ;
        RECT 14.070 14.665 14.240 15.365 ;
        RECT 14.410 15.005 14.580 15.785 ;
        RECT 14.900 15.735 15.270 16.235 ;
        RECT 15.450 15.785 15.855 15.955 ;
        RECT 16.025 15.785 16.810 15.955 ;
        RECT 15.450 15.555 15.620 15.785 ;
        RECT 14.790 15.255 15.620 15.555 ;
        RECT 16.005 15.285 16.470 15.615 ;
        RECT 14.790 15.225 14.990 15.255 ;
        RECT 15.110 15.005 15.280 15.075 ;
        RECT 14.410 14.835 15.280 15.005 ;
        RECT 14.770 14.745 15.280 14.835 ;
        RECT 13.320 14.280 13.625 14.410 ;
        RECT 14.070 14.300 14.600 14.665 ;
        RECT 12.940 13.685 13.205 14.145 ;
        RECT 13.375 13.855 13.625 14.280 ;
        RECT 14.770 14.130 14.940 14.745 ;
        RECT 13.835 13.960 14.940 14.130 ;
        RECT 15.110 13.685 15.280 14.485 ;
        RECT 15.450 14.185 15.620 15.255 ;
        RECT 15.790 14.355 15.980 15.075 ;
        RECT 16.150 14.325 16.470 15.285 ;
        RECT 16.640 15.325 16.810 15.785 ;
        RECT 17.085 15.705 17.295 16.235 ;
        RECT 17.555 15.495 17.885 16.020 ;
        RECT 18.055 15.625 18.225 16.235 ;
        RECT 18.395 15.580 18.725 16.015 ;
        RECT 19.110 15.725 19.350 16.235 ;
        RECT 19.530 15.725 19.810 16.055 ;
        RECT 20.040 15.725 20.255 16.235 ;
        RECT 18.395 15.495 18.775 15.580 ;
        RECT 17.685 15.325 17.885 15.495 ;
        RECT 18.550 15.455 18.775 15.495 ;
        RECT 16.640 14.995 17.515 15.325 ;
        RECT 17.685 14.995 18.435 15.325 ;
        RECT 15.450 13.855 15.700 14.185 ;
        RECT 16.640 14.155 16.810 14.995 ;
        RECT 17.685 14.790 17.875 14.995 ;
        RECT 18.605 14.875 18.775 15.455 ;
        RECT 19.005 14.995 19.360 15.555 ;
        RECT 18.560 14.825 18.775 14.875 ;
        RECT 19.530 14.825 19.700 15.725 ;
        RECT 19.870 14.995 20.135 15.555 ;
        RECT 20.425 15.495 21.040 16.065 ;
        RECT 21.335 15.685 21.505 15.975 ;
        RECT 21.675 15.855 22.005 16.235 ;
        RECT 21.335 15.515 22.000 15.685 ;
        RECT 20.385 14.825 20.555 15.325 ;
        RECT 16.980 14.415 17.875 14.790 ;
        RECT 18.385 14.745 18.775 14.825 ;
        RECT 15.925 13.985 16.810 14.155 ;
        RECT 16.990 13.685 17.305 14.185 ;
        RECT 17.535 13.855 17.875 14.415 ;
        RECT 18.045 13.685 18.215 14.695 ;
        RECT 18.385 13.900 18.715 14.745 ;
        RECT 19.130 14.655 20.555 14.825 ;
        RECT 19.130 14.480 19.520 14.655 ;
        RECT 20.005 13.685 20.335 14.485 ;
        RECT 20.725 14.475 21.040 15.495 ;
        RECT 21.250 14.695 21.600 15.345 ;
        RECT 21.770 14.525 22.000 15.515 ;
        RECT 20.505 13.855 21.040 14.475 ;
        RECT 21.335 14.355 22.000 14.525 ;
        RECT 21.335 13.855 21.505 14.355 ;
        RECT 21.675 13.685 22.005 14.185 ;
        RECT 22.175 13.855 22.360 15.975 ;
        RECT 22.615 15.775 22.865 16.235 ;
        RECT 23.035 15.785 23.370 15.955 ;
        RECT 23.565 15.785 24.240 15.955 ;
        RECT 23.035 15.645 23.205 15.785 ;
        RECT 22.530 14.655 22.810 15.605 ;
        RECT 22.980 15.515 23.205 15.645 ;
        RECT 22.980 14.410 23.150 15.515 ;
        RECT 23.375 15.365 23.900 15.585 ;
        RECT 23.320 14.600 23.560 15.195 ;
        RECT 23.730 14.665 23.900 15.365 ;
        RECT 24.070 15.005 24.240 15.785 ;
        RECT 24.560 15.735 24.930 16.235 ;
        RECT 25.110 15.785 25.515 15.955 ;
        RECT 25.685 15.785 26.470 15.955 ;
        RECT 25.110 15.555 25.280 15.785 ;
        RECT 24.450 15.255 25.280 15.555 ;
        RECT 25.665 15.285 26.130 15.615 ;
        RECT 24.450 15.225 24.650 15.255 ;
        RECT 24.770 15.005 24.940 15.075 ;
        RECT 24.070 14.835 24.940 15.005 ;
        RECT 24.430 14.745 24.940 14.835 ;
        RECT 22.980 14.280 23.285 14.410 ;
        RECT 23.730 14.300 24.260 14.665 ;
        RECT 22.600 13.685 22.865 14.145 ;
        RECT 23.035 13.855 23.285 14.280 ;
        RECT 24.430 14.130 24.600 14.745 ;
        RECT 23.495 13.960 24.600 14.130 ;
        RECT 24.770 13.685 24.940 14.485 ;
        RECT 25.110 14.185 25.280 15.255 ;
        RECT 25.450 14.355 25.640 15.075 ;
        RECT 25.810 14.325 26.130 15.285 ;
        RECT 26.300 15.325 26.470 15.785 ;
        RECT 26.745 15.705 26.955 16.235 ;
        RECT 27.215 15.495 27.545 16.020 ;
        RECT 27.715 15.625 27.885 16.235 ;
        RECT 28.055 15.580 28.385 16.015 ;
        RECT 28.055 15.495 28.435 15.580 ;
        RECT 27.345 15.325 27.545 15.495 ;
        RECT 28.210 15.455 28.435 15.495 ;
        RECT 26.300 14.995 27.175 15.325 ;
        RECT 27.345 14.995 28.095 15.325 ;
        RECT 25.110 13.855 25.360 14.185 ;
        RECT 26.300 14.155 26.470 14.995 ;
        RECT 27.345 14.790 27.535 14.995 ;
        RECT 28.265 14.875 28.435 15.455 ;
        RECT 28.220 14.825 28.435 14.875 ;
        RECT 26.640 14.415 27.535 14.790 ;
        RECT 28.045 14.745 28.435 14.825 ;
        RECT 28.640 15.495 29.255 16.065 ;
        RECT 29.425 15.725 29.640 16.235 ;
        RECT 29.870 15.725 30.150 16.055 ;
        RECT 30.330 15.725 30.570 16.235 ;
        RECT 25.585 13.985 26.470 14.155 ;
        RECT 26.650 13.685 26.965 14.185 ;
        RECT 27.195 13.855 27.535 14.415 ;
        RECT 27.705 13.685 27.875 14.695 ;
        RECT 28.045 13.900 28.375 14.745 ;
        RECT 28.640 14.475 28.955 15.495 ;
        RECT 29.125 14.825 29.295 15.325 ;
        RECT 29.545 14.995 29.810 15.555 ;
        RECT 29.980 14.825 30.150 15.725 ;
        RECT 30.320 14.995 30.675 15.555 ;
        RECT 31.365 15.510 31.655 16.235 ;
        RECT 32.335 15.580 32.665 16.015 ;
        RECT 32.835 15.625 33.005 16.235 ;
        RECT 32.285 15.495 32.665 15.580 ;
        RECT 33.175 15.495 33.505 16.020 ;
        RECT 33.765 15.705 33.975 16.235 ;
        RECT 34.250 15.785 35.035 15.955 ;
        RECT 35.205 15.785 35.610 15.955 ;
        RECT 32.285 15.455 32.510 15.495 ;
        RECT 32.285 14.875 32.455 15.455 ;
        RECT 33.175 15.325 33.375 15.495 ;
        RECT 34.250 15.325 34.420 15.785 ;
        RECT 32.625 14.995 33.375 15.325 ;
        RECT 33.545 14.995 34.420 15.325 ;
        RECT 29.125 14.655 30.550 14.825 ;
        RECT 28.640 13.855 29.175 14.475 ;
        RECT 29.345 13.685 29.675 14.485 ;
        RECT 30.160 14.480 30.550 14.655 ;
        RECT 31.365 13.685 31.655 14.850 ;
        RECT 32.285 14.825 32.500 14.875 ;
        RECT 32.285 14.745 32.675 14.825 ;
        RECT 32.345 13.900 32.675 14.745 ;
        RECT 33.185 14.790 33.375 14.995 ;
        RECT 32.845 13.685 33.015 14.695 ;
        RECT 33.185 14.415 34.080 14.790 ;
        RECT 33.185 13.855 33.525 14.415 ;
        RECT 33.755 13.685 34.070 14.185 ;
        RECT 34.250 14.155 34.420 14.995 ;
        RECT 34.590 15.285 35.055 15.615 ;
        RECT 35.440 15.555 35.610 15.785 ;
        RECT 35.790 15.735 36.160 16.235 ;
        RECT 36.480 15.785 37.155 15.955 ;
        RECT 37.350 15.785 37.685 15.955 ;
        RECT 34.590 14.325 34.910 15.285 ;
        RECT 35.440 15.255 36.270 15.555 ;
        RECT 35.080 14.355 35.270 15.075 ;
        RECT 35.440 14.185 35.610 15.255 ;
        RECT 36.070 15.225 36.270 15.255 ;
        RECT 35.780 15.005 35.950 15.075 ;
        RECT 36.480 15.005 36.650 15.785 ;
        RECT 37.515 15.645 37.685 15.785 ;
        RECT 37.855 15.775 38.105 16.235 ;
        RECT 35.780 14.835 36.650 15.005 ;
        RECT 36.820 15.365 37.345 15.585 ;
        RECT 37.515 15.515 37.740 15.645 ;
        RECT 35.780 14.745 36.290 14.835 ;
        RECT 34.250 13.985 35.135 14.155 ;
        RECT 35.360 13.855 35.610 14.185 ;
        RECT 35.780 13.685 35.950 14.485 ;
        RECT 36.120 14.130 36.290 14.745 ;
        RECT 36.820 14.665 36.990 15.365 ;
        RECT 36.460 14.300 36.990 14.665 ;
        RECT 37.160 14.600 37.400 15.195 ;
        RECT 37.570 14.410 37.740 15.515 ;
        RECT 37.910 14.655 38.190 15.605 ;
        RECT 37.435 14.280 37.740 14.410 ;
        RECT 36.120 13.960 37.225 14.130 ;
        RECT 37.435 13.855 37.685 14.280 ;
        RECT 37.855 13.685 38.120 14.145 ;
        RECT 38.360 13.855 38.545 15.975 ;
        RECT 38.715 15.855 39.045 16.235 ;
        RECT 39.215 15.685 39.385 15.975 ;
        RECT 38.720 15.515 39.385 15.685 ;
        RECT 40.195 15.685 40.365 15.975 ;
        RECT 40.535 15.855 40.865 16.235 ;
        RECT 40.195 15.515 40.860 15.685 ;
        RECT 38.720 14.525 38.950 15.515 ;
        RECT 39.120 14.695 39.470 15.345 ;
        RECT 40.110 14.695 40.460 15.345 ;
        RECT 40.630 14.525 40.860 15.515 ;
        RECT 38.720 14.355 39.385 14.525 ;
        RECT 38.715 13.685 39.045 14.185 ;
        RECT 39.215 13.855 39.385 14.355 ;
        RECT 40.195 14.355 40.860 14.525 ;
        RECT 40.195 13.855 40.365 14.355 ;
        RECT 40.535 13.685 40.865 14.185 ;
        RECT 41.035 13.855 41.220 15.975 ;
        RECT 41.475 15.775 41.725 16.235 ;
        RECT 41.895 15.785 42.230 15.955 ;
        RECT 42.425 15.785 43.100 15.955 ;
        RECT 41.895 15.645 42.065 15.785 ;
        RECT 41.390 14.655 41.670 15.605 ;
        RECT 41.840 15.515 42.065 15.645 ;
        RECT 41.840 14.410 42.010 15.515 ;
        RECT 42.235 15.365 42.760 15.585 ;
        RECT 42.180 14.600 42.420 15.195 ;
        RECT 42.590 14.665 42.760 15.365 ;
        RECT 42.930 15.005 43.100 15.785 ;
        RECT 43.420 15.735 43.790 16.235 ;
        RECT 43.970 15.785 44.375 15.955 ;
        RECT 44.545 15.785 45.330 15.955 ;
        RECT 43.970 15.555 44.140 15.785 ;
        RECT 43.310 15.255 44.140 15.555 ;
        RECT 44.525 15.285 44.990 15.615 ;
        RECT 43.310 15.225 43.510 15.255 ;
        RECT 43.630 15.005 43.800 15.075 ;
        RECT 42.930 14.835 43.800 15.005 ;
        RECT 43.290 14.745 43.800 14.835 ;
        RECT 41.840 14.280 42.145 14.410 ;
        RECT 42.590 14.300 43.120 14.665 ;
        RECT 41.460 13.685 41.725 14.145 ;
        RECT 41.895 13.855 42.145 14.280 ;
        RECT 43.290 14.130 43.460 14.745 ;
        RECT 42.355 13.960 43.460 14.130 ;
        RECT 43.630 13.685 43.800 14.485 ;
        RECT 43.970 14.185 44.140 15.255 ;
        RECT 44.310 14.355 44.500 15.075 ;
        RECT 44.670 14.325 44.990 15.285 ;
        RECT 45.160 15.325 45.330 15.785 ;
        RECT 45.605 15.705 45.815 16.235 ;
        RECT 46.075 15.495 46.405 16.020 ;
        RECT 46.575 15.625 46.745 16.235 ;
        RECT 46.915 15.580 47.245 16.015 ;
        RECT 47.555 15.685 47.725 15.975 ;
        RECT 47.895 15.855 48.225 16.235 ;
        RECT 46.915 15.495 47.295 15.580 ;
        RECT 47.555 15.515 48.220 15.685 ;
        RECT 46.205 15.325 46.405 15.495 ;
        RECT 47.070 15.455 47.295 15.495 ;
        RECT 45.160 14.995 46.035 15.325 ;
        RECT 46.205 14.995 46.955 15.325 ;
        RECT 43.970 13.855 44.220 14.185 ;
        RECT 45.160 14.155 45.330 14.995 ;
        RECT 46.205 14.790 46.395 14.995 ;
        RECT 47.125 14.875 47.295 15.455 ;
        RECT 47.080 14.825 47.295 14.875 ;
        RECT 45.500 14.415 46.395 14.790 ;
        RECT 46.905 14.745 47.295 14.825 ;
        RECT 44.445 13.985 45.330 14.155 ;
        RECT 45.510 13.685 45.825 14.185 ;
        RECT 46.055 13.855 46.395 14.415 ;
        RECT 46.565 13.685 46.735 14.695 ;
        RECT 46.905 13.900 47.235 14.745 ;
        RECT 47.470 14.695 47.820 15.345 ;
        RECT 47.990 14.525 48.220 15.515 ;
        RECT 47.555 14.355 48.220 14.525 ;
        RECT 47.555 13.855 47.725 14.355 ;
        RECT 47.895 13.685 48.225 14.185 ;
        RECT 48.395 13.855 48.580 15.975 ;
        RECT 48.835 15.775 49.085 16.235 ;
        RECT 49.255 15.785 49.590 15.955 ;
        RECT 49.785 15.785 50.460 15.955 ;
        RECT 49.255 15.645 49.425 15.785 ;
        RECT 48.750 14.655 49.030 15.605 ;
        RECT 49.200 15.515 49.425 15.645 ;
        RECT 49.200 14.410 49.370 15.515 ;
        RECT 49.595 15.365 50.120 15.585 ;
        RECT 49.540 14.600 49.780 15.195 ;
        RECT 49.950 14.665 50.120 15.365 ;
        RECT 50.290 15.005 50.460 15.785 ;
        RECT 50.780 15.735 51.150 16.235 ;
        RECT 51.330 15.785 51.735 15.955 ;
        RECT 51.905 15.785 52.690 15.955 ;
        RECT 51.330 15.555 51.500 15.785 ;
        RECT 50.670 15.255 51.500 15.555 ;
        RECT 51.885 15.285 52.350 15.615 ;
        RECT 50.670 15.225 50.870 15.255 ;
        RECT 50.990 15.005 51.160 15.075 ;
        RECT 50.290 14.835 51.160 15.005 ;
        RECT 50.650 14.745 51.160 14.835 ;
        RECT 49.200 14.280 49.505 14.410 ;
        RECT 49.950 14.300 50.480 14.665 ;
        RECT 48.820 13.685 49.085 14.145 ;
        RECT 49.255 13.855 49.505 14.280 ;
        RECT 50.650 14.130 50.820 14.745 ;
        RECT 49.715 13.960 50.820 14.130 ;
        RECT 50.990 13.685 51.160 14.485 ;
        RECT 51.330 14.185 51.500 15.255 ;
        RECT 51.670 14.355 51.860 15.075 ;
        RECT 52.030 14.325 52.350 15.285 ;
        RECT 52.520 15.325 52.690 15.785 ;
        RECT 52.965 15.705 53.175 16.235 ;
        RECT 53.435 15.495 53.765 16.020 ;
        RECT 53.935 15.625 54.105 16.235 ;
        RECT 54.275 15.580 54.605 16.015 ;
        RECT 54.275 15.495 54.655 15.580 ;
        RECT 53.565 15.325 53.765 15.495 ;
        RECT 54.430 15.455 54.655 15.495 ;
        RECT 52.520 14.995 53.395 15.325 ;
        RECT 53.565 14.995 54.315 15.325 ;
        RECT 51.330 13.855 51.580 14.185 ;
        RECT 52.520 14.155 52.690 14.995 ;
        RECT 53.565 14.790 53.755 14.995 ;
        RECT 54.485 14.875 54.655 15.455 ;
        RECT 54.440 14.825 54.655 14.875 ;
        RECT 52.860 14.415 53.755 14.790 ;
        RECT 54.265 14.745 54.655 14.825 ;
        RECT 54.860 15.495 55.475 16.065 ;
        RECT 55.645 15.725 55.860 16.235 ;
        RECT 56.090 15.725 56.370 16.055 ;
        RECT 56.550 15.725 56.790 16.235 ;
        RECT 51.805 13.985 52.690 14.155 ;
        RECT 52.870 13.685 53.185 14.185 ;
        RECT 53.415 13.855 53.755 14.415 ;
        RECT 53.925 13.685 54.095 14.695 ;
        RECT 54.265 13.900 54.595 14.745 ;
        RECT 54.860 14.475 55.175 15.495 ;
        RECT 55.345 14.825 55.515 15.325 ;
        RECT 55.765 14.995 56.030 15.555 ;
        RECT 56.200 14.825 56.370 15.725 ;
        RECT 56.540 14.995 56.895 15.555 ;
        RECT 57.125 15.510 57.415 16.235 ;
        RECT 57.585 15.735 57.845 16.065 ;
        RECT 58.015 15.875 58.345 16.235 ;
        RECT 58.600 15.855 59.900 16.065 ;
        RECT 55.345 14.655 56.770 14.825 ;
        RECT 54.860 13.855 55.395 14.475 ;
        RECT 55.565 13.685 55.895 14.485 ;
        RECT 56.380 14.480 56.770 14.655 ;
        RECT 57.125 13.685 57.415 14.850 ;
        RECT 57.585 14.535 57.755 15.735 ;
        RECT 58.600 15.705 58.770 15.855 ;
        RECT 58.015 15.580 58.770 15.705 ;
        RECT 57.925 15.535 58.770 15.580 ;
        RECT 57.925 15.415 58.195 15.535 ;
        RECT 57.925 14.840 58.095 15.415 ;
        RECT 58.325 14.975 58.735 15.280 ;
        RECT 59.025 15.245 59.235 15.645 ;
        RECT 58.905 15.035 59.235 15.245 ;
        RECT 59.480 15.245 59.700 15.645 ;
        RECT 60.175 15.470 60.630 16.235 ;
        RECT 60.805 15.485 62.015 16.235 ;
        RECT 62.275 15.685 62.445 15.975 ;
        RECT 62.615 15.855 62.945 16.235 ;
        RECT 62.275 15.515 62.940 15.685 ;
        RECT 59.480 15.035 59.955 15.245 ;
        RECT 60.145 15.045 60.635 15.245 ;
        RECT 60.805 14.945 61.325 15.485 ;
        RECT 57.925 14.805 58.125 14.840 ;
        RECT 59.455 14.805 60.630 14.865 ;
        RECT 57.925 14.695 60.630 14.805 ;
        RECT 61.495 14.775 62.015 15.315 ;
        RECT 57.985 14.635 59.785 14.695 ;
        RECT 59.455 14.605 59.785 14.635 ;
        RECT 57.585 13.855 57.845 14.535 ;
        RECT 58.015 13.685 58.265 14.465 ;
        RECT 58.515 14.435 59.350 14.445 ;
        RECT 59.940 14.435 60.125 14.525 ;
        RECT 58.515 14.235 60.125 14.435 ;
        RECT 58.515 13.855 58.765 14.235 ;
        RECT 59.895 14.195 60.125 14.235 ;
        RECT 60.375 14.075 60.630 14.695 ;
        RECT 58.935 13.685 59.290 14.065 ;
        RECT 60.295 13.855 60.630 14.075 ;
        RECT 60.805 13.685 62.015 14.775 ;
        RECT 62.190 14.695 62.540 15.345 ;
        RECT 62.710 14.525 62.940 15.515 ;
        RECT 62.275 14.355 62.940 14.525 ;
        RECT 62.275 13.855 62.445 14.355 ;
        RECT 62.615 13.685 62.945 14.185 ;
        RECT 63.115 13.855 63.300 15.975 ;
        RECT 63.555 15.775 63.805 16.235 ;
        RECT 63.975 15.785 64.310 15.955 ;
        RECT 64.505 15.785 65.180 15.955 ;
        RECT 63.975 15.645 64.145 15.785 ;
        RECT 63.470 14.655 63.750 15.605 ;
        RECT 63.920 15.515 64.145 15.645 ;
        RECT 63.920 14.410 64.090 15.515 ;
        RECT 64.315 15.365 64.840 15.585 ;
        RECT 64.260 14.600 64.500 15.195 ;
        RECT 64.670 14.665 64.840 15.365 ;
        RECT 65.010 15.005 65.180 15.785 ;
        RECT 65.500 15.735 65.870 16.235 ;
        RECT 66.050 15.785 66.455 15.955 ;
        RECT 66.625 15.785 67.410 15.955 ;
        RECT 66.050 15.555 66.220 15.785 ;
        RECT 65.390 15.255 66.220 15.555 ;
        RECT 66.605 15.285 67.070 15.615 ;
        RECT 65.390 15.225 65.590 15.255 ;
        RECT 65.710 15.005 65.880 15.075 ;
        RECT 65.010 14.835 65.880 15.005 ;
        RECT 65.370 14.745 65.880 14.835 ;
        RECT 63.920 14.280 64.225 14.410 ;
        RECT 64.670 14.300 65.200 14.665 ;
        RECT 63.540 13.685 63.805 14.145 ;
        RECT 63.975 13.855 64.225 14.280 ;
        RECT 65.370 14.130 65.540 14.745 ;
        RECT 64.435 13.960 65.540 14.130 ;
        RECT 65.710 13.685 65.880 14.485 ;
        RECT 66.050 14.185 66.220 15.255 ;
        RECT 66.390 14.355 66.580 15.075 ;
        RECT 66.750 14.325 67.070 15.285 ;
        RECT 67.240 15.325 67.410 15.785 ;
        RECT 67.685 15.705 67.895 16.235 ;
        RECT 68.155 15.495 68.485 16.020 ;
        RECT 68.655 15.625 68.825 16.235 ;
        RECT 68.995 15.580 69.325 16.015 ;
        RECT 69.710 15.725 69.950 16.235 ;
        RECT 70.130 15.725 70.410 16.055 ;
        RECT 70.640 15.725 70.855 16.235 ;
        RECT 68.995 15.495 69.375 15.580 ;
        RECT 68.285 15.325 68.485 15.495 ;
        RECT 69.150 15.455 69.375 15.495 ;
        RECT 67.240 14.995 68.115 15.325 ;
        RECT 68.285 14.995 69.035 15.325 ;
        RECT 66.050 13.855 66.300 14.185 ;
        RECT 67.240 14.155 67.410 14.995 ;
        RECT 68.285 14.790 68.475 14.995 ;
        RECT 69.205 14.875 69.375 15.455 ;
        RECT 69.605 14.995 69.960 15.555 ;
        RECT 69.160 14.825 69.375 14.875 ;
        RECT 70.130 14.825 70.300 15.725 ;
        RECT 70.470 14.995 70.735 15.555 ;
        RECT 71.025 15.495 71.640 16.065 ;
        RECT 70.985 14.825 71.155 15.325 ;
        RECT 67.580 14.415 68.475 14.790 ;
        RECT 68.985 14.745 69.375 14.825 ;
        RECT 66.525 13.985 67.410 14.155 ;
        RECT 67.590 13.685 67.905 14.185 ;
        RECT 68.135 13.855 68.475 14.415 ;
        RECT 68.645 13.685 68.815 14.695 ;
        RECT 68.985 13.900 69.315 14.745 ;
        RECT 69.730 14.655 71.155 14.825 ;
        RECT 69.730 14.480 70.120 14.655 ;
        RECT 70.605 13.685 70.935 14.485 ;
        RECT 71.325 14.475 71.640 15.495 ;
        RECT 71.845 15.485 73.055 16.235 ;
        RECT 73.315 15.685 73.485 15.975 ;
        RECT 73.655 15.855 73.985 16.235 ;
        RECT 73.315 15.515 73.980 15.685 ;
        RECT 71.845 14.945 72.365 15.485 ;
        RECT 72.535 14.775 73.055 15.315 ;
        RECT 71.105 13.855 71.640 14.475 ;
        RECT 71.845 13.685 73.055 14.775 ;
        RECT 73.230 14.695 73.580 15.345 ;
        RECT 73.750 14.525 73.980 15.515 ;
        RECT 73.315 14.355 73.980 14.525 ;
        RECT 73.315 13.855 73.485 14.355 ;
        RECT 73.655 13.685 73.985 14.185 ;
        RECT 74.155 13.855 74.340 15.975 ;
        RECT 74.595 15.775 74.845 16.235 ;
        RECT 75.015 15.785 75.350 15.955 ;
        RECT 75.545 15.785 76.220 15.955 ;
        RECT 75.015 15.645 75.185 15.785 ;
        RECT 74.510 14.655 74.790 15.605 ;
        RECT 74.960 15.515 75.185 15.645 ;
        RECT 74.960 14.410 75.130 15.515 ;
        RECT 75.355 15.365 75.880 15.585 ;
        RECT 75.300 14.600 75.540 15.195 ;
        RECT 75.710 14.665 75.880 15.365 ;
        RECT 76.050 15.005 76.220 15.785 ;
        RECT 76.540 15.735 76.910 16.235 ;
        RECT 77.090 15.785 77.495 15.955 ;
        RECT 77.665 15.785 78.450 15.955 ;
        RECT 77.090 15.555 77.260 15.785 ;
        RECT 76.430 15.255 77.260 15.555 ;
        RECT 77.645 15.285 78.110 15.615 ;
        RECT 76.430 15.225 76.630 15.255 ;
        RECT 76.750 15.005 76.920 15.075 ;
        RECT 76.050 14.835 76.920 15.005 ;
        RECT 76.410 14.745 76.920 14.835 ;
        RECT 74.960 14.280 75.265 14.410 ;
        RECT 75.710 14.300 76.240 14.665 ;
        RECT 74.580 13.685 74.845 14.145 ;
        RECT 75.015 13.855 75.265 14.280 ;
        RECT 76.410 14.130 76.580 14.745 ;
        RECT 75.475 13.960 76.580 14.130 ;
        RECT 76.750 13.685 76.920 14.485 ;
        RECT 77.090 14.185 77.260 15.255 ;
        RECT 77.430 14.355 77.620 15.075 ;
        RECT 77.790 14.325 78.110 15.285 ;
        RECT 78.280 15.325 78.450 15.785 ;
        RECT 78.725 15.705 78.935 16.235 ;
        RECT 79.195 15.495 79.525 16.020 ;
        RECT 79.695 15.625 79.865 16.235 ;
        RECT 80.035 15.580 80.365 16.015 ;
        RECT 80.675 15.685 80.845 16.065 ;
        RECT 81.060 15.855 81.390 16.235 ;
        RECT 80.035 15.495 80.415 15.580 ;
        RECT 80.675 15.515 81.390 15.685 ;
        RECT 79.325 15.325 79.525 15.495 ;
        RECT 80.190 15.455 80.415 15.495 ;
        RECT 78.280 14.995 79.155 15.325 ;
        RECT 79.325 14.995 80.075 15.325 ;
        RECT 77.090 13.855 77.340 14.185 ;
        RECT 78.280 14.155 78.450 14.995 ;
        RECT 79.325 14.790 79.515 14.995 ;
        RECT 80.245 14.875 80.415 15.455 ;
        RECT 80.585 14.965 80.940 15.335 ;
        RECT 81.220 15.325 81.390 15.515 ;
        RECT 81.560 15.490 81.815 16.065 ;
        RECT 81.220 14.995 81.475 15.325 ;
        RECT 80.200 14.825 80.415 14.875 ;
        RECT 78.620 14.415 79.515 14.790 ;
        RECT 80.025 14.745 80.415 14.825 ;
        RECT 81.220 14.785 81.390 14.995 ;
        RECT 77.565 13.985 78.450 14.155 ;
        RECT 78.630 13.685 78.945 14.185 ;
        RECT 79.175 13.855 79.515 14.415 ;
        RECT 79.685 13.685 79.855 14.695 ;
        RECT 80.025 13.900 80.355 14.745 ;
        RECT 80.675 14.615 81.390 14.785 ;
        RECT 81.645 14.760 81.815 15.490 ;
        RECT 81.990 15.395 82.250 16.235 ;
        RECT 82.885 15.485 84.095 16.235 ;
        RECT 80.675 13.855 80.845 14.615 ;
        RECT 81.060 13.685 81.390 14.445 ;
        RECT 81.560 13.855 81.815 14.760 ;
        RECT 81.990 13.685 82.250 14.835 ;
        RECT 82.885 14.775 83.405 15.315 ;
        RECT 83.575 14.945 84.095 15.485 ;
        RECT 82.885 13.685 84.095 14.775 ;
        RECT 5.520 13.515 84.180 13.685 ;
        RECT 5.605 12.425 6.815 13.515 ;
        RECT 7.075 12.845 7.245 13.345 ;
        RECT 7.415 13.015 7.745 13.515 ;
        RECT 7.075 12.675 7.740 12.845 ;
        RECT 5.605 11.715 6.125 12.255 ;
        RECT 6.295 11.885 6.815 12.425 ;
        RECT 6.990 11.855 7.340 12.505 ;
        RECT 5.605 10.965 6.815 11.715 ;
        RECT 7.510 11.685 7.740 12.675 ;
        RECT 7.075 11.515 7.740 11.685 ;
        RECT 7.075 11.225 7.245 11.515 ;
        RECT 7.415 10.965 7.745 11.345 ;
        RECT 7.915 11.225 8.100 13.345 ;
        RECT 8.340 13.055 8.605 13.515 ;
        RECT 8.775 12.920 9.025 13.345 ;
        RECT 9.235 13.070 10.340 13.240 ;
        RECT 8.720 12.790 9.025 12.920 ;
        RECT 8.270 11.595 8.550 12.545 ;
        RECT 8.720 11.685 8.890 12.790 ;
        RECT 9.060 12.005 9.300 12.600 ;
        RECT 9.470 12.535 10.000 12.900 ;
        RECT 9.470 11.835 9.640 12.535 ;
        RECT 10.170 12.455 10.340 13.070 ;
        RECT 10.510 12.715 10.680 13.515 ;
        RECT 10.850 13.015 11.100 13.345 ;
        RECT 11.325 13.045 12.210 13.215 ;
        RECT 10.170 12.365 10.680 12.455 ;
        RECT 8.720 11.555 8.945 11.685 ;
        RECT 9.115 11.615 9.640 11.835 ;
        RECT 9.810 12.195 10.680 12.365 ;
        RECT 8.355 10.965 8.605 11.425 ;
        RECT 8.775 11.415 8.945 11.555 ;
        RECT 9.810 11.415 9.980 12.195 ;
        RECT 10.510 12.125 10.680 12.195 ;
        RECT 10.190 11.945 10.390 11.975 ;
        RECT 10.850 11.945 11.020 13.015 ;
        RECT 11.190 12.125 11.380 12.845 ;
        RECT 10.190 11.645 11.020 11.945 ;
        RECT 11.550 11.915 11.870 12.875 ;
        RECT 8.775 11.245 9.110 11.415 ;
        RECT 9.305 11.245 9.980 11.415 ;
        RECT 10.300 10.965 10.670 11.465 ;
        RECT 10.850 11.415 11.020 11.645 ;
        RECT 11.405 11.585 11.870 11.915 ;
        RECT 12.040 12.205 12.210 13.045 ;
        RECT 12.390 13.015 12.705 13.515 ;
        RECT 12.935 12.785 13.275 13.345 ;
        RECT 12.380 12.410 13.275 12.785 ;
        RECT 13.445 12.505 13.615 13.515 ;
        RECT 13.085 12.205 13.275 12.410 ;
        RECT 13.785 12.455 14.115 13.300 ;
        RECT 15.300 12.725 15.835 13.345 ;
        RECT 13.785 12.375 14.175 12.455 ;
        RECT 13.960 12.325 14.175 12.375 ;
        RECT 12.040 11.875 12.915 12.205 ;
        RECT 13.085 11.875 13.835 12.205 ;
        RECT 12.040 11.415 12.210 11.875 ;
        RECT 13.085 11.705 13.285 11.875 ;
        RECT 14.005 11.745 14.175 12.325 ;
        RECT 13.950 11.705 14.175 11.745 ;
        RECT 10.850 11.245 11.255 11.415 ;
        RECT 11.425 11.245 12.210 11.415 ;
        RECT 12.485 10.965 12.695 11.495 ;
        RECT 12.955 11.180 13.285 11.705 ;
        RECT 13.795 11.620 14.175 11.705 ;
        RECT 15.300 11.705 15.615 12.725 ;
        RECT 16.005 12.715 16.335 13.515 ;
        RECT 16.820 12.545 17.210 12.720 ;
        RECT 15.785 12.375 17.210 12.545 ;
        RECT 15.785 11.875 15.955 12.375 ;
        RECT 13.455 10.965 13.625 11.575 ;
        RECT 13.795 11.185 14.125 11.620 ;
        RECT 15.300 11.135 15.915 11.705 ;
        RECT 16.205 11.645 16.470 12.205 ;
        RECT 16.640 11.475 16.810 12.375 ;
        RECT 18.485 12.350 18.775 13.515 ;
        RECT 19.870 12.365 20.130 13.515 ;
        RECT 20.305 12.440 20.560 13.345 ;
        RECT 20.730 12.755 21.060 13.515 ;
        RECT 21.275 12.585 21.445 13.345 ;
        RECT 16.980 11.645 17.335 12.205 ;
        RECT 16.085 10.965 16.300 11.475 ;
        RECT 16.530 11.145 16.810 11.475 ;
        RECT 16.990 10.965 17.230 11.475 ;
        RECT 18.485 10.965 18.775 11.690 ;
        RECT 19.870 10.965 20.130 11.805 ;
        RECT 20.305 11.710 20.475 12.440 ;
        RECT 20.730 12.415 21.445 12.585 ;
        RECT 20.730 12.205 20.900 12.415 ;
        RECT 22.170 12.365 22.430 13.515 ;
        RECT 22.605 12.440 22.860 13.345 ;
        RECT 23.030 12.755 23.360 13.515 ;
        RECT 23.575 12.585 23.745 13.345 ;
        RECT 20.645 11.875 20.900 12.205 ;
        RECT 20.305 11.135 20.560 11.710 ;
        RECT 20.730 11.685 20.900 11.875 ;
        RECT 21.180 11.865 21.535 12.235 ;
        RECT 20.730 11.515 21.445 11.685 ;
        RECT 20.730 10.965 21.060 11.345 ;
        RECT 21.275 11.135 21.445 11.515 ;
        RECT 22.170 10.965 22.430 11.805 ;
        RECT 22.605 11.710 22.775 12.440 ;
        RECT 23.030 12.415 23.745 12.585 ;
        RECT 23.030 12.205 23.200 12.415 ;
        RECT 24.010 12.365 24.270 13.515 ;
        RECT 24.445 12.440 24.700 13.345 ;
        RECT 24.870 12.755 25.200 13.515 ;
        RECT 25.415 12.585 25.585 13.345 ;
        RECT 22.945 11.875 23.200 12.205 ;
        RECT 22.605 11.135 22.860 11.710 ;
        RECT 23.030 11.685 23.200 11.875 ;
        RECT 23.480 11.865 23.835 12.235 ;
        RECT 23.030 11.515 23.745 11.685 ;
        RECT 23.030 10.965 23.360 11.345 ;
        RECT 23.575 11.135 23.745 11.515 ;
        RECT 24.010 10.965 24.270 11.805 ;
        RECT 24.445 11.710 24.615 12.440 ;
        RECT 24.870 12.415 25.585 12.585 ;
        RECT 24.870 12.205 25.040 12.415 ;
        RECT 25.850 12.365 26.110 13.515 ;
        RECT 26.285 12.440 26.540 13.345 ;
        RECT 26.710 12.755 27.040 13.515 ;
        RECT 27.255 12.585 27.425 13.345 ;
        RECT 24.785 11.875 25.040 12.205 ;
        RECT 24.445 11.135 24.700 11.710 ;
        RECT 24.870 11.685 25.040 11.875 ;
        RECT 25.320 11.865 25.675 12.235 ;
        RECT 24.870 11.515 25.585 11.685 ;
        RECT 24.870 10.965 25.200 11.345 ;
        RECT 25.415 11.135 25.585 11.515 ;
        RECT 25.850 10.965 26.110 11.805 ;
        RECT 26.285 11.710 26.455 12.440 ;
        RECT 26.710 12.415 27.425 12.585 ;
        RECT 26.710 12.205 26.880 12.415 ;
        RECT 27.690 12.365 27.950 13.515 ;
        RECT 28.125 12.440 28.380 13.345 ;
        RECT 28.550 12.755 28.880 13.515 ;
        RECT 29.095 12.585 29.265 13.345 ;
        RECT 26.625 11.875 26.880 12.205 ;
        RECT 26.285 11.135 26.540 11.710 ;
        RECT 26.710 11.685 26.880 11.875 ;
        RECT 27.160 11.865 27.515 12.235 ;
        RECT 26.710 11.515 27.425 11.685 ;
        RECT 26.710 10.965 27.040 11.345 ;
        RECT 27.255 11.135 27.425 11.515 ;
        RECT 27.690 10.965 27.950 11.805 ;
        RECT 28.125 11.710 28.295 12.440 ;
        RECT 28.550 12.415 29.265 12.585 ;
        RECT 28.550 12.205 28.720 12.415 ;
        RECT 29.530 12.365 29.790 13.515 ;
        RECT 29.965 12.440 30.220 13.345 ;
        RECT 30.390 12.755 30.720 13.515 ;
        RECT 30.935 12.585 31.105 13.345 ;
        RECT 28.465 11.875 28.720 12.205 ;
        RECT 28.125 11.135 28.380 11.710 ;
        RECT 28.550 11.685 28.720 11.875 ;
        RECT 29.000 11.865 29.355 12.235 ;
        RECT 28.550 11.515 29.265 11.685 ;
        RECT 28.550 10.965 28.880 11.345 ;
        RECT 29.095 11.135 29.265 11.515 ;
        RECT 29.530 10.965 29.790 11.805 ;
        RECT 29.965 11.710 30.135 12.440 ;
        RECT 30.390 12.415 31.105 12.585 ;
        RECT 30.390 12.205 30.560 12.415 ;
        RECT 31.365 12.350 31.655 13.515 ;
        RECT 32.750 13.125 33.085 13.345 ;
        RECT 34.090 13.135 34.445 13.515 ;
        RECT 32.750 12.505 33.005 13.125 ;
        RECT 33.255 12.965 33.485 13.005 ;
        RECT 34.615 12.965 34.865 13.345 ;
        RECT 33.255 12.765 34.865 12.965 ;
        RECT 33.255 12.675 33.440 12.765 ;
        RECT 34.030 12.755 34.865 12.765 ;
        RECT 35.115 12.735 35.365 13.515 ;
        RECT 35.535 12.665 35.795 13.345 ;
        RECT 33.595 12.565 33.925 12.595 ;
        RECT 33.595 12.505 35.395 12.565 ;
        RECT 32.750 12.395 35.455 12.505 ;
        RECT 32.750 12.335 33.925 12.395 ;
        RECT 35.255 12.360 35.455 12.395 ;
        RECT 30.305 11.875 30.560 12.205 ;
        RECT 29.965 11.135 30.220 11.710 ;
        RECT 30.390 11.685 30.560 11.875 ;
        RECT 30.840 11.865 31.195 12.235 ;
        RECT 32.745 11.955 33.235 12.155 ;
        RECT 33.425 11.955 33.900 12.165 ;
        RECT 30.390 11.515 31.105 11.685 ;
        RECT 30.390 10.965 30.720 11.345 ;
        RECT 30.935 11.135 31.105 11.515 ;
        RECT 31.365 10.965 31.655 11.690 ;
        RECT 32.750 10.965 33.205 11.730 ;
        RECT 33.680 11.555 33.900 11.955 ;
        RECT 34.145 11.955 34.475 12.165 ;
        RECT 34.145 11.555 34.355 11.955 ;
        RECT 34.645 11.920 35.055 12.225 ;
        RECT 35.285 11.785 35.455 12.360 ;
        RECT 35.185 11.665 35.455 11.785 ;
        RECT 34.610 11.620 35.455 11.665 ;
        RECT 34.610 11.495 35.365 11.620 ;
        RECT 34.610 11.345 34.780 11.495 ;
        RECT 35.625 11.465 35.795 12.665 ;
        RECT 36.150 12.545 36.540 12.720 ;
        RECT 37.025 12.715 37.355 13.515 ;
        RECT 37.525 12.725 38.060 13.345 ;
        RECT 36.150 12.375 37.575 12.545 ;
        RECT 36.025 11.645 36.380 12.205 ;
        RECT 36.550 11.475 36.720 12.375 ;
        RECT 36.890 11.645 37.155 12.205 ;
        RECT 37.405 11.875 37.575 12.375 ;
        RECT 37.745 11.705 38.060 12.725 ;
        RECT 38.270 12.365 38.530 13.515 ;
        RECT 38.705 12.440 38.960 13.345 ;
        RECT 39.130 12.755 39.460 13.515 ;
        RECT 39.675 12.585 39.845 13.345 ;
        RECT 33.480 11.135 34.780 11.345 ;
        RECT 35.035 10.965 35.365 11.325 ;
        RECT 35.535 11.135 35.795 11.465 ;
        RECT 36.130 10.965 36.370 11.475 ;
        RECT 36.550 11.145 36.830 11.475 ;
        RECT 37.060 10.965 37.275 11.475 ;
        RECT 37.445 11.135 38.060 11.705 ;
        RECT 38.270 10.965 38.530 11.805 ;
        RECT 38.705 11.710 38.875 12.440 ;
        RECT 39.130 12.415 39.845 12.585 ;
        RECT 40.195 12.585 40.365 13.345 ;
        RECT 40.580 12.755 40.910 13.515 ;
        RECT 40.195 12.415 40.910 12.585 ;
        RECT 41.080 12.440 41.335 13.345 ;
        RECT 39.130 12.205 39.300 12.415 ;
        RECT 39.045 11.875 39.300 12.205 ;
        RECT 38.705 11.135 38.960 11.710 ;
        RECT 39.130 11.685 39.300 11.875 ;
        RECT 39.580 11.865 39.935 12.235 ;
        RECT 40.105 11.865 40.460 12.235 ;
        RECT 40.740 12.205 40.910 12.415 ;
        RECT 40.740 11.875 40.995 12.205 ;
        RECT 40.740 11.685 40.910 11.875 ;
        RECT 41.165 11.710 41.335 12.440 ;
        RECT 41.510 12.365 41.770 13.515 ;
        RECT 42.130 12.545 42.520 12.720 ;
        RECT 43.005 12.715 43.335 13.515 ;
        RECT 43.505 12.725 44.040 13.345 ;
        RECT 42.130 12.375 43.555 12.545 ;
        RECT 39.130 11.515 39.845 11.685 ;
        RECT 39.130 10.965 39.460 11.345 ;
        RECT 39.675 11.135 39.845 11.515 ;
        RECT 40.195 11.515 40.910 11.685 ;
        RECT 40.195 11.135 40.365 11.515 ;
        RECT 40.580 10.965 40.910 11.345 ;
        RECT 41.080 11.135 41.335 11.710 ;
        RECT 41.510 10.965 41.770 11.805 ;
        RECT 42.005 11.645 42.360 12.205 ;
        RECT 42.530 11.475 42.700 12.375 ;
        RECT 42.870 11.645 43.135 12.205 ;
        RECT 43.385 11.875 43.555 12.375 ;
        RECT 43.725 11.705 44.040 12.725 ;
        RECT 44.245 12.350 44.535 13.515 ;
        RECT 45.630 12.365 45.890 13.515 ;
        RECT 46.065 12.440 46.320 13.345 ;
        RECT 46.490 12.755 46.820 13.515 ;
        RECT 47.035 12.585 47.205 13.345 ;
        RECT 42.110 10.965 42.350 11.475 ;
        RECT 42.530 11.145 42.810 11.475 ;
        RECT 43.040 10.965 43.255 11.475 ;
        RECT 43.425 11.135 44.040 11.705 ;
        RECT 44.245 10.965 44.535 11.690 ;
        RECT 45.630 10.965 45.890 11.805 ;
        RECT 46.065 11.710 46.235 12.440 ;
        RECT 46.490 12.415 47.205 12.585 ;
        RECT 47.465 12.425 48.675 13.515 ;
        RECT 46.490 12.205 46.660 12.415 ;
        RECT 46.405 11.875 46.660 12.205 ;
        RECT 46.065 11.135 46.320 11.710 ;
        RECT 46.490 11.685 46.660 11.875 ;
        RECT 46.940 11.865 47.295 12.235 ;
        RECT 47.465 11.715 47.985 12.255 ;
        RECT 48.155 11.885 48.675 12.425 ;
        RECT 48.850 12.365 49.110 13.515 ;
        RECT 49.285 12.440 49.540 13.345 ;
        RECT 49.710 12.755 50.040 13.515 ;
        RECT 50.255 12.585 50.425 13.345 ;
        RECT 46.490 11.515 47.205 11.685 ;
        RECT 46.490 10.965 46.820 11.345 ;
        RECT 47.035 11.135 47.205 11.515 ;
        RECT 47.465 10.965 48.675 11.715 ;
        RECT 48.850 10.965 49.110 11.805 ;
        RECT 49.285 11.710 49.455 12.440 ;
        RECT 49.710 12.415 50.425 12.585 ;
        RECT 50.685 12.425 51.895 13.515 ;
        RECT 49.710 12.205 49.880 12.415 ;
        RECT 49.625 11.875 49.880 12.205 ;
        RECT 49.285 11.135 49.540 11.710 ;
        RECT 49.710 11.685 49.880 11.875 ;
        RECT 50.160 11.865 50.515 12.235 ;
        RECT 50.685 11.715 51.205 12.255 ;
        RECT 51.375 11.885 51.895 12.425 ;
        RECT 52.155 12.585 52.325 13.345 ;
        RECT 52.540 12.755 52.870 13.515 ;
        RECT 52.155 12.415 52.870 12.585 ;
        RECT 53.040 12.440 53.295 13.345 ;
        RECT 52.065 11.865 52.420 12.235 ;
        RECT 52.700 12.205 52.870 12.415 ;
        RECT 52.700 11.875 52.955 12.205 ;
        RECT 49.710 11.515 50.425 11.685 ;
        RECT 49.710 10.965 50.040 11.345 ;
        RECT 50.255 11.135 50.425 11.515 ;
        RECT 50.685 10.965 51.895 11.715 ;
        RECT 52.700 11.685 52.870 11.875 ;
        RECT 53.125 11.710 53.295 12.440 ;
        RECT 53.470 12.365 53.730 13.515 ;
        RECT 53.905 12.425 55.115 13.515 ;
        RECT 52.155 11.515 52.870 11.685 ;
        RECT 52.155 11.135 52.325 11.515 ;
        RECT 52.540 10.965 52.870 11.345 ;
        RECT 53.040 11.135 53.295 11.710 ;
        RECT 53.470 10.965 53.730 11.805 ;
        RECT 53.905 11.715 54.425 12.255 ;
        RECT 54.595 11.885 55.115 12.425 ;
        RECT 55.290 12.365 55.550 13.515 ;
        RECT 55.725 12.440 55.980 13.345 ;
        RECT 56.150 12.755 56.480 13.515 ;
        RECT 56.695 12.585 56.865 13.345 ;
        RECT 53.905 10.965 55.115 11.715 ;
        RECT 55.290 10.965 55.550 11.805 ;
        RECT 55.725 11.710 55.895 12.440 ;
        RECT 56.150 12.415 56.865 12.585 ;
        RECT 56.150 12.205 56.320 12.415 ;
        RECT 57.125 12.350 57.415 13.515 ;
        RECT 58.510 12.365 58.770 13.515 ;
        RECT 58.945 12.440 59.200 13.345 ;
        RECT 59.370 12.755 59.700 13.515 ;
        RECT 59.915 12.585 60.085 13.345 ;
        RECT 56.065 11.875 56.320 12.205 ;
        RECT 55.725 11.135 55.980 11.710 ;
        RECT 56.150 11.685 56.320 11.875 ;
        RECT 56.600 11.865 56.955 12.235 ;
        RECT 56.150 11.515 56.865 11.685 ;
        RECT 56.150 10.965 56.480 11.345 ;
        RECT 56.695 11.135 56.865 11.515 ;
        RECT 57.125 10.965 57.415 11.690 ;
        RECT 58.510 10.965 58.770 11.805 ;
        RECT 58.945 11.710 59.115 12.440 ;
        RECT 59.370 12.415 60.085 12.585 ;
        RECT 60.345 12.425 61.555 13.515 ;
        RECT 59.370 12.205 59.540 12.415 ;
        RECT 59.285 11.875 59.540 12.205 ;
        RECT 58.945 11.135 59.200 11.710 ;
        RECT 59.370 11.685 59.540 11.875 ;
        RECT 59.820 11.865 60.175 12.235 ;
        RECT 60.345 11.715 60.865 12.255 ;
        RECT 61.035 11.885 61.555 12.425 ;
        RECT 61.730 12.365 61.990 13.515 ;
        RECT 62.165 12.440 62.420 13.345 ;
        RECT 62.590 12.755 62.920 13.515 ;
        RECT 63.135 12.585 63.305 13.345 ;
        RECT 59.370 11.515 60.085 11.685 ;
        RECT 59.370 10.965 59.700 11.345 ;
        RECT 59.915 11.135 60.085 11.515 ;
        RECT 60.345 10.965 61.555 11.715 ;
        RECT 61.730 10.965 61.990 11.805 ;
        RECT 62.165 11.710 62.335 12.440 ;
        RECT 62.590 12.415 63.305 12.585 ;
        RECT 63.565 12.425 64.775 13.515 ;
        RECT 62.590 12.205 62.760 12.415 ;
        RECT 62.505 11.875 62.760 12.205 ;
        RECT 62.165 11.135 62.420 11.710 ;
        RECT 62.590 11.685 62.760 11.875 ;
        RECT 63.040 11.865 63.395 12.235 ;
        RECT 63.565 11.715 64.085 12.255 ;
        RECT 64.255 11.885 64.775 12.425 ;
        RECT 65.035 12.585 65.205 13.345 ;
        RECT 65.420 12.755 65.750 13.515 ;
        RECT 65.035 12.415 65.750 12.585 ;
        RECT 65.920 12.440 66.175 13.345 ;
        RECT 64.945 11.865 65.300 12.235 ;
        RECT 65.580 12.205 65.750 12.415 ;
        RECT 65.580 11.875 65.835 12.205 ;
        RECT 62.590 11.515 63.305 11.685 ;
        RECT 62.590 10.965 62.920 11.345 ;
        RECT 63.135 11.135 63.305 11.515 ;
        RECT 63.565 10.965 64.775 11.715 ;
        RECT 65.580 11.685 65.750 11.875 ;
        RECT 66.005 11.710 66.175 12.440 ;
        RECT 66.350 12.365 66.610 13.515 ;
        RECT 66.785 12.425 67.995 13.515 ;
        RECT 65.035 11.515 65.750 11.685 ;
        RECT 65.035 11.135 65.205 11.515 ;
        RECT 65.420 10.965 65.750 11.345 ;
        RECT 65.920 11.135 66.175 11.710 ;
        RECT 66.350 10.965 66.610 11.805 ;
        RECT 66.785 11.715 67.305 12.255 ;
        RECT 67.475 11.885 67.995 12.425 ;
        RECT 68.170 12.365 68.430 13.515 ;
        RECT 68.605 12.440 68.860 13.345 ;
        RECT 69.030 12.755 69.360 13.515 ;
        RECT 69.575 12.585 69.745 13.345 ;
        RECT 66.785 10.965 67.995 11.715 ;
        RECT 68.170 10.965 68.430 11.805 ;
        RECT 68.605 11.710 68.775 12.440 ;
        RECT 69.030 12.415 69.745 12.585 ;
        RECT 69.030 12.205 69.200 12.415 ;
        RECT 70.005 12.350 70.295 13.515 ;
        RECT 70.650 12.545 71.040 12.720 ;
        RECT 71.525 12.715 71.855 13.515 ;
        RECT 72.025 12.725 72.560 13.345 ;
        RECT 70.650 12.375 72.075 12.545 ;
        RECT 68.945 11.875 69.200 12.205 ;
        RECT 68.605 11.135 68.860 11.710 ;
        RECT 69.030 11.685 69.200 11.875 ;
        RECT 69.480 11.865 69.835 12.235 ;
        RECT 69.030 11.515 69.745 11.685 ;
        RECT 69.030 10.965 69.360 11.345 ;
        RECT 69.575 11.135 69.745 11.515 ;
        RECT 70.005 10.965 70.295 11.690 ;
        RECT 70.525 11.645 70.880 12.205 ;
        RECT 71.050 11.475 71.220 12.375 ;
        RECT 71.390 11.645 71.655 12.205 ;
        RECT 71.905 11.875 72.075 12.375 ;
        RECT 72.245 11.705 72.560 12.725 ;
        RECT 72.950 12.545 73.340 12.720 ;
        RECT 73.825 12.715 74.155 13.515 ;
        RECT 74.325 12.725 74.860 13.345 ;
        RECT 72.950 12.375 74.375 12.545 ;
        RECT 70.630 10.965 70.870 11.475 ;
        RECT 71.050 11.145 71.330 11.475 ;
        RECT 71.560 10.965 71.775 11.475 ;
        RECT 71.945 11.135 72.560 11.705 ;
        RECT 72.825 11.645 73.180 12.205 ;
        RECT 73.350 11.475 73.520 12.375 ;
        RECT 73.690 11.645 73.955 12.205 ;
        RECT 74.205 11.875 74.375 12.375 ;
        RECT 74.545 11.705 74.860 12.725 ;
        RECT 75.615 12.845 75.785 13.345 ;
        RECT 75.955 13.015 76.285 13.515 ;
        RECT 75.615 12.675 76.280 12.845 ;
        RECT 75.530 11.855 75.880 12.505 ;
        RECT 72.930 10.965 73.170 11.475 ;
        RECT 73.350 11.145 73.630 11.475 ;
        RECT 73.860 10.965 74.075 11.475 ;
        RECT 74.245 11.135 74.860 11.705 ;
        RECT 76.050 11.685 76.280 12.675 ;
        RECT 75.615 11.515 76.280 11.685 ;
        RECT 75.615 11.225 75.785 11.515 ;
        RECT 75.955 10.965 76.285 11.345 ;
        RECT 76.455 11.225 76.640 13.345 ;
        RECT 76.880 13.055 77.145 13.515 ;
        RECT 77.315 12.920 77.565 13.345 ;
        RECT 77.775 13.070 78.880 13.240 ;
        RECT 77.260 12.790 77.565 12.920 ;
        RECT 76.810 11.595 77.090 12.545 ;
        RECT 77.260 11.685 77.430 12.790 ;
        RECT 77.600 12.005 77.840 12.600 ;
        RECT 78.010 12.535 78.540 12.900 ;
        RECT 78.010 11.835 78.180 12.535 ;
        RECT 78.710 12.455 78.880 13.070 ;
        RECT 79.050 12.715 79.220 13.515 ;
        RECT 79.390 13.015 79.640 13.345 ;
        RECT 79.865 13.045 80.750 13.215 ;
        RECT 78.710 12.365 79.220 12.455 ;
        RECT 77.260 11.555 77.485 11.685 ;
        RECT 77.655 11.615 78.180 11.835 ;
        RECT 78.350 12.195 79.220 12.365 ;
        RECT 76.895 10.965 77.145 11.425 ;
        RECT 77.315 11.415 77.485 11.555 ;
        RECT 78.350 11.415 78.520 12.195 ;
        RECT 79.050 12.125 79.220 12.195 ;
        RECT 78.730 11.945 78.930 11.975 ;
        RECT 79.390 11.945 79.560 13.015 ;
        RECT 79.730 12.125 79.920 12.845 ;
        RECT 78.730 11.645 79.560 11.945 ;
        RECT 80.090 11.915 80.410 12.875 ;
        RECT 77.315 11.245 77.650 11.415 ;
        RECT 77.845 11.245 78.520 11.415 ;
        RECT 78.840 10.965 79.210 11.465 ;
        RECT 79.390 11.415 79.560 11.645 ;
        RECT 79.945 11.585 80.410 11.915 ;
        RECT 80.580 12.205 80.750 13.045 ;
        RECT 80.930 13.015 81.245 13.515 ;
        RECT 81.475 12.785 81.815 13.345 ;
        RECT 80.920 12.410 81.815 12.785 ;
        RECT 81.985 12.505 82.155 13.515 ;
        RECT 81.625 12.205 81.815 12.410 ;
        RECT 82.325 12.455 82.655 13.300 ;
        RECT 82.325 12.375 82.715 12.455 ;
        RECT 82.500 12.325 82.715 12.375 ;
        RECT 80.580 11.875 81.455 12.205 ;
        RECT 81.625 11.875 82.375 12.205 ;
        RECT 80.580 11.415 80.750 11.875 ;
        RECT 81.625 11.705 81.825 11.875 ;
        RECT 82.545 11.745 82.715 12.325 ;
        RECT 82.885 12.425 84.095 13.515 ;
        RECT 82.885 11.885 83.405 12.425 ;
        RECT 82.490 11.705 82.715 11.745 ;
        RECT 83.575 11.715 84.095 12.255 ;
        RECT 79.390 11.245 79.795 11.415 ;
        RECT 79.965 11.245 80.750 11.415 ;
        RECT 81.025 10.965 81.235 11.495 ;
        RECT 81.495 11.180 81.825 11.705 ;
        RECT 82.335 11.620 82.715 11.705 ;
        RECT 81.995 10.965 82.165 11.575 ;
        RECT 82.335 11.185 82.665 11.620 ;
        RECT 82.885 10.965 84.095 11.715 ;
        RECT 5.520 10.795 84.180 10.965 ;
      LAYER met1 ;
        RECT 5.520 198.320 84.180 198.800 ;
        RECT 43.310 198.120 43.630 198.180 ;
        RECT 51.145 198.120 51.435 198.165 ;
        RECT 43.310 197.980 51.435 198.120 ;
        RECT 43.310 197.920 43.630 197.980 ;
        RECT 51.145 197.935 51.435 197.980 ;
        RECT 54.810 197.100 55.130 197.160 ;
        RECT 55.285 197.100 55.575 197.145 ;
        RECT 54.810 196.960 55.575 197.100 ;
        RECT 54.810 196.900 55.130 196.960 ;
        RECT 55.285 196.915 55.575 196.960 ;
        RECT 64.470 197.100 64.790 197.160 ;
        RECT 65.865 197.100 66.155 197.145 ;
        RECT 64.470 196.960 66.155 197.100 ;
        RECT 64.470 196.900 64.790 196.960 ;
        RECT 65.865 196.915 66.155 196.960 ;
        RECT 41.010 196.760 41.330 196.820 ;
        RECT 52.065 196.760 52.355 196.805 ;
        RECT 41.010 196.620 52.355 196.760 ;
        RECT 41.010 196.560 41.330 196.620 ;
        RECT 52.065 196.575 52.355 196.620 ;
        RECT 50.210 196.220 50.530 196.480 ;
        RECT 51.065 196.420 51.355 196.465 ;
        RECT 53.890 196.420 54.210 196.480 ;
        RECT 51.065 196.280 54.210 196.420 ;
        RECT 51.065 196.235 51.355 196.280 ;
        RECT 53.890 196.220 54.210 196.280 ;
        RECT 56.205 196.420 56.495 196.465 ;
        RECT 56.650 196.420 56.970 196.480 ;
        RECT 56.205 196.280 56.970 196.420 ;
        RECT 56.205 196.235 56.495 196.280 ;
        RECT 56.650 196.220 56.970 196.280 ;
        RECT 63.090 196.420 63.410 196.480 ;
        RECT 64.945 196.420 65.235 196.465 ;
        RECT 63.090 196.280 65.235 196.420 ;
        RECT 63.090 196.220 63.410 196.280 ;
        RECT 64.945 196.235 65.235 196.280 ;
        RECT 5.520 195.600 84.180 196.080 ;
        RECT 37.805 195.215 38.095 195.445 ;
        RECT 50.210 195.400 50.530 195.460 ;
        RECT 50.210 195.260 50.900 195.400 ;
        RECT 35.030 195.060 35.350 195.120 ;
        RECT 36.870 195.105 37.190 195.120 ;
        RECT 35.965 195.060 36.255 195.105 ;
        RECT 35.030 194.920 36.255 195.060 ;
        RECT 35.030 194.860 35.350 194.920 ;
        RECT 35.965 194.875 36.255 194.920 ;
        RECT 36.870 194.875 37.255 195.105 ;
        RECT 37.880 195.060 38.020 195.215 ;
        RECT 50.210 195.200 50.530 195.260 ;
        RECT 50.760 195.105 50.900 195.260 ;
        RECT 39.490 195.060 39.780 195.105 ;
        RECT 37.880 194.920 39.780 195.060 ;
        RECT 39.490 194.875 39.780 194.920 ;
        RECT 50.640 194.875 50.930 195.105 ;
        RECT 34.570 194.520 34.890 194.780 ;
        RECT 35.490 194.520 35.810 194.780 ;
        RECT 36.040 194.720 36.180 194.875 ;
        RECT 36.870 194.860 37.190 194.875 ;
        RECT 41.010 194.720 41.330 194.780 ;
        RECT 36.040 194.580 41.330 194.720 ;
        RECT 41.010 194.520 41.330 194.580 ;
        RECT 63.550 194.720 63.870 194.780 ;
        RECT 65.450 194.720 65.740 194.765 ;
        RECT 63.550 194.580 65.740 194.720 ;
        RECT 63.550 194.520 63.870 194.580 ;
        RECT 65.450 194.535 65.740 194.580 ;
        RECT 30.430 194.380 30.750 194.440 ;
        RECT 38.265 194.380 38.555 194.425 ;
        RECT 30.430 194.240 38.555 194.380 ;
        RECT 30.430 194.180 30.750 194.240 ;
        RECT 38.265 194.195 38.555 194.240 ;
        RECT 39.145 194.380 39.435 194.425 ;
        RECT 40.335 194.380 40.625 194.425 ;
        RECT 42.855 194.380 43.145 194.425 ;
        RECT 39.145 194.240 43.145 194.380 ;
        RECT 39.145 194.195 39.435 194.240 ;
        RECT 40.335 194.195 40.625 194.240 ;
        RECT 42.855 194.195 43.145 194.240 ;
        RECT 48.830 194.380 49.150 194.440 ;
        RECT 49.305 194.380 49.595 194.425 ;
        RECT 48.830 194.240 49.595 194.380 ;
        RECT 48.830 194.180 49.150 194.240 ;
        RECT 49.305 194.195 49.595 194.240 ;
        RECT 50.185 194.380 50.475 194.425 ;
        RECT 51.375 194.380 51.665 194.425 ;
        RECT 53.895 194.380 54.185 194.425 ;
        RECT 50.185 194.240 54.185 194.380 ;
        RECT 50.185 194.195 50.475 194.240 ;
        RECT 51.375 194.195 51.665 194.240 ;
        RECT 53.895 194.195 54.185 194.240 ;
        RECT 62.195 194.380 62.485 194.425 ;
        RECT 64.715 194.380 65.005 194.425 ;
        RECT 65.905 194.380 66.195 194.425 ;
        RECT 62.195 194.240 66.195 194.380 ;
        RECT 62.195 194.195 62.485 194.240 ;
        RECT 64.715 194.195 65.005 194.240 ;
        RECT 65.905 194.195 66.195 194.240 ;
        RECT 66.785 194.380 67.075 194.425 ;
        RECT 69.530 194.380 69.850 194.440 ;
        RECT 66.785 194.240 69.850 194.380 ;
        RECT 66.785 194.195 67.075 194.240 ;
        RECT 69.530 194.180 69.850 194.240 ;
        RECT 38.750 194.040 39.040 194.085 ;
        RECT 40.850 194.040 41.140 194.085 ;
        RECT 42.420 194.040 42.710 194.085 ;
        RECT 38.750 193.900 42.710 194.040 ;
        RECT 38.750 193.855 39.040 193.900 ;
        RECT 40.850 193.855 41.140 193.900 ;
        RECT 42.420 193.855 42.710 193.900 ;
        RECT 49.790 194.040 50.080 194.085 ;
        RECT 51.890 194.040 52.180 194.085 ;
        RECT 53.460 194.040 53.750 194.085 ;
        RECT 49.790 193.900 53.750 194.040 ;
        RECT 49.790 193.855 50.080 193.900 ;
        RECT 51.890 193.855 52.180 193.900 ;
        RECT 53.460 193.855 53.750 193.900 ;
        RECT 62.630 194.040 62.920 194.085 ;
        RECT 64.200 194.040 64.490 194.085 ;
        RECT 66.300 194.040 66.590 194.085 ;
        RECT 62.630 193.900 66.590 194.040 ;
        RECT 62.630 193.855 62.920 193.900 ;
        RECT 64.200 193.855 64.490 193.900 ;
        RECT 66.300 193.855 66.590 193.900 ;
        RECT 35.490 193.500 35.810 193.760 ;
        RECT 36.885 193.700 37.175 193.745 ;
        RECT 39.630 193.700 39.950 193.760 ;
        RECT 36.885 193.560 39.950 193.700 ;
        RECT 36.885 193.515 37.175 193.560 ;
        RECT 39.630 193.500 39.950 193.560 ;
        RECT 41.470 193.700 41.790 193.760 ;
        RECT 45.165 193.700 45.455 193.745 ;
        RECT 41.470 193.560 45.455 193.700 ;
        RECT 41.470 193.500 41.790 193.560 ;
        RECT 45.165 193.515 45.455 193.560 ;
        RECT 55.270 193.700 55.590 193.760 ;
        RECT 56.205 193.700 56.495 193.745 ;
        RECT 55.270 193.560 56.495 193.700 ;
        RECT 55.270 193.500 55.590 193.560 ;
        RECT 56.205 193.515 56.495 193.560 ;
        RECT 59.885 193.700 60.175 193.745 ;
        RECT 60.330 193.700 60.650 193.760 ;
        RECT 59.885 193.560 60.650 193.700 ;
        RECT 59.885 193.515 60.175 193.560 ;
        RECT 60.330 193.500 60.650 193.560 ;
        RECT 5.520 192.880 84.180 193.360 ;
        RECT 38.710 192.680 39.030 192.740 ;
        RECT 39.185 192.680 39.475 192.725 ;
        RECT 38.710 192.540 39.475 192.680 ;
        RECT 38.710 192.480 39.030 192.540 ;
        RECT 39.185 192.495 39.475 192.540 ;
        RECT 39.630 192.680 39.950 192.740 ;
        RECT 42.865 192.680 43.155 192.725 ;
        RECT 43.310 192.680 43.630 192.740 ;
        RECT 39.630 192.540 43.630 192.680 ;
        RECT 39.630 192.480 39.950 192.540 ;
        RECT 42.865 192.495 43.155 192.540 ;
        RECT 43.310 192.480 43.630 192.540 ;
        RECT 53.890 192.480 54.210 192.740 ;
        RECT 60.345 192.680 60.635 192.725 ;
        RECT 60.790 192.680 61.110 192.740 ;
        RECT 60.345 192.540 61.110 192.680 ;
        RECT 60.345 192.495 60.635 192.540 ;
        RECT 60.790 192.480 61.110 192.540 ;
        RECT 61.265 192.680 61.555 192.725 ;
        RECT 63.550 192.680 63.870 192.740 ;
        RECT 61.265 192.540 63.870 192.680 ;
        RECT 61.265 192.495 61.555 192.540 ;
        RECT 63.550 192.480 63.870 192.540 ;
        RECT 30.930 192.340 31.220 192.385 ;
        RECT 33.030 192.340 33.320 192.385 ;
        RECT 34.600 192.340 34.890 192.385 ;
        RECT 30.930 192.200 34.890 192.340 ;
        RECT 30.930 192.155 31.220 192.200 ;
        RECT 33.030 192.155 33.320 192.200 ;
        RECT 34.600 192.155 34.890 192.200 ;
        RECT 36.870 192.340 37.190 192.400 ;
        RECT 40.565 192.340 40.855 192.385 ;
        RECT 36.870 192.200 40.855 192.340 ;
        RECT 36.870 192.140 37.190 192.200 ;
        RECT 40.565 192.155 40.855 192.200 ;
        RECT 45.190 192.340 45.480 192.385 ;
        RECT 47.290 192.340 47.580 192.385 ;
        RECT 48.860 192.340 49.150 192.385 ;
        RECT 45.190 192.200 49.150 192.340 ;
        RECT 45.190 192.155 45.480 192.200 ;
        RECT 47.290 192.155 47.580 192.200 ;
        RECT 48.860 192.155 49.150 192.200 ;
        RECT 65.390 192.340 65.680 192.385 ;
        RECT 66.960 192.340 67.250 192.385 ;
        RECT 69.060 192.340 69.350 192.385 ;
        RECT 65.390 192.200 69.350 192.340 ;
        RECT 65.390 192.155 65.680 192.200 ;
        RECT 66.960 192.155 67.250 192.200 ;
        RECT 69.060 192.155 69.350 192.200 ;
        RECT 30.430 191.800 30.750 192.060 ;
        RECT 31.325 192.000 31.615 192.045 ;
        RECT 32.515 192.000 32.805 192.045 ;
        RECT 35.035 192.000 35.325 192.045 ;
        RECT 45.585 192.000 45.875 192.045 ;
        RECT 46.775 192.000 47.065 192.045 ;
        RECT 49.295 192.000 49.585 192.045 ;
        RECT 55.745 192.000 56.035 192.045 ;
        RECT 31.325 191.860 35.325 192.000 ;
        RECT 31.325 191.815 31.615 191.860 ;
        RECT 32.515 191.815 32.805 191.860 ;
        RECT 35.035 191.815 35.325 191.860 ;
        RECT 38.340 191.860 41.700 192.000 ;
        RECT 31.780 191.320 32.070 191.365 ;
        RECT 33.190 191.320 33.510 191.380 ;
        RECT 31.780 191.180 33.510 191.320 ;
        RECT 31.780 191.135 32.070 191.180 ;
        RECT 33.190 191.120 33.510 191.180 ;
        RECT 38.340 191.040 38.480 191.860 ;
        RECT 40.550 191.460 40.870 191.720 ;
        RECT 41.560 191.705 41.700 191.860 ;
        RECT 45.585 191.860 49.585 192.000 ;
        RECT 45.585 191.815 45.875 191.860 ;
        RECT 46.775 191.815 47.065 191.860 ;
        RECT 49.295 191.815 49.585 191.860 ;
        RECT 53.980 191.860 56.035 192.000 ;
        RECT 41.485 191.475 41.775 191.705 ;
        RECT 42.390 191.660 42.710 191.720 ;
        RECT 44.705 191.660 44.995 191.705 ;
        RECT 48.830 191.660 49.150 191.720 ;
        RECT 42.390 191.520 49.150 191.660 ;
        RECT 42.390 191.460 42.710 191.520 ;
        RECT 44.705 191.475 44.995 191.520 ;
        RECT 48.830 191.460 49.150 191.520 ;
        RECT 52.970 191.460 53.290 191.720 ;
        RECT 53.980 191.705 54.120 191.860 ;
        RECT 55.745 191.815 56.035 191.860 ;
        RECT 64.955 192.000 65.245 192.045 ;
        RECT 67.475 192.000 67.765 192.045 ;
        RECT 68.665 192.000 68.955 192.045 ;
        RECT 64.955 191.860 68.955 192.000 ;
        RECT 64.955 191.815 65.245 191.860 ;
        RECT 67.475 191.815 67.765 191.860 ;
        RECT 68.665 191.815 68.955 191.860 ;
        RECT 69.530 191.800 69.850 192.060 ;
        RECT 53.905 191.475 54.195 191.705 ;
        RECT 55.270 191.460 55.590 191.720 ;
        RECT 56.205 191.660 56.495 191.705 ;
        RECT 57.570 191.660 57.890 191.720 ;
        RECT 58.045 191.660 58.335 191.705 ;
        RECT 56.205 191.520 58.335 191.660 ;
        RECT 56.205 191.475 56.495 191.520 ;
        RECT 57.570 191.460 57.890 191.520 ;
        RECT 58.045 191.475 58.335 191.520 ;
        RECT 58.965 191.660 59.255 191.705 ;
        RECT 60.790 191.660 61.110 191.720 ;
        RECT 58.965 191.520 61.110 191.660 ;
        RECT 58.965 191.475 59.255 191.520 ;
        RECT 60.790 191.460 61.110 191.520 ;
        RECT 40.105 191.135 40.395 191.365 ;
        RECT 41.010 191.320 41.330 191.380 ;
        RECT 41.945 191.320 42.235 191.365 ;
        RECT 45.930 191.320 46.220 191.365 ;
        RECT 41.010 191.180 42.235 191.320 ;
        RECT 37.345 190.980 37.635 191.025 ;
        RECT 37.790 190.980 38.110 191.040 ;
        RECT 37.345 190.840 38.110 190.980 ;
        RECT 37.345 190.795 37.635 190.840 ;
        RECT 37.790 190.780 38.110 190.840 ;
        RECT 38.250 190.780 38.570 191.040 ;
        RECT 39.170 191.025 39.490 191.040 ;
        RECT 39.105 190.795 39.490 191.025 ;
        RECT 40.180 190.980 40.320 191.135 ;
        RECT 41.010 191.120 41.330 191.180 ;
        RECT 41.945 191.135 42.235 191.180 ;
        RECT 43.860 191.180 46.220 191.320 ;
        RECT 41.470 190.980 41.790 191.040 ;
        RECT 40.180 190.840 41.790 190.980 ;
        RECT 39.170 190.780 39.490 190.795 ;
        RECT 41.470 190.780 41.790 190.840 ;
        RECT 42.850 191.025 43.170 191.040 ;
        RECT 43.860 191.025 44.000 191.180 ;
        RECT 45.930 191.135 46.220 191.180 ;
        RECT 59.410 191.120 59.730 191.380 ;
        RECT 65.390 191.320 65.710 191.380 ;
        RECT 68.210 191.320 68.500 191.365 ;
        RECT 65.390 191.180 68.500 191.320 ;
        RECT 65.390 191.120 65.710 191.180 ;
        RECT 68.210 191.135 68.500 191.180 ;
        RECT 42.850 190.795 43.235 191.025 ;
        RECT 43.785 190.795 44.075 191.025 ;
        RECT 42.850 190.780 43.170 190.795 ;
        RECT 51.590 190.780 51.910 191.040 ;
        RECT 58.505 190.980 58.795 191.025 ;
        RECT 60.425 190.980 60.715 191.025 ;
        RECT 58.505 190.840 60.715 190.980 ;
        RECT 58.505 190.795 58.795 190.840 ;
        RECT 60.425 190.795 60.715 190.840 ;
        RECT 61.710 190.980 62.030 191.040 ;
        RECT 62.645 190.980 62.935 191.025 ;
        RECT 61.710 190.840 62.935 190.980 ;
        RECT 61.710 190.780 62.030 190.840 ;
        RECT 62.645 190.795 62.935 190.840 ;
        RECT 5.520 190.160 84.180 190.640 ;
        RECT 33.190 189.760 33.510 190.020 ;
        RECT 34.045 189.960 34.335 190.005 ;
        RECT 35.490 189.960 35.810 190.020 ;
        RECT 34.045 189.820 35.810 189.960 ;
        RECT 34.045 189.775 34.335 189.820 ;
        RECT 35.490 189.760 35.810 189.820 ;
        RECT 35.950 189.760 36.270 190.020 ;
        RECT 38.250 189.760 38.570 190.020 ;
        RECT 40.550 190.005 40.870 190.020 ;
        RECT 40.550 189.960 40.885 190.005 ;
        RECT 40.385 189.820 40.885 189.960 ;
        RECT 40.550 189.775 40.885 189.820 ;
        RECT 41.025 189.960 41.315 190.005 ;
        RECT 43.770 189.960 44.090 190.020 ;
        RECT 49.750 189.960 50.070 190.020 ;
        RECT 51.590 189.960 51.910 190.020 ;
        RECT 41.025 189.820 51.910 189.960 ;
        RECT 41.025 189.775 41.315 189.820 ;
        RECT 40.550 189.760 40.870 189.775 ;
        RECT 43.770 189.760 44.090 189.820 ;
        RECT 49.750 189.760 50.070 189.820 ;
        RECT 51.590 189.760 51.910 189.820 ;
        RECT 52.970 189.960 53.290 190.020 ;
        RECT 60.345 189.960 60.635 190.005 ;
        RECT 52.970 189.820 60.635 189.960 ;
        RECT 52.970 189.760 53.290 189.820 ;
        RECT 60.345 189.775 60.635 189.820 ;
        RECT 61.250 189.960 61.570 190.020 ;
        RECT 63.565 189.960 63.855 190.005 ;
        RECT 61.250 189.820 63.855 189.960 ;
        RECT 61.250 189.760 61.570 189.820 ;
        RECT 63.565 189.775 63.855 189.820 ;
        RECT 65.390 189.760 65.710 190.020 ;
        RECT 35.030 189.420 35.350 189.680 ;
        RECT 38.340 189.620 38.480 189.760 ;
        RECT 35.580 189.480 38.480 189.620 ;
        RECT 38.725 189.620 39.015 189.665 ;
        RECT 39.170 189.620 39.490 189.680 ;
        RECT 38.725 189.480 41.700 189.620 ;
        RECT 35.580 189.325 35.720 189.480 ;
        RECT 38.725 189.435 39.015 189.480 ;
        RECT 39.170 189.420 39.490 189.480 ;
        RECT 35.505 189.095 35.795 189.325 ;
        RECT 36.425 189.280 36.715 189.325 ;
        RECT 37.790 189.280 38.110 189.340 ;
        RECT 36.425 189.140 38.110 189.280 ;
        RECT 36.425 189.095 36.715 189.140 ;
        RECT 37.790 189.080 38.110 189.140 ;
        RECT 38.250 189.080 38.570 189.340 ;
        RECT 41.560 189.325 41.700 189.480 ;
        RECT 43.770 189.325 44.090 189.340 ;
        RECT 40.105 189.280 40.395 189.325 ;
        RECT 41.485 189.280 41.775 189.325 ;
        RECT 43.770 189.280 44.110 189.325 ;
        RECT 40.105 189.140 40.780 189.280 ;
        RECT 40.105 189.095 40.395 189.140 ;
        RECT 36.885 188.600 37.175 188.645 ;
        RECT 40.640 188.600 40.780 189.140 ;
        RECT 41.485 189.140 43.495 189.280 ;
        RECT 41.485 189.095 41.775 189.140 ;
        RECT 41.945 188.940 42.235 188.985 ;
        RECT 42.850 188.940 43.170 189.000 ;
        RECT 41.945 188.800 43.170 188.940 ;
        RECT 43.355 188.940 43.495 189.140 ;
        RECT 43.770 189.140 44.285 189.280 ;
        RECT 43.770 189.095 44.110 189.140 ;
        RECT 43.770 189.080 44.090 189.095 ;
        RECT 44.245 188.940 44.535 188.985 ;
        RECT 53.060 188.940 53.200 189.760 ;
        RECT 56.205 189.620 56.495 189.665 ;
        RECT 63.090 189.620 63.410 189.680 ;
        RECT 56.205 189.480 63.410 189.620 ;
        RECT 56.205 189.435 56.495 189.480 ;
        RECT 63.090 189.420 63.410 189.480 ;
        RECT 64.485 189.620 64.775 189.665 ;
        RECT 67.705 189.620 67.995 189.665 ;
        RECT 64.485 189.480 67.995 189.620 ;
        RECT 64.485 189.435 64.775 189.480 ;
        RECT 67.705 189.435 67.995 189.480 ;
        RECT 55.270 189.280 55.590 189.340 ;
        RECT 57.585 189.280 57.875 189.325 ;
        RECT 58.505 189.280 58.795 189.325 ;
        RECT 55.270 189.140 57.875 189.280 ;
        RECT 55.270 189.080 55.590 189.140 ;
        RECT 57.585 189.095 57.875 189.140 ;
        RECT 58.120 189.140 58.795 189.280 ;
        RECT 43.355 188.800 53.200 188.940 ;
        RECT 56.190 188.940 56.510 189.000 ;
        RECT 58.120 188.940 58.260 189.140 ;
        RECT 58.505 189.095 58.795 189.140 ;
        RECT 58.965 189.095 59.255 189.325 ;
        RECT 59.425 189.095 59.715 189.325 ;
        RECT 60.330 189.280 60.650 189.340 ;
        RECT 60.805 189.280 61.095 189.325 ;
        RECT 60.330 189.140 61.095 189.280 ;
        RECT 59.040 188.940 59.180 189.095 ;
        RECT 56.190 188.800 58.260 188.940 ;
        RECT 58.580 188.800 59.180 188.940 ;
        RECT 59.500 188.940 59.640 189.095 ;
        RECT 60.330 189.080 60.650 189.140 ;
        RECT 60.805 189.095 61.095 189.140 ;
        RECT 61.710 189.080 62.030 189.340 ;
        RECT 62.185 189.280 62.475 189.325 ;
        RECT 62.185 189.140 62.860 189.280 ;
        RECT 62.185 189.095 62.475 189.140 ;
        RECT 62.720 188.940 62.860 189.140 ;
        RECT 64.010 189.080 64.330 189.340 ;
        RECT 65.865 189.095 66.155 189.325 ;
        RECT 63.090 188.940 63.410 189.000 ;
        RECT 65.940 188.940 66.080 189.095 ;
        RECT 66.770 189.080 67.090 189.340 ;
        RECT 59.500 188.800 66.080 188.940 ;
        RECT 41.945 188.755 42.235 188.800 ;
        RECT 42.850 188.740 43.170 188.800 ;
        RECT 44.245 188.755 44.535 188.800 ;
        RECT 56.190 188.740 56.510 188.800 ;
        RECT 58.580 188.660 58.720 188.800 ;
        RECT 63.090 188.740 63.410 188.800 ;
        RECT 41.470 188.600 41.790 188.660 ;
        RECT 36.885 188.460 41.790 188.600 ;
        RECT 36.885 188.415 37.175 188.460 ;
        RECT 41.470 188.400 41.790 188.460 ;
        RECT 58.490 188.400 58.810 188.660 ;
        RECT 60.790 188.400 61.110 188.660 ;
        RECT 62.645 188.600 62.935 188.645 ;
        RECT 62.030 188.460 62.935 188.600 ;
        RECT 34.110 188.060 34.430 188.320 ;
        RECT 34.570 188.260 34.890 188.320 ;
        RECT 39.645 188.260 39.935 188.305 ;
        RECT 34.570 188.120 39.935 188.260 ;
        RECT 34.570 188.060 34.890 188.120 ;
        RECT 39.645 188.075 39.935 188.120 ;
        RECT 54.350 188.260 54.670 188.320 ;
        RECT 54.825 188.260 55.115 188.305 ;
        RECT 54.350 188.120 55.115 188.260 ;
        RECT 54.350 188.060 54.670 188.120 ;
        RECT 54.825 188.075 55.115 188.120 ;
        RECT 55.730 188.260 56.050 188.320 ;
        RECT 59.410 188.260 59.730 188.320 ;
        RECT 62.030 188.260 62.170 188.460 ;
        RECT 62.645 188.415 62.935 188.460 ;
        RECT 55.730 188.120 62.170 188.260 ;
        RECT 55.730 188.060 56.050 188.120 ;
        RECT 59.410 188.060 59.730 188.120 ;
        RECT 5.520 187.440 84.180 187.920 ;
        RECT 34.110 187.240 34.430 187.300 ;
        RECT 34.585 187.240 34.875 187.285 ;
        RECT 43.310 187.240 43.630 187.300 ;
        RECT 34.110 187.100 43.630 187.240 ;
        RECT 34.110 187.040 34.430 187.100 ;
        RECT 34.585 187.055 34.875 187.100 ;
        RECT 43.310 187.040 43.630 187.100 ;
        RECT 57.570 187.040 57.890 187.300 ;
        RECT 58.490 187.040 58.810 187.300 ;
        RECT 63.565 187.240 63.855 187.285 ;
        RECT 64.010 187.240 64.330 187.300 ;
        RECT 63.565 187.100 64.330 187.240 ;
        RECT 63.565 187.055 63.855 187.100 ;
        RECT 64.010 187.040 64.330 187.100 ;
        RECT 50.685 186.900 50.975 186.945 ;
        RECT 52.970 186.900 53.290 186.960 ;
        RECT 50.685 186.760 53.290 186.900 ;
        RECT 50.685 186.715 50.975 186.760 ;
        RECT 52.970 186.700 53.290 186.760 ;
        RECT 54.350 186.900 54.670 186.960 ;
        RECT 54.350 186.760 56.880 186.900 ;
        RECT 54.350 186.700 54.670 186.760 ;
        RECT 56.740 186.605 56.880 186.760 ;
        RECT 53.445 186.560 53.735 186.605 ;
        RECT 49.840 186.420 52.740 186.560 ;
        RECT 49.840 186.280 49.980 186.420 ;
        RECT 35.030 186.020 35.350 186.280 ;
        RECT 49.290 186.020 49.610 186.280 ;
        RECT 49.750 186.020 50.070 186.280 ;
        RECT 52.600 186.265 52.740 186.420 ;
        RECT 53.445 186.420 55.500 186.560 ;
        RECT 53.445 186.375 53.735 186.420 ;
        RECT 55.360 186.280 55.500 186.420 ;
        RECT 56.665 186.375 56.955 186.605 ;
        RECT 58.490 186.560 58.810 186.620 ;
        RECT 61.710 186.560 62.030 186.620 ;
        RECT 58.490 186.420 64.240 186.560 ;
        RECT 58.490 186.360 58.810 186.420 ;
        RECT 61.710 186.360 62.030 186.420 ;
        RECT 52.065 186.220 52.355 186.265 ;
        RECT 50.300 186.080 52.355 186.220 ;
        RECT 35.120 185.880 35.260 186.020 ;
        RECT 35.505 185.880 35.795 185.925 ;
        RECT 35.120 185.740 35.795 185.880 ;
        RECT 49.380 185.880 49.520 186.020 ;
        RECT 50.300 185.880 50.440 186.080 ;
        RECT 52.065 186.035 52.355 186.080 ;
        RECT 52.525 186.035 52.815 186.265 ;
        RECT 53.890 186.020 54.210 186.280 ;
        RECT 55.270 186.020 55.590 186.280 ;
        RECT 56.190 186.020 56.510 186.280 ;
        RECT 63.090 186.220 63.410 186.280 ;
        RECT 64.100 186.265 64.240 186.420 ;
        RECT 59.040 186.080 63.410 186.220 ;
        RECT 49.380 185.740 50.440 185.880 ;
        RECT 50.685 185.880 50.975 185.925 ;
        RECT 54.365 185.880 54.655 185.925 ;
        RECT 50.685 185.740 54.655 185.880 ;
        RECT 35.505 185.695 35.795 185.740 ;
        RECT 50.685 185.695 50.975 185.740 ;
        RECT 54.365 185.695 54.655 185.740 ;
        RECT 58.425 185.880 58.715 185.925 ;
        RECT 59.040 185.880 59.180 186.080 ;
        RECT 63.090 186.020 63.410 186.080 ;
        RECT 64.025 186.220 64.315 186.265 ;
        RECT 66.770 186.220 67.090 186.280 ;
        RECT 64.025 186.080 67.090 186.220 ;
        RECT 64.025 186.035 64.315 186.080 ;
        RECT 66.770 186.020 67.090 186.080 ;
        RECT 58.425 185.740 59.180 185.880 ;
        RECT 59.425 185.880 59.715 185.925 ;
        RECT 60.330 185.880 60.650 185.940 ;
        RECT 59.425 185.740 60.650 185.880 ;
        RECT 63.180 185.880 63.320 186.020 ;
        RECT 64.930 185.880 65.250 185.940 ;
        RECT 63.180 185.740 65.250 185.880 ;
        RECT 58.425 185.695 58.715 185.740 ;
        RECT 59.425 185.695 59.715 185.740 ;
        RECT 33.650 185.340 33.970 185.600 ;
        RECT 34.505 185.540 34.795 185.585 ;
        RECT 35.030 185.540 35.350 185.600 ;
        RECT 34.505 185.400 35.350 185.540 ;
        RECT 34.505 185.355 34.795 185.400 ;
        RECT 35.030 185.340 35.350 185.400 ;
        RECT 50.210 185.540 50.530 185.600 ;
        RECT 51.145 185.540 51.435 185.585 ;
        RECT 50.210 185.400 51.435 185.540 ;
        RECT 50.210 185.340 50.530 185.400 ;
        RECT 51.145 185.355 51.435 185.400 ;
        RECT 56.190 185.540 56.510 185.600 ;
        RECT 59.500 185.540 59.640 185.695 ;
        RECT 60.330 185.680 60.650 185.740 ;
        RECT 64.930 185.680 65.250 185.740 ;
        RECT 56.190 185.400 59.640 185.540 ;
        RECT 56.190 185.340 56.510 185.400 ;
        RECT 5.520 184.720 84.180 185.200 ;
        RECT 49.305 184.520 49.595 184.565 ;
        RECT 49.750 184.520 50.070 184.580 ;
        RECT 49.305 184.380 50.070 184.520 ;
        RECT 49.305 184.335 49.595 184.380 ;
        RECT 49.750 184.320 50.070 184.380 ;
        RECT 14.790 184.225 15.110 184.240 ;
        RECT 14.725 183.995 15.110 184.225 ;
        RECT 15.725 183.995 16.015 184.225 ;
        RECT 33.160 184.180 33.450 184.225 ;
        RECT 33.650 184.180 33.970 184.240 ;
        RECT 33.160 184.040 33.970 184.180 ;
        RECT 33.160 183.995 33.450 184.040 ;
        RECT 14.790 183.980 15.110 183.995 ;
        RECT 10.190 183.500 10.510 183.560 ;
        RECT 15.800 183.500 15.940 183.995 ;
        RECT 33.650 183.980 33.970 184.040 ;
        RECT 45.150 184.180 45.470 184.240 ;
        RECT 55.730 184.180 56.050 184.240 ;
        RECT 45.150 184.040 56.050 184.180 ;
        RECT 45.150 183.980 45.470 184.040 ;
        RECT 55.730 183.980 56.050 184.040 ;
        RECT 20.310 183.840 20.630 183.900 ;
        RECT 21.145 183.840 21.435 183.885 ;
        RECT 20.310 183.700 21.435 183.840 ;
        RECT 20.310 183.640 20.630 183.700 ;
        RECT 21.145 183.655 21.435 183.700 ;
        RECT 30.430 183.840 30.750 183.900 ;
        RECT 31.825 183.840 32.115 183.885 ;
        RECT 30.430 183.700 32.115 183.840 ;
        RECT 30.430 183.640 30.750 183.700 ;
        RECT 31.825 183.655 32.115 183.700 ;
        RECT 48.845 183.655 49.135 183.885 ;
        RECT 10.190 183.360 15.940 183.500 ;
        RECT 18.010 183.500 18.330 183.560 ;
        RECT 19.865 183.500 20.155 183.545 ;
        RECT 18.010 183.360 20.155 183.500 ;
        RECT 10.190 183.300 10.510 183.360 ;
        RECT 18.010 183.300 18.330 183.360 ;
        RECT 19.865 183.315 20.155 183.360 ;
        RECT 20.745 183.500 21.035 183.545 ;
        RECT 21.935 183.500 22.225 183.545 ;
        RECT 24.455 183.500 24.745 183.545 ;
        RECT 20.745 183.360 24.745 183.500 ;
        RECT 20.745 183.315 21.035 183.360 ;
        RECT 21.935 183.315 22.225 183.360 ;
        RECT 24.455 183.315 24.745 183.360 ;
        RECT 32.705 183.500 32.995 183.545 ;
        RECT 33.895 183.500 34.185 183.545 ;
        RECT 36.415 183.500 36.705 183.545 ;
        RECT 32.705 183.360 36.705 183.500 ;
        RECT 48.920 183.500 49.060 183.655 ;
        RECT 50.210 183.640 50.530 183.900 ;
        RECT 52.050 183.840 52.370 183.900 ;
        RECT 52.985 183.840 53.275 183.885 ;
        RECT 52.050 183.700 53.275 183.840 ;
        RECT 52.050 183.640 52.370 183.700 ;
        RECT 52.985 183.655 53.275 183.700 ;
        RECT 53.445 183.840 53.735 183.885 ;
        RECT 56.190 183.840 56.510 183.900 ;
        RECT 53.445 183.700 56.510 183.840 ;
        RECT 53.445 183.655 53.735 183.700 ;
        RECT 56.190 183.640 56.510 183.700 ;
        RECT 49.290 183.500 49.610 183.560 ;
        RECT 51.130 183.500 51.450 183.560 ;
        RECT 48.920 183.360 51.450 183.500 ;
        RECT 32.705 183.315 32.995 183.360 ;
        RECT 33.895 183.315 34.185 183.360 ;
        RECT 36.415 183.315 36.705 183.360 ;
        RECT 49.290 183.300 49.610 183.360 ;
        RECT 51.130 183.300 51.450 183.360 ;
        RECT 54.365 183.500 54.655 183.545 ;
        RECT 58.490 183.500 58.810 183.560 ;
        RECT 54.365 183.360 58.810 183.500 ;
        RECT 54.365 183.315 54.655 183.360 ;
        RECT 58.490 183.300 58.810 183.360 ;
        RECT 20.350 183.160 20.640 183.205 ;
        RECT 22.450 183.160 22.740 183.205 ;
        RECT 24.020 183.160 24.310 183.205 ;
        RECT 20.350 183.020 24.310 183.160 ;
        RECT 20.350 182.975 20.640 183.020 ;
        RECT 22.450 182.975 22.740 183.020 ;
        RECT 24.020 182.975 24.310 183.020 ;
        RECT 32.310 183.160 32.600 183.205 ;
        RECT 34.410 183.160 34.700 183.205 ;
        RECT 35.980 183.160 36.270 183.205 ;
        RECT 32.310 183.020 36.270 183.160 ;
        RECT 32.310 182.975 32.600 183.020 ;
        RECT 34.410 182.975 34.700 183.020 ;
        RECT 35.980 182.975 36.270 183.020 ;
        RECT 39.630 183.160 39.950 183.220 ;
        RECT 41.010 183.160 41.330 183.220 ;
        RECT 60.790 183.160 61.110 183.220 ;
        RECT 39.630 183.020 61.110 183.160 ;
        RECT 39.630 182.960 39.950 183.020 ;
        RECT 41.010 182.960 41.330 183.020 ;
        RECT 60.790 182.960 61.110 183.020 ;
        RECT 13.870 182.620 14.190 182.880 ;
        RECT 14.805 182.820 15.095 182.865 ;
        RECT 19.850 182.820 20.170 182.880 ;
        RECT 14.805 182.680 20.170 182.820 ;
        RECT 14.805 182.635 15.095 182.680 ;
        RECT 19.850 182.620 20.170 182.680 ;
        RECT 26.750 182.620 27.070 182.880 ;
        RECT 36.410 182.820 36.730 182.880 ;
        RECT 38.725 182.820 39.015 182.865 ;
        RECT 36.410 182.680 39.015 182.820 ;
        RECT 36.410 182.620 36.730 182.680 ;
        RECT 38.725 182.635 39.015 182.680 ;
        RECT 50.225 182.820 50.515 182.865 ;
        RECT 52.510 182.820 52.830 182.880 ;
        RECT 50.225 182.680 52.830 182.820 ;
        RECT 50.225 182.635 50.515 182.680 ;
        RECT 52.510 182.620 52.830 182.680 ;
        RECT 53.890 182.620 54.210 182.880 ;
        RECT 5.520 182.000 84.180 182.480 ;
        RECT 10.190 181.600 10.510 181.860 ;
        RECT 19.865 181.800 20.155 181.845 ;
        RECT 20.310 181.800 20.630 181.860 ;
        RECT 19.865 181.660 20.630 181.800 ;
        RECT 19.865 181.615 20.155 181.660 ;
        RECT 20.310 181.600 20.630 181.660 ;
        RECT 20.770 181.600 21.090 181.860 ;
        RECT 30.445 181.800 30.735 181.845 ;
        RECT 21.320 181.660 30.735 181.800 ;
        RECT 13.870 181.460 14.160 181.505 ;
        RECT 15.440 181.460 15.730 181.505 ;
        RECT 17.540 181.460 17.830 181.505 ;
        RECT 13.870 181.320 17.830 181.460 ;
        RECT 13.870 181.275 14.160 181.320 ;
        RECT 15.440 181.275 15.730 181.320 ;
        RECT 17.540 181.275 17.830 181.320 ;
        RECT 13.435 181.120 13.725 181.165 ;
        RECT 15.955 181.120 16.245 181.165 ;
        RECT 17.145 181.120 17.435 181.165 ;
        RECT 13.435 180.980 17.435 181.120 ;
        RECT 13.435 180.935 13.725 180.980 ;
        RECT 15.955 180.935 16.245 180.980 ;
        RECT 17.145 180.935 17.435 180.980 ;
        RECT 9.745 180.595 10.035 180.825 ;
        RECT 9.820 180.440 9.960 180.595 ;
        RECT 10.650 180.580 10.970 180.840 ;
        RECT 13.870 180.780 14.190 180.840 ;
        RECT 16.690 180.780 16.980 180.825 ;
        RECT 13.870 180.640 16.980 180.780 ;
        RECT 13.870 180.580 14.190 180.640 ;
        RECT 16.690 180.595 16.980 180.640 ;
        RECT 18.010 180.580 18.330 180.840 ;
        RECT 20.705 180.440 20.995 180.485 ;
        RECT 21.320 180.440 21.460 181.660 ;
        RECT 30.445 181.615 30.735 181.660 ;
        RECT 35.030 181.600 35.350 181.860 ;
        RECT 50.210 181.800 50.530 181.860 ;
        RECT 57.110 181.800 57.430 181.860 ;
        RECT 50.210 181.660 57.430 181.800 ;
        RECT 50.210 181.600 50.530 181.660 ;
        RECT 23.160 181.320 28.820 181.460 ;
        RECT 22.610 180.780 22.930 180.840 ;
        RECT 23.160 180.825 23.300 181.320 ;
        RECT 23.530 181.120 23.850 181.180 ;
        RECT 23.530 180.980 26.520 181.120 ;
        RECT 23.530 180.920 23.850 180.980 ;
        RECT 23.085 180.780 23.375 180.825 ;
        RECT 22.610 180.640 23.375 180.780 ;
        RECT 22.610 180.580 22.930 180.640 ;
        RECT 23.085 180.595 23.375 180.640 ;
        RECT 23.990 180.580 24.310 180.840 ;
        RECT 24.450 180.580 24.770 180.840 ;
        RECT 26.380 180.825 26.520 180.980 ;
        RECT 26.305 180.780 26.595 180.825 ;
        RECT 26.750 180.780 27.070 180.840 ;
        RECT 26.305 180.640 27.070 180.780 ;
        RECT 27.300 180.790 27.440 181.320 ;
        RECT 28.680 181.120 28.820 181.320 ;
        RECT 33.665 181.120 33.955 181.165 ;
        RECT 34.570 181.120 34.890 181.180 ;
        RECT 28.680 180.980 32.040 181.120 ;
        RECT 27.685 180.790 27.975 180.825 ;
        RECT 27.300 180.650 27.975 180.790 ;
        RECT 26.305 180.595 26.595 180.640 ;
        RECT 26.750 180.580 27.070 180.640 ;
        RECT 27.685 180.595 27.975 180.650 ;
        RECT 28.130 180.580 28.450 180.840 ;
        RECT 28.680 180.780 28.820 180.980 ;
        RECT 29.065 180.780 29.355 180.825 ;
        RECT 28.680 180.640 29.355 180.780 ;
        RECT 29.065 180.595 29.355 180.640 ;
        RECT 29.510 180.580 29.830 180.840 ;
        RECT 31.900 180.825 32.040 180.980 ;
        RECT 33.665 180.980 34.890 181.120 ;
        RECT 33.665 180.935 33.955 180.980 ;
        RECT 34.570 180.920 34.890 180.980 ;
        RECT 30.445 180.780 30.735 180.825 ;
        RECT 30.445 180.640 31.580 180.780 ;
        RECT 30.445 180.595 30.735 180.640 ;
        RECT 9.820 180.300 11.340 180.440 ;
        RECT 11.200 180.145 11.340 180.300 ;
        RECT 20.705 180.300 21.460 180.440 ;
        RECT 21.705 180.440 21.995 180.485 ;
        RECT 25.385 180.440 25.675 180.485 ;
        RECT 25.830 180.440 26.150 180.500 ;
        RECT 21.705 180.300 26.150 180.440 ;
        RECT 26.840 180.440 26.980 180.580 ;
        RECT 30.905 180.440 31.195 180.485 ;
        RECT 26.840 180.300 31.195 180.440 ;
        RECT 20.705 180.255 20.995 180.300 ;
        RECT 21.705 180.255 21.995 180.300 ;
        RECT 25.385 180.255 25.675 180.300 ;
        RECT 25.830 180.240 26.150 180.300 ;
        RECT 30.905 180.255 31.195 180.300 ;
        RECT 11.125 180.100 11.415 180.145 ;
        RECT 16.170 180.100 16.490 180.160 ;
        RECT 11.125 179.960 16.490 180.100 ;
        RECT 11.125 179.915 11.415 179.960 ;
        RECT 16.170 179.900 16.490 179.960 ;
        RECT 22.165 180.100 22.455 180.145 ;
        RECT 23.070 180.100 23.390 180.160 ;
        RECT 22.165 179.960 23.390 180.100 ;
        RECT 22.165 179.915 22.455 179.960 ;
        RECT 23.070 179.900 23.390 179.960 ;
        RECT 24.910 180.100 25.230 180.160 ;
        RECT 26.750 180.100 27.070 180.160 ;
        RECT 27.225 180.100 27.515 180.145 ;
        RECT 31.440 180.100 31.580 180.640 ;
        RECT 31.825 180.595 32.115 180.825 ;
        RECT 33.205 180.780 33.495 180.825 ;
        RECT 35.950 180.780 36.270 180.840 ;
        RECT 33.205 180.640 36.270 180.780 ;
        RECT 33.205 180.595 33.495 180.640 ;
        RECT 35.950 180.580 36.270 180.640 ;
        RECT 45.610 180.580 45.930 180.840 ;
        RECT 47.005 180.780 47.295 180.825 ;
        RECT 49.750 180.780 50.070 180.840 ;
        RECT 51.680 180.825 51.820 181.660 ;
        RECT 57.110 181.600 57.430 181.660 ;
        RECT 60.790 181.800 61.110 181.860 ;
        RECT 61.265 181.800 61.555 181.845 ;
        RECT 60.790 181.660 61.555 181.800 ;
        RECT 60.790 181.600 61.110 181.660 ;
        RECT 61.265 181.615 61.555 181.660 ;
        RECT 52.985 181.460 53.275 181.505 ;
        RECT 53.890 181.460 54.210 181.520 ;
        RECT 52.985 181.320 54.210 181.460 ;
        RECT 52.985 181.275 53.275 181.320 ;
        RECT 53.890 181.260 54.210 181.320 ;
        RECT 60.330 181.460 60.650 181.520 ;
        RECT 62.645 181.460 62.935 181.505 ;
        RECT 60.330 181.320 62.935 181.460 ;
        RECT 60.330 181.260 60.650 181.320 ;
        RECT 62.645 181.275 62.935 181.320 ;
        RECT 65.390 181.460 65.680 181.505 ;
        RECT 66.960 181.460 67.250 181.505 ;
        RECT 69.060 181.460 69.350 181.505 ;
        RECT 65.390 181.320 69.350 181.460 ;
        RECT 65.390 181.275 65.680 181.320 ;
        RECT 66.960 181.275 67.250 181.320 ;
        RECT 69.060 181.275 69.350 181.320 ;
        RECT 54.900 180.980 56.880 181.120 ;
        RECT 47.005 180.640 50.070 180.780 ;
        RECT 47.005 180.595 47.295 180.640 ;
        RECT 49.750 180.580 50.070 180.640 ;
        RECT 51.605 180.595 51.895 180.825 ;
        RECT 52.525 180.780 52.815 180.825 ;
        RECT 52.970 180.780 53.290 180.840 ;
        RECT 52.525 180.640 53.290 180.780 ;
        RECT 52.525 180.595 52.815 180.640 ;
        RECT 52.970 180.580 53.290 180.640 ;
        RECT 53.445 180.595 53.735 180.825 ;
        RECT 53.905 180.790 54.195 180.825 ;
        RECT 54.900 180.790 55.040 180.980 ;
        RECT 53.905 180.650 55.040 180.790 ;
        RECT 55.730 180.780 56.050 180.840 ;
        RECT 56.205 180.780 56.495 180.825 ;
        RECT 53.905 180.595 54.195 180.650 ;
        RECT 55.730 180.640 56.495 180.780 ;
        RECT 56.740 180.780 56.880 180.980 ;
        RECT 57.110 180.920 57.430 181.180 ;
        RECT 64.955 181.120 65.245 181.165 ;
        RECT 67.475 181.120 67.765 181.165 ;
        RECT 68.665 181.120 68.955 181.165 ;
        RECT 64.955 180.980 68.955 181.120 ;
        RECT 64.955 180.935 65.245 180.980 ;
        RECT 67.475 180.935 67.765 180.980 ;
        RECT 68.665 180.935 68.955 180.980 ;
        RECT 69.530 180.920 69.850 181.180 ;
        RECT 56.740 180.640 57.340 180.780 ;
        RECT 35.490 180.440 35.810 180.500 ;
        RECT 40.105 180.440 40.395 180.485 ;
        RECT 35.490 180.300 40.395 180.440 ;
        RECT 35.490 180.240 35.810 180.300 ;
        RECT 40.105 180.255 40.395 180.300 ;
        RECT 42.850 180.440 43.170 180.500 ;
        RECT 46.545 180.440 46.835 180.485 ;
        RECT 42.850 180.300 46.835 180.440 ;
        RECT 53.520 180.440 53.660 180.595 ;
        RECT 55.730 180.580 56.050 180.640 ;
        RECT 56.205 180.595 56.495 180.640 ;
        RECT 56.650 180.440 56.970 180.500 ;
        RECT 53.520 180.300 56.970 180.440 ;
        RECT 57.200 180.440 57.340 180.640 ;
        RECT 57.570 180.580 57.890 180.840 ;
        RECT 59.425 180.780 59.715 180.825 ;
        RECT 65.390 180.780 65.710 180.840 ;
        RECT 59.425 180.640 65.710 180.780 ;
        RECT 59.425 180.595 59.715 180.640 ;
        RECT 65.390 180.580 65.710 180.640 ;
        RECT 58.045 180.440 58.335 180.485 ;
        RECT 57.200 180.300 58.335 180.440 ;
        RECT 42.850 180.240 43.170 180.300 ;
        RECT 46.545 180.255 46.835 180.300 ;
        RECT 56.650 180.240 56.970 180.300 ;
        RECT 58.045 180.255 58.335 180.300 ;
        RECT 64.010 180.440 64.330 180.500 ;
        RECT 68.210 180.440 68.500 180.485 ;
        RECT 64.010 180.300 68.500 180.440 ;
        RECT 64.010 180.240 64.330 180.300 ;
        RECT 68.210 180.255 68.500 180.300 ;
        RECT 24.910 179.960 31.580 180.100 ;
        RECT 37.330 180.100 37.650 180.160 ;
        RECT 39.645 180.100 39.935 180.145 ;
        RECT 41.010 180.100 41.330 180.160 ;
        RECT 37.330 179.960 41.330 180.100 ;
        RECT 24.910 179.900 25.230 179.960 ;
        RECT 26.750 179.900 27.070 179.960 ;
        RECT 27.225 179.915 27.515 179.960 ;
        RECT 37.330 179.900 37.650 179.960 ;
        RECT 39.645 179.915 39.935 179.960 ;
        RECT 41.010 179.900 41.330 179.960 ;
        RECT 44.705 180.100 44.995 180.145 ;
        RECT 45.150 180.100 45.470 180.160 ;
        RECT 44.705 179.960 45.470 180.100 ;
        RECT 44.705 179.915 44.995 179.960 ;
        RECT 45.150 179.900 45.470 179.960 ;
        RECT 52.970 180.100 53.290 180.160 ;
        RECT 54.825 180.100 55.115 180.145 ;
        RECT 52.970 179.960 55.115 180.100 ;
        RECT 52.970 179.900 53.290 179.960 ;
        RECT 54.825 179.915 55.115 179.960 ;
        RECT 55.270 179.900 55.590 180.160 ;
        RECT 61.250 179.900 61.570 180.160 ;
        RECT 62.170 179.900 62.490 180.160 ;
        RECT 5.520 179.280 84.180 179.760 ;
        RECT 14.345 179.080 14.635 179.125 ;
        RECT 14.790 179.080 15.110 179.140 ;
        RECT 14.345 178.940 15.110 179.080 ;
        RECT 14.345 178.895 14.635 178.940 ;
        RECT 14.790 178.880 15.110 178.940 ;
        RECT 23.990 179.080 24.310 179.140 ;
        RECT 26.290 179.080 26.610 179.140 ;
        RECT 27.670 179.080 27.990 179.140 ;
        RECT 23.990 178.940 24.680 179.080 ;
        RECT 23.990 178.880 24.310 178.940 ;
        RECT 16.170 178.740 16.490 178.800 ;
        RECT 22.610 178.740 22.930 178.800 ;
        RECT 24.540 178.785 24.680 178.940 ;
        RECT 26.290 178.940 27.990 179.080 ;
        RECT 26.290 178.880 26.610 178.940 ;
        RECT 27.670 178.880 27.990 178.940 ;
        RECT 35.505 179.080 35.795 179.125 ;
        RECT 41.485 179.080 41.775 179.125 ;
        RECT 35.505 178.940 41.775 179.080 ;
        RECT 35.505 178.895 35.795 178.940 ;
        RECT 41.485 178.895 41.775 178.940 ;
        RECT 42.850 178.880 43.170 179.140 ;
        RECT 44.705 179.080 44.995 179.125 ;
        RECT 45.610 179.080 45.930 179.140 ;
        RECT 44.705 178.940 45.930 179.080 ;
        RECT 44.705 178.895 44.995 178.940 ;
        RECT 45.610 178.880 45.930 178.940 ;
        RECT 49.750 178.880 50.070 179.140 ;
        RECT 51.130 179.080 51.450 179.140 ;
        RECT 56.665 179.080 56.955 179.125 ;
        RECT 57.570 179.080 57.890 179.140 ;
        RECT 51.130 178.940 55.960 179.080 ;
        RECT 51.130 178.880 51.450 178.940 ;
        RECT 23.545 178.740 23.835 178.785 ;
        RECT 16.170 178.600 23.835 178.740 ;
        RECT 16.170 178.540 16.490 178.600 ;
        RECT 22.610 178.540 22.930 178.600 ;
        RECT 23.545 178.555 23.835 178.600 ;
        RECT 24.465 178.740 24.755 178.785 ;
        RECT 36.425 178.740 36.715 178.785 ;
        RECT 42.070 178.740 42.360 178.785 ;
        RECT 24.465 178.600 28.820 178.740 ;
        RECT 24.465 178.555 24.755 178.600 ;
        RECT 28.680 178.460 28.820 178.600 ;
        RECT 36.425 178.600 42.360 178.740 ;
        RECT 42.940 178.740 43.080 178.880 ;
        RECT 51.590 178.740 51.910 178.800 ;
        RECT 55.270 178.740 55.590 178.800 ;
        RECT 42.940 178.600 48.140 178.740 ;
        RECT 36.425 178.555 36.715 178.600 ;
        RECT 42.070 178.555 42.360 178.600 ;
        RECT 10.650 178.400 10.970 178.460 ;
        RECT 15.265 178.400 15.555 178.445 ;
        RECT 10.650 178.260 15.555 178.400 ;
        RECT 10.650 178.200 10.970 178.260 ;
        RECT 15.265 178.215 15.555 178.260 ;
        RECT 15.340 178.060 15.480 178.215 ;
        RECT 23.990 178.200 24.310 178.460 ;
        RECT 27.225 178.215 27.515 178.445 ;
        RECT 25.385 178.060 25.675 178.105 ;
        RECT 26.750 178.060 27.070 178.120 ;
        RECT 15.340 177.920 27.070 178.060 ;
        RECT 27.300 178.060 27.440 178.215 ;
        RECT 27.670 178.200 27.990 178.460 ;
        RECT 28.130 178.200 28.450 178.460 ;
        RECT 28.590 178.200 28.910 178.460 ;
        RECT 33.650 178.200 33.970 178.460 ;
        RECT 35.950 178.200 36.270 178.460 ;
        RECT 36.885 178.400 37.175 178.445 ;
        RECT 37.330 178.400 37.650 178.460 ;
        RECT 36.885 178.260 37.650 178.400 ;
        RECT 36.885 178.215 37.175 178.260 ;
        RECT 37.330 178.200 37.650 178.260 ;
        RECT 38.265 178.215 38.555 178.445 ;
        RECT 39.185 178.400 39.475 178.445 ;
        RECT 41.025 178.400 41.315 178.445 ;
        RECT 39.185 178.260 41.315 178.400 ;
        RECT 39.185 178.215 39.475 178.260 ;
        RECT 41.025 178.215 41.315 178.260 ;
        RECT 43.325 178.400 43.615 178.445 ;
        RECT 43.325 178.260 44.460 178.400 ;
        RECT 43.325 178.215 43.615 178.260 ;
        RECT 29.970 178.060 30.290 178.120 ;
        RECT 33.205 178.060 33.495 178.105 ;
        RECT 27.300 177.920 33.495 178.060 ;
        RECT 36.040 178.060 36.180 178.200 ;
        RECT 38.340 178.060 38.480 178.215 ;
        RECT 36.040 177.920 38.480 178.060 ;
        RECT 25.385 177.875 25.675 177.920 ;
        RECT 26.750 177.860 27.070 177.920 ;
        RECT 29.970 177.860 30.290 177.920 ;
        RECT 33.205 177.875 33.495 177.920 ;
        RECT 20.770 177.380 21.090 177.440 ;
        RECT 22.625 177.380 22.915 177.425 ;
        RECT 23.530 177.380 23.850 177.440 ;
        RECT 20.770 177.240 23.850 177.380 ;
        RECT 20.770 177.180 21.090 177.240 ;
        RECT 22.625 177.195 22.915 177.240 ;
        RECT 23.530 177.180 23.850 177.240 ;
        RECT 26.305 177.380 26.595 177.425 ;
        RECT 26.750 177.380 27.070 177.440 ;
        RECT 26.305 177.240 27.070 177.380 ;
        RECT 38.340 177.380 38.480 177.920 ;
        RECT 39.645 178.060 39.935 178.105 ;
        RECT 40.090 178.060 40.410 178.120 ;
        RECT 39.645 177.920 40.410 178.060 ;
        RECT 41.100 178.060 41.240 178.215 ;
        RECT 43.785 178.060 44.075 178.105 ;
        RECT 41.100 177.920 44.075 178.060 ;
        RECT 39.645 177.875 39.935 177.920 ;
        RECT 40.090 177.860 40.410 177.920 ;
        RECT 43.785 177.875 44.075 177.920 ;
        RECT 39.170 177.720 39.490 177.780 ;
        RECT 44.320 177.720 44.460 178.260 ;
        RECT 46.085 178.215 46.375 178.445 ;
        RECT 47.005 178.400 47.295 178.445 ;
        RECT 47.450 178.400 47.770 178.460 ;
        RECT 48.000 178.445 48.140 178.600 ;
        RECT 51.590 178.600 55.590 178.740 ;
        RECT 55.820 178.740 55.960 178.940 ;
        RECT 56.665 178.940 57.890 179.080 ;
        RECT 56.665 178.895 56.955 178.940 ;
        RECT 57.570 178.880 57.890 178.940 ;
        RECT 65.390 179.080 65.710 179.140 ;
        RECT 70.005 179.080 70.295 179.125 ;
        RECT 65.390 178.940 70.295 179.080 ;
        RECT 65.390 178.880 65.710 178.940 ;
        RECT 70.005 178.895 70.295 178.940 ;
        RECT 57.110 178.740 57.430 178.800 ;
        RECT 58.505 178.740 58.795 178.785 ;
        RECT 55.820 178.600 58.795 178.740 ;
        RECT 51.590 178.540 51.910 178.600 ;
        RECT 55.270 178.540 55.590 178.600 ;
        RECT 57.110 178.540 57.430 178.600 ;
        RECT 58.505 178.555 58.795 178.600 ;
        RECT 60.790 178.540 61.110 178.800 ;
        RECT 61.710 178.785 62.030 178.800 ;
        RECT 61.710 178.555 62.095 178.785 ;
        RECT 62.630 178.740 62.950 178.800 ;
        RECT 64.330 178.740 64.620 178.785 ;
        RECT 62.630 178.600 64.620 178.740 ;
        RECT 61.710 178.540 62.030 178.555 ;
        RECT 62.630 178.540 62.950 178.600 ;
        RECT 64.330 178.555 64.620 178.600 ;
        RECT 47.005 178.260 47.770 178.400 ;
        RECT 47.005 178.215 47.295 178.260 ;
        RECT 44.690 177.860 45.010 178.120 ;
        RECT 46.160 178.060 46.300 178.215 ;
        RECT 47.450 178.200 47.770 178.260 ;
        RECT 47.925 178.215 48.215 178.445 ;
        RECT 49.305 178.400 49.595 178.445 ;
        RECT 49.750 178.400 50.070 178.460 ;
        RECT 49.305 178.260 50.070 178.400 ;
        RECT 49.305 178.215 49.595 178.260 ;
        RECT 49.750 178.200 50.070 178.260 ;
        RECT 50.685 178.215 50.975 178.445 ;
        RECT 48.370 178.060 48.690 178.120 ;
        RECT 46.160 177.920 48.690 178.060 ;
        RECT 39.170 177.580 44.460 177.720 ;
        RECT 39.170 177.520 39.490 177.580 ;
        RECT 40.550 177.380 40.870 177.440 ;
        RECT 38.340 177.240 40.870 177.380 ;
        RECT 26.305 177.195 26.595 177.240 ;
        RECT 26.750 177.180 27.070 177.240 ;
        RECT 40.550 177.180 40.870 177.240 ;
        RECT 41.010 177.380 41.330 177.440 ;
        RECT 46.160 177.380 46.300 177.920 ;
        RECT 48.370 177.860 48.690 177.920 ;
        RECT 48.830 178.060 49.150 178.120 ;
        RECT 50.760 178.060 50.900 178.215 ;
        RECT 51.130 178.200 51.450 178.460 ;
        RECT 52.510 178.200 52.830 178.460 ;
        RECT 52.970 178.200 53.290 178.460 ;
        RECT 53.905 178.400 54.195 178.445 ;
        RECT 60.330 178.400 60.650 178.460 ;
        RECT 53.905 178.260 55.040 178.400 ;
        RECT 53.905 178.215 54.195 178.260 ;
        RECT 54.900 178.120 55.040 178.260 ;
        RECT 55.820 178.260 60.650 178.400 ;
        RECT 48.830 177.920 50.900 178.060 ;
        RECT 48.830 177.860 49.150 177.920 ;
        RECT 54.810 177.860 55.130 178.120 ;
        RECT 55.285 177.875 55.575 178.105 ;
        RECT 54.350 177.720 54.670 177.780 ;
        RECT 55.360 177.720 55.500 177.875 ;
        RECT 54.350 177.580 55.500 177.720 ;
        RECT 54.350 177.520 54.670 177.580 ;
        RECT 41.010 177.240 46.300 177.380 ;
        RECT 41.010 177.180 41.330 177.240 ;
        RECT 49.290 177.180 49.610 177.440 ;
        RECT 55.820 177.425 55.960 178.260 ;
        RECT 60.330 178.200 60.650 178.260 ;
        RECT 62.170 178.060 62.490 178.120 ;
        RECT 58.580 177.920 62.490 178.060 ;
        RECT 56.650 177.720 56.970 177.780 ;
        RECT 57.585 177.720 57.875 177.765 ;
        RECT 56.650 177.580 57.875 177.720 ;
        RECT 56.650 177.520 56.970 177.580 ;
        RECT 57.585 177.535 57.875 177.580 ;
        RECT 58.580 177.425 58.720 177.920 ;
        RECT 62.170 177.860 62.490 177.920 ;
        RECT 63.090 177.860 63.410 178.120 ;
        RECT 63.985 178.060 64.275 178.105 ;
        RECT 65.175 178.060 65.465 178.105 ;
        RECT 67.695 178.060 67.985 178.105 ;
        RECT 63.985 177.920 67.985 178.060 ;
        RECT 63.985 177.875 64.275 177.920 ;
        RECT 65.175 177.875 65.465 177.920 ;
        RECT 67.695 177.875 67.985 177.920 ;
        RECT 63.590 177.720 63.880 177.765 ;
        RECT 65.690 177.720 65.980 177.765 ;
        RECT 67.260 177.720 67.550 177.765 ;
        RECT 63.590 177.580 67.550 177.720 ;
        RECT 63.590 177.535 63.880 177.580 ;
        RECT 65.690 177.535 65.980 177.580 ;
        RECT 67.260 177.535 67.550 177.580 ;
        RECT 55.745 177.195 56.035 177.425 ;
        RECT 58.505 177.195 58.795 177.425 ;
        RECT 61.250 177.380 61.570 177.440 ;
        RECT 61.725 177.380 62.015 177.425 ;
        RECT 61.250 177.240 62.015 177.380 ;
        RECT 61.250 177.180 61.570 177.240 ;
        RECT 61.725 177.195 62.015 177.240 ;
        RECT 62.645 177.380 62.935 177.425 ;
        RECT 64.010 177.380 64.330 177.440 ;
        RECT 62.645 177.240 64.330 177.380 ;
        RECT 62.645 177.195 62.935 177.240 ;
        RECT 64.010 177.180 64.330 177.240 ;
        RECT 5.520 176.560 84.180 177.040 ;
        RECT 10.650 176.360 10.970 176.420 ;
        RECT 11.125 176.360 11.415 176.405 ;
        RECT 10.650 176.220 11.415 176.360 ;
        RECT 10.650 176.160 10.970 176.220 ;
        RECT 11.125 176.175 11.415 176.220 ;
        RECT 20.785 176.360 21.075 176.405 ;
        RECT 23.070 176.360 23.390 176.420 ;
        RECT 20.785 176.220 23.390 176.360 ;
        RECT 20.785 176.175 21.075 176.220 ;
        RECT 23.070 176.160 23.390 176.220 ;
        RECT 28.590 176.360 28.910 176.420 ;
        RECT 29.065 176.360 29.355 176.405 ;
        RECT 28.590 176.220 29.355 176.360 ;
        RECT 28.590 176.160 28.910 176.220 ;
        RECT 29.065 176.175 29.355 176.220 ;
        RECT 29.970 176.160 30.290 176.420 ;
        RECT 40.090 176.160 40.410 176.420 ;
        RECT 41.930 176.160 42.250 176.420 ;
        RECT 42.940 176.220 44.000 176.360 ;
        RECT 13.870 176.020 14.160 176.065 ;
        RECT 15.440 176.020 15.730 176.065 ;
        RECT 17.540 176.020 17.830 176.065 ;
        RECT 13.870 175.880 17.830 176.020 ;
        RECT 13.870 175.835 14.160 175.880 ;
        RECT 15.440 175.835 15.730 175.880 ;
        RECT 17.540 175.835 17.830 175.880 ;
        RECT 18.945 176.020 19.235 176.065 ;
        RECT 20.310 176.020 20.630 176.080 ;
        RECT 18.945 175.880 20.630 176.020 ;
        RECT 18.945 175.835 19.235 175.880 ;
        RECT 20.310 175.820 20.630 175.880 ;
        RECT 22.650 176.020 22.940 176.065 ;
        RECT 24.750 176.020 25.040 176.065 ;
        RECT 26.320 176.020 26.610 176.065 ;
        RECT 22.650 175.880 26.610 176.020 ;
        RECT 22.650 175.835 22.940 175.880 ;
        RECT 24.750 175.835 25.040 175.880 ;
        RECT 26.320 175.835 26.610 175.880 ;
        RECT 29.510 176.020 29.830 176.080 ;
        RECT 30.905 176.020 31.195 176.065 ;
        RECT 34.110 176.020 34.430 176.080 ;
        RECT 29.510 175.880 34.430 176.020 ;
        RECT 29.510 175.820 29.830 175.880 ;
        RECT 30.905 175.835 31.195 175.880 ;
        RECT 34.110 175.820 34.430 175.880 ;
        RECT 13.435 175.680 13.725 175.725 ;
        RECT 15.955 175.680 16.245 175.725 ;
        RECT 17.145 175.680 17.435 175.725 ;
        RECT 13.435 175.540 17.435 175.680 ;
        RECT 13.435 175.495 13.725 175.540 ;
        RECT 15.955 175.495 16.245 175.540 ;
        RECT 17.145 175.495 17.435 175.540 ;
        RECT 23.045 175.680 23.335 175.725 ;
        RECT 24.235 175.680 24.525 175.725 ;
        RECT 26.755 175.680 27.045 175.725 ;
        RECT 23.045 175.540 27.045 175.680 ;
        RECT 23.045 175.495 23.335 175.540 ;
        RECT 24.235 175.495 24.525 175.540 ;
        RECT 26.755 175.495 27.045 175.540 ;
        RECT 18.010 175.140 18.330 175.400 ;
        RECT 22.165 175.340 22.455 175.385 ;
        RECT 30.430 175.340 30.750 175.400 ;
        RECT 22.165 175.200 30.750 175.340 ;
        RECT 22.165 175.155 22.455 175.200 ;
        RECT 30.430 175.140 30.750 175.200 ;
        RECT 37.790 175.340 38.110 175.400 ;
        RECT 38.265 175.340 38.555 175.385 ;
        RECT 37.790 175.200 38.555 175.340 ;
        RECT 37.790 175.140 38.110 175.200 ;
        RECT 38.265 175.155 38.555 175.200 ;
        RECT 39.170 175.140 39.490 175.400 ;
        RECT 40.180 175.340 40.320 176.160 ;
        RECT 40.550 175.680 40.870 175.740 ;
        RECT 41.485 175.680 41.775 175.725 ;
        RECT 40.550 175.540 41.775 175.680 ;
        RECT 40.550 175.480 40.870 175.540 ;
        RECT 41.485 175.495 41.775 175.540 ;
        RECT 41.025 175.340 41.315 175.385 ;
        RECT 40.180 175.200 41.315 175.340 ;
        RECT 41.025 175.155 41.315 175.200 ;
        RECT 42.405 175.340 42.695 175.385 ;
        RECT 42.940 175.340 43.080 176.220 ;
        RECT 43.325 175.835 43.615 176.065 ;
        RECT 43.860 176.020 44.000 176.220 ;
        RECT 44.690 176.160 45.010 176.420 ;
        RECT 48.830 176.160 49.150 176.420 ;
        RECT 49.750 176.160 50.070 176.420 ;
        RECT 50.685 176.360 50.975 176.405 ;
        RECT 51.130 176.360 51.450 176.420 ;
        RECT 54.825 176.360 55.115 176.405 ;
        RECT 50.685 176.220 55.115 176.360 ;
        RECT 50.685 176.175 50.975 176.220 ;
        RECT 51.130 176.160 51.450 176.220 ;
        RECT 54.825 176.175 55.115 176.220 ;
        RECT 61.710 176.360 62.030 176.420 ;
        RECT 61.710 176.220 64.240 176.360 ;
        RECT 61.710 176.160 62.030 176.220 ;
        RECT 46.530 176.020 46.850 176.080 ;
        RECT 52.050 176.020 52.370 176.080 ;
        RECT 43.860 175.880 52.370 176.020 ;
        RECT 42.405 175.200 43.080 175.340 ;
        RECT 43.400 175.340 43.540 175.835 ;
        RECT 46.530 175.820 46.850 175.880 ;
        RECT 52.050 175.820 52.370 175.880 ;
        RECT 52.985 176.020 53.275 176.065 ;
        RECT 53.890 176.020 54.210 176.080 ;
        RECT 52.985 175.880 54.210 176.020 ;
        RECT 52.985 175.835 53.275 175.880 ;
        RECT 53.890 175.820 54.210 175.880 ;
        RECT 47.005 175.680 47.295 175.725 ;
        RECT 49.750 175.680 50.070 175.740 ;
        RECT 61.250 175.680 61.570 175.740 ;
        RECT 64.100 175.725 64.240 176.220 ;
        RECT 47.005 175.540 48.370 175.680 ;
        RECT 47.005 175.495 47.295 175.540 ;
        RECT 48.230 175.400 48.370 175.540 ;
        RECT 49.750 175.540 61.570 175.680 ;
        RECT 49.750 175.480 50.070 175.540 ;
        RECT 61.250 175.480 61.570 175.540 ;
        RECT 62.645 175.680 62.935 175.725 ;
        RECT 62.645 175.540 63.780 175.680 ;
        RECT 62.645 175.495 62.935 175.540 ;
        RECT 45.625 175.340 45.915 175.385 ;
        RECT 43.400 175.200 45.915 175.340 ;
        RECT 42.405 175.155 42.695 175.200 ;
        RECT 45.625 175.155 45.915 175.200 ;
        RECT 46.085 175.155 46.375 175.385 ;
        RECT 15.250 175.000 15.570 175.060 ;
        RECT 16.690 175.000 16.980 175.045 ;
        RECT 23.390 175.000 23.680 175.045 ;
        RECT 15.250 174.860 16.980 175.000 ;
        RECT 15.250 174.800 15.570 174.860 ;
        RECT 16.690 174.815 16.980 174.860 ;
        RECT 21.780 174.860 23.680 175.000 ;
        RECT 20.770 174.460 21.090 174.720 ;
        RECT 21.780 174.705 21.920 174.860 ;
        RECT 23.390 174.815 23.680 174.860 ;
        RECT 27.670 175.000 27.990 175.060 ;
        RECT 32.285 175.000 32.575 175.045 ;
        RECT 27.670 174.860 32.575 175.000 ;
        RECT 27.670 174.800 27.990 174.860 ;
        RECT 32.285 174.815 32.575 174.860 ;
        RECT 33.650 175.000 33.970 175.060 ;
        RECT 41.470 175.000 41.790 175.060 ;
        RECT 46.160 175.000 46.300 175.155 ;
        RECT 47.450 175.140 47.770 175.400 ;
        RECT 48.230 175.200 48.690 175.400 ;
        RECT 48.370 175.140 48.690 175.200 ;
        RECT 49.305 175.340 49.595 175.385 ;
        RECT 52.510 175.340 52.830 175.400 ;
        RECT 53.445 175.340 53.735 175.385 ;
        RECT 49.305 175.200 52.280 175.340 ;
        RECT 49.305 175.155 49.595 175.200 ;
        RECT 33.650 174.860 46.300 175.000 ;
        RECT 48.460 175.000 48.600 175.140 ;
        RECT 52.140 175.060 52.280 175.200 ;
        RECT 52.510 175.200 53.735 175.340 ;
        RECT 52.510 175.140 52.830 175.200 ;
        RECT 53.445 175.155 53.735 175.200 ;
        RECT 56.205 175.155 56.495 175.385 ;
        RECT 51.130 175.000 51.450 175.060 ;
        RECT 48.460 174.860 51.450 175.000 ;
        RECT 33.650 174.800 33.970 174.860 ;
        RECT 41.470 174.800 41.790 174.860 ;
        RECT 51.130 174.800 51.450 174.860 ;
        RECT 51.590 174.800 51.910 175.060 ;
        RECT 52.050 174.800 52.370 175.060 ;
        RECT 21.705 174.475 21.995 174.705 ;
        RECT 50.605 174.660 50.895 174.705 ;
        RECT 53.445 174.660 53.735 174.705 ;
        RECT 50.605 174.520 53.735 174.660 ;
        RECT 56.280 174.660 56.420 175.155 ;
        RECT 56.650 175.140 56.970 175.400 ;
        RECT 57.125 175.340 57.415 175.385 ;
        RECT 57.570 175.340 57.890 175.400 ;
        RECT 57.125 175.200 57.890 175.340 ;
        RECT 57.125 175.155 57.415 175.200 ;
        RECT 57.570 175.140 57.890 175.200 ;
        RECT 58.030 175.140 58.350 175.400 ;
        RECT 63.640 175.385 63.780 175.540 ;
        RECT 64.025 175.495 64.315 175.725 ;
        RECT 62.215 175.155 62.505 175.385 ;
        RECT 63.105 175.155 63.395 175.385 ;
        RECT 63.565 175.155 63.855 175.385 ;
        RECT 64.485 175.340 64.775 175.385 ;
        RECT 64.930 175.340 65.250 175.400 ;
        RECT 64.485 175.200 65.250 175.340 ;
        RECT 64.485 175.155 64.775 175.200 ;
        RECT 60.330 175.000 60.650 175.060 ;
        RECT 62.260 175.000 62.400 175.155 ;
        RECT 60.330 174.860 62.400 175.000 ;
        RECT 60.330 174.800 60.650 174.860 ;
        RECT 62.170 174.660 62.490 174.720 ;
        RECT 56.280 174.520 62.490 174.660 ;
        RECT 63.180 174.660 63.320 175.155 ;
        RECT 64.930 175.140 65.250 175.200 ;
        RECT 63.550 174.660 63.870 174.720 ;
        RECT 63.180 174.520 63.870 174.660 ;
        RECT 50.605 174.475 50.895 174.520 ;
        RECT 53.445 174.475 53.735 174.520 ;
        RECT 62.170 174.460 62.490 174.520 ;
        RECT 63.550 174.460 63.870 174.520 ;
        RECT 5.520 173.840 84.180 174.320 ;
        RECT 15.250 173.440 15.570 173.700 ;
        RECT 41.930 173.640 42.250 173.700 ;
        RECT 55.730 173.640 56.050 173.700 ;
        RECT 41.930 173.500 56.050 173.640 ;
        RECT 41.930 173.440 42.250 173.500 ;
        RECT 55.730 173.440 56.050 173.500 ;
        RECT 10.650 173.300 10.970 173.360 ;
        RECT 12.965 173.300 13.255 173.345 ;
        RECT 10.650 173.160 13.255 173.300 ;
        RECT 10.650 173.100 10.970 173.160 ;
        RECT 12.965 173.115 13.255 173.160 ;
        RECT 53.430 173.300 53.750 173.360 ;
        RECT 56.650 173.300 56.970 173.360 ;
        RECT 64.485 173.300 64.775 173.345 ;
        RECT 65.850 173.300 66.170 173.360 ;
        RECT 53.430 173.160 56.970 173.300 ;
        RECT 53.430 173.100 53.750 173.160 ;
        RECT 56.650 173.100 56.970 173.160 ;
        RECT 63.640 173.160 64.775 173.300 ;
        RECT 63.640 173.020 63.780 173.160 ;
        RECT 64.485 173.115 64.775 173.160 ;
        RECT 65.020 173.160 66.170 173.300 ;
        RECT 36.885 172.960 37.175 173.005 ;
        RECT 37.330 172.960 37.650 173.020 ;
        RECT 36.885 172.820 37.650 172.960 ;
        RECT 36.885 172.775 37.175 172.820 ;
        RECT 37.330 172.760 37.650 172.820 ;
        RECT 37.805 172.960 38.095 173.005 ;
        RECT 41.010 172.960 41.330 173.020 ;
        RECT 37.805 172.820 41.330 172.960 ;
        RECT 37.805 172.775 38.095 172.820 ;
        RECT 41.010 172.760 41.330 172.820 ;
        RECT 61.250 172.760 61.570 173.020 ;
        RECT 62.630 172.760 62.950 173.020 ;
        RECT 63.550 172.760 63.870 173.020 ;
        RECT 64.010 172.760 64.330 173.020 ;
        RECT 65.020 173.005 65.160 173.160 ;
        RECT 65.850 173.100 66.170 173.160 ;
        RECT 64.945 172.775 65.235 173.005 ;
        RECT 65.390 172.760 65.710 173.020 ;
        RECT 66.325 172.960 66.615 173.005 ;
        RECT 66.770 172.960 67.090 173.020 ;
        RECT 66.325 172.820 67.090 172.960 ;
        RECT 66.325 172.775 66.615 172.820 ;
        RECT 66.770 172.760 67.090 172.820 ;
        RECT 60.805 172.620 61.095 172.665 ;
        RECT 62.170 172.620 62.490 172.680 ;
        RECT 60.805 172.480 62.490 172.620 ;
        RECT 60.805 172.435 61.095 172.480 ;
        RECT 14.330 172.280 14.650 172.340 ;
        RECT 20.770 172.280 21.090 172.340 ;
        RECT 14.330 172.140 21.090 172.280 ;
        RECT 14.330 172.080 14.650 172.140 ;
        RECT 20.770 172.080 21.090 172.140 ;
        RECT 36.410 172.280 36.730 172.340 ;
        RECT 43.310 172.280 43.630 172.340 ;
        RECT 46.070 172.280 46.390 172.340 ;
        RECT 36.410 172.140 46.390 172.280 ;
        RECT 61.800 172.280 61.940 172.480 ;
        RECT 62.170 172.420 62.490 172.480 ;
        RECT 63.105 172.620 63.395 172.665 ;
        RECT 64.470 172.620 64.790 172.680 ;
        RECT 63.105 172.480 64.790 172.620 ;
        RECT 63.105 172.435 63.395 172.480 ;
        RECT 64.470 172.420 64.790 172.480 ;
        RECT 64.010 172.280 64.330 172.340 ;
        RECT 61.800 172.140 64.330 172.280 ;
        RECT 36.410 172.080 36.730 172.140 ;
        RECT 43.310 172.080 43.630 172.140 ;
        RECT 46.070 172.080 46.390 172.140 ;
        RECT 64.010 172.080 64.330 172.140 ;
        RECT 35.950 171.940 36.270 172.000 ;
        RECT 36.885 171.940 37.175 171.985 ;
        RECT 35.950 171.800 37.175 171.940 ;
        RECT 35.950 171.740 36.270 171.800 ;
        RECT 36.885 171.755 37.175 171.800 ;
        RECT 45.150 171.940 45.470 172.000 ;
        RECT 61.710 171.940 62.030 172.000 ;
        RECT 45.150 171.800 62.030 171.940 ;
        RECT 45.150 171.740 45.470 171.800 ;
        RECT 61.710 171.740 62.030 171.800 ;
        RECT 63.550 171.940 63.870 172.000 ;
        RECT 64.930 171.940 65.250 172.000 ;
        RECT 63.550 171.800 65.250 171.940 ;
        RECT 63.550 171.740 63.870 171.800 ;
        RECT 64.930 171.740 65.250 171.800 ;
        RECT 5.520 171.120 84.180 171.600 ;
        RECT 22.610 170.920 22.930 170.980 ;
        RECT 23.085 170.920 23.375 170.965 ;
        RECT 22.610 170.780 23.375 170.920 ;
        RECT 22.610 170.720 22.930 170.780 ;
        RECT 23.085 170.735 23.375 170.780 ;
        RECT 25.385 170.920 25.675 170.965 ;
        RECT 29.510 170.920 29.830 170.980 ;
        RECT 25.385 170.780 29.830 170.920 ;
        RECT 25.385 170.735 25.675 170.780 ;
        RECT 20.770 170.580 21.090 170.640 ;
        RECT 24.465 170.580 24.755 170.625 ;
        RECT 20.770 170.440 24.755 170.580 ;
        RECT 20.770 170.380 21.090 170.440 ;
        RECT 24.465 170.395 24.755 170.440 ;
        RECT 22.150 170.240 22.470 170.300 ;
        RECT 25.460 170.240 25.600 170.735 ;
        RECT 29.510 170.720 29.830 170.780 ;
        RECT 35.965 170.920 36.255 170.965 ;
        RECT 36.410 170.920 36.730 170.980 ;
        RECT 35.965 170.780 36.730 170.920 ;
        RECT 35.965 170.735 36.255 170.780 ;
        RECT 36.410 170.720 36.730 170.780 ;
        RECT 38.265 170.920 38.555 170.965 ;
        RECT 39.170 170.920 39.490 170.980 ;
        RECT 38.265 170.780 39.490 170.920 ;
        RECT 38.265 170.735 38.555 170.780 ;
        RECT 39.170 170.720 39.490 170.780 ;
        RECT 41.010 170.720 41.330 170.980 ;
        RECT 51.145 170.920 51.435 170.965 ;
        RECT 52.050 170.920 52.370 170.980 ;
        RECT 51.145 170.780 52.370 170.920 ;
        RECT 51.145 170.735 51.435 170.780 ;
        RECT 52.050 170.720 52.370 170.780 ;
        RECT 62.185 170.920 62.475 170.965 ;
        RECT 62.630 170.920 62.950 170.980 ;
        RECT 62.185 170.780 62.950 170.920 ;
        RECT 62.185 170.735 62.475 170.780 ;
        RECT 62.630 170.720 62.950 170.780 ;
        RECT 65.390 170.920 65.710 170.980 ;
        RECT 68.610 170.920 68.930 170.980 ;
        RECT 65.390 170.780 68.930 170.920 ;
        RECT 65.390 170.720 65.710 170.780 ;
        RECT 68.610 170.720 68.930 170.780 ;
        RECT 36.870 170.580 37.190 170.640 ;
        RECT 39.630 170.580 39.950 170.640 ;
        RECT 46.085 170.580 46.375 170.625 ;
        RECT 36.870 170.440 46.375 170.580 ;
        RECT 36.870 170.380 37.190 170.440 ;
        RECT 39.630 170.380 39.950 170.440 ;
        RECT 46.085 170.395 46.375 170.440 ;
        RECT 50.685 170.395 50.975 170.625 ;
        RECT 58.965 170.580 59.255 170.625 ;
        RECT 63.550 170.580 63.870 170.640 ;
        RECT 58.965 170.440 63.870 170.580 ;
        RECT 58.965 170.395 59.255 170.440 ;
        RECT 22.150 170.100 25.600 170.240 ;
        RECT 22.150 170.040 22.470 170.100 ;
        RECT 30.430 170.040 30.750 170.300 ;
        RECT 50.210 170.240 50.530 170.300 ;
        RECT 34.660 170.100 50.530 170.240 ;
        RECT 50.760 170.240 50.900 170.395 ;
        RECT 63.550 170.380 63.870 170.440 ;
        RECT 64.930 170.580 65.250 170.640 ;
        RECT 66.770 170.580 67.090 170.640 ;
        RECT 64.930 170.440 67.090 170.580 ;
        RECT 64.930 170.380 65.250 170.440 ;
        RECT 66.770 170.380 67.090 170.440 ;
        RECT 70.950 170.580 71.240 170.625 ;
        RECT 73.050 170.580 73.340 170.625 ;
        RECT 74.620 170.580 74.910 170.625 ;
        RECT 70.950 170.440 74.910 170.580 ;
        RECT 70.950 170.395 71.240 170.440 ;
        RECT 73.050 170.395 73.340 170.440 ;
        RECT 74.620 170.395 74.910 170.440 ;
        RECT 61.725 170.240 62.015 170.285 ;
        RECT 62.170 170.240 62.490 170.300 ;
        RECT 69.530 170.240 69.850 170.300 ;
        RECT 70.465 170.240 70.755 170.285 ;
        RECT 50.760 170.100 54.120 170.240 ;
        RECT 21.690 169.900 22.010 169.960 ;
        RECT 23.530 169.900 23.850 169.960 ;
        RECT 34.660 169.945 34.800 170.100 ;
        RECT 50.210 170.040 50.530 170.100 ;
        RECT 21.690 169.760 23.850 169.900 ;
        RECT 21.690 169.700 22.010 169.760 ;
        RECT 23.530 169.700 23.850 169.760 ;
        RECT 34.585 169.715 34.875 169.945 ;
        RECT 35.030 169.900 35.350 169.960 ;
        RECT 39.645 169.900 39.935 169.945 ;
        RECT 35.030 169.760 39.935 169.900 ;
        RECT 35.030 169.700 35.350 169.760 ;
        RECT 19.850 169.560 20.170 169.620 ;
        RECT 22.165 169.560 22.455 169.605 ;
        RECT 19.850 169.420 22.455 169.560 ;
        RECT 23.620 169.560 23.760 169.700 ;
        RECT 25.225 169.560 25.515 169.605 ;
        RECT 23.620 169.420 25.515 169.560 ;
        RECT 19.850 169.360 20.170 169.420 ;
        RECT 22.165 169.375 22.455 169.420 ;
        RECT 25.225 169.375 25.515 169.420 ;
        RECT 26.305 169.560 26.595 169.605 ;
        RECT 27.210 169.560 27.530 169.620 ;
        RECT 35.950 169.605 36.270 169.620 ;
        RECT 26.305 169.420 27.530 169.560 ;
        RECT 26.305 169.375 26.595 169.420 ;
        RECT 27.210 169.360 27.530 169.420 ;
        RECT 35.885 169.375 36.270 169.605 ;
        RECT 35.950 169.360 36.270 169.375 ;
        RECT 36.870 169.360 37.190 169.620 ;
        RECT 38.340 169.605 38.480 169.760 ;
        RECT 39.645 169.715 39.935 169.760 ;
        RECT 40.090 169.900 40.410 169.960 ;
        RECT 41.025 169.900 41.315 169.945 ;
        RECT 40.090 169.760 41.315 169.900 ;
        RECT 40.090 169.700 40.410 169.760 ;
        RECT 41.025 169.715 41.315 169.760 ;
        RECT 45.150 169.700 45.470 169.960 ;
        RECT 47.465 169.900 47.755 169.945 ;
        RECT 49.290 169.900 49.610 169.960 ;
        RECT 47.465 169.760 49.610 169.900 ;
        RECT 47.465 169.715 47.755 169.760 ;
        RECT 49.290 169.700 49.610 169.760 ;
        RECT 49.750 169.700 50.070 169.960 ;
        RECT 50.685 169.715 50.975 169.945 ;
        RECT 38.185 169.420 38.480 169.605 ;
        RECT 38.185 169.375 38.475 169.420 ;
        RECT 39.185 169.375 39.475 169.605 ;
        RECT 46.070 169.560 46.390 169.620 ;
        RECT 46.545 169.560 46.835 169.605 ;
        RECT 46.070 169.420 46.835 169.560 ;
        RECT 50.760 169.560 50.900 169.715 ;
        RECT 52.050 169.700 52.370 169.960 ;
        RECT 53.980 169.945 54.120 170.100 ;
        RECT 56.280 170.100 62.490 170.240 ;
        RECT 56.280 169.960 56.420 170.100 ;
        RECT 61.725 170.055 62.015 170.100 ;
        RECT 62.170 170.040 62.490 170.100 ;
        RECT 63.180 170.100 66.080 170.240 ;
        RECT 53.905 169.715 54.195 169.945 ;
        RECT 55.730 169.900 56.050 169.960 ;
        RECT 55.535 169.760 56.050 169.900 ;
        RECT 55.730 169.700 56.050 169.760 ;
        RECT 56.190 169.700 56.510 169.960 ;
        RECT 60.345 169.900 60.635 169.945 ;
        RECT 61.250 169.900 61.570 169.960 ;
        RECT 63.180 169.945 63.320 170.100 ;
        RECT 65.940 169.960 66.080 170.100 ;
        RECT 69.530 170.100 70.755 170.240 ;
        RECT 69.530 170.040 69.850 170.100 ;
        RECT 70.465 170.055 70.755 170.100 ;
        RECT 71.345 170.240 71.635 170.285 ;
        RECT 72.535 170.240 72.825 170.285 ;
        RECT 75.055 170.240 75.345 170.285 ;
        RECT 71.345 170.100 75.345 170.240 ;
        RECT 71.345 170.055 71.635 170.100 ;
        RECT 72.535 170.055 72.825 170.100 ;
        RECT 75.055 170.055 75.345 170.100 ;
        RECT 60.345 169.760 61.570 169.900 ;
        RECT 60.345 169.715 60.635 169.760 ;
        RECT 61.250 169.700 61.570 169.760 ;
        RECT 63.105 169.715 63.395 169.945 ;
        RECT 64.010 169.700 64.330 169.960 ;
        RECT 65.850 169.700 66.170 169.960 ;
        RECT 67.245 169.900 67.535 169.945 ;
        RECT 71.745 169.900 72.035 169.945 ;
        RECT 67.245 169.760 72.035 169.900 ;
        RECT 67.245 169.715 67.535 169.760 ;
        RECT 71.745 169.715 72.035 169.760 ;
        RECT 52.525 169.560 52.815 169.605 ;
        RECT 50.760 169.420 52.815 169.560 ;
        RECT 23.070 169.265 23.390 169.280 ;
        RECT 23.070 169.035 23.455 169.265 ;
        RECT 23.070 169.020 23.390 169.035 ;
        RECT 23.990 169.020 24.310 169.280 ;
        RECT 34.570 169.220 34.890 169.280 ;
        RECT 35.045 169.220 35.335 169.265 ;
        RECT 34.570 169.080 35.335 169.220 ;
        RECT 34.570 169.020 34.890 169.080 ;
        RECT 35.045 169.035 35.335 169.080 ;
        RECT 37.330 169.020 37.650 169.280 ;
        RECT 39.260 169.220 39.400 169.375 ;
        RECT 46.070 169.360 46.390 169.420 ;
        RECT 46.545 169.375 46.835 169.420 ;
        RECT 52.525 169.375 52.815 169.420 ;
        RECT 52.985 169.560 53.275 169.605 ;
        RECT 54.365 169.560 54.655 169.605 ;
        RECT 52.985 169.420 54.655 169.560 ;
        RECT 52.985 169.375 53.275 169.420 ;
        RECT 54.365 169.375 54.655 169.420 ;
        RECT 59.885 169.560 60.175 169.605 ;
        RECT 61.710 169.560 62.030 169.620 ;
        RECT 64.485 169.560 64.775 169.605 ;
        RECT 66.325 169.560 66.615 169.605 ;
        RECT 67.705 169.560 67.995 169.605 ;
        RECT 59.885 169.420 61.480 169.560 ;
        RECT 59.885 169.375 60.175 169.420 ;
        RECT 40.105 169.220 40.395 169.265 ;
        RECT 40.550 169.220 40.870 169.280 ;
        RECT 39.260 169.080 40.870 169.220 ;
        RECT 52.600 169.220 52.740 169.375 ;
        RECT 59.960 169.220 60.100 169.375 ;
        RECT 52.600 169.080 60.100 169.220 ;
        RECT 60.330 169.220 60.650 169.280 ;
        RECT 60.805 169.220 61.095 169.265 ;
        RECT 60.330 169.080 61.095 169.220 ;
        RECT 61.340 169.220 61.480 169.420 ;
        RECT 61.710 169.420 66.080 169.560 ;
        RECT 61.710 169.360 62.030 169.420 ;
        RECT 64.485 169.375 64.775 169.420 ;
        RECT 65.940 169.280 66.080 169.420 ;
        RECT 66.325 169.420 67.995 169.560 ;
        RECT 66.325 169.375 66.615 169.420 ;
        RECT 67.705 169.375 67.995 169.420 ;
        RECT 68.610 169.360 68.930 169.620 ;
        RECT 69.545 169.375 69.835 169.605 ;
        RECT 64.930 169.220 65.250 169.280 ;
        RECT 61.340 169.080 65.250 169.220 ;
        RECT 40.105 169.035 40.395 169.080 ;
        RECT 40.550 169.020 40.870 169.080 ;
        RECT 60.330 169.020 60.650 169.080 ;
        RECT 60.805 169.035 61.095 169.080 ;
        RECT 64.930 169.020 65.250 169.080 ;
        RECT 65.390 169.020 65.710 169.280 ;
        RECT 65.850 169.020 66.170 169.280 ;
        RECT 66.770 169.220 67.090 169.280 ;
        RECT 69.620 169.220 69.760 169.375 ;
        RECT 77.365 169.220 77.655 169.265 ;
        RECT 66.770 169.080 77.655 169.220 ;
        RECT 66.770 169.020 67.090 169.080 ;
        RECT 77.365 169.035 77.655 169.080 ;
        RECT 5.520 168.400 84.180 168.880 ;
        RECT 22.610 168.000 22.930 168.260 ;
        RECT 49.750 168.200 50.070 168.260 ;
        RECT 53.890 168.200 54.210 168.260 ;
        RECT 34.660 168.060 54.210 168.200 ;
        RECT 18.010 167.860 18.330 167.920 ;
        RECT 23.070 167.860 23.390 167.920 ;
        RECT 30.430 167.860 30.750 167.920 ;
        RECT 14.420 167.720 23.390 167.860 ;
        RECT 14.420 167.565 14.560 167.720 ;
        RECT 18.010 167.660 18.330 167.720 ;
        RECT 23.070 167.660 23.390 167.720 ;
        RECT 24.080 167.720 30.750 167.860 ;
        RECT 14.345 167.335 14.635 167.565 ;
        RECT 14.790 167.520 15.110 167.580 ;
        RECT 15.625 167.520 15.915 167.565 ;
        RECT 14.790 167.380 15.915 167.520 ;
        RECT 14.790 167.320 15.110 167.380 ;
        RECT 15.625 167.335 15.915 167.380 ;
        RECT 21.690 167.320 22.010 167.580 ;
        RECT 22.150 167.520 22.470 167.580 ;
        RECT 22.625 167.520 22.915 167.565 ;
        RECT 24.080 167.520 24.220 167.720 ;
        RECT 30.430 167.660 30.750 167.720 ;
        RECT 24.450 167.565 24.770 167.580 ;
        RECT 22.150 167.380 22.915 167.520 ;
        RECT 22.150 167.320 22.470 167.380 ;
        RECT 22.625 167.335 22.915 167.380 ;
        RECT 23.160 167.380 24.220 167.520 ;
        RECT 24.420 167.520 24.770 167.565 ;
        RECT 34.110 167.520 34.430 167.580 ;
        RECT 34.660 167.565 34.800 168.060 ;
        RECT 49.750 168.000 50.070 168.060 ;
        RECT 53.890 168.000 54.210 168.060 ;
        RECT 57.585 168.200 57.875 168.245 ;
        RECT 58.030 168.200 58.350 168.260 ;
        RECT 57.585 168.060 58.350 168.200 ;
        RECT 57.585 168.015 57.875 168.060 ;
        RECT 58.030 168.000 58.350 168.060 ;
        RECT 58.490 168.000 58.810 168.260 ;
        RECT 50.670 167.860 50.990 167.920 ;
        RECT 63.090 167.860 63.410 167.920 ;
        RECT 42.480 167.720 63.410 167.860 ;
        RECT 42.480 167.580 42.620 167.720 ;
        RECT 50.670 167.660 50.990 167.720 ;
        RECT 63.090 167.660 63.410 167.720 ;
        RECT 34.585 167.520 34.875 167.565 ;
        RECT 24.420 167.380 24.920 167.520 ;
        RECT 34.110 167.380 34.875 167.520 ;
        RECT 23.160 167.225 23.300 167.380 ;
        RECT 24.420 167.335 24.770 167.380 ;
        RECT 24.450 167.320 24.770 167.335 ;
        RECT 34.110 167.320 34.430 167.380 ;
        RECT 34.585 167.335 34.875 167.380 ;
        RECT 38.725 167.520 39.015 167.565 ;
        RECT 41.470 167.520 41.790 167.580 ;
        RECT 38.725 167.380 41.790 167.520 ;
        RECT 38.725 167.335 39.015 167.380 ;
        RECT 41.470 167.320 41.790 167.380 ;
        RECT 41.945 167.520 42.235 167.565 ;
        RECT 42.390 167.520 42.710 167.580 ;
        RECT 43.310 167.565 43.630 167.580 ;
        RECT 41.945 167.380 42.710 167.520 ;
        RECT 41.945 167.335 42.235 167.380 ;
        RECT 42.390 167.320 42.710 167.380 ;
        RECT 43.280 167.335 43.630 167.565 ;
        RECT 49.305 167.520 49.595 167.565 ;
        RECT 43.310 167.320 43.630 167.335 ;
        RECT 48.920 167.380 49.595 167.520 ;
        RECT 15.225 167.180 15.515 167.225 ;
        RECT 16.415 167.180 16.705 167.225 ;
        RECT 18.935 167.180 19.225 167.225 ;
        RECT 15.225 167.040 19.225 167.180 ;
        RECT 15.225 166.995 15.515 167.040 ;
        RECT 16.415 166.995 16.705 167.040 ;
        RECT 18.935 166.995 19.225 167.040 ;
        RECT 23.085 166.995 23.375 167.225 ;
        RECT 23.965 167.180 24.255 167.225 ;
        RECT 25.155 167.180 25.445 167.225 ;
        RECT 27.675 167.180 27.965 167.225 ;
        RECT 23.965 167.040 27.965 167.180 ;
        RECT 23.965 166.995 24.255 167.040 ;
        RECT 25.155 166.995 25.445 167.040 ;
        RECT 27.675 166.995 27.965 167.040 ;
        RECT 32.745 167.180 33.035 167.225 ;
        RECT 37.805 167.180 38.095 167.225 ;
        RECT 32.745 167.040 38.095 167.180 ;
        RECT 32.745 166.995 33.035 167.040 ;
        RECT 37.805 166.995 38.095 167.040 ;
        RECT 42.825 167.180 43.115 167.225 ;
        RECT 44.015 167.180 44.305 167.225 ;
        RECT 46.535 167.180 46.825 167.225 ;
        RECT 42.825 167.040 46.825 167.180 ;
        RECT 42.825 166.995 43.115 167.040 ;
        RECT 44.015 166.995 44.305 167.040 ;
        RECT 46.535 166.995 46.825 167.040 ;
        RECT 14.830 166.840 15.120 166.885 ;
        RECT 16.930 166.840 17.220 166.885 ;
        RECT 18.500 166.840 18.790 166.885 ;
        RECT 14.830 166.700 18.790 166.840 ;
        RECT 14.830 166.655 15.120 166.700 ;
        RECT 16.930 166.655 17.220 166.700 ;
        RECT 18.500 166.655 18.790 166.700 ;
        RECT 23.570 166.840 23.860 166.885 ;
        RECT 25.670 166.840 25.960 166.885 ;
        RECT 27.240 166.840 27.530 166.885 ;
        RECT 23.570 166.700 27.530 166.840 ;
        RECT 23.570 166.655 23.860 166.700 ;
        RECT 25.670 166.655 25.960 166.700 ;
        RECT 27.240 166.655 27.530 166.700 ;
        RECT 38.250 166.640 38.570 166.900 ;
        RECT 42.430 166.840 42.720 166.885 ;
        RECT 44.530 166.840 44.820 166.885 ;
        RECT 46.100 166.840 46.390 166.885 ;
        RECT 42.430 166.700 46.390 166.840 ;
        RECT 42.430 166.655 42.720 166.700 ;
        RECT 44.530 166.655 44.820 166.700 ;
        RECT 46.100 166.655 46.390 166.700 ;
        RECT 19.390 166.500 19.710 166.560 ;
        RECT 21.245 166.500 21.535 166.545 ;
        RECT 19.390 166.360 21.535 166.500 ;
        RECT 19.390 166.300 19.710 166.360 ;
        RECT 21.245 166.315 21.535 166.360 ;
        RECT 21.690 166.500 22.010 166.560 ;
        RECT 23.990 166.500 24.310 166.560 ;
        RECT 21.690 166.360 24.310 166.500 ;
        RECT 21.690 166.300 22.010 166.360 ;
        RECT 23.990 166.300 24.310 166.360 ;
        RECT 29.510 166.500 29.830 166.560 ;
        RECT 29.985 166.500 30.275 166.545 ;
        RECT 29.510 166.360 30.275 166.500 ;
        RECT 29.510 166.300 29.830 166.360 ;
        RECT 29.985 166.315 30.275 166.360 ;
        RECT 43.770 166.500 44.090 166.560 ;
        RECT 47.450 166.500 47.770 166.560 ;
        RECT 48.920 166.545 49.060 167.380 ;
        RECT 49.305 167.335 49.595 167.380 ;
        RECT 49.750 167.520 50.070 167.580 ;
        RECT 51.145 167.520 51.435 167.565 ;
        RECT 49.750 167.380 51.435 167.520 ;
        RECT 49.750 167.320 50.070 167.380 ;
        RECT 51.145 167.335 51.435 167.380 ;
        RECT 53.890 167.320 54.210 167.580 ;
        RECT 58.490 167.520 58.780 167.565 ;
        RECT 59.870 167.520 60.190 167.580 ;
        RECT 58.490 167.380 60.190 167.520 ;
        RECT 58.490 167.335 58.780 167.380 ;
        RECT 59.870 167.320 60.190 167.380 ;
        RECT 60.345 167.520 60.635 167.565 ;
        RECT 61.250 167.520 61.570 167.580 ;
        RECT 64.010 167.520 64.330 167.580 ;
        RECT 68.670 167.520 68.960 167.565 ;
        RECT 60.345 167.380 62.170 167.520 ;
        RECT 60.345 167.335 60.635 167.380 ;
        RECT 61.250 167.320 61.570 167.380 ;
        RECT 50.225 167.180 50.515 167.225 ;
        RECT 56.190 167.180 56.510 167.240 ;
        RECT 50.225 167.040 56.510 167.180 ;
        RECT 50.225 166.995 50.515 167.040 ;
        RECT 56.190 166.980 56.510 167.040 ;
        RECT 60.790 166.980 61.110 167.240 ;
        RECT 49.765 166.840 50.055 166.885 ;
        RECT 52.050 166.840 52.370 166.900 ;
        RECT 49.765 166.700 52.370 166.840 ;
        RECT 62.030 166.840 62.170 167.380 ;
        RECT 64.010 167.380 68.960 167.520 ;
        RECT 64.010 167.320 64.330 167.380 ;
        RECT 68.670 167.335 68.960 167.380 ;
        RECT 69.530 167.520 69.850 167.580 ;
        RECT 70.005 167.520 70.295 167.565 ;
        RECT 69.530 167.380 70.295 167.520 ;
        RECT 69.530 167.320 69.850 167.380 ;
        RECT 70.005 167.335 70.295 167.380 ;
        RECT 65.415 167.180 65.705 167.225 ;
        RECT 67.935 167.180 68.225 167.225 ;
        RECT 69.125 167.180 69.415 167.225 ;
        RECT 65.415 167.040 69.415 167.180 ;
        RECT 65.415 166.995 65.705 167.040 ;
        RECT 67.935 166.995 68.225 167.040 ;
        RECT 69.125 166.995 69.415 167.040 ;
        RECT 63.105 166.840 63.395 166.885 ;
        RECT 62.030 166.700 63.395 166.840 ;
        RECT 49.765 166.655 50.055 166.700 ;
        RECT 52.050 166.640 52.370 166.700 ;
        RECT 63.105 166.655 63.395 166.700 ;
        RECT 65.850 166.840 66.140 166.885 ;
        RECT 67.420 166.840 67.710 166.885 ;
        RECT 69.520 166.840 69.810 166.885 ;
        RECT 65.850 166.700 69.810 166.840 ;
        RECT 65.850 166.655 66.140 166.700 ;
        RECT 67.420 166.655 67.710 166.700 ;
        RECT 69.520 166.655 69.810 166.700 ;
        RECT 48.845 166.500 49.135 166.545 ;
        RECT 43.770 166.360 49.135 166.500 ;
        RECT 43.770 166.300 44.090 166.360 ;
        RECT 47.450 166.300 47.770 166.360 ;
        RECT 48.845 166.315 49.135 166.360 ;
        RECT 50.225 166.500 50.515 166.545 ;
        RECT 52.510 166.500 52.830 166.560 ;
        RECT 50.225 166.360 52.830 166.500 ;
        RECT 50.225 166.315 50.515 166.360 ;
        RECT 52.510 166.300 52.830 166.360 ;
        RECT 52.970 166.300 53.290 166.560 ;
        RECT 53.890 166.500 54.210 166.560 ;
        RECT 63.550 166.500 63.870 166.560 ;
        RECT 53.890 166.360 63.870 166.500 ;
        RECT 53.890 166.300 54.210 166.360 ;
        RECT 63.550 166.300 63.870 166.360 ;
        RECT 5.520 165.680 84.180 166.160 ;
        RECT 14.790 165.280 15.110 165.540 ;
        RECT 15.725 165.480 16.015 165.525 ;
        RECT 18.945 165.480 19.235 165.525 ;
        RECT 34.110 165.480 34.430 165.540 ;
        RECT 15.725 165.340 19.235 165.480 ;
        RECT 15.725 165.295 16.015 165.340 ;
        RECT 18.945 165.295 19.235 165.340 ;
        RECT 28.680 165.340 34.430 165.480 ;
        RECT 17.565 165.140 17.855 165.185 ;
        RECT 20.310 165.140 20.630 165.200 ;
        RECT 17.565 165.000 20.630 165.140 ;
        RECT 17.565 164.955 17.855 165.000 ;
        RECT 20.310 164.940 20.630 165.000 ;
        RECT 23.990 164.800 24.310 164.860 ;
        RECT 21.320 164.660 24.310 164.800 ;
        RECT 21.320 164.520 21.460 164.660 ;
        RECT 23.990 164.600 24.310 164.660 ;
        RECT 19.390 164.460 19.710 164.520 ;
        RECT 19.865 164.460 20.155 164.505 ;
        RECT 19.390 164.320 20.155 164.460 ;
        RECT 19.390 164.260 19.710 164.320 ;
        RECT 19.865 164.275 20.155 164.320 ;
        RECT 19.940 164.120 20.080 164.275 ;
        RECT 21.230 164.260 21.550 164.520 ;
        RECT 23.070 164.260 23.390 164.520 ;
        RECT 27.670 164.260 27.990 164.520 ;
        RECT 28.680 164.505 28.820 165.340 ;
        RECT 34.110 165.280 34.430 165.340 ;
        RECT 40.090 165.280 40.410 165.540 ;
        RECT 43.310 165.480 43.630 165.540 ;
        RECT 43.785 165.480 44.075 165.525 ;
        RECT 43.310 165.340 44.075 165.480 ;
        RECT 43.310 165.280 43.630 165.340 ;
        RECT 43.785 165.295 44.075 165.340 ;
        RECT 46.530 165.480 46.850 165.540 ;
        RECT 49.290 165.480 49.610 165.540 ;
        RECT 46.530 165.340 49.610 165.480 ;
        RECT 46.530 165.280 46.850 165.340 ;
        RECT 49.290 165.280 49.610 165.340 ;
        RECT 64.010 165.280 64.330 165.540 ;
        RECT 64.945 165.480 65.235 165.525 ;
        RECT 65.390 165.480 65.710 165.540 ;
        RECT 64.945 165.340 65.710 165.480 ;
        RECT 64.945 165.295 65.235 165.340 ;
        RECT 33.690 165.140 33.980 165.185 ;
        RECT 35.790 165.140 36.080 165.185 ;
        RECT 37.360 165.140 37.650 165.185 ;
        RECT 33.690 165.000 37.650 165.140 ;
        RECT 33.690 164.955 33.980 165.000 ;
        RECT 35.790 164.955 36.080 165.000 ;
        RECT 37.360 164.955 37.650 165.000 ;
        RECT 41.470 165.140 41.790 165.200 ;
        RECT 46.990 165.140 47.310 165.200 ;
        RECT 48.845 165.140 49.135 165.185 ;
        RECT 41.470 165.000 55.960 165.140 ;
        RECT 41.470 164.940 41.790 165.000 ;
        RECT 46.990 164.940 47.310 165.000 ;
        RECT 48.845 164.955 49.135 165.000 ;
        RECT 55.820 164.860 55.960 165.000 ;
        RECT 34.085 164.800 34.375 164.845 ;
        RECT 35.275 164.800 35.565 164.845 ;
        RECT 37.795 164.800 38.085 164.845 ;
        RECT 34.085 164.660 38.085 164.800 ;
        RECT 34.085 164.615 34.375 164.660 ;
        RECT 35.275 164.615 35.565 164.660 ;
        RECT 37.795 164.615 38.085 164.660 ;
        RECT 40.640 164.660 45.840 164.800 ;
        RECT 28.605 164.275 28.895 164.505 ;
        RECT 29.985 164.460 30.275 164.505 ;
        RECT 30.430 164.460 30.750 164.520 ;
        RECT 32.270 164.460 32.590 164.520 ;
        RECT 34.570 164.505 34.890 164.520 ;
        RECT 33.205 164.460 33.495 164.505 ;
        RECT 34.540 164.460 34.890 164.505 ;
        RECT 29.985 164.320 33.495 164.460 ;
        RECT 34.375 164.320 34.890 164.460 ;
        RECT 29.985 164.275 30.275 164.320 ;
        RECT 30.430 164.260 30.750 164.320 ;
        RECT 32.270 164.260 32.590 164.320 ;
        RECT 33.205 164.275 33.495 164.320 ;
        RECT 34.540 164.275 34.890 164.320 ;
        RECT 34.570 164.260 34.890 164.275 ;
        RECT 36.870 164.460 37.190 164.520 ;
        RECT 40.640 164.505 40.780 164.660 ;
        RECT 40.565 164.460 40.855 164.505 ;
        RECT 36.870 164.320 40.855 164.460 ;
        RECT 36.870 164.260 37.190 164.320 ;
        RECT 40.565 164.275 40.855 164.320 ;
        RECT 41.470 164.260 41.790 164.520 ;
        RECT 41.945 164.275 42.235 164.505 ;
        RECT 42.405 164.460 42.695 164.505 ;
        RECT 43.770 164.460 44.090 164.520 ;
        RECT 42.405 164.320 44.090 164.460 ;
        RECT 42.405 164.275 42.695 164.320 ;
        RECT 21.690 164.120 22.010 164.180 ;
        RECT 19.940 163.980 22.010 164.120 ;
        RECT 21.690 163.920 22.010 163.980 ;
        RECT 29.525 164.120 29.815 164.165 ;
        RECT 35.030 164.120 35.350 164.180 ;
        RECT 29.525 163.980 35.350 164.120 ;
        RECT 29.525 163.935 29.815 163.980 ;
        RECT 35.030 163.920 35.350 163.980 ;
        RECT 37.330 164.120 37.650 164.180 ;
        RECT 42.020 164.120 42.160 164.275 ;
        RECT 43.770 164.260 44.090 164.320 ;
        RECT 44.705 164.460 44.995 164.505 ;
        RECT 45.150 164.460 45.470 164.520 ;
        RECT 45.700 164.505 45.840 164.660 ;
        RECT 49.750 164.600 50.070 164.860 ;
        RECT 50.670 164.800 50.990 164.860 ;
        RECT 53.905 164.800 54.195 164.845 ;
        RECT 54.350 164.800 54.670 164.860 ;
        RECT 50.670 164.660 54.670 164.800 ;
        RECT 50.670 164.600 50.990 164.660 ;
        RECT 53.905 164.615 54.195 164.660 ;
        RECT 54.350 164.600 54.670 164.660 ;
        RECT 55.730 164.600 56.050 164.860 ;
        RECT 58.045 164.800 58.335 164.845 ;
        RECT 60.790 164.800 61.110 164.860 ;
        RECT 65.020 164.800 65.160 165.295 ;
        RECT 65.390 165.280 65.710 165.340 ;
        RECT 58.045 164.660 61.110 164.800 ;
        RECT 58.045 164.615 58.335 164.660 ;
        RECT 60.790 164.600 61.110 164.660 ;
        RECT 62.030 164.660 65.160 164.800 ;
        RECT 44.705 164.320 45.470 164.460 ;
        RECT 44.705 164.275 44.995 164.320 ;
        RECT 37.330 163.980 42.160 164.120 ;
        RECT 42.850 164.120 43.170 164.180 ;
        RECT 44.780 164.120 44.920 164.275 ;
        RECT 45.150 164.260 45.470 164.320 ;
        RECT 45.625 164.275 45.915 164.505 ;
        RECT 46.085 164.275 46.375 164.505 ;
        RECT 46.160 164.120 46.300 164.275 ;
        RECT 50.210 164.260 50.530 164.520 ;
        RECT 52.970 164.460 53.290 164.520 ;
        RECT 56.205 164.460 56.495 164.505 ;
        RECT 51.220 164.320 56.495 164.460 ;
        RECT 51.220 164.180 51.360 164.320 ;
        RECT 52.970 164.260 53.290 164.320 ;
        RECT 56.205 164.275 56.495 164.320 ;
        RECT 47.465 164.120 47.755 164.165 ;
        RECT 51.130 164.120 51.450 164.180 ;
        RECT 42.850 163.980 44.920 164.120 ;
        RECT 45.240 163.980 51.450 164.120 ;
        RECT 37.330 163.920 37.650 163.980 ;
        RECT 42.850 163.920 43.170 163.980 ;
        RECT 15.725 163.780 16.015 163.825 ;
        RECT 17.550 163.780 17.870 163.840 ;
        RECT 19.850 163.780 20.170 163.840 ;
        RECT 15.725 163.640 20.170 163.780 ;
        RECT 15.725 163.595 16.015 163.640 ;
        RECT 17.550 163.580 17.870 163.640 ;
        RECT 19.850 163.580 20.170 163.640 ;
        RECT 20.310 163.780 20.630 163.840 ;
        RECT 20.785 163.780 21.075 163.825 ;
        RECT 29.050 163.780 29.370 163.840 ;
        RECT 20.310 163.640 29.370 163.780 ;
        RECT 20.310 163.580 20.630 163.640 ;
        RECT 20.785 163.595 21.075 163.640 ;
        RECT 29.050 163.580 29.370 163.640 ;
        RECT 31.350 163.780 31.670 163.840 ;
        RECT 45.240 163.780 45.380 163.980 ;
        RECT 47.465 163.935 47.755 163.980 ;
        RECT 51.130 163.920 51.450 163.980 ;
        RECT 31.350 163.640 45.380 163.780 ;
        RECT 31.350 163.580 31.670 163.640 ;
        RECT 45.610 163.580 45.930 163.840 ;
        RECT 46.070 163.780 46.390 163.840 ;
        RECT 62.030 163.780 62.170 164.660 ;
        RECT 63.105 164.460 63.395 164.505 ;
        RECT 69.530 164.460 69.850 164.520 ;
        RECT 63.105 164.320 69.850 164.460 ;
        RECT 63.105 164.275 63.395 164.320 ;
        RECT 69.530 164.260 69.850 164.320 ;
        RECT 64.470 164.165 64.790 164.180 ;
        RECT 64.470 163.935 65.075 164.165 ;
        RECT 64.470 163.920 64.790 163.935 ;
        RECT 65.850 163.920 66.170 164.180 ;
        RECT 46.070 163.640 62.170 163.780 ;
        RECT 46.070 163.580 46.390 163.640 ;
        RECT 5.520 162.960 84.180 163.440 ;
        RECT 19.405 162.760 19.695 162.805 ;
        RECT 21.230 162.760 21.550 162.820 ;
        RECT 19.405 162.620 21.550 162.760 ;
        RECT 19.405 162.575 19.695 162.620 ;
        RECT 21.230 162.560 21.550 162.620 ;
        RECT 25.830 162.760 26.150 162.820 ;
        RECT 38.250 162.760 38.570 162.820 ;
        RECT 52.510 162.760 52.830 162.820 ;
        RECT 25.830 162.620 52.830 162.760 ;
        RECT 25.830 162.560 26.150 162.620 ;
        RECT 38.250 162.560 38.570 162.620 ;
        RECT 52.510 162.560 52.830 162.620 ;
        RECT 56.665 162.760 56.955 162.805 ;
        RECT 58.490 162.760 58.810 162.820 ;
        RECT 56.665 162.620 58.810 162.760 ;
        RECT 56.665 162.575 56.955 162.620 ;
        RECT 58.490 162.560 58.810 162.620 ;
        RECT 16.185 162.420 16.475 162.465 ;
        RECT 20.770 162.420 21.090 162.480 ;
        RECT 16.185 162.280 21.090 162.420 ;
        RECT 16.185 162.235 16.475 162.280 ;
        RECT 20.770 162.220 21.090 162.280 ;
        RECT 28.605 162.420 28.895 162.465 ;
        RECT 31.350 162.420 31.670 162.480 ;
        RECT 28.605 162.280 31.670 162.420 ;
        RECT 28.605 162.235 28.895 162.280 ;
        RECT 31.350 162.220 31.670 162.280 ;
        RECT 50.210 162.420 50.530 162.480 ;
        RECT 59.410 162.420 59.730 162.480 ;
        RECT 60.805 162.420 61.095 162.465 ;
        RECT 50.210 162.280 61.095 162.420 ;
        RECT 50.210 162.220 50.530 162.280 ;
        RECT 59.410 162.220 59.730 162.280 ;
        RECT 60.805 162.235 61.095 162.280 ;
        RECT 64.945 162.420 65.235 162.465 ;
        RECT 69.530 162.420 69.850 162.480 ;
        RECT 64.945 162.280 69.850 162.420 ;
        RECT 64.945 162.235 65.235 162.280 ;
        RECT 69.530 162.220 69.850 162.280 ;
        RECT 17.105 161.895 17.395 162.125 ;
        RECT 17.180 161.740 17.320 161.895 ;
        RECT 19.850 161.880 20.170 162.140 ;
        RECT 20.325 162.080 20.615 162.125 ;
        RECT 21.690 162.080 22.010 162.140 ;
        RECT 20.325 161.940 24.220 162.080 ;
        RECT 20.325 161.895 20.615 161.940 ;
        RECT 21.690 161.880 22.010 161.940 ;
        RECT 22.625 161.740 22.915 161.785 ;
        RECT 23.070 161.740 23.390 161.800 ;
        RECT 17.180 161.600 21.460 161.740 ;
        RECT 21.320 161.445 21.460 161.600 ;
        RECT 22.625 161.600 23.390 161.740 ;
        RECT 24.080 161.740 24.220 161.940 ;
        RECT 26.290 161.880 26.610 162.140 ;
        RECT 27.685 161.895 27.975 162.125 ;
        RECT 29.065 162.080 29.355 162.125 ;
        RECT 29.510 162.080 29.830 162.140 ;
        RECT 29.065 161.940 29.830 162.080 ;
        RECT 29.065 161.895 29.355 161.940 ;
        RECT 27.210 161.740 27.530 161.800 ;
        RECT 27.760 161.740 27.900 161.895 ;
        RECT 29.510 161.880 29.830 161.940 ;
        RECT 50.670 161.880 50.990 162.140 ;
        RECT 51.130 162.080 51.450 162.140 ;
        RECT 55.730 162.125 56.050 162.140 ;
        RECT 54.825 162.080 55.115 162.125 ;
        RECT 51.130 161.940 55.115 162.080 ;
        RECT 51.130 161.880 51.450 161.940 ;
        RECT 54.825 161.895 55.115 161.940 ;
        RECT 55.595 161.895 56.050 162.125 ;
        RECT 55.730 161.880 56.050 161.895 ;
        RECT 56.190 162.080 56.510 162.140 ;
        RECT 58.045 162.080 58.335 162.125 ;
        RECT 56.190 161.940 58.335 162.080 ;
        RECT 56.190 161.880 56.510 161.940 ;
        RECT 58.045 161.895 58.335 161.940 ;
        RECT 29.970 161.740 30.290 161.800 ;
        RECT 24.080 161.600 30.290 161.740 ;
        RECT 22.625 161.555 22.915 161.600 ;
        RECT 23.070 161.540 23.390 161.600 ;
        RECT 27.210 161.540 27.530 161.600 ;
        RECT 29.970 161.540 30.290 161.600 ;
        RECT 21.245 161.400 21.535 161.445 ;
        RECT 23.990 161.400 24.310 161.460 ;
        RECT 21.245 161.260 24.310 161.400 ;
        RECT 21.245 161.215 21.535 161.260 ;
        RECT 23.990 161.200 24.310 161.260 ;
        RECT 18.010 160.860 18.330 161.120 ;
        RECT 18.470 160.860 18.790 161.120 ;
        RECT 24.910 161.060 25.230 161.120 ;
        RECT 26.765 161.060 27.055 161.105 ;
        RECT 24.910 160.920 27.055 161.060 ;
        RECT 55.820 161.060 55.960 161.880 ;
        RECT 57.110 161.060 57.430 161.120 ;
        RECT 58.505 161.060 58.795 161.105 ;
        RECT 55.820 160.920 58.795 161.060 ;
        RECT 24.910 160.860 25.230 160.920 ;
        RECT 26.765 160.875 27.055 160.920 ;
        RECT 57.110 160.860 57.430 160.920 ;
        RECT 58.505 160.875 58.795 160.920 ;
        RECT 5.520 160.240 84.180 160.720 ;
        RECT 18.010 160.040 18.330 160.100 ;
        RECT 20.785 160.040 21.075 160.085 ;
        RECT 18.010 159.900 21.075 160.040 ;
        RECT 18.010 159.840 18.330 159.900 ;
        RECT 20.785 159.855 21.075 159.900 ;
        RECT 23.530 160.040 23.850 160.100 ;
        RECT 24.005 160.040 24.295 160.085 ;
        RECT 29.510 160.040 29.830 160.100 ;
        RECT 23.530 159.900 24.295 160.040 ;
        RECT 23.530 159.840 23.850 159.900 ;
        RECT 24.005 159.855 24.295 159.900 ;
        RECT 24.540 159.900 29.830 160.040 ;
        RECT 18.470 159.700 18.790 159.760 ;
        RECT 18.945 159.700 19.235 159.745 ;
        RECT 18.470 159.560 19.235 159.700 ;
        RECT 18.470 159.500 18.790 159.560 ;
        RECT 18.945 159.515 19.235 159.560 ;
        RECT 24.540 159.360 24.680 159.900 ;
        RECT 29.510 159.840 29.830 159.900 ;
        RECT 35.030 160.040 35.350 160.100 ;
        RECT 35.030 159.900 48.600 160.040 ;
        RECT 35.030 159.840 35.350 159.900 ;
        RECT 25.830 159.700 26.150 159.760 ;
        RECT 27.210 159.700 27.530 159.760 ;
        RECT 28.605 159.700 28.895 159.745 ;
        RECT 25.830 159.560 26.520 159.700 ;
        RECT 25.830 159.500 26.150 159.560 ;
        RECT 21.780 159.220 24.680 159.360 ;
        RECT 14.790 159.020 15.110 159.080 ;
        RECT 14.790 158.880 19.620 159.020 ;
        RECT 14.790 158.820 15.110 158.880 ;
        RECT 19.480 158.680 19.620 158.880 ;
        RECT 20.785 158.680 21.075 158.725 ;
        RECT 19.480 158.540 21.075 158.680 ;
        RECT 21.780 158.680 21.920 159.220 ;
        RECT 22.165 159.020 22.455 159.065 ;
        RECT 24.450 159.020 24.770 159.080 ;
        RECT 22.165 158.880 24.770 159.020 ;
        RECT 22.165 158.835 22.455 158.880 ;
        RECT 24.450 158.820 24.770 158.880 ;
        RECT 24.910 158.820 25.230 159.080 ;
        RECT 26.380 159.065 26.520 159.560 ;
        RECT 27.210 159.560 28.895 159.700 ;
        RECT 27.210 159.500 27.530 159.560 ;
        RECT 28.605 159.515 28.895 159.560 ;
        RECT 30.890 159.700 31.210 159.760 ;
        RECT 30.890 159.560 43.080 159.700 ;
        RECT 30.890 159.500 31.210 159.560 ;
        RECT 26.750 159.160 27.070 159.420 ;
        RECT 29.065 159.360 29.355 159.405 ;
        RECT 27.760 159.220 29.355 159.360 ;
        RECT 27.760 159.065 27.900 159.220 ;
        RECT 29.065 159.175 29.355 159.220 ;
        RECT 29.510 159.360 29.830 159.420 ;
        RECT 29.510 159.220 31.120 159.360 ;
        RECT 29.510 159.160 29.830 159.220 ;
        RECT 25.845 159.020 26.135 159.065 ;
        RECT 25.735 158.880 26.135 159.020 ;
        RECT 25.845 158.835 26.135 158.880 ;
        RECT 26.305 159.020 26.595 159.065 ;
        RECT 26.305 158.880 26.705 159.020 ;
        RECT 26.305 158.835 26.595 158.880 ;
        RECT 27.685 158.835 27.975 159.065 ;
        RECT 23.085 158.680 23.375 158.725 ;
        RECT 21.780 158.540 23.375 158.680 ;
        RECT 20.785 158.495 21.075 158.540 ;
        RECT 23.085 158.495 23.375 158.540 ;
        RECT 23.990 158.680 24.310 158.740 ;
        RECT 25.920 158.680 26.060 158.835 ;
        RECT 23.990 158.540 26.060 158.680 ;
        RECT 26.380 158.680 26.520 158.835 ;
        RECT 29.970 158.820 30.290 159.080 ;
        RECT 30.980 159.065 31.120 159.220 ;
        RECT 35.030 159.160 35.350 159.420 ;
        RECT 42.940 159.405 43.080 159.560 ;
        RECT 42.865 159.175 43.155 159.405 ;
        RECT 30.905 158.835 31.195 159.065 ;
        RECT 31.350 158.820 31.670 159.080 ;
        RECT 34.570 158.820 34.890 159.080 ;
        RECT 41.945 159.020 42.235 159.065 ;
        RECT 35.120 158.880 42.235 159.020 ;
        RECT 26.750 158.680 27.070 158.740 ;
        RECT 26.380 158.540 27.070 158.680 ;
        RECT 23.990 158.480 24.310 158.540 ;
        RECT 26.750 158.480 27.070 158.540 ;
        RECT 34.110 158.680 34.430 158.740 ;
        RECT 35.120 158.680 35.260 158.880 ;
        RECT 41.945 158.835 42.235 158.880 ;
        RECT 42.390 158.820 42.710 159.080 ;
        RECT 43.325 159.020 43.615 159.065 ;
        RECT 46.530 159.020 46.850 159.080 ;
        RECT 48.460 159.065 48.600 159.900 ;
        RECT 53.060 159.560 61.020 159.700 ;
        RECT 51.605 159.360 51.895 159.405 ;
        RECT 51.605 159.220 52.740 159.360 ;
        RECT 51.605 159.175 51.895 159.220 ;
        RECT 47.005 159.020 47.295 159.065 ;
        RECT 43.325 158.880 47.295 159.020 ;
        RECT 43.325 158.835 43.615 158.880 ;
        RECT 46.530 158.820 46.850 158.880 ;
        RECT 47.005 158.835 47.295 158.880 ;
        RECT 48.385 158.835 48.675 159.065 ;
        RECT 51.130 158.820 51.450 159.080 ;
        RECT 52.600 159.065 52.740 159.220 ;
        RECT 52.065 159.020 52.355 159.065 ;
        RECT 51.955 158.880 52.355 159.020 ;
        RECT 52.600 158.880 52.915 159.065 ;
        RECT 52.065 158.835 52.355 158.880 ;
        RECT 52.625 158.835 52.915 158.880 ;
        RECT 34.110 158.540 35.260 158.680 ;
        RECT 40.105 158.680 40.395 158.725 ;
        RECT 40.105 158.540 47.220 158.680 ;
        RECT 34.110 158.480 34.430 158.540 ;
        RECT 40.105 158.495 40.395 158.540 ;
        RECT 47.080 158.400 47.220 158.540 ;
        RECT 47.925 158.495 48.215 158.725 ;
        RECT 52.140 158.680 52.280 158.835 ;
        RECT 53.060 158.680 53.200 159.560 ;
        RECT 55.745 159.360 56.035 159.405 ;
        RECT 53.520 159.220 56.035 159.360 ;
        RECT 53.520 159.065 53.660 159.220 ;
        RECT 55.745 159.175 56.035 159.220 ;
        RECT 60.345 159.175 60.635 159.405 ;
        RECT 53.445 158.835 53.735 159.065 ;
        RECT 53.905 158.835 54.195 159.065 ;
        RECT 54.485 159.020 54.775 159.065 ;
        RECT 57.110 159.020 57.430 159.080 ;
        RECT 54.440 158.835 54.775 159.020 ;
        RECT 56.915 158.880 57.430 159.020 ;
        RECT 53.980 158.680 54.120 158.835 ;
        RECT 52.140 158.540 54.120 158.680 ;
        RECT 21.690 158.140 22.010 158.400 ;
        RECT 32.730 158.140 33.050 158.400 ;
        RECT 39.630 158.140 39.950 158.400 ;
        RECT 40.550 158.340 40.870 158.400 ;
        RECT 41.025 158.340 41.315 158.385 ;
        RECT 40.550 158.200 41.315 158.340 ;
        RECT 40.550 158.140 40.870 158.200 ;
        RECT 41.025 158.155 41.315 158.200 ;
        RECT 45.610 158.340 45.930 158.400 ;
        RECT 46.085 158.340 46.375 158.385 ;
        RECT 45.610 158.200 46.375 158.340 ;
        RECT 45.610 158.140 45.930 158.200 ;
        RECT 46.085 158.155 46.375 158.200 ;
        RECT 46.990 158.140 47.310 158.400 ;
        RECT 47.450 158.340 47.770 158.400 ;
        RECT 48.000 158.340 48.140 158.495 ;
        RECT 49.305 158.340 49.595 158.385 ;
        RECT 54.440 158.340 54.580 158.835 ;
        RECT 57.110 158.820 57.430 158.880 ;
        RECT 57.570 159.020 57.890 159.080 ;
        RECT 60.420 159.020 60.560 159.175 ;
        RECT 60.880 159.065 61.020 159.560 ;
        RECT 62.645 159.360 62.935 159.405 ;
        RECT 65.530 159.360 65.820 159.405 ;
        RECT 62.645 159.220 65.820 159.360 ;
        RECT 62.645 159.175 62.935 159.220 ;
        RECT 65.530 159.175 65.820 159.220 ;
        RECT 57.570 158.880 60.560 159.020 ;
        RECT 60.805 159.020 61.095 159.065 ;
        RECT 62.170 159.020 62.490 159.080 ;
        RECT 60.805 158.880 62.490 159.020 ;
        RECT 57.570 158.820 57.890 158.880 ;
        RECT 60.805 158.835 61.095 158.880 ;
        RECT 62.170 158.820 62.490 158.880 ;
        RECT 63.090 158.820 63.410 159.080 ;
        RECT 64.470 158.820 64.790 159.080 ;
        RECT 64.930 158.820 65.250 159.080 ;
        RECT 47.450 158.200 54.580 158.340 ;
        RECT 47.450 158.140 47.770 158.200 ;
        RECT 49.305 158.155 49.595 158.200 ;
        RECT 55.270 158.140 55.590 158.400 ;
        RECT 66.325 158.340 66.615 158.385 ;
        RECT 66.770 158.340 67.090 158.400 ;
        RECT 66.325 158.200 67.090 158.340 ;
        RECT 66.325 158.155 66.615 158.200 ;
        RECT 66.770 158.140 67.090 158.200 ;
        RECT 5.520 157.520 84.180 158.000 ;
        RECT 16.645 157.135 16.935 157.365 ;
        RECT 16.720 156.640 16.860 157.135 ;
        RECT 23.530 157.120 23.850 157.380 ;
        RECT 23.990 157.320 24.310 157.380 ;
        RECT 24.925 157.320 25.215 157.365 ;
        RECT 23.990 157.180 25.215 157.320 ;
        RECT 23.990 157.120 24.310 157.180 ;
        RECT 24.925 157.135 25.215 157.180 ;
        RECT 30.905 157.320 31.195 157.365 ;
        RECT 35.030 157.320 35.350 157.380 ;
        RECT 39.185 157.320 39.475 157.365 ;
        RECT 42.390 157.320 42.710 157.380 ;
        RECT 30.905 157.180 35.350 157.320 ;
        RECT 38.975 157.180 42.710 157.320 ;
        RECT 30.905 157.135 31.195 157.180 ;
        RECT 35.030 157.120 35.350 157.180 ;
        RECT 39.185 157.135 39.475 157.180 ;
        RECT 21.690 156.980 22.010 157.040 ;
        RECT 22.210 156.980 22.500 157.025 ;
        RECT 21.690 156.840 22.500 156.980 ;
        RECT 21.690 156.780 22.010 156.840 ;
        RECT 22.210 156.795 22.500 156.840 ;
        RECT 23.620 156.640 23.760 157.120 ;
        RECT 34.110 156.980 34.430 157.040 ;
        RECT 30.060 156.840 34.430 156.980 ;
        RECT 25.830 156.640 26.150 156.700 ;
        RECT 30.060 156.685 30.200 156.840 ;
        RECT 34.110 156.780 34.430 156.840 ;
        RECT 34.570 156.980 34.890 157.040 ;
        RECT 39.260 156.980 39.400 157.135 ;
        RECT 42.390 157.120 42.710 157.180 ;
        RECT 46.530 157.120 46.850 157.380 ;
        RECT 54.350 156.980 54.670 157.040 ;
        RECT 65.850 156.980 66.170 157.040 ;
        RECT 66.770 157.025 67.090 157.040 ;
        RECT 34.570 156.840 39.400 156.980 ;
        RECT 39.720 156.840 54.670 156.980 ;
        RECT 34.570 156.780 34.890 156.840 ;
        RECT 16.720 156.500 26.150 156.640 ;
        RECT 25.830 156.440 26.150 156.500 ;
        RECT 29.985 156.455 30.275 156.685 ;
        RECT 30.890 156.640 31.210 156.700 ;
        RECT 31.810 156.640 32.130 156.700 ;
        RECT 30.890 156.500 32.130 156.640 ;
        RECT 30.890 156.440 31.210 156.500 ;
        RECT 31.810 156.440 32.130 156.500 ;
        RECT 32.270 156.440 32.590 156.700 ;
        RECT 33.650 156.685 33.970 156.700 ;
        RECT 39.720 156.685 39.860 156.840 ;
        RECT 54.350 156.780 54.670 156.840 ;
        RECT 62.030 156.840 66.170 156.980 ;
        RECT 41.010 156.685 41.330 156.700 ;
        RECT 33.620 156.455 33.970 156.685 ;
        RECT 39.645 156.455 39.935 156.685 ;
        RECT 40.980 156.455 41.330 156.685 ;
        RECT 33.650 156.440 33.970 156.455 ;
        RECT 41.010 156.440 41.330 156.455 ;
        RECT 45.610 156.640 45.930 156.700 ;
        RECT 49.305 156.640 49.595 156.685 ;
        RECT 45.610 156.500 49.595 156.640 ;
        RECT 45.610 156.440 45.930 156.500 ;
        RECT 49.305 156.455 49.595 156.500 ;
        RECT 49.750 156.640 50.070 156.700 ;
        RECT 50.225 156.640 50.515 156.685 ;
        RECT 49.750 156.500 50.515 156.640 ;
        RECT 49.750 156.440 50.070 156.500 ;
        RECT 50.225 156.455 50.515 156.500 ;
        RECT 50.685 156.640 50.975 156.685 ;
        RECT 57.570 156.640 57.890 156.700 ;
        RECT 62.030 156.640 62.170 156.840 ;
        RECT 65.850 156.780 66.170 156.840 ;
        RECT 66.740 156.795 67.090 157.025 ;
        RECT 66.770 156.780 67.090 156.795 ;
        RECT 67.690 156.780 68.010 157.040 ;
        RECT 67.780 156.640 67.920 156.780 ;
        RECT 50.685 156.500 62.170 156.640 ;
        RECT 65.020 156.500 67.920 156.640 ;
        RECT 50.685 156.455 50.975 156.500 ;
        RECT 57.570 156.440 57.890 156.500 ;
        RECT 65.020 156.360 65.160 156.500 ;
        RECT 18.955 156.300 19.245 156.345 ;
        RECT 21.475 156.300 21.765 156.345 ;
        RECT 22.665 156.300 22.955 156.345 ;
        RECT 18.955 156.160 22.955 156.300 ;
        RECT 18.955 156.115 19.245 156.160 ;
        RECT 21.475 156.115 21.765 156.160 ;
        RECT 22.665 156.115 22.955 156.160 ;
        RECT 23.530 156.100 23.850 156.360 ;
        RECT 27.225 156.300 27.515 156.345 ;
        RECT 28.130 156.300 28.450 156.360 ;
        RECT 27.225 156.160 28.450 156.300 ;
        RECT 27.225 156.115 27.515 156.160 ;
        RECT 28.130 156.100 28.450 156.160 ;
        RECT 33.165 156.300 33.455 156.345 ;
        RECT 34.355 156.300 34.645 156.345 ;
        RECT 36.875 156.300 37.165 156.345 ;
        RECT 33.165 156.160 37.165 156.300 ;
        RECT 33.165 156.115 33.455 156.160 ;
        RECT 34.355 156.115 34.645 156.160 ;
        RECT 36.875 156.115 37.165 156.160 ;
        RECT 40.525 156.300 40.815 156.345 ;
        RECT 41.715 156.300 42.005 156.345 ;
        RECT 44.235 156.300 44.525 156.345 ;
        RECT 40.525 156.160 44.525 156.300 ;
        RECT 40.525 156.115 40.815 156.160 ;
        RECT 41.715 156.115 42.005 156.160 ;
        RECT 44.235 156.115 44.525 156.160 ;
        RECT 46.990 156.300 47.310 156.360 ;
        RECT 64.930 156.300 65.250 156.360 ;
        RECT 46.990 156.160 65.250 156.300 ;
        RECT 46.990 156.100 47.310 156.160 ;
        RECT 64.930 156.100 65.250 156.160 ;
        RECT 65.405 156.300 65.695 156.345 ;
        RECT 66.285 156.300 66.575 156.345 ;
        RECT 67.475 156.300 67.765 156.345 ;
        RECT 69.995 156.300 70.285 156.345 ;
        RECT 65.405 156.115 65.745 156.300 ;
        RECT 66.285 156.160 70.285 156.300 ;
        RECT 66.285 156.115 66.575 156.160 ;
        RECT 67.475 156.115 67.765 156.160 ;
        RECT 69.995 156.115 70.285 156.160 ;
        RECT 19.390 155.960 19.680 156.005 ;
        RECT 20.960 155.960 21.250 156.005 ;
        RECT 23.060 155.960 23.350 156.005 ;
        RECT 19.390 155.820 23.350 155.960 ;
        RECT 19.390 155.775 19.680 155.820 ;
        RECT 20.960 155.775 21.250 155.820 ;
        RECT 23.060 155.775 23.350 155.820 ;
        RECT 32.770 155.960 33.060 156.005 ;
        RECT 34.870 155.960 35.160 156.005 ;
        RECT 36.440 155.960 36.730 156.005 ;
        RECT 32.770 155.820 36.730 155.960 ;
        RECT 32.770 155.775 33.060 155.820 ;
        RECT 34.870 155.775 35.160 155.820 ;
        RECT 36.440 155.775 36.730 155.820 ;
        RECT 40.130 155.960 40.420 156.005 ;
        RECT 42.230 155.960 42.520 156.005 ;
        RECT 43.800 155.960 44.090 156.005 ;
        RECT 40.130 155.820 44.090 155.960 ;
        RECT 40.130 155.775 40.420 155.820 ;
        RECT 42.230 155.775 42.520 155.820 ;
        RECT 43.800 155.775 44.090 155.820 ;
        RECT 44.690 155.960 45.010 156.020 ;
        RECT 63.090 155.960 63.410 156.020 ;
        RECT 64.010 155.960 64.330 156.020 ;
        RECT 44.690 155.820 64.330 155.960 ;
        RECT 44.690 155.760 45.010 155.820 ;
        RECT 63.090 155.760 63.410 155.820 ;
        RECT 64.010 155.760 64.330 155.820 ;
        RECT 26.765 155.620 27.055 155.665 ;
        RECT 27.670 155.620 27.990 155.680 ;
        RECT 26.765 155.480 27.990 155.620 ;
        RECT 26.765 155.435 27.055 155.480 ;
        RECT 27.670 155.420 27.990 155.480 ;
        RECT 48.385 155.620 48.675 155.665 ;
        RECT 53.430 155.620 53.750 155.680 ;
        RECT 48.385 155.480 53.750 155.620 ;
        RECT 48.385 155.435 48.675 155.480 ;
        RECT 53.430 155.420 53.750 155.480 ;
        RECT 53.890 155.620 54.210 155.680 ;
        RECT 64.930 155.620 65.250 155.680 ;
        RECT 53.890 155.480 65.250 155.620 ;
        RECT 65.605 155.620 65.745 156.115 ;
        RECT 65.890 155.960 66.180 156.005 ;
        RECT 67.990 155.960 68.280 156.005 ;
        RECT 69.560 155.960 69.850 156.005 ;
        RECT 65.890 155.820 69.850 155.960 ;
        RECT 65.890 155.775 66.180 155.820 ;
        RECT 67.990 155.775 68.280 155.820 ;
        RECT 69.560 155.775 69.850 155.820 ;
        RECT 70.450 155.620 70.770 155.680 ;
        RECT 65.605 155.480 70.770 155.620 ;
        RECT 53.890 155.420 54.210 155.480 ;
        RECT 64.930 155.420 65.250 155.480 ;
        RECT 70.450 155.420 70.770 155.480 ;
        RECT 72.290 155.420 72.610 155.680 ;
        RECT 5.520 154.800 84.180 155.280 ;
        RECT 32.745 154.600 33.035 154.645 ;
        RECT 33.650 154.600 33.970 154.660 ;
        RECT 32.745 154.460 33.970 154.600 ;
        RECT 32.745 154.415 33.035 154.460 ;
        RECT 33.650 154.400 33.970 154.460 ;
        RECT 41.010 154.400 41.330 154.660 ;
        RECT 46.545 154.600 46.835 154.645 ;
        RECT 46.990 154.600 47.310 154.660 ;
        RECT 46.545 154.460 47.310 154.600 ;
        RECT 46.545 154.415 46.835 154.460 ;
        RECT 46.990 154.400 47.310 154.460 ;
        RECT 52.985 154.600 53.275 154.645 ;
        RECT 55.270 154.600 55.590 154.660 ;
        RECT 52.985 154.460 55.590 154.600 ;
        RECT 52.985 154.415 53.275 154.460 ;
        RECT 55.270 154.400 55.590 154.460 ;
        RECT 64.010 154.600 64.330 154.660 ;
        RECT 66.310 154.600 66.630 154.660 ;
        RECT 64.010 154.460 66.630 154.600 ;
        RECT 64.010 154.400 64.330 154.460 ;
        RECT 66.310 154.400 66.630 154.460 ;
        RECT 44.690 154.260 45.010 154.320 ;
        RECT 37.880 154.120 45.010 154.260 ;
        RECT 18.470 153.920 18.790 153.980 ;
        RECT 25.830 153.920 26.150 153.980 ;
        RECT 27.225 153.920 27.515 153.965 ;
        RECT 18.470 153.780 20.080 153.920 ;
        RECT 18.470 153.720 18.790 153.780 ;
        RECT 18.945 153.580 19.235 153.625 ;
        RECT 19.390 153.580 19.710 153.640 ;
        RECT 19.940 153.625 20.080 153.780 ;
        RECT 25.830 153.780 27.515 153.920 ;
        RECT 25.830 153.720 26.150 153.780 ;
        RECT 27.225 153.735 27.515 153.780 ;
        RECT 32.730 153.920 33.050 153.980 ;
        RECT 37.880 153.965 38.020 154.120 ;
        RECT 44.690 154.060 45.010 154.120 ;
        RECT 49.305 154.260 49.595 154.305 ;
        RECT 50.225 154.260 50.515 154.305 ;
        RECT 53.890 154.260 54.210 154.320 ;
        RECT 60.345 154.260 60.635 154.305 ;
        RECT 49.305 154.120 50.515 154.260 ;
        RECT 49.305 154.075 49.595 154.120 ;
        RECT 50.225 154.075 50.515 154.120 ;
        RECT 50.760 154.120 54.210 154.260 ;
        RECT 33.540 153.920 33.830 153.965 ;
        RECT 32.730 153.780 33.830 153.920 ;
        RECT 32.730 153.720 33.050 153.780 ;
        RECT 33.540 153.735 33.830 153.780 ;
        RECT 35.965 153.920 36.255 153.965 ;
        RECT 37.805 153.920 38.095 153.965 ;
        RECT 50.760 153.920 50.900 154.120 ;
        RECT 53.890 154.060 54.210 154.120 ;
        RECT 56.740 154.120 60.635 154.260 ;
        RECT 35.965 153.780 38.095 153.920 ;
        RECT 35.965 153.735 36.255 153.780 ;
        RECT 37.805 153.735 38.095 153.780 ;
        RECT 43.400 153.780 50.900 153.920 ;
        RECT 52.065 153.920 52.355 153.965 ;
        RECT 55.730 153.920 56.050 153.980 ;
        RECT 52.065 153.780 56.050 153.920 ;
        RECT 18.945 153.440 19.710 153.580 ;
        RECT 18.945 153.395 19.235 153.440 ;
        RECT 19.390 153.380 19.710 153.440 ;
        RECT 19.865 153.395 20.155 153.625 ;
        RECT 26.305 153.580 26.595 153.625 ;
        RECT 26.750 153.580 27.070 153.640 ;
        RECT 26.305 153.440 27.070 153.580 ;
        RECT 26.305 153.395 26.595 153.440 ;
        RECT 26.750 153.380 27.070 153.440 ;
        RECT 40.090 153.625 40.410 153.640 ;
        RECT 40.090 153.395 40.520 153.625 ;
        RECT 40.090 153.380 40.410 153.395 ;
        RECT 34.585 153.240 34.875 153.285 ;
        RECT 39.185 153.240 39.475 153.285 ;
        RECT 41.930 153.240 42.250 153.300 ;
        RECT 34.585 153.100 42.250 153.240 ;
        RECT 34.585 153.055 34.875 153.100 ;
        RECT 39.185 153.055 39.475 153.100 ;
        RECT 41.930 153.040 42.250 153.100 ;
        RECT 15.710 152.900 16.030 152.960 ;
        RECT 18.945 152.900 19.235 152.945 ;
        RECT 15.710 152.760 19.235 152.900 ;
        RECT 15.710 152.700 16.030 152.760 ;
        RECT 18.945 152.715 19.235 152.760 ;
        RECT 23.990 152.900 24.310 152.960 ;
        RECT 25.385 152.900 25.675 152.945 ;
        RECT 23.990 152.760 25.675 152.900 ;
        RECT 23.990 152.700 24.310 152.760 ;
        RECT 25.385 152.715 25.675 152.760 ;
        RECT 34.125 152.900 34.415 152.945 ;
        RECT 35.030 152.900 35.350 152.960 ;
        RECT 39.630 152.900 39.950 152.960 ;
        RECT 43.400 152.900 43.540 153.780 ;
        RECT 52.065 153.735 52.355 153.780 ;
        RECT 55.730 153.720 56.050 153.780 ;
        RECT 56.740 153.640 56.880 154.120 ;
        RECT 60.345 154.075 60.635 154.120 ;
        RECT 64.930 154.260 65.250 154.320 ;
        RECT 67.230 154.260 67.550 154.320 ;
        RECT 64.930 154.120 67.550 154.260 ;
        RECT 64.930 154.060 65.250 154.120 ;
        RECT 67.230 154.060 67.550 154.120 ;
        RECT 70.950 154.260 71.240 154.305 ;
        RECT 73.050 154.260 73.340 154.305 ;
        RECT 74.620 154.260 74.910 154.305 ;
        RECT 70.950 154.120 74.910 154.260 ;
        RECT 70.950 154.075 71.240 154.120 ;
        RECT 73.050 154.075 73.340 154.120 ;
        RECT 74.620 154.075 74.910 154.120 ;
        RECT 58.490 153.720 58.810 153.980 ;
        RECT 60.790 153.920 61.110 153.980 ;
        RECT 62.645 153.920 62.935 153.965 ;
        RECT 69.990 153.920 70.310 153.980 ;
        RECT 60.790 153.780 62.935 153.920 ;
        RECT 60.790 153.720 61.110 153.780 ;
        RECT 62.645 153.735 62.935 153.780 ;
        RECT 65.020 153.780 70.310 153.920 ;
        RECT 46.530 153.580 46.850 153.640 ;
        RECT 47.170 153.580 47.460 153.625 ;
        RECT 46.530 153.440 47.460 153.580 ;
        RECT 46.530 153.380 46.850 153.440 ;
        RECT 47.170 153.395 47.460 153.440 ;
        RECT 49.750 153.380 50.070 153.640 ;
        RECT 51.130 153.380 51.450 153.640 ;
        RECT 53.430 153.380 53.750 153.640 ;
        RECT 54.810 153.380 55.130 153.640 ;
        RECT 55.285 153.395 55.575 153.625 ;
        RECT 56.205 153.580 56.495 153.625 ;
        RECT 55.820 153.440 56.495 153.580 ;
        RECT 55.360 153.240 55.500 153.395 ;
        RECT 48.230 153.100 55.500 153.240 ;
        RECT 34.125 152.760 43.540 152.900 ;
        RECT 46.530 152.900 46.850 152.960 ;
        RECT 47.450 152.900 47.770 152.960 ;
        RECT 48.230 152.900 48.370 153.100 ;
        RECT 46.530 152.760 48.370 152.900 ;
        RECT 34.125 152.715 34.415 152.760 ;
        RECT 35.030 152.700 35.350 152.760 ;
        RECT 39.630 152.700 39.950 152.760 ;
        RECT 46.530 152.700 46.850 152.760 ;
        RECT 47.450 152.700 47.770 152.760 ;
        RECT 53.890 152.700 54.210 152.960 ;
        RECT 55.820 152.900 55.960 153.440 ;
        RECT 56.205 153.395 56.495 153.440 ;
        RECT 56.650 153.380 56.970 153.640 ;
        RECT 58.950 153.380 59.270 153.640 ;
        RECT 62.170 153.380 62.490 153.640 ;
        RECT 64.010 153.380 64.330 153.640 ;
        RECT 65.020 153.625 65.160 153.780 ;
        RECT 69.990 153.720 70.310 153.780 ;
        RECT 70.450 153.720 70.770 153.980 ;
        RECT 71.345 153.920 71.635 153.965 ;
        RECT 72.535 153.920 72.825 153.965 ;
        RECT 75.055 153.920 75.345 153.965 ;
        RECT 71.345 153.780 75.345 153.920 ;
        RECT 71.345 153.735 71.635 153.780 ;
        RECT 72.535 153.735 72.825 153.780 ;
        RECT 75.055 153.735 75.345 153.780 ;
        RECT 64.945 153.395 65.235 153.625 ;
        RECT 65.405 153.580 65.695 153.625 ;
        RECT 66.310 153.580 66.630 153.640 ;
        RECT 65.405 153.440 66.630 153.580 ;
        RECT 65.405 153.395 65.695 153.440 ;
        RECT 66.310 153.380 66.630 153.440 ;
        RECT 67.230 153.380 67.550 153.640 ;
        RECT 64.485 153.240 64.775 153.285 ;
        RECT 67.830 153.240 68.120 153.285 ;
        RECT 71.690 153.240 71.980 153.285 ;
        RECT 64.485 153.100 68.120 153.240 ;
        RECT 64.485 153.055 64.775 153.100 ;
        RECT 67.830 153.055 68.120 153.100 ;
        RECT 68.700 153.100 71.980 153.240 ;
        RECT 56.190 152.900 56.510 152.960 ;
        RECT 57.125 152.900 57.415 152.945 ;
        RECT 55.820 152.760 57.415 152.900 ;
        RECT 56.190 152.700 56.510 152.760 ;
        RECT 57.125 152.715 57.415 152.760 ;
        RECT 65.390 152.900 65.710 152.960 ;
        RECT 68.700 152.945 68.840 153.100 ;
        RECT 71.690 153.055 71.980 153.100 ;
        RECT 66.785 152.900 67.075 152.945 ;
        RECT 65.390 152.760 67.075 152.900 ;
        RECT 65.390 152.700 65.710 152.760 ;
        RECT 66.785 152.715 67.075 152.760 ;
        RECT 68.625 152.715 68.915 152.945 ;
        RECT 70.450 152.900 70.770 152.960 ;
        RECT 77.365 152.900 77.655 152.945 ;
        RECT 70.450 152.760 77.655 152.900 ;
        RECT 70.450 152.700 70.770 152.760 ;
        RECT 77.365 152.715 77.655 152.760 ;
        RECT 5.520 152.080 84.180 152.560 ;
        RECT 19.390 151.880 19.710 151.940 ;
        RECT 18.100 151.740 19.710 151.880 ;
        RECT 14.790 151.340 15.110 151.600 ;
        RECT 18.100 151.585 18.240 151.740 ;
        RECT 19.390 151.680 19.710 151.740 ;
        RECT 26.305 151.880 26.595 151.925 ;
        RECT 26.750 151.880 27.070 151.940 ;
        RECT 27.670 151.880 27.990 151.940 ;
        RECT 26.305 151.740 27.990 151.880 ;
        RECT 26.305 151.695 26.595 151.740 ;
        RECT 26.750 151.680 27.070 151.740 ;
        RECT 27.670 151.680 27.990 151.740 ;
        RECT 42.390 151.880 42.710 151.940 ;
        RECT 49.750 151.880 50.070 151.940 ;
        RECT 54.365 151.880 54.655 151.925 ;
        RECT 64.010 151.880 64.330 151.940 ;
        RECT 66.770 151.880 67.090 151.940 ;
        RECT 42.390 151.740 45.380 151.880 ;
        RECT 42.390 151.680 42.710 151.740 ;
        RECT 15.885 151.540 16.175 151.585 ;
        RECT 17.105 151.540 17.395 151.585 ;
        RECT 15.885 151.400 17.395 151.540 ;
        RECT 15.885 151.355 16.175 151.400 ;
        RECT 17.105 151.355 17.395 151.400 ;
        RECT 18.025 151.355 18.315 151.585 ;
        RECT 18.470 151.540 18.790 151.600 ;
        RECT 18.945 151.540 19.235 151.585 ;
        RECT 23.530 151.540 23.850 151.600 ;
        RECT 18.470 151.400 19.235 151.540 ;
        RECT 18.470 151.340 18.790 151.400 ;
        RECT 18.945 151.355 19.235 151.400 ;
        RECT 19.480 151.400 23.850 151.540 ;
        RECT 19.480 151.245 19.620 151.400 ;
        RECT 23.530 151.340 23.850 151.400 ;
        RECT 31.810 151.540 32.130 151.600 ;
        RECT 31.810 151.400 43.540 151.540 ;
        RECT 31.810 151.340 32.130 151.400 ;
        RECT 19.405 151.015 19.695 151.245 ;
        RECT 20.685 151.200 20.975 151.245 ;
        RECT 19.940 151.060 20.975 151.200 ;
        RECT 19.940 150.860 20.080 151.060 ;
        RECT 20.685 151.015 20.975 151.060 ;
        RECT 41.470 151.200 41.790 151.260 ;
        RECT 43.400 151.245 43.540 151.400 ;
        RECT 45.240 151.245 45.380 151.740 ;
        RECT 49.750 151.740 54.655 151.880 ;
        RECT 49.750 151.680 50.070 151.740 ;
        RECT 54.365 151.695 54.655 151.740 ;
        RECT 62.720 151.740 63.780 151.880 ;
        RECT 62.720 151.585 62.860 151.740 ;
        RECT 62.645 151.355 62.935 151.585 ;
        RECT 63.090 151.340 63.410 151.600 ;
        RECT 63.640 151.540 63.780 151.740 ;
        RECT 64.010 151.740 67.090 151.880 ;
        RECT 64.010 151.680 64.330 151.740 ;
        RECT 66.770 151.680 67.090 151.740 ;
        RECT 65.850 151.540 66.170 151.600 ;
        RECT 67.545 151.540 67.835 151.585 ;
        RECT 63.640 151.400 67.835 151.540 ;
        RECT 65.850 151.340 66.170 151.400 ;
        RECT 67.545 151.355 67.835 151.400 ;
        RECT 68.625 151.540 68.915 151.585 ;
        RECT 70.450 151.540 70.770 151.600 ;
        RECT 68.625 151.400 70.770 151.540 ;
        RECT 68.625 151.355 68.915 151.400 ;
        RECT 42.405 151.200 42.695 151.245 ;
        RECT 41.470 151.060 42.695 151.200 ;
        RECT 41.470 151.000 41.790 151.060 ;
        RECT 42.405 151.015 42.695 151.060 ;
        RECT 43.325 151.200 43.615 151.245 ;
        RECT 44.705 151.200 44.995 151.245 ;
        RECT 43.325 151.060 44.995 151.200 ;
        RECT 43.325 151.015 43.615 151.060 ;
        RECT 44.705 151.015 44.995 151.060 ;
        RECT 45.165 151.015 45.455 151.245 ;
        RECT 45.610 151.200 45.930 151.260 ;
        RECT 46.085 151.200 46.375 151.245 ;
        RECT 45.610 151.060 46.375 151.200 ;
        RECT 16.720 150.720 20.080 150.860 ;
        RECT 20.285 150.860 20.575 150.905 ;
        RECT 21.475 150.860 21.765 150.905 ;
        RECT 23.995 150.860 24.285 150.905 ;
        RECT 20.285 150.720 24.285 150.860 ;
        RECT 42.480 150.860 42.620 151.015 ;
        RECT 45.240 150.860 45.380 151.015 ;
        RECT 45.610 151.000 45.930 151.060 ;
        RECT 46.085 151.015 46.375 151.060 ;
        RECT 46.990 151.000 47.310 151.260 ;
        RECT 48.385 151.200 48.675 151.245 ;
        RECT 49.290 151.200 49.610 151.260 ;
        RECT 48.385 151.060 49.610 151.200 ;
        RECT 48.385 151.015 48.675 151.060 ;
        RECT 49.290 151.000 49.610 151.060 ;
        RECT 55.270 151.000 55.590 151.260 ;
        RECT 56.205 151.200 56.495 151.245 ;
        RECT 56.650 151.200 56.970 151.260 ;
        RECT 56.205 151.060 56.970 151.200 ;
        RECT 56.205 151.015 56.495 151.060 ;
        RECT 56.650 151.000 56.970 151.060 ;
        RECT 58.950 151.200 59.270 151.260 ;
        RECT 59.425 151.200 59.715 151.245 ;
        RECT 58.950 151.060 59.715 151.200 ;
        RECT 58.950 151.000 59.270 151.060 ;
        RECT 59.425 151.015 59.715 151.060 ;
        RECT 60.345 151.200 60.635 151.245 ;
        RECT 60.790 151.200 61.110 151.260 ;
        RECT 60.345 151.060 61.110 151.200 ;
        RECT 60.345 151.015 60.635 151.060 ;
        RECT 47.465 150.860 47.755 150.905 ;
        RECT 42.480 150.720 44.920 150.860 ;
        RECT 45.240 150.720 47.755 150.860 ;
        RECT 59.500 150.860 59.640 151.015 ;
        RECT 60.790 151.000 61.110 151.060 ;
        RECT 62.170 151.200 62.490 151.260 ;
        RECT 63.565 151.200 63.855 151.245 ;
        RECT 68.700 151.200 68.840 151.355 ;
        RECT 70.450 151.340 70.770 151.400 ;
        RECT 62.170 151.060 68.840 151.200 ;
        RECT 62.170 151.000 62.490 151.060 ;
        RECT 63.565 151.015 63.855 151.060 ;
        RECT 69.085 151.015 69.375 151.245 ;
        RECT 69.545 151.200 69.835 151.245 ;
        RECT 72.290 151.200 72.610 151.260 ;
        RECT 69.545 151.060 72.610 151.200 ;
        RECT 69.545 151.015 69.835 151.060 ;
        RECT 65.850 150.860 66.170 150.920 ;
        RECT 68.610 150.860 68.930 150.920 ;
        RECT 69.160 150.860 69.300 151.015 ;
        RECT 59.500 150.720 64.700 150.860 ;
        RECT 16.720 150.565 16.860 150.720 ;
        RECT 20.285 150.675 20.575 150.720 ;
        RECT 21.475 150.675 21.765 150.720 ;
        RECT 23.995 150.675 24.285 150.720 ;
        RECT 16.645 150.335 16.935 150.565 ;
        RECT 19.890 150.520 20.180 150.565 ;
        RECT 21.990 150.520 22.280 150.565 ;
        RECT 23.560 150.520 23.850 150.565 ;
        RECT 19.890 150.380 23.850 150.520 ;
        RECT 19.890 150.335 20.180 150.380 ;
        RECT 21.990 150.335 22.280 150.380 ;
        RECT 23.560 150.335 23.850 150.380 ;
        RECT 28.130 150.520 28.450 150.580 ;
        RECT 31.350 150.520 31.670 150.580 ;
        RECT 44.780 150.520 44.920 150.720 ;
        RECT 47.465 150.675 47.755 150.720 ;
        RECT 45.625 150.520 45.915 150.565 ;
        RECT 46.530 150.520 46.850 150.580 ;
        RECT 47.910 150.520 48.230 150.580 ;
        RECT 62.170 150.520 62.490 150.580 ;
        RECT 64.560 150.565 64.700 150.720 ;
        RECT 65.850 150.720 69.300 150.860 ;
        RECT 65.850 150.660 66.170 150.720 ;
        RECT 68.610 150.660 68.930 150.720 ;
        RECT 28.130 150.380 44.460 150.520 ;
        RECT 44.780 150.380 46.850 150.520 ;
        RECT 28.130 150.320 28.450 150.380 ;
        RECT 31.350 150.320 31.670 150.380 ;
        RECT 15.710 149.980 16.030 150.240 ;
        RECT 42.390 149.980 42.710 150.240 ;
        RECT 43.770 149.980 44.090 150.240 ;
        RECT 44.320 150.180 44.460 150.380 ;
        RECT 45.625 150.335 45.915 150.380 ;
        RECT 46.530 150.320 46.850 150.380 ;
        RECT 47.080 150.380 48.230 150.520 ;
        RECT 47.080 150.225 47.220 150.380 ;
        RECT 47.910 150.320 48.230 150.380 ;
        RECT 60.420 150.380 62.490 150.520 ;
        RECT 47.005 150.180 47.295 150.225 ;
        RECT 44.320 150.040 47.295 150.180 ;
        RECT 47.005 149.995 47.295 150.040 ;
        RECT 47.450 150.180 47.770 150.240 ;
        RECT 49.305 150.180 49.595 150.225 ;
        RECT 47.450 150.040 49.595 150.180 ;
        RECT 47.450 149.980 47.770 150.040 ;
        RECT 49.305 149.995 49.595 150.040 ;
        RECT 56.190 149.980 56.510 150.240 ;
        RECT 57.110 150.180 57.430 150.240 ;
        RECT 60.420 150.225 60.560 150.380 ;
        RECT 62.170 150.320 62.490 150.380 ;
        RECT 64.485 150.520 64.775 150.565 ;
        RECT 68.150 150.520 68.470 150.580 ;
        RECT 64.485 150.380 68.470 150.520 ;
        RECT 64.485 150.335 64.775 150.380 ;
        RECT 68.150 150.320 68.470 150.380 ;
        RECT 58.505 150.180 58.795 150.225 ;
        RECT 57.110 150.040 58.795 150.180 ;
        RECT 57.110 149.980 57.430 150.040 ;
        RECT 58.505 149.995 58.795 150.040 ;
        RECT 60.345 149.995 60.635 150.225 ;
        RECT 61.710 149.980 62.030 150.240 ;
        RECT 63.090 150.180 63.410 150.240 ;
        RECT 67.705 150.180 67.995 150.225 ;
        RECT 69.620 150.180 69.760 151.015 ;
        RECT 72.290 151.000 72.610 151.060 ;
        RECT 69.990 150.520 70.310 150.580 ;
        RECT 70.465 150.520 70.755 150.565 ;
        RECT 69.990 150.380 70.755 150.520 ;
        RECT 69.990 150.320 70.310 150.380 ;
        RECT 70.465 150.335 70.755 150.380 ;
        RECT 63.090 150.040 69.760 150.180 ;
        RECT 63.090 149.980 63.410 150.040 ;
        RECT 67.705 149.995 67.995 150.040 ;
        RECT 5.520 149.360 84.180 149.840 ;
        RECT 42.390 148.960 42.710 149.220 ;
        RECT 52.050 149.160 52.370 149.220 ;
        RECT 56.190 149.160 56.510 149.220 ;
        RECT 56.665 149.160 56.955 149.205 ;
        RECT 52.050 149.020 55.960 149.160 ;
        RECT 52.050 148.960 52.370 149.020 ;
        RECT 11.610 148.820 11.900 148.865 ;
        RECT 13.710 148.820 14.000 148.865 ;
        RECT 15.280 148.820 15.570 148.865 ;
        RECT 11.610 148.680 15.570 148.820 ;
        RECT 11.610 148.635 11.900 148.680 ;
        RECT 13.710 148.635 14.000 148.680 ;
        RECT 15.280 148.635 15.570 148.680 ;
        RECT 29.525 148.820 29.815 148.865 ;
        RECT 46.990 148.820 47.310 148.880 ;
        RECT 55.820 148.820 55.960 149.020 ;
        RECT 56.190 149.020 56.955 149.160 ;
        RECT 56.190 148.960 56.510 149.020 ;
        RECT 56.665 148.975 56.955 149.020 ;
        RECT 64.470 148.820 64.790 148.880 ;
        RECT 65.850 148.820 66.170 148.880 ;
        RECT 29.525 148.680 37.560 148.820 ;
        RECT 29.525 148.635 29.815 148.680 ;
        RECT 12.005 148.480 12.295 148.525 ;
        RECT 13.195 148.480 13.485 148.525 ;
        RECT 15.715 148.480 16.005 148.525 ;
        RECT 12.005 148.340 16.005 148.480 ;
        RECT 12.005 148.295 12.295 148.340 ;
        RECT 13.195 148.295 13.485 148.340 ;
        RECT 15.715 148.295 16.005 148.340 ;
        RECT 18.470 148.480 18.790 148.540 ;
        RECT 23.530 148.480 23.850 148.540 ;
        RECT 29.050 148.480 29.370 148.540 ;
        RECT 18.470 148.340 21.460 148.480 ;
        RECT 18.470 148.280 18.790 148.340 ;
        RECT 11.110 147.940 11.430 148.200 ;
        RECT 21.320 148.185 21.460 148.340 ;
        RECT 23.530 148.340 25.145 148.480 ;
        RECT 23.530 148.280 23.850 148.340 ;
        RECT 25.005 148.185 25.145 148.340 ;
        RECT 25.920 148.340 29.370 148.480 ;
        RECT 25.920 148.185 26.060 148.340 ;
        RECT 29.050 148.280 29.370 148.340 ;
        RECT 19.865 147.955 20.155 148.185 ;
        RECT 21.245 147.955 21.535 148.185 ;
        RECT 24.465 147.955 24.755 148.185 ;
        RECT 24.930 147.955 25.220 148.185 ;
        RECT 25.845 147.955 26.135 148.185 ;
        RECT 26.995 148.140 27.285 148.185 ;
        RECT 29.600 148.140 29.740 148.635 ;
        RECT 33.665 148.295 33.955 148.525 ;
        RECT 26.995 148.000 29.740 148.140 ;
        RECT 26.995 147.955 27.285 148.000 ;
        RECT 12.490 147.845 12.810 147.860 ;
        RECT 12.460 147.615 12.810 147.845 ;
        RECT 19.940 147.800 20.080 147.955 ;
        RECT 24.540 147.800 24.680 147.955 ;
        RECT 30.890 147.940 31.210 148.200 ;
        RECT 31.350 147.940 31.670 148.200 ;
        RECT 31.810 148.140 32.130 148.200 ;
        RECT 33.205 148.140 33.495 148.185 ;
        RECT 31.810 148.000 33.495 148.140 ;
        RECT 33.740 148.140 33.880 148.295 ;
        RECT 35.030 148.280 35.350 148.540 ;
        RECT 37.420 148.525 37.560 148.680 ;
        RECT 42.480 148.680 47.310 148.820 ;
        RECT 42.480 148.525 42.620 148.680 ;
        RECT 46.990 148.620 47.310 148.680 ;
        RECT 51.680 148.680 55.500 148.820 ;
        RECT 55.820 148.680 66.170 148.820 ;
        RECT 37.345 148.295 37.635 148.525 ;
        RECT 42.405 148.295 42.695 148.525 ;
        RECT 43.770 148.480 44.090 148.540 ;
        RECT 48.845 148.480 49.135 148.525 ;
        RECT 43.770 148.340 49.135 148.480 ;
        RECT 43.770 148.280 44.090 148.340 ;
        RECT 48.845 148.295 49.135 148.340 ;
        RECT 34.110 148.140 34.430 148.200 ;
        RECT 36.870 148.140 37.190 148.200 ;
        RECT 33.740 148.000 37.190 148.140 ;
        RECT 31.810 147.940 32.130 148.000 ;
        RECT 33.205 147.955 33.495 148.000 ;
        RECT 34.110 147.940 34.430 148.000 ;
        RECT 36.870 147.940 37.190 148.000 ;
        RECT 37.805 148.140 38.095 148.185 ;
        RECT 37.805 148.000 42.620 148.140 ;
        RECT 37.805 147.955 38.095 148.000 ;
        RECT 12.490 147.600 12.810 147.615 ;
        RECT 18.100 147.660 24.680 147.800 ;
        RECT 26.305 147.800 26.595 147.845 ;
        RECT 26.305 147.660 26.980 147.800 ;
        RECT 18.100 147.520 18.240 147.660 ;
        RECT 26.305 147.615 26.595 147.660 ;
        RECT 26.840 147.520 26.980 147.660 ;
        RECT 41.485 147.615 41.775 147.845 ;
        RECT 42.480 147.800 42.620 148.000 ;
        RECT 42.850 147.940 43.170 148.200 ;
        RECT 45.165 148.140 45.455 148.185 ;
        RECT 43.400 148.000 45.455 148.140 ;
        RECT 43.400 147.860 43.540 148.000 ;
        RECT 45.165 147.955 45.455 148.000 ;
        RECT 47.450 147.940 47.770 148.200 ;
        RECT 50.685 148.140 50.975 148.185 ;
        RECT 51.680 148.140 51.820 148.680 ;
        RECT 52.050 148.280 52.370 148.540 ;
        RECT 53.430 148.185 53.750 148.200 ;
        RECT 50.685 148.000 51.820 148.140 ;
        RECT 50.685 147.955 50.975 148.000 ;
        RECT 52.525 147.955 52.815 148.185 ;
        RECT 53.265 147.955 53.750 148.185 ;
        RECT 43.310 147.800 43.630 147.860 ;
        RECT 51.130 147.800 51.450 147.860 ;
        RECT 52.600 147.800 52.740 147.955 ;
        RECT 53.430 147.940 53.750 147.955 ;
        RECT 53.890 147.940 54.210 148.200 ;
        RECT 54.850 147.955 55.140 148.185 ;
        RECT 55.360 148.140 55.500 148.680 ;
        RECT 64.470 148.620 64.790 148.680 ;
        RECT 65.850 148.620 66.170 148.680 ;
        RECT 67.705 148.480 67.995 148.525 ;
        RECT 66.860 148.340 67.995 148.480 ;
        RECT 55.360 148.000 55.960 148.140 ;
        RECT 42.480 147.660 43.630 147.800 ;
        RECT 18.010 147.260 18.330 147.520 ;
        RECT 18.930 147.260 19.250 147.520 ;
        RECT 19.390 147.460 19.710 147.520 ;
        RECT 20.785 147.460 21.075 147.505 ;
        RECT 26.750 147.460 27.070 147.520 ;
        RECT 19.390 147.320 27.070 147.460 ;
        RECT 19.390 147.260 19.710 147.320 ;
        RECT 20.785 147.275 21.075 147.320 ;
        RECT 26.750 147.260 27.070 147.320 ;
        RECT 27.670 147.260 27.990 147.520 ;
        RECT 39.645 147.460 39.935 147.505 ;
        RECT 41.560 147.460 41.700 147.615 ;
        RECT 43.310 147.600 43.630 147.660 ;
        RECT 43.860 147.660 52.740 147.800 ;
        RECT 43.860 147.505 44.000 147.660 ;
        RECT 51.130 147.600 51.450 147.660 ;
        RECT 54.350 147.600 54.670 147.860 ;
        RECT 39.645 147.320 41.700 147.460 ;
        RECT 39.645 147.275 39.935 147.320 ;
        RECT 43.785 147.275 44.075 147.505 ;
        RECT 45.630 147.460 45.920 147.505 ;
        RECT 52.070 147.460 52.360 147.505 ;
        RECT 45.630 147.320 52.360 147.460 ;
        RECT 45.630 147.275 45.920 147.320 ;
        RECT 52.070 147.275 52.360 147.320 ;
        RECT 52.970 147.460 53.290 147.520 ;
        RECT 54.900 147.460 55.040 147.955 ;
        RECT 55.820 147.505 55.960 148.000 ;
        RECT 56.205 147.955 56.495 148.185 ;
        RECT 57.125 148.140 57.415 148.185 ;
        RECT 59.870 148.140 60.190 148.200 ;
        RECT 57.125 148.000 60.190 148.140 ;
        RECT 57.125 147.955 57.415 148.000 ;
        RECT 56.280 147.800 56.420 147.955 ;
        RECT 59.870 147.940 60.190 148.000 ;
        RECT 61.710 148.140 62.030 148.200 ;
        RECT 66.860 148.185 67.000 148.340 ;
        RECT 67.705 148.295 67.995 148.340 ;
        RECT 65.865 148.140 66.155 148.185 ;
        RECT 61.710 148.000 66.155 148.140 ;
        RECT 61.710 147.940 62.030 148.000 ;
        RECT 65.865 147.955 66.155 148.000 ;
        RECT 66.785 147.955 67.075 148.185 ;
        RECT 67.230 147.940 67.550 148.200 ;
        RECT 68.150 148.140 68.470 148.200 ;
        RECT 74.130 148.140 74.450 148.200 ;
        RECT 68.150 148.000 74.450 148.140 ;
        RECT 68.150 147.940 68.470 148.000 ;
        RECT 74.130 147.940 74.450 148.000 ;
        RECT 58.030 147.800 58.350 147.860 ;
        RECT 60.790 147.800 61.110 147.860 ;
        RECT 56.280 147.660 61.110 147.800 ;
        RECT 58.030 147.600 58.350 147.660 ;
        RECT 60.790 147.600 61.110 147.660 ;
        RECT 52.970 147.320 55.040 147.460 ;
        RECT 52.970 147.260 53.290 147.320 ;
        RECT 55.745 147.275 56.035 147.505 ;
        RECT 64.470 147.460 64.790 147.520 ;
        RECT 66.325 147.460 66.615 147.505 ;
        RECT 64.470 147.320 66.615 147.460 ;
        RECT 64.470 147.260 64.790 147.320 ;
        RECT 66.325 147.275 66.615 147.320 ;
        RECT 5.520 146.640 84.180 147.120 ;
        RECT 12.490 146.240 12.810 146.500 ;
        RECT 13.425 146.440 13.715 146.485 ;
        RECT 14.790 146.440 15.110 146.500 ;
        RECT 13.425 146.300 15.110 146.440 ;
        RECT 13.425 146.255 13.715 146.300 ;
        RECT 14.790 146.240 15.110 146.300 ;
        RECT 17.025 146.440 17.315 146.485 ;
        RECT 18.470 146.440 18.790 146.500 ;
        RECT 17.025 146.300 18.790 146.440 ;
        RECT 17.025 146.255 17.315 146.300 ;
        RECT 18.470 146.240 18.790 146.300 ;
        RECT 23.530 146.440 23.850 146.500 ;
        RECT 31.810 146.440 32.130 146.500 ;
        RECT 41.945 146.440 42.235 146.485 ;
        RECT 23.530 146.300 31.580 146.440 ;
        RECT 23.530 146.240 23.850 146.300 ;
        RECT 18.010 145.900 18.330 146.160 ;
        RECT 27.670 146.100 27.990 146.160 ;
        RECT 25.460 145.960 27.990 146.100 ;
        RECT 31.440 146.100 31.580 146.300 ;
        RECT 31.810 146.300 42.235 146.440 ;
        RECT 31.810 146.240 32.130 146.300 ;
        RECT 41.945 146.255 42.235 146.300 ;
        RECT 43.785 146.440 44.075 146.485 ;
        RECT 46.990 146.440 47.310 146.500 ;
        RECT 43.785 146.300 47.310 146.440 ;
        RECT 43.785 146.255 44.075 146.300 ;
        RECT 46.990 146.240 47.310 146.300 ;
        RECT 52.970 146.240 53.290 146.500 ;
        RECT 53.430 146.240 53.750 146.500 ;
        RECT 64.930 146.440 65.250 146.500 ;
        RECT 65.405 146.440 65.695 146.485 ;
        RECT 64.930 146.300 65.695 146.440 ;
        RECT 64.930 146.240 65.250 146.300 ;
        RECT 65.405 146.255 65.695 146.300 ;
        RECT 66.785 146.255 67.075 146.485 ;
        RECT 57.110 146.100 57.430 146.160 ;
        RECT 31.440 145.960 41.240 146.100 ;
        RECT 23.990 145.560 24.310 145.820 ;
        RECT 24.450 145.760 24.770 145.820 ;
        RECT 25.460 145.805 25.600 145.960 ;
        RECT 27.670 145.900 27.990 145.960 ;
        RECT 24.925 145.760 25.215 145.805 ;
        RECT 24.450 145.620 25.215 145.760 ;
        RECT 24.450 145.560 24.770 145.620 ;
        RECT 24.925 145.575 25.215 145.620 ;
        RECT 25.385 145.575 25.675 145.805 ;
        RECT 26.750 145.560 27.070 145.820 ;
        RECT 35.950 145.760 36.270 145.820 ;
        RECT 37.390 145.760 37.680 145.805 ;
        RECT 35.950 145.620 37.680 145.760 ;
        RECT 41.100 145.760 41.240 145.960 ;
        RECT 55.820 145.960 57.430 146.100 ;
        RECT 41.470 145.760 41.790 145.820 ;
        RECT 41.100 145.620 41.790 145.760 ;
        RECT 35.950 145.560 36.270 145.620 ;
        RECT 37.390 145.575 37.680 145.620 ;
        RECT 41.470 145.560 41.790 145.620 ;
        RECT 42.390 145.760 42.710 145.820 ;
        RECT 42.865 145.760 43.155 145.805 ;
        RECT 42.390 145.620 43.155 145.760 ;
        RECT 42.390 145.560 42.710 145.620 ;
        RECT 42.865 145.575 43.155 145.620 ;
        RECT 51.130 145.560 51.450 145.820 ;
        RECT 52.065 145.760 52.355 145.805 ;
        RECT 52.970 145.760 53.290 145.820 ;
        RECT 55.820 145.805 55.960 145.960 ;
        RECT 57.110 145.900 57.430 145.960 ;
        RECT 57.585 145.915 57.875 146.145 ;
        RECT 58.490 146.100 58.810 146.160 ;
        RECT 61.265 146.100 61.555 146.145 ;
        RECT 63.550 146.100 63.870 146.160 ;
        RECT 58.490 145.960 59.640 146.100 ;
        RECT 54.825 145.760 55.115 145.805 ;
        RECT 52.065 145.620 55.115 145.760 ;
        RECT 52.065 145.575 52.355 145.620 ;
        RECT 52.970 145.560 53.290 145.620 ;
        RECT 54.825 145.575 55.115 145.620 ;
        RECT 55.285 145.575 55.575 145.805 ;
        RECT 55.745 145.575 56.035 145.805 ;
        RECT 56.665 145.760 56.955 145.805 ;
        RECT 57.660 145.760 57.800 145.915 ;
        RECT 58.490 145.900 58.810 145.960 ;
        RECT 56.665 145.620 57.800 145.760 ;
        RECT 56.665 145.575 56.955 145.620 ;
        RECT 25.940 145.420 26.230 145.465 ;
        RECT 27.210 145.420 27.530 145.480 ;
        RECT 25.940 145.280 27.530 145.420 ;
        RECT 25.940 145.235 26.230 145.280 ;
        RECT 27.210 145.220 27.530 145.280 ;
        RECT 34.135 145.420 34.425 145.465 ;
        RECT 36.655 145.420 36.945 145.465 ;
        RECT 37.845 145.420 38.135 145.465 ;
        RECT 34.135 145.280 38.135 145.420 ;
        RECT 34.135 145.235 34.425 145.280 ;
        RECT 36.655 145.235 36.945 145.280 ;
        RECT 37.845 145.235 38.135 145.280 ;
        RECT 38.710 145.220 39.030 145.480 ;
        RECT 51.220 145.420 51.360 145.560 ;
        RECT 55.360 145.420 55.500 145.575 ;
        RECT 58.950 145.560 59.270 145.820 ;
        RECT 59.500 145.805 59.640 145.960 ;
        RECT 59.960 145.960 61.555 146.100 ;
        RECT 59.960 145.820 60.100 145.960 ;
        RECT 61.265 145.915 61.555 145.960 ;
        RECT 62.720 145.960 63.870 146.100 ;
        RECT 66.860 146.100 67.000 146.255 ;
        RECT 74.130 146.240 74.450 146.500 ;
        RECT 68.470 146.100 68.760 146.145 ;
        RECT 66.860 145.960 68.760 146.100 ;
        RECT 59.425 145.575 59.715 145.805 ;
        RECT 59.870 145.560 60.190 145.820 ;
        RECT 60.790 145.560 61.110 145.820 ;
        RECT 62.720 145.805 62.860 145.960 ;
        RECT 63.550 145.900 63.870 145.960 ;
        RECT 68.470 145.915 68.760 145.960 ;
        RECT 62.640 145.575 62.930 145.805 ;
        RECT 63.105 145.575 63.395 145.805 ;
        RECT 64.010 145.760 64.330 145.820 ;
        RECT 64.945 145.760 65.235 145.805 ;
        RECT 65.390 145.760 65.710 145.820 ;
        RECT 64.010 145.620 65.710 145.760 ;
        RECT 51.220 145.280 55.500 145.420 ;
        RECT 60.330 145.420 60.650 145.480 ;
        RECT 63.180 145.420 63.320 145.575 ;
        RECT 64.010 145.560 64.330 145.620 ;
        RECT 64.945 145.575 65.235 145.620 ;
        RECT 65.390 145.560 65.710 145.620 ;
        RECT 60.330 145.280 63.320 145.420 ;
        RECT 60.330 145.220 60.650 145.280 ;
        RECT 63.550 145.220 63.870 145.480 ;
        RECT 64.470 145.420 64.790 145.480 ;
        RECT 65.990 145.420 66.280 145.465 ;
        RECT 64.470 145.280 66.280 145.420 ;
        RECT 64.470 145.220 64.790 145.280 ;
        RECT 65.990 145.235 66.280 145.280 ;
        RECT 67.230 145.220 67.550 145.480 ;
        RECT 68.125 145.420 68.415 145.465 ;
        RECT 69.315 145.420 69.605 145.465 ;
        RECT 71.835 145.420 72.125 145.465 ;
        RECT 68.125 145.280 72.125 145.420 ;
        RECT 68.125 145.235 68.415 145.280 ;
        RECT 69.315 145.235 69.605 145.280 ;
        RECT 71.835 145.235 72.125 145.280 ;
        RECT 15.265 145.080 15.555 145.125 ;
        RECT 16.170 145.080 16.490 145.140 ;
        RECT 18.930 145.080 19.250 145.140 ;
        RECT 15.265 144.940 16.490 145.080 ;
        RECT 15.265 144.895 15.555 144.940 ;
        RECT 16.170 144.880 16.490 144.940 ;
        RECT 16.720 144.940 19.250 145.080 ;
        RECT 13.425 144.740 13.715 144.785 ;
        RECT 16.720 144.740 16.860 144.940 ;
        RECT 18.930 144.880 19.250 144.940 ;
        RECT 24.465 145.080 24.755 145.125 ;
        RECT 33.650 145.080 33.970 145.140 ;
        RECT 24.465 144.940 33.970 145.080 ;
        RECT 24.465 144.895 24.755 144.940 ;
        RECT 33.650 144.880 33.970 144.940 ;
        RECT 34.570 145.080 34.860 145.125 ;
        RECT 36.140 145.080 36.430 145.125 ;
        RECT 38.240 145.080 38.530 145.125 ;
        RECT 34.570 144.940 38.530 145.080 ;
        RECT 34.570 144.895 34.860 144.940 ;
        RECT 36.140 144.895 36.430 144.940 ;
        RECT 38.240 144.895 38.530 144.940 ;
        RECT 67.730 145.080 68.020 145.125 ;
        RECT 69.830 145.080 70.120 145.125 ;
        RECT 71.400 145.080 71.690 145.125 ;
        RECT 67.730 144.940 71.690 145.080 ;
        RECT 67.730 144.895 68.020 144.940 ;
        RECT 69.830 144.895 70.120 144.940 ;
        RECT 71.400 144.895 71.690 144.940 ;
        RECT 13.425 144.600 16.860 144.740 ;
        RECT 17.105 144.740 17.395 144.785 ;
        RECT 19.390 144.740 19.710 144.800 ;
        RECT 17.105 144.600 19.710 144.740 ;
        RECT 13.425 144.555 13.715 144.600 ;
        RECT 17.105 144.555 17.395 144.600 ;
        RECT 19.390 144.540 19.710 144.600 ;
        RECT 5.520 143.920 84.180 144.400 ;
        RECT 22.625 143.720 22.915 143.765 ;
        RECT 23.990 143.720 24.310 143.780 ;
        RECT 22.625 143.580 24.310 143.720 ;
        RECT 22.625 143.535 22.915 143.580 ;
        RECT 23.990 143.520 24.310 143.580 ;
        RECT 29.050 143.720 29.370 143.780 ;
        RECT 30.905 143.720 31.195 143.765 ;
        RECT 29.050 143.580 31.195 143.720 ;
        RECT 29.050 143.520 29.370 143.580 ;
        RECT 30.905 143.535 31.195 143.580 ;
        RECT 35.950 143.520 36.270 143.780 ;
        RECT 51.130 143.720 51.450 143.780 ;
        RECT 52.525 143.720 52.815 143.765 ;
        RECT 53.445 143.720 53.735 143.765 ;
        RECT 51.130 143.580 53.735 143.720 ;
        RECT 51.130 143.520 51.450 143.580 ;
        RECT 52.525 143.535 52.815 143.580 ;
        RECT 53.445 143.535 53.735 143.580 ;
        RECT 55.270 143.720 55.590 143.780 ;
        RECT 55.745 143.720 56.035 143.765 ;
        RECT 55.270 143.580 56.035 143.720 ;
        RECT 55.270 143.520 55.590 143.580 ;
        RECT 55.745 143.535 56.035 143.580 ;
        RECT 21.230 143.380 21.550 143.440 ;
        RECT 26.750 143.380 27.070 143.440 ;
        RECT 39.170 143.380 39.490 143.440 ;
        RECT 21.230 143.240 27.070 143.380 ;
        RECT 21.230 143.180 21.550 143.240 ;
        RECT 26.750 143.180 27.070 143.240 ;
        RECT 34.660 143.240 39.490 143.380 ;
        RECT 34.660 143.100 34.800 143.240 ;
        RECT 39.170 143.180 39.490 143.240 ;
        RECT 66.770 143.380 67.090 143.440 ;
        RECT 68.165 143.380 68.455 143.425 ;
        RECT 70.465 143.380 70.755 143.425 ;
        RECT 66.770 143.240 70.755 143.380 ;
        RECT 66.770 143.180 67.090 143.240 ;
        RECT 68.165 143.195 68.455 143.240 ;
        RECT 70.465 143.195 70.755 143.240 ;
        RECT 19.850 143.040 20.170 143.100 ;
        RECT 19.850 142.900 26.060 143.040 ;
        RECT 19.850 142.840 20.170 142.900 ;
        RECT 20.310 142.500 20.630 142.760 ;
        RECT 21.230 142.500 21.550 142.760 ;
        RECT 21.690 142.700 22.010 142.760 ;
        RECT 23.530 142.700 23.850 142.760 ;
        RECT 25.000 142.745 25.140 142.900 ;
        RECT 21.690 142.560 23.850 142.700 ;
        RECT 21.690 142.500 22.010 142.560 ;
        RECT 23.530 142.500 23.850 142.560 ;
        RECT 24.925 142.515 25.215 142.745 ;
        RECT 25.385 142.515 25.675 142.745 ;
        RECT 25.460 142.360 25.600 142.515 ;
        RECT 24.540 142.220 25.600 142.360 ;
        RECT 25.920 142.360 26.060 142.900 ;
        RECT 34.570 142.840 34.890 143.100 ;
        RECT 35.030 143.085 35.350 143.100 ;
        RECT 35.030 142.855 35.460 143.085 ;
        RECT 63.565 143.040 63.855 143.085 ;
        RECT 67.230 143.040 67.550 143.100 ;
        RECT 63.565 142.900 67.550 143.040 ;
        RECT 63.565 142.855 63.855 142.900 ;
        RECT 35.030 142.840 35.350 142.855 ;
        RECT 28.605 142.700 28.895 142.745 ;
        RECT 31.365 142.700 31.655 142.745 ;
        RECT 28.605 142.560 31.655 142.700 ;
        RECT 28.605 142.515 28.895 142.560 ;
        RECT 31.365 142.515 31.655 142.560 ;
        RECT 32.745 142.700 33.035 142.745 ;
        RECT 41.010 142.700 41.330 142.760 ;
        RECT 32.745 142.560 41.330 142.700 ;
        RECT 32.745 142.515 33.035 142.560 ;
        RECT 41.010 142.500 41.330 142.560 ;
        RECT 51.145 142.515 51.435 142.745 ;
        RECT 51.605 142.700 51.895 142.745 ;
        RECT 52.510 142.700 52.830 142.760 ;
        RECT 51.605 142.560 52.830 142.700 ;
        RECT 51.605 142.515 51.895 142.560 ;
        RECT 29.065 142.360 29.355 142.405 ;
        RECT 25.920 142.220 29.355 142.360 ;
        RECT 18.470 142.020 18.790 142.080 ;
        RECT 20.785 142.020 21.075 142.065 ;
        RECT 18.470 141.880 21.075 142.020 ;
        RECT 18.470 141.820 18.790 141.880 ;
        RECT 20.785 141.835 21.075 141.880 ;
        RECT 23.990 142.020 24.310 142.080 ;
        RECT 24.540 142.065 24.680 142.220 ;
        RECT 29.065 142.175 29.355 142.220 ;
        RECT 29.985 142.175 30.275 142.405 ;
        RECT 34.125 142.360 34.415 142.405 ;
        RECT 39.630 142.360 39.950 142.420 ;
        RECT 41.930 142.360 42.250 142.420 ;
        RECT 34.125 142.220 42.250 142.360 ;
        RECT 51.220 142.360 51.360 142.515 ;
        RECT 52.510 142.500 52.830 142.560 ;
        RECT 52.970 142.500 53.290 142.760 ;
        RECT 54.825 142.700 55.115 142.745 ;
        RECT 57.570 142.700 57.890 142.760 ;
        RECT 54.825 142.560 57.890 142.700 ;
        RECT 54.825 142.515 55.115 142.560 ;
        RECT 57.570 142.500 57.890 142.560 ;
        RECT 58.965 142.700 59.255 142.745 ;
        RECT 63.640 142.700 63.780 142.855 ;
        RECT 67.230 142.840 67.550 142.900 ;
        RECT 58.965 142.560 62.170 142.700 ;
        RECT 58.965 142.515 59.255 142.560 ;
        RECT 62.030 142.420 62.170 142.560 ;
        RECT 53.430 142.360 53.750 142.420 ;
        RECT 51.220 142.220 53.750 142.360 ;
        RECT 34.125 142.175 34.415 142.220 ;
        RECT 24.465 142.020 24.755 142.065 ;
        RECT 30.060 142.020 30.200 142.175 ;
        RECT 39.630 142.160 39.950 142.220 ;
        RECT 41.930 142.160 42.250 142.220 ;
        RECT 53.430 142.160 53.750 142.220 ;
        RECT 57.110 142.360 57.430 142.420 ;
        RECT 59.410 142.360 59.730 142.420 ;
        RECT 57.110 142.220 59.730 142.360 ;
        RECT 57.110 142.160 57.430 142.220 ;
        RECT 59.410 142.160 59.730 142.220 ;
        RECT 61.710 142.360 62.170 142.420 ;
        RECT 62.720 142.560 63.780 142.700 ;
        RECT 62.720 142.360 62.860 142.560 ;
        RECT 65.850 142.500 66.170 142.760 ;
        RECT 69.070 142.700 69.390 142.760 ;
        RECT 71.385 142.700 71.675 142.745 ;
        RECT 69.070 142.560 71.675 142.700 ;
        RECT 69.070 142.500 69.390 142.560 ;
        RECT 71.385 142.515 71.675 142.560 ;
        RECT 61.710 142.220 62.860 142.360 ;
        RECT 63.090 142.360 63.410 142.420 ;
        RECT 65.405 142.360 65.695 142.405 ;
        RECT 67.690 142.360 68.010 142.420 ;
        RECT 63.090 142.220 68.010 142.360 ;
        RECT 61.710 142.160 62.030 142.220 ;
        RECT 63.090 142.160 63.410 142.220 ;
        RECT 65.405 142.175 65.695 142.220 ;
        RECT 67.690 142.160 68.010 142.220 ;
        RECT 68.165 142.360 68.455 142.405 ;
        RECT 68.610 142.360 68.930 142.420 ;
        RECT 68.165 142.220 68.930 142.360 ;
        RECT 68.165 142.175 68.455 142.220 ;
        RECT 68.610 142.160 68.930 142.220 ;
        RECT 23.990 141.880 30.200 142.020 ;
        RECT 31.350 142.020 31.670 142.080 ;
        RECT 31.825 142.020 32.115 142.065 ;
        RECT 31.350 141.880 32.115 142.020 ;
        RECT 23.990 141.820 24.310 141.880 ;
        RECT 24.465 141.835 24.755 141.880 ;
        RECT 31.350 141.820 31.670 141.880 ;
        RECT 31.825 141.835 32.115 141.880 ;
        RECT 64.470 141.820 64.790 142.080 ;
        RECT 5.520 141.200 84.180 141.680 ;
        RECT 15.265 141.000 15.555 141.045 ;
        RECT 18.010 141.000 18.330 141.060 ;
        RECT 20.310 141.000 20.630 141.060 ;
        RECT 15.265 140.860 20.630 141.000 ;
        RECT 15.265 140.815 15.555 140.860 ;
        RECT 18.010 140.800 18.330 140.860 ;
        RECT 20.310 140.800 20.630 140.860 ;
        RECT 43.310 141.000 43.630 141.060 ;
        RECT 43.785 141.000 44.075 141.045 ;
        RECT 43.310 140.860 44.075 141.000 ;
        RECT 43.310 140.800 43.630 140.860 ;
        RECT 43.785 140.815 44.075 140.860 ;
        RECT 52.065 141.000 52.355 141.045 ;
        RECT 52.970 141.000 53.290 141.060 ;
        RECT 52.065 140.860 53.290 141.000 ;
        RECT 52.065 140.815 52.355 140.860 ;
        RECT 52.970 140.800 53.290 140.860 ;
        RECT 57.570 140.800 57.890 141.060 ;
        RECT 68.610 141.000 68.930 141.060 ;
        RECT 69.085 141.000 69.375 141.045 ;
        RECT 68.610 140.860 69.375 141.000 ;
        RECT 68.610 140.800 68.930 140.860 ;
        RECT 69.085 140.815 69.375 140.860 ;
        RECT 21.230 140.660 21.550 140.720 ;
        RECT 19.940 140.520 21.550 140.660 ;
        RECT 16.170 140.320 16.490 140.380 ;
        RECT 17.565 140.320 17.855 140.365 ;
        RECT 16.170 140.180 17.855 140.320 ;
        RECT 16.170 140.120 16.490 140.180 ;
        RECT 17.565 140.135 17.855 140.180 ;
        RECT 18.485 140.320 18.775 140.365 ;
        RECT 19.390 140.320 19.710 140.380 ;
        RECT 19.940 140.365 20.080 140.520 ;
        RECT 21.230 140.460 21.550 140.520 ;
        RECT 23.545 140.660 23.835 140.705 ;
        RECT 26.290 140.660 26.610 140.720 ;
        RECT 31.350 140.660 31.670 140.720 ;
        RECT 38.710 140.660 39.030 140.720 ;
        RECT 42.390 140.660 42.710 140.720 ;
        RECT 23.545 140.520 26.610 140.660 ;
        RECT 23.545 140.475 23.835 140.520 ;
        RECT 26.290 140.460 26.610 140.520 ;
        RECT 30.520 140.520 31.670 140.660 ;
        RECT 18.485 140.180 19.710 140.320 ;
        RECT 18.485 140.135 18.775 140.180 ;
        RECT 17.105 139.980 17.395 140.025 ;
        RECT 18.560 139.980 18.700 140.135 ;
        RECT 19.390 140.120 19.710 140.180 ;
        RECT 19.865 140.135 20.155 140.365 ;
        RECT 17.105 139.840 18.700 139.980 ;
        RECT 18.930 139.980 19.250 140.040 ;
        RECT 19.940 139.980 20.080 140.135 ;
        RECT 21.690 140.120 22.010 140.380 ;
        RECT 30.520 140.365 30.660 140.520 ;
        RECT 31.350 140.460 31.670 140.520 ;
        RECT 31.900 140.520 39.030 140.660 ;
        RECT 31.900 140.380 32.040 140.520 ;
        RECT 38.710 140.460 39.030 140.520 ;
        RECT 40.640 140.520 42.710 140.660 ;
        RECT 22.165 140.320 22.455 140.365 ;
        RECT 30.445 140.320 30.735 140.365 ;
        RECT 22.165 140.180 30.735 140.320 ;
        RECT 22.165 140.135 22.455 140.180 ;
        RECT 30.445 140.135 30.735 140.180 ;
        RECT 30.905 140.135 31.195 140.365 ;
        RECT 18.930 139.840 20.080 139.980 ;
        RECT 23.070 139.980 23.390 140.040 ;
        RECT 27.225 139.980 27.515 140.025 ;
        RECT 23.070 139.840 27.515 139.980 ;
        RECT 17.105 139.795 17.395 139.840 ;
        RECT 18.930 139.780 19.250 139.840 ;
        RECT 23.070 139.780 23.390 139.840 ;
        RECT 27.225 139.795 27.515 139.840 ;
        RECT 28.590 139.780 28.910 140.040 ;
        RECT 18.470 139.640 18.790 139.700 ;
        RECT 30.980 139.640 31.120 140.135 ;
        RECT 31.810 140.120 32.130 140.380 ;
        RECT 33.650 140.320 33.970 140.380 ;
        RECT 35.505 140.320 35.795 140.365 ;
        RECT 33.650 140.180 35.795 140.320 ;
        RECT 33.650 140.120 33.970 140.180 ;
        RECT 35.505 140.135 35.795 140.180 ;
        RECT 36.870 140.320 37.190 140.380 ;
        RECT 40.640 140.365 40.780 140.520 ;
        RECT 42.390 140.460 42.710 140.520 ;
        RECT 42.865 140.660 43.155 140.705 ;
        RECT 51.590 140.660 51.910 140.720 ;
        RECT 63.520 140.660 63.810 140.705 ;
        RECT 64.470 140.660 64.790 140.720 ;
        RECT 42.865 140.520 51.360 140.660 ;
        RECT 42.865 140.475 43.155 140.520 ;
        RECT 36.870 140.180 37.560 140.320 ;
        RECT 36.870 140.120 37.190 140.180 ;
        RECT 18.470 139.500 31.120 139.640 ;
        RECT 37.420 139.640 37.560 140.180 ;
        RECT 37.805 140.135 38.095 140.365 ;
        RECT 40.565 140.135 40.855 140.365 ;
        RECT 37.880 139.980 38.020 140.135 ;
        RECT 41.470 140.120 41.790 140.380 ;
        RECT 49.290 140.365 49.610 140.380 ;
        RECT 49.290 140.135 49.640 140.365 ;
        RECT 51.220 140.320 51.360 140.520 ;
        RECT 51.590 140.520 59.180 140.660 ;
        RECT 51.590 140.460 51.910 140.520 ;
        RECT 52.050 140.320 52.370 140.380 ;
        RECT 51.220 140.180 52.370 140.320 ;
        RECT 49.290 140.120 49.610 140.135 ;
        RECT 52.050 140.120 52.370 140.180 ;
        RECT 52.510 140.320 52.830 140.380 ;
        RECT 52.985 140.320 53.275 140.365 ;
        RECT 52.510 140.180 53.275 140.320 ;
        RECT 52.510 140.120 52.830 140.180 ;
        RECT 52.985 140.135 53.275 140.180 ;
        RECT 53.430 140.120 53.750 140.380 ;
        RECT 54.900 140.365 55.040 140.520 ;
        RECT 54.825 140.135 55.115 140.365 ;
        RECT 58.490 140.120 58.810 140.380 ;
        RECT 41.025 139.980 41.315 140.025 ;
        RECT 37.880 139.840 41.315 139.980 ;
        RECT 41.025 139.795 41.315 139.840 ;
        RECT 46.095 139.980 46.385 140.025 ;
        RECT 48.615 139.980 48.905 140.025 ;
        RECT 49.805 139.980 50.095 140.025 ;
        RECT 46.095 139.840 50.095 139.980 ;
        RECT 46.095 139.795 46.385 139.840 ;
        RECT 48.615 139.795 48.905 139.840 ;
        RECT 49.805 139.795 50.095 139.840 ;
        RECT 50.670 139.780 50.990 140.040 ;
        RECT 54.365 139.980 54.655 140.025 ;
        RECT 58.580 139.980 58.720 140.120 ;
        RECT 54.365 139.840 58.720 139.980 ;
        RECT 59.040 139.980 59.180 140.520 ;
        RECT 63.520 140.520 64.790 140.660 ;
        RECT 63.520 140.475 63.810 140.520 ;
        RECT 64.470 140.460 64.790 140.520 ;
        RECT 59.425 140.320 59.715 140.365 ;
        RECT 60.330 140.320 60.650 140.380 ;
        RECT 59.425 140.180 60.650 140.320 ;
        RECT 59.425 140.135 59.715 140.180 ;
        RECT 60.330 140.120 60.650 140.180 ;
        RECT 59.885 139.980 60.175 140.025 ;
        RECT 59.040 139.840 60.175 139.980 ;
        RECT 54.365 139.795 54.655 139.840 ;
        RECT 59.885 139.795 60.175 139.840 ;
        RECT 61.710 139.980 62.030 140.040 ;
        RECT 62.185 139.980 62.475 140.025 ;
        RECT 61.710 139.840 62.475 139.980 ;
        RECT 61.710 139.780 62.030 139.840 ;
        RECT 62.185 139.795 62.475 139.840 ;
        RECT 63.065 139.980 63.355 140.025 ;
        RECT 64.255 139.980 64.545 140.025 ;
        RECT 66.775 139.980 67.065 140.025 ;
        RECT 63.065 139.840 67.065 139.980 ;
        RECT 63.065 139.795 63.355 139.840 ;
        RECT 64.255 139.795 64.545 139.840 ;
        RECT 66.775 139.795 67.065 139.840 ;
        RECT 41.930 139.640 42.250 139.700 ;
        RECT 37.420 139.500 42.250 139.640 ;
        RECT 18.470 139.440 18.790 139.500 ;
        RECT 41.930 139.440 42.250 139.500 ;
        RECT 46.530 139.640 46.820 139.685 ;
        RECT 48.100 139.640 48.390 139.685 ;
        RECT 50.200 139.640 50.490 139.685 ;
        RECT 46.530 139.500 50.490 139.640 ;
        RECT 46.530 139.455 46.820 139.500 ;
        RECT 48.100 139.455 48.390 139.500 ;
        RECT 50.200 139.455 50.490 139.500 ;
        RECT 62.670 139.640 62.960 139.685 ;
        RECT 64.770 139.640 65.060 139.685 ;
        RECT 66.340 139.640 66.630 139.685 ;
        RECT 62.670 139.500 66.630 139.640 ;
        RECT 62.670 139.455 62.960 139.500 ;
        RECT 64.770 139.455 65.060 139.500 ;
        RECT 66.340 139.455 66.630 139.500 ;
        RECT 19.390 139.100 19.710 139.360 ;
        RECT 19.850 139.300 20.170 139.360 ;
        RECT 20.325 139.300 20.615 139.345 ;
        RECT 19.850 139.160 20.615 139.300 ;
        RECT 19.850 139.100 20.170 139.160 ;
        RECT 20.325 139.115 20.615 139.160 ;
        RECT 23.085 139.300 23.375 139.345 ;
        RECT 23.530 139.300 23.850 139.360 ;
        RECT 23.085 139.160 23.850 139.300 ;
        RECT 23.085 139.115 23.375 139.160 ;
        RECT 23.530 139.100 23.850 139.160 ;
        RECT 29.525 139.300 29.815 139.345 ;
        RECT 31.350 139.300 31.670 139.360 ;
        RECT 29.525 139.160 31.670 139.300 ;
        RECT 29.525 139.115 29.815 139.160 ;
        RECT 31.350 139.100 31.670 139.160 ;
        RECT 34.570 139.100 34.890 139.360 ;
        RECT 37.790 139.100 38.110 139.360 ;
        RECT 39.630 139.300 39.950 139.360 ;
        RECT 42.405 139.300 42.695 139.345 ;
        RECT 45.610 139.300 45.930 139.360 ;
        RECT 39.630 139.160 45.930 139.300 ;
        RECT 39.630 139.100 39.950 139.160 ;
        RECT 42.405 139.115 42.695 139.160 ;
        RECT 45.610 139.100 45.930 139.160 ;
        RECT 5.520 138.480 84.180 138.960 ;
        RECT 18.025 138.280 18.315 138.325 ;
        RECT 19.850 138.280 20.170 138.340 ;
        RECT 28.590 138.280 28.910 138.340 ;
        RECT 18.025 138.140 20.170 138.280 ;
        RECT 18.025 138.095 18.315 138.140 ;
        RECT 19.850 138.080 20.170 138.140 ;
        RECT 20.400 138.140 28.910 138.280 ;
        RECT 20.400 138.000 20.540 138.140 ;
        RECT 28.590 138.080 28.910 138.140 ;
        RECT 41.025 138.280 41.315 138.325 ;
        RECT 42.390 138.280 42.710 138.340 ;
        RECT 41.025 138.140 42.710 138.280 ;
        RECT 41.025 138.095 41.315 138.140 ;
        RECT 42.390 138.080 42.710 138.140 ;
        RECT 42.865 138.280 43.155 138.325 ;
        RECT 47.450 138.280 47.770 138.340 ;
        RECT 49.290 138.280 49.610 138.340 ;
        RECT 42.865 138.140 47.770 138.280 ;
        RECT 42.865 138.095 43.155 138.140 ;
        RECT 47.450 138.080 47.770 138.140 ;
        RECT 48.000 138.140 49.610 138.280 ;
        RECT 11.610 137.940 11.900 137.985 ;
        RECT 13.710 137.940 14.000 137.985 ;
        RECT 15.280 137.940 15.570 137.985 ;
        RECT 11.610 137.800 15.570 137.940 ;
        RECT 11.610 137.755 11.900 137.800 ;
        RECT 13.710 137.755 14.000 137.800 ;
        RECT 15.280 137.755 15.570 137.800 ;
        RECT 20.310 137.740 20.630 138.000 ;
        RECT 23.990 137.940 24.280 137.985 ;
        RECT 25.560 137.940 25.850 137.985 ;
        RECT 27.660 137.940 27.950 137.985 ;
        RECT 23.990 137.800 27.950 137.940 ;
        RECT 23.990 137.755 24.280 137.800 ;
        RECT 25.560 137.755 25.850 137.800 ;
        RECT 27.660 137.755 27.950 137.800 ;
        RECT 34.610 137.940 34.900 137.985 ;
        RECT 36.710 137.940 37.000 137.985 ;
        RECT 38.280 137.940 38.570 137.985 ;
        RECT 34.610 137.800 38.570 137.940 ;
        RECT 34.610 137.755 34.900 137.800 ;
        RECT 36.710 137.755 37.000 137.800 ;
        RECT 38.280 137.755 38.570 137.800 ;
        RECT 41.470 137.940 41.790 138.000 ;
        RECT 43.785 137.940 44.075 137.985 ;
        RECT 44.690 137.940 45.010 138.000 ;
        RECT 48.000 137.985 48.140 138.140 ;
        RECT 49.290 138.080 49.610 138.140 ;
        RECT 41.470 137.800 45.010 137.940 ;
        RECT 41.470 137.740 41.790 137.800 ;
        RECT 43.785 137.755 44.075 137.800 ;
        RECT 44.690 137.740 45.010 137.800 ;
        RECT 45.240 137.800 47.680 137.940 ;
        RECT 11.110 137.400 11.430 137.660 ;
        RECT 12.005 137.600 12.295 137.645 ;
        RECT 13.195 137.600 13.485 137.645 ;
        RECT 15.715 137.600 16.005 137.645 ;
        RECT 12.005 137.460 16.005 137.600 ;
        RECT 12.005 137.415 12.295 137.460 ;
        RECT 13.195 137.415 13.485 137.460 ;
        RECT 15.715 137.415 16.005 137.460 ;
        RECT 23.555 137.600 23.845 137.645 ;
        RECT 26.075 137.600 26.365 137.645 ;
        RECT 27.265 137.600 27.555 137.645 ;
        RECT 31.810 137.600 32.130 137.660 ;
        RECT 34.125 137.600 34.415 137.645 ;
        RECT 23.555 137.460 27.555 137.600 ;
        RECT 23.555 137.415 23.845 137.460 ;
        RECT 26.075 137.415 26.365 137.460 ;
        RECT 27.265 137.415 27.555 137.460 ;
        RECT 29.140 137.460 34.415 137.600 ;
        RECT 11.200 137.260 11.340 137.400 ;
        RECT 29.140 137.320 29.280 137.460 ;
        RECT 31.810 137.400 32.130 137.460 ;
        RECT 34.125 137.415 34.415 137.460 ;
        RECT 35.005 137.600 35.295 137.645 ;
        RECT 36.195 137.600 36.485 137.645 ;
        RECT 38.715 137.600 39.005 137.645 ;
        RECT 43.310 137.600 43.630 137.660 ;
        RECT 45.240 137.600 45.380 137.800 ;
        RECT 35.005 137.460 39.005 137.600 ;
        RECT 35.005 137.415 35.295 137.460 ;
        RECT 36.195 137.415 36.485 137.460 ;
        RECT 38.715 137.415 39.005 137.460 ;
        RECT 42.020 137.460 43.630 137.600 ;
        RECT 15.250 137.260 15.570 137.320 ;
        RECT 23.070 137.260 23.390 137.320 ;
        RECT 11.200 137.120 23.390 137.260 ;
        RECT 15.250 137.060 15.570 137.120 ;
        RECT 23.070 137.060 23.390 137.120 ;
        RECT 28.145 137.260 28.435 137.305 ;
        RECT 29.050 137.260 29.370 137.320 ;
        RECT 28.145 137.120 29.370 137.260 ;
        RECT 28.145 137.075 28.435 137.120 ;
        RECT 29.050 137.060 29.370 137.120 ;
        RECT 31.350 137.060 31.670 137.320 ;
        RECT 12.460 136.920 12.750 136.965 ;
        RECT 13.410 136.920 13.730 136.980 ;
        RECT 12.460 136.780 13.730 136.920 ;
        RECT 12.460 136.735 12.750 136.780 ;
        RECT 13.410 136.720 13.730 136.780 ;
        RECT 17.550 136.920 17.870 136.980 ;
        RECT 19.865 136.920 20.155 136.965 ;
        RECT 17.550 136.780 20.155 136.920 ;
        RECT 17.550 136.720 17.870 136.780 ;
        RECT 19.865 136.735 20.155 136.780 ;
        RECT 26.920 136.920 27.210 136.965 ;
        RECT 28.605 136.920 28.895 136.965 ;
        RECT 26.920 136.780 28.895 136.920 ;
        RECT 26.920 136.735 27.210 136.780 ;
        RECT 28.605 136.735 28.895 136.780 ;
        RECT 35.460 136.920 35.750 136.965 ;
        RECT 37.330 136.920 37.650 136.980 ;
        RECT 42.020 136.965 42.160 137.460 ;
        RECT 43.310 137.400 43.630 137.460 ;
        RECT 44.320 137.460 45.380 137.600 ;
        RECT 47.540 137.600 47.680 137.800 ;
        RECT 47.925 137.755 48.215 137.985 ;
        RECT 48.370 137.740 48.690 138.000 ;
        RECT 47.540 137.460 49.980 137.600 ;
        RECT 42.850 136.965 43.170 136.980 ;
        RECT 35.460 136.780 37.650 136.920 ;
        RECT 35.460 136.735 35.750 136.780 ;
        RECT 37.330 136.720 37.650 136.780 ;
        RECT 41.945 136.735 42.235 136.965 ;
        RECT 42.850 136.920 43.315 136.965 ;
        RECT 44.320 136.920 44.460 137.460 ;
        RECT 44.705 137.075 44.995 137.305 ;
        RECT 45.610 137.260 45.930 137.320 ;
        RECT 46.085 137.260 46.375 137.305 ;
        RECT 46.530 137.260 46.850 137.320 ;
        RECT 49.840 137.305 49.980 137.460 ;
        RECT 50.670 137.400 50.990 137.660 ;
        RECT 53.890 137.600 54.210 137.660 ;
        RECT 56.665 137.600 56.955 137.645 ;
        RECT 51.220 137.460 56.955 137.600 ;
        RECT 45.610 137.120 46.850 137.260 ;
        RECT 42.850 136.780 44.460 136.920 ;
        RECT 42.850 136.735 43.315 136.780 ;
        RECT 42.850 136.720 43.170 136.735 ;
        RECT 14.790 136.580 15.110 136.640 ;
        RECT 20.310 136.580 20.630 136.640 ;
        RECT 14.790 136.440 20.630 136.580 ;
        RECT 14.790 136.380 15.110 136.440 ;
        RECT 20.310 136.380 20.630 136.440 ;
        RECT 21.245 136.580 21.535 136.625 ;
        RECT 23.990 136.580 24.310 136.640 ;
        RECT 21.245 136.440 24.310 136.580 ;
        RECT 21.245 136.395 21.535 136.440 ;
        RECT 23.990 136.380 24.310 136.440 ;
        RECT 41.010 136.580 41.330 136.640 ;
        RECT 44.780 136.580 44.920 137.075 ;
        RECT 45.610 137.060 45.930 137.120 ;
        RECT 46.085 137.075 46.375 137.120 ;
        RECT 46.530 137.060 46.850 137.120 ;
        RECT 49.765 137.260 50.055 137.305 ;
        RECT 51.220 137.260 51.360 137.460 ;
        RECT 53.890 137.400 54.210 137.460 ;
        RECT 56.665 137.415 56.955 137.460 ;
        RECT 49.765 137.120 51.360 137.260 ;
        RECT 55.730 137.260 56.050 137.320 ;
        RECT 58.490 137.260 58.810 137.320 ;
        RECT 59.425 137.260 59.715 137.305 ;
        RECT 55.730 137.120 59.715 137.260 ;
        RECT 49.765 137.075 50.055 137.120 ;
        RECT 55.730 137.060 56.050 137.120 ;
        RECT 58.490 137.060 58.810 137.120 ;
        RECT 59.425 137.075 59.715 137.120 ;
        RECT 45.150 136.920 45.470 136.980 ;
        RECT 47.130 136.920 47.420 136.965 ;
        RECT 45.150 136.780 47.420 136.920 ;
        RECT 45.150 136.720 45.470 136.780 ;
        RECT 47.130 136.735 47.420 136.780 ;
        RECT 47.910 136.920 48.230 136.980 ;
        RECT 48.385 136.920 48.675 136.965 ;
        RECT 47.910 136.780 48.675 136.920 ;
        RECT 47.910 136.720 48.230 136.780 ;
        RECT 48.385 136.735 48.675 136.780 ;
        RECT 51.130 136.920 51.450 136.980 ;
        RECT 54.825 136.920 55.115 136.965 ;
        RECT 57.110 136.920 57.430 136.980 ;
        RECT 51.130 136.780 57.430 136.920 ;
        RECT 51.130 136.720 51.450 136.780 ;
        RECT 54.825 136.735 55.115 136.780 ;
        RECT 57.110 136.720 57.430 136.780 ;
        RECT 57.585 136.920 57.875 136.965 ;
        RECT 58.950 136.920 59.270 136.980 ;
        RECT 61.250 136.920 61.570 136.980 ;
        RECT 57.585 136.780 61.570 136.920 ;
        RECT 57.585 136.735 57.875 136.780 ;
        RECT 58.950 136.720 59.270 136.780 ;
        RECT 61.250 136.720 61.570 136.780 ;
        RECT 41.010 136.440 44.920 136.580 ;
        RECT 41.010 136.380 41.330 136.440 ;
        RECT 46.530 136.380 46.850 136.640 ;
        RECT 48.830 136.580 49.150 136.640 ;
        RECT 49.305 136.580 49.595 136.625 ;
        RECT 52.970 136.580 53.290 136.640 ;
        RECT 48.830 136.440 53.290 136.580 ;
        RECT 48.830 136.380 49.150 136.440 ;
        RECT 49.305 136.395 49.595 136.440 ;
        RECT 52.970 136.380 53.290 136.440 ;
        RECT 58.030 136.380 58.350 136.640 ;
        RECT 58.505 136.580 58.795 136.625 ;
        RECT 60.330 136.580 60.650 136.640 ;
        RECT 58.505 136.440 60.650 136.580 ;
        RECT 58.505 136.395 58.795 136.440 ;
        RECT 60.330 136.380 60.650 136.440 ;
        RECT 5.520 135.760 84.180 136.240 ;
        RECT 13.410 135.360 13.730 135.620 ;
        RECT 14.345 135.560 14.635 135.605 ;
        RECT 14.790 135.560 15.110 135.620 ;
        RECT 14.345 135.420 15.110 135.560 ;
        RECT 14.345 135.375 14.635 135.420 ;
        RECT 14.790 135.360 15.110 135.420 ;
        RECT 19.865 135.560 20.155 135.605 ;
        RECT 21.325 135.560 21.615 135.605 ;
        RECT 19.865 135.420 21.615 135.560 ;
        RECT 19.865 135.375 20.155 135.420 ;
        RECT 21.325 135.375 21.615 135.420 ;
        RECT 22.165 135.375 22.455 135.605 ;
        RECT 37.330 135.560 37.650 135.620 ;
        RECT 37.805 135.560 38.095 135.605 ;
        RECT 37.330 135.420 38.095 135.560 ;
        RECT 18.010 135.220 18.330 135.280 ;
        RECT 16.260 135.080 18.330 135.220 ;
        RECT 16.260 134.925 16.400 135.080 ;
        RECT 18.010 135.020 18.330 135.080 ;
        RECT 20.310 135.020 20.630 135.280 ;
        RECT 22.240 135.220 22.380 135.375 ;
        RECT 37.330 135.360 37.650 135.420 ;
        RECT 37.805 135.375 38.095 135.420 ;
        RECT 39.170 135.360 39.490 135.620 ;
        RECT 39.630 135.360 39.950 135.620 ;
        RECT 41.485 135.560 41.775 135.605 ;
        RECT 41.930 135.560 42.250 135.620 ;
        RECT 41.485 135.420 42.250 135.560 ;
        RECT 41.485 135.375 41.775 135.420 ;
        RECT 41.930 135.360 42.250 135.420 ;
        RECT 42.390 135.560 42.710 135.620 ;
        RECT 43.325 135.560 43.615 135.605 ;
        RECT 42.390 135.420 43.615 135.560 ;
        RECT 42.390 135.360 42.710 135.420 ;
        RECT 43.325 135.375 43.615 135.420 ;
        RECT 45.150 135.360 45.470 135.620 ;
        RECT 52.050 135.560 52.370 135.620 ;
        RECT 63.090 135.560 63.410 135.620 ;
        RECT 64.025 135.560 64.315 135.605 ;
        RECT 52.050 135.420 64.315 135.560 ;
        RECT 52.050 135.360 52.370 135.420 ;
        RECT 63.090 135.360 63.410 135.420 ;
        RECT 64.025 135.375 64.315 135.420 ;
        RECT 65.405 135.375 65.695 135.605 ;
        RECT 23.850 135.220 24.140 135.265 ;
        RECT 22.240 135.080 24.140 135.220 ;
        RECT 23.850 135.035 24.140 135.080 ;
        RECT 27.670 135.220 27.990 135.280 ;
        RECT 32.745 135.220 33.035 135.265 ;
        RECT 51.130 135.220 51.450 135.280 ;
        RECT 27.670 135.080 51.450 135.220 ;
        RECT 27.670 135.020 27.990 135.080 ;
        RECT 32.745 135.035 33.035 135.080 ;
        RECT 51.130 135.020 51.450 135.080 ;
        RECT 53.430 135.220 53.750 135.280 ;
        RECT 62.170 135.220 62.490 135.280 ;
        RECT 63.550 135.220 63.870 135.280 ;
        RECT 53.430 135.080 63.870 135.220 ;
        RECT 65.480 135.220 65.620 135.375 ;
        RECT 71.430 135.220 71.720 135.265 ;
        RECT 65.480 135.080 71.720 135.220 ;
        RECT 53.430 135.020 53.750 135.080 ;
        RECT 62.170 135.020 62.490 135.080 ;
        RECT 63.550 135.020 63.870 135.080 ;
        RECT 71.430 135.035 71.720 135.080 ;
        RECT 8.365 134.880 8.655 134.925 ;
        RECT 8.365 134.740 13.870 134.880 ;
        RECT 8.365 134.695 8.655 134.740 ;
        RECT 13.730 134.540 13.870 134.740 ;
        RECT 16.185 134.695 16.475 134.925 ;
        RECT 18.930 134.880 19.250 134.940 ;
        RECT 22.625 134.880 22.915 134.925 ;
        RECT 23.070 134.880 23.390 134.940 ;
        RECT 18.930 134.740 22.380 134.880 ;
        RECT 18.930 134.680 19.250 134.740 ;
        RECT 20.310 134.540 20.630 134.600 ;
        RECT 13.730 134.400 20.630 134.540 ;
        RECT 20.310 134.340 20.630 134.400 ;
        RECT 18.470 134.200 18.790 134.260 ;
        RECT 18.470 134.060 21.460 134.200 ;
        RECT 18.470 134.000 18.790 134.060 ;
        RECT 4.210 133.860 4.530 133.920 ;
        RECT 7.445 133.860 7.735 133.905 ;
        RECT 4.210 133.720 7.735 133.860 ;
        RECT 4.210 133.660 4.530 133.720 ;
        RECT 7.445 133.675 7.735 133.720 ;
        RECT 14.345 133.860 14.635 133.905 ;
        RECT 19.390 133.860 19.710 133.920 ;
        RECT 21.320 133.905 21.460 134.060 ;
        RECT 14.345 133.720 19.710 133.860 ;
        RECT 14.345 133.675 14.635 133.720 ;
        RECT 19.390 133.660 19.710 133.720 ;
        RECT 21.245 133.675 21.535 133.905 ;
        RECT 22.240 133.860 22.380 134.740 ;
        RECT 22.625 134.740 23.390 134.880 ;
        RECT 22.625 134.695 22.915 134.740 ;
        RECT 23.070 134.680 23.390 134.740 ;
        RECT 37.790 134.880 38.110 134.940 ;
        RECT 38.600 134.880 38.890 134.925 ;
        RECT 37.790 134.740 38.890 134.880 ;
        RECT 37.790 134.680 38.110 134.740 ;
        RECT 38.600 134.695 38.890 134.740 ;
        RECT 42.390 134.680 42.710 134.940 ;
        RECT 42.865 134.695 43.155 134.925 ;
        RECT 43.310 134.880 43.630 134.940 ;
        RECT 44.245 134.880 44.535 134.925 ;
        RECT 43.310 134.740 44.535 134.880 ;
        RECT 23.505 134.540 23.795 134.585 ;
        RECT 24.695 134.540 24.985 134.585 ;
        RECT 27.215 134.540 27.505 134.585 ;
        RECT 23.505 134.400 27.505 134.540 ;
        RECT 23.505 134.355 23.795 134.400 ;
        RECT 24.695 134.355 24.985 134.400 ;
        RECT 27.215 134.355 27.505 134.400 ;
        RECT 29.050 134.540 29.370 134.600 ;
        RECT 36.425 134.540 36.715 134.585 ;
        RECT 29.050 134.400 36.715 134.540 ;
        RECT 29.050 134.340 29.370 134.400 ;
        RECT 36.425 134.355 36.715 134.400 ;
        RECT 41.010 134.340 41.330 134.600 ;
        RECT 42.940 134.540 43.080 134.695 ;
        RECT 43.310 134.680 43.630 134.740 ;
        RECT 44.245 134.695 44.535 134.740 ;
        RECT 44.320 134.540 44.460 134.695 ;
        RECT 44.690 134.680 45.010 134.940 ;
        RECT 45.625 134.880 45.915 134.925 ;
        RECT 48.370 134.880 48.690 134.940 ;
        RECT 45.625 134.740 48.690 134.880 ;
        RECT 45.625 134.695 45.915 134.740 ;
        RECT 48.370 134.680 48.690 134.740 ;
        RECT 50.670 134.680 50.990 134.940 ;
        RECT 58.030 134.880 58.350 134.940 ;
        RECT 59.425 134.880 59.715 134.925 ;
        RECT 58.030 134.740 59.715 134.880 ;
        RECT 58.030 134.680 58.350 134.740 ;
        RECT 59.425 134.695 59.715 134.740 ;
        RECT 60.330 134.680 60.650 134.940 ;
        RECT 69.070 134.880 69.390 134.940 ;
        RECT 60.880 134.740 69.390 134.880 ;
        RECT 47.910 134.540 48.230 134.600 ;
        RECT 60.880 134.540 61.020 134.740 ;
        RECT 69.070 134.680 69.390 134.740 ;
        RECT 69.530 134.880 69.850 134.940 ;
        RECT 72.765 134.880 73.055 134.925 ;
        RECT 69.530 134.740 73.055 134.880 ;
        RECT 69.530 134.680 69.850 134.740 ;
        RECT 72.765 134.695 73.055 134.740 ;
        RECT 42.940 134.400 43.540 134.540 ;
        RECT 44.320 134.400 48.230 134.540 ;
        RECT 23.110 134.200 23.400 134.245 ;
        RECT 25.210 134.200 25.500 134.245 ;
        RECT 26.780 134.200 27.070 134.245 ;
        RECT 23.110 134.060 27.070 134.200 ;
        RECT 23.110 134.015 23.400 134.060 ;
        RECT 25.210 134.015 25.500 134.060 ;
        RECT 26.780 134.015 27.070 134.060 ;
        RECT 29.525 133.860 29.815 133.905 ;
        RECT 22.240 133.720 29.815 133.860 ;
        RECT 29.525 133.675 29.815 133.720 ;
        RECT 41.930 133.860 42.250 133.920 ;
        RECT 43.400 133.860 43.540 134.400 ;
        RECT 47.910 134.340 48.230 134.400 ;
        RECT 48.460 134.400 61.020 134.540 ;
        RECT 45.610 134.200 45.930 134.260 ;
        RECT 48.460 134.200 48.600 134.400 ;
        RECT 62.170 134.340 62.490 134.600 ;
        RECT 63.550 134.340 63.870 134.600 ;
        RECT 64.610 134.540 64.900 134.585 ;
        RECT 65.390 134.540 65.710 134.600 ;
        RECT 64.610 134.400 65.710 134.540 ;
        RECT 64.610 134.355 64.900 134.400 ;
        RECT 65.390 134.340 65.710 134.400 ;
        RECT 68.175 134.540 68.465 134.585 ;
        RECT 70.695 134.540 70.985 134.585 ;
        RECT 71.885 134.540 72.175 134.585 ;
        RECT 68.175 134.400 72.175 134.540 ;
        RECT 68.175 134.355 68.465 134.400 ;
        RECT 70.695 134.355 70.985 134.400 ;
        RECT 71.885 134.355 72.175 134.400 ;
        RECT 45.610 134.060 48.600 134.200 ;
        RECT 58.490 134.200 58.810 134.260 ;
        RECT 65.865 134.200 66.155 134.245 ;
        RECT 58.490 134.060 66.155 134.200 ;
        RECT 45.610 134.000 45.930 134.060 ;
        RECT 58.490 134.000 58.810 134.060 ;
        RECT 65.865 134.015 66.155 134.060 ;
        RECT 68.610 134.200 68.900 134.245 ;
        RECT 70.180 134.200 70.470 134.245 ;
        RECT 72.280 134.200 72.570 134.245 ;
        RECT 68.610 134.060 72.570 134.200 ;
        RECT 68.610 134.015 68.900 134.060 ;
        RECT 70.180 134.015 70.470 134.060 ;
        RECT 72.280 134.015 72.570 134.060 ;
        RECT 48.830 133.860 49.150 133.920 ;
        RECT 41.930 133.720 49.150 133.860 ;
        RECT 41.930 133.660 42.250 133.720 ;
        RECT 48.830 133.660 49.150 133.720 ;
        RECT 60.345 133.860 60.635 133.905 ;
        RECT 60.790 133.860 61.110 133.920 ;
        RECT 60.345 133.720 61.110 133.860 ;
        RECT 60.345 133.675 60.635 133.720 ;
        RECT 60.790 133.660 61.110 133.720 ;
        RECT 5.520 133.040 84.180 133.520 ;
        RECT 35.030 132.840 35.350 132.900 ;
        RECT 39.170 132.840 39.490 132.900 ;
        RECT 46.530 132.840 46.850 132.900 ;
        RECT 35.030 132.700 46.850 132.840 ;
        RECT 35.030 132.640 35.350 132.700 ;
        RECT 39.170 132.640 39.490 132.700 ;
        RECT 46.530 132.640 46.850 132.700 ;
        RECT 58.030 132.640 58.350 132.900 ;
        RECT 58.490 132.840 58.810 132.900 ;
        RECT 58.965 132.840 59.255 132.885 ;
        RECT 58.490 132.700 59.255 132.840 ;
        RECT 58.490 132.640 58.810 132.700 ;
        RECT 58.965 132.655 59.255 132.700 ;
        RECT 26.290 132.300 26.610 132.560 ;
        RECT 30.930 132.500 31.220 132.545 ;
        RECT 33.030 132.500 33.320 132.545 ;
        RECT 34.600 132.500 34.890 132.545 ;
        RECT 57.110 132.500 57.430 132.560 ;
        RECT 30.930 132.360 34.890 132.500 ;
        RECT 30.930 132.315 31.220 132.360 ;
        RECT 33.030 132.315 33.320 132.360 ;
        RECT 34.600 132.315 34.890 132.360 ;
        RECT 51.680 132.360 57.430 132.500 ;
        RECT 51.680 132.220 51.820 132.360 ;
        RECT 57.110 132.300 57.430 132.360 ;
        RECT 31.325 132.160 31.615 132.205 ;
        RECT 32.515 132.160 32.805 132.205 ;
        RECT 35.035 132.160 35.325 132.205 ;
        RECT 31.325 132.020 35.325 132.160 ;
        RECT 31.325 131.975 31.615 132.020 ;
        RECT 32.515 131.975 32.805 132.020 ;
        RECT 35.035 131.975 35.325 132.020 ;
        RECT 41.010 132.160 41.330 132.220 ;
        RECT 44.705 132.160 44.995 132.205 ;
        RECT 41.010 132.020 50.440 132.160 ;
        RECT 41.010 131.960 41.330 132.020 ;
        RECT 44.705 131.975 44.995 132.020 ;
        RECT 23.070 131.820 23.390 131.880 ;
        RECT 23.545 131.820 23.835 131.865 ;
        RECT 23.070 131.680 23.835 131.820 ;
        RECT 23.070 131.620 23.390 131.680 ;
        RECT 23.545 131.635 23.835 131.680 ;
        RECT 23.990 131.820 24.310 131.880 ;
        RECT 27.685 131.820 27.975 131.865 ;
        RECT 23.990 131.680 27.975 131.820 ;
        RECT 23.990 131.620 24.310 131.680 ;
        RECT 27.685 131.635 27.975 131.680 ;
        RECT 29.050 131.820 29.370 131.880 ;
        RECT 30.445 131.820 30.735 131.865 ;
        RECT 34.570 131.820 34.890 131.880 ;
        RECT 29.050 131.680 30.735 131.820 ;
        RECT 29.050 131.620 29.370 131.680 ;
        RECT 30.445 131.635 30.735 131.680 ;
        RECT 30.980 131.680 34.890 131.820 ;
        RECT 26.305 131.480 26.595 131.525 ;
        RECT 26.750 131.480 27.070 131.540 ;
        RECT 26.305 131.340 27.070 131.480 ;
        RECT 26.305 131.295 26.595 131.340 ;
        RECT 26.750 131.280 27.070 131.340 ;
        RECT 27.225 131.480 27.515 131.525 ;
        RECT 30.980 131.480 31.120 131.680 ;
        RECT 34.570 131.620 34.890 131.680 ;
        RECT 45.610 131.620 45.930 131.880 ;
        RECT 50.300 131.865 50.440 132.020 ;
        RECT 51.590 131.960 51.910 132.220 ;
        RECT 52.050 131.960 52.370 132.220 ;
        RECT 50.225 131.820 50.515 131.865 ;
        RECT 53.430 131.820 53.750 131.880 ;
        RECT 50.225 131.680 53.750 131.820 ;
        RECT 50.225 131.635 50.515 131.680 ;
        RECT 53.430 131.620 53.750 131.680 ;
        RECT 53.890 131.620 54.210 131.880 ;
        RECT 54.825 131.635 55.115 131.865 ;
        RECT 31.810 131.525 32.130 131.540 ;
        RECT 27.225 131.340 31.120 131.480 ;
        RECT 27.225 131.295 27.515 131.340 ;
        RECT 31.780 131.295 32.130 131.525 ;
        RECT 52.650 131.480 52.940 131.525 ;
        RECT 54.365 131.480 54.655 131.525 ;
        RECT 52.650 131.340 54.655 131.480 ;
        RECT 54.900 131.480 55.040 131.635 ;
        RECT 55.730 131.620 56.050 131.880 ;
        RECT 56.665 131.820 56.955 131.865 ;
        RECT 58.120 131.820 58.260 132.640 ;
        RECT 59.040 132.160 59.180 132.655 ;
        RECT 60.330 132.640 60.650 132.900 ;
        RECT 61.250 132.840 61.570 132.900 ;
        RECT 65.390 132.840 65.710 132.900 ;
        RECT 65.865 132.840 66.155 132.885 ;
        RECT 61.250 132.700 62.170 132.840 ;
        RECT 61.250 132.640 61.570 132.700 ;
        RECT 62.030 132.160 62.170 132.700 ;
        RECT 65.390 132.700 66.155 132.840 ;
        RECT 65.390 132.640 65.710 132.700 ;
        RECT 65.865 132.655 66.155 132.700 ;
        RECT 63.565 132.160 63.855 132.205 ;
        RECT 59.040 132.020 61.020 132.160 ;
        RECT 56.665 131.680 58.260 131.820 ;
        RECT 60.880 131.820 61.020 132.020 ;
        RECT 61.800 132.020 63.855 132.160 ;
        RECT 61.800 131.865 61.940 132.020 ;
        RECT 63.565 131.975 63.855 132.020 ;
        RECT 61.265 131.820 61.555 131.865 ;
        RECT 60.880 131.680 61.555 131.820 ;
        RECT 56.665 131.635 56.955 131.680 ;
        RECT 61.265 131.635 61.555 131.680 ;
        RECT 61.725 131.635 62.015 131.865 ;
        RECT 64.025 131.635 64.315 131.865 ;
        RECT 58.950 131.525 59.270 131.540 ;
        RECT 56.205 131.480 56.495 131.525 ;
        RECT 54.900 131.340 56.495 131.480 ;
        RECT 52.650 131.295 52.940 131.340 ;
        RECT 54.365 131.295 54.655 131.340 ;
        RECT 56.205 131.295 56.495 131.340 ;
        RECT 58.885 131.295 59.270 131.525 ;
        RECT 21.230 131.140 21.550 131.200 ;
        RECT 27.300 131.140 27.440 131.295 ;
        RECT 31.810 131.280 32.130 131.295 ;
        RECT 58.950 131.280 59.270 131.295 ;
        RECT 59.870 131.480 60.190 131.540 ;
        RECT 60.345 131.480 60.635 131.525 ;
        RECT 59.870 131.340 60.635 131.480 ;
        RECT 61.340 131.480 61.480 131.635 ;
        RECT 64.100 131.480 64.240 131.635 ;
        RECT 61.340 131.340 64.240 131.480 ;
        RECT 59.870 131.280 60.190 131.340 ;
        RECT 60.345 131.295 60.635 131.340 ;
        RECT 21.230 131.000 27.440 131.140 ;
        RECT 37.345 131.140 37.635 131.185 ;
        RECT 39.630 131.140 39.950 131.200 ;
        RECT 37.345 131.000 39.950 131.140 ;
        RECT 21.230 130.940 21.550 131.000 ;
        RECT 37.345 130.955 37.635 131.000 ;
        RECT 39.630 130.940 39.950 131.000 ;
        RECT 53.430 130.940 53.750 131.200 ;
        RECT 5.520 130.320 84.180 130.800 ;
        RECT 17.550 130.120 17.870 130.180 ;
        RECT 19.405 130.120 19.695 130.165 ;
        RECT 17.550 129.980 19.695 130.120 ;
        RECT 17.550 129.920 17.870 129.980 ;
        RECT 19.405 129.935 19.695 129.980 ;
        RECT 20.325 130.120 20.615 130.165 ;
        RECT 23.530 130.120 23.850 130.180 ;
        RECT 20.325 129.980 23.850 130.120 ;
        RECT 20.325 129.935 20.615 129.980 ;
        RECT 23.530 129.920 23.850 129.980 ;
        RECT 32.745 130.120 33.035 130.165 ;
        RECT 46.085 130.120 46.375 130.165 ;
        RECT 46.530 130.120 46.850 130.180 ;
        RECT 32.745 129.980 42.160 130.120 ;
        RECT 32.745 129.935 33.035 129.980 ;
        RECT 31.825 129.780 32.115 129.825 ;
        RECT 41.010 129.780 41.330 129.840 ;
        RECT 31.825 129.640 41.330 129.780 ;
        RECT 42.020 129.780 42.160 129.980 ;
        RECT 46.085 129.980 46.850 130.120 ;
        RECT 46.085 129.935 46.375 129.980 ;
        RECT 46.530 129.920 46.850 129.980 ;
        RECT 55.730 130.120 56.050 130.180 ;
        RECT 56.665 130.120 56.955 130.165 ;
        RECT 55.730 129.980 56.955 130.120 ;
        RECT 55.730 129.920 56.050 129.980 ;
        RECT 56.665 129.935 56.955 129.980 ;
        RECT 59.870 130.120 60.190 130.180 ;
        RECT 65.405 130.120 65.695 130.165 ;
        RECT 59.870 129.980 65.695 130.120 ;
        RECT 59.870 129.920 60.190 129.980 ;
        RECT 65.405 129.935 65.695 129.980 ;
        RECT 45.150 129.780 45.470 129.840 ;
        RECT 45.625 129.780 45.915 129.825 ;
        RECT 42.020 129.640 45.915 129.780 ;
        RECT 31.825 129.595 32.115 129.640 ;
        RECT 41.010 129.580 41.330 129.640 ;
        RECT 45.150 129.580 45.470 129.640 ;
        RECT 45.625 129.595 45.915 129.640 ;
        RECT 51.100 129.780 51.390 129.825 ;
        RECT 53.430 129.780 53.750 129.840 ;
        RECT 61.710 129.780 62.030 129.840 ;
        RECT 66.310 129.780 66.630 129.840 ;
        RECT 68.610 129.780 68.930 129.840 ;
        RECT 51.100 129.640 53.750 129.780 ;
        RECT 51.100 129.595 51.390 129.640 ;
        RECT 53.430 129.580 53.750 129.640 ;
        RECT 58.580 129.640 68.930 129.780 ;
        RECT 33.205 129.440 33.495 129.485 ;
        RECT 35.030 129.440 35.350 129.500 ;
        RECT 33.205 129.300 35.350 129.440 ;
        RECT 33.205 129.255 33.495 129.300 ;
        RECT 35.030 129.240 35.350 129.300 ;
        RECT 38.725 129.440 39.015 129.485 ;
        RECT 39.170 129.440 39.490 129.500 ;
        RECT 38.725 129.300 39.490 129.440 ;
        RECT 38.725 129.255 39.015 129.300 ;
        RECT 39.170 129.240 39.490 129.300 ;
        RECT 39.630 129.240 39.950 129.500 ;
        RECT 41.930 129.240 42.250 129.500 ;
        RECT 46.670 129.440 46.960 129.485 ;
        RECT 43.860 129.300 46.960 129.440 ;
        RECT 22.165 129.100 22.455 129.145 ;
        RECT 23.070 129.100 23.390 129.160 ;
        RECT 22.165 128.960 23.390 129.100 ;
        RECT 22.165 128.915 22.455 128.960 ;
        RECT 23.070 128.900 23.390 128.960 ;
        RECT 28.130 128.900 28.450 129.160 ;
        RECT 38.265 129.100 38.555 129.145 ;
        RECT 39.720 129.100 39.860 129.240 ;
        RECT 38.265 128.960 39.860 129.100 ;
        RECT 38.265 128.915 38.555 128.960 ;
        RECT 42.390 128.900 42.710 129.160 ;
        RECT 43.860 129.145 44.000 129.300 ;
        RECT 46.670 129.255 46.960 129.300 ;
        RECT 49.765 129.440 50.055 129.485 ;
        RECT 50.210 129.440 50.530 129.500 ;
        RECT 58.580 129.485 58.720 129.640 ;
        RECT 61.710 129.580 62.030 129.640 ;
        RECT 66.310 129.580 66.630 129.640 ;
        RECT 68.610 129.580 68.930 129.640 ;
        RECT 59.870 129.485 60.190 129.500 ;
        RECT 49.765 129.300 50.530 129.440 ;
        RECT 49.765 129.255 50.055 129.300 ;
        RECT 50.210 129.240 50.530 129.300 ;
        RECT 58.505 129.255 58.795 129.485 ;
        RECT 59.840 129.255 60.190 129.485 ;
        RECT 59.870 129.240 60.190 129.255 ;
        RECT 43.785 128.915 44.075 129.145 ;
        RECT 44.245 128.915 44.535 129.145 ;
        RECT 50.645 129.100 50.935 129.145 ;
        RECT 51.835 129.100 52.125 129.145 ;
        RECT 54.355 129.100 54.645 129.145 ;
        RECT 50.645 128.960 54.645 129.100 ;
        RECT 50.645 128.915 50.935 128.960 ;
        RECT 51.835 128.915 52.125 128.960 ;
        RECT 54.355 128.915 54.645 128.960 ;
        RECT 59.385 129.100 59.675 129.145 ;
        RECT 60.575 129.100 60.865 129.145 ;
        RECT 63.095 129.100 63.385 129.145 ;
        RECT 59.385 128.960 63.385 129.100 ;
        RECT 59.385 128.915 59.675 128.960 ;
        RECT 60.575 128.915 60.865 128.960 ;
        RECT 63.095 128.915 63.385 128.960 ;
        RECT 31.810 128.560 32.130 128.820 ;
        RECT 41.010 128.760 41.330 128.820 ;
        RECT 44.320 128.760 44.460 128.915 ;
        RECT 41.010 128.620 44.460 128.760 ;
        RECT 50.250 128.760 50.540 128.805 ;
        RECT 52.350 128.760 52.640 128.805 ;
        RECT 53.920 128.760 54.210 128.805 ;
        RECT 50.250 128.620 54.210 128.760 ;
        RECT 41.010 128.560 41.330 128.620 ;
        RECT 50.250 128.575 50.540 128.620 ;
        RECT 52.350 128.575 52.640 128.620 ;
        RECT 53.920 128.575 54.210 128.620 ;
        RECT 58.990 128.760 59.280 128.805 ;
        RECT 61.090 128.760 61.380 128.805 ;
        RECT 62.660 128.760 62.950 128.805 ;
        RECT 58.990 128.620 62.950 128.760 ;
        RECT 58.990 128.575 59.280 128.620 ;
        RECT 61.090 128.575 61.380 128.620 ;
        RECT 62.660 128.575 62.950 128.620 ;
        RECT 20.325 128.420 20.615 128.465 ;
        RECT 21.230 128.420 21.550 128.480 ;
        RECT 20.325 128.280 21.550 128.420 ;
        RECT 20.325 128.235 20.615 128.280 ;
        RECT 21.230 128.220 21.550 128.280 ;
        RECT 23.530 128.420 23.850 128.480 ;
        RECT 26.305 128.420 26.595 128.465 ;
        RECT 26.750 128.420 27.070 128.480 ;
        RECT 23.530 128.280 27.070 128.420 ;
        RECT 23.530 128.220 23.850 128.280 ;
        RECT 26.305 128.235 26.595 128.280 ;
        RECT 26.750 128.220 27.070 128.280 ;
        RECT 29.970 128.420 30.290 128.480 ;
        RECT 30.905 128.420 31.195 128.465 ;
        RECT 29.970 128.280 31.195 128.420 ;
        RECT 29.970 128.220 30.290 128.280 ;
        RECT 30.905 128.235 31.195 128.280 ;
        RECT 35.030 128.220 35.350 128.480 ;
        RECT 37.790 128.420 38.110 128.480 ;
        RECT 39.185 128.420 39.475 128.465 ;
        RECT 37.790 128.280 39.475 128.420 ;
        RECT 37.790 128.220 38.110 128.280 ;
        RECT 39.185 128.235 39.475 128.280 ;
        RECT 47.450 128.220 47.770 128.480 ;
        RECT 5.520 127.600 84.180 128.080 ;
        RECT 52.970 127.200 53.290 127.460 ;
        RECT 59.870 127.400 60.190 127.460 ;
        RECT 60.805 127.400 61.095 127.445 ;
        RECT 59.870 127.260 61.095 127.400 ;
        RECT 59.870 127.200 60.190 127.260 ;
        RECT 60.805 127.215 61.095 127.260 ;
        RECT 21.690 127.060 21.980 127.105 ;
        RECT 23.260 127.060 23.550 127.105 ;
        RECT 25.360 127.060 25.650 127.105 ;
        RECT 21.690 126.920 25.650 127.060 ;
        RECT 21.690 126.875 21.980 126.920 ;
        RECT 23.260 126.875 23.550 126.920 ;
        RECT 25.360 126.875 25.650 126.920 ;
        RECT 29.090 127.060 29.380 127.105 ;
        RECT 31.190 127.060 31.480 127.105 ;
        RECT 32.760 127.060 33.050 127.105 ;
        RECT 29.090 126.920 33.050 127.060 ;
        RECT 29.090 126.875 29.380 126.920 ;
        RECT 31.190 126.875 31.480 126.920 ;
        RECT 32.760 126.875 33.050 126.920 ;
        RECT 34.570 127.060 34.890 127.120 ;
        RECT 39.185 127.060 39.475 127.105 ;
        RECT 34.570 126.920 39.475 127.060 ;
        RECT 34.570 126.860 34.890 126.920 ;
        RECT 39.185 126.875 39.475 126.920 ;
        RECT 46.570 127.060 46.860 127.105 ;
        RECT 48.670 127.060 48.960 127.105 ;
        RECT 50.240 127.060 50.530 127.105 ;
        RECT 62.170 127.060 62.490 127.120 ;
        RECT 46.570 126.920 50.530 127.060 ;
        RECT 46.570 126.875 46.860 126.920 ;
        RECT 48.670 126.875 48.960 126.920 ;
        RECT 50.240 126.875 50.530 126.920 ;
        RECT 57.660 126.920 62.490 127.060 ;
        RECT 21.255 126.720 21.545 126.765 ;
        RECT 23.775 126.720 24.065 126.765 ;
        RECT 24.965 126.720 25.255 126.765 ;
        RECT 26.290 126.720 26.610 126.780 ;
        RECT 21.255 126.580 25.255 126.720 ;
        RECT 21.255 126.535 21.545 126.580 ;
        RECT 23.775 126.535 24.065 126.580 ;
        RECT 24.965 126.535 25.255 126.580 ;
        RECT 25.460 126.580 26.610 126.720 ;
        RECT 24.565 126.380 24.855 126.425 ;
        RECT 25.460 126.380 25.600 126.580 ;
        RECT 26.290 126.520 26.610 126.580 ;
        RECT 29.485 126.720 29.775 126.765 ;
        RECT 30.675 126.720 30.965 126.765 ;
        RECT 33.195 126.720 33.485 126.765 ;
        RECT 38.265 126.720 38.555 126.765 ;
        RECT 29.485 126.580 33.485 126.720 ;
        RECT 29.485 126.535 29.775 126.580 ;
        RECT 30.675 126.535 30.965 126.580 ;
        RECT 33.195 126.535 33.485 126.580 ;
        RECT 36.960 126.580 38.555 126.720 ;
        RECT 24.565 126.240 25.600 126.380 ;
        RECT 25.845 126.380 26.135 126.425 ;
        RECT 28.605 126.380 28.895 126.425 ;
        RECT 29.050 126.380 29.370 126.440 ;
        RECT 29.970 126.425 30.290 126.440 ;
        RECT 29.940 126.380 30.290 126.425 ;
        RECT 32.730 126.380 33.050 126.440 ;
        RECT 25.845 126.240 29.370 126.380 ;
        RECT 29.775 126.240 30.290 126.380 ;
        RECT 24.565 126.195 24.855 126.240 ;
        RECT 25.845 126.195 26.135 126.240 ;
        RECT 28.605 126.195 28.895 126.240 ;
        RECT 29.050 126.180 29.370 126.240 ;
        RECT 29.940 126.195 30.290 126.240 ;
        RECT 29.970 126.180 30.290 126.195 ;
        RECT 30.980 126.240 33.050 126.380 ;
        RECT 20.770 126.040 21.090 126.100 ;
        RECT 27.225 126.040 27.515 126.085 ;
        RECT 20.770 125.900 27.515 126.040 ;
        RECT 20.770 125.840 21.090 125.900 ;
        RECT 27.225 125.855 27.515 125.900 ;
        RECT 28.145 126.040 28.435 126.085 ;
        RECT 30.980 126.040 31.120 126.240 ;
        RECT 32.730 126.180 33.050 126.240 ;
        RECT 35.490 126.380 35.810 126.440 ;
        RECT 36.425 126.380 36.715 126.425 ;
        RECT 35.490 126.240 36.715 126.380 ;
        RECT 35.490 126.180 35.810 126.240 ;
        RECT 36.425 126.195 36.715 126.240 ;
        RECT 35.965 126.040 36.255 126.085 ;
        RECT 28.145 125.900 31.120 126.040 ;
        RECT 31.440 125.900 36.255 126.040 ;
        RECT 28.145 125.855 28.435 125.900 ;
        RECT 18.930 125.500 19.250 125.760 ;
        RECT 26.305 125.700 26.595 125.745 ;
        RECT 31.440 125.700 31.580 125.900 ;
        RECT 35.965 125.855 36.255 125.900 ;
        RECT 26.305 125.560 31.580 125.700 ;
        RECT 32.730 125.700 33.050 125.760 ;
        RECT 35.505 125.700 35.795 125.745 ;
        RECT 36.960 125.700 37.100 126.580 ;
        RECT 38.265 126.535 38.555 126.580 ;
        RECT 39.630 126.720 39.950 126.780 ;
        RECT 57.660 126.765 57.800 126.920 ;
        RECT 62.170 126.860 62.490 126.920 ;
        RECT 46.965 126.720 47.255 126.765 ;
        RECT 48.155 126.720 48.445 126.765 ;
        RECT 50.675 126.720 50.965 126.765 ;
        RECT 39.630 126.580 45.840 126.720 ;
        RECT 37.790 126.180 38.110 126.440 ;
        RECT 38.340 126.380 38.480 126.535 ;
        RECT 39.630 126.520 39.950 126.580 ;
        RECT 41.470 126.380 41.790 126.440 ;
        RECT 45.700 126.425 45.840 126.580 ;
        RECT 46.965 126.580 50.965 126.720 ;
        RECT 46.965 126.535 47.255 126.580 ;
        RECT 48.155 126.535 48.445 126.580 ;
        RECT 50.675 126.535 50.965 126.580 ;
        RECT 57.585 126.535 57.875 126.765 ;
        RECT 60.010 126.720 60.300 126.765 ;
        RECT 60.790 126.720 61.110 126.780 ;
        RECT 60.010 126.580 61.110 126.720 ;
        RECT 60.010 126.535 60.300 126.580 ;
        RECT 60.790 126.520 61.110 126.580 ;
        RECT 42.405 126.380 42.695 126.425 ;
        RECT 44.705 126.380 44.995 126.425 ;
        RECT 38.340 126.240 44.995 126.380 ;
        RECT 41.470 126.180 41.790 126.240 ;
        RECT 42.405 126.195 42.695 126.240 ;
        RECT 44.705 126.195 44.995 126.240 ;
        RECT 45.625 126.195 45.915 126.425 ;
        RECT 46.085 126.380 46.375 126.425 ;
        RECT 50.210 126.380 50.530 126.440 ;
        RECT 46.085 126.240 50.530 126.380 ;
        RECT 46.085 126.195 46.375 126.240 ;
        RECT 50.210 126.180 50.530 126.240 ;
        RECT 57.110 126.380 57.430 126.440 ;
        RECT 58.965 126.380 59.255 126.425 ;
        RECT 57.110 126.240 59.255 126.380 ;
        RECT 57.110 126.180 57.430 126.240 ;
        RECT 58.965 126.195 59.255 126.240 ;
        RECT 37.330 126.040 37.650 126.100 ;
        RECT 47.450 126.085 47.770 126.100 ;
        RECT 39.645 126.040 39.935 126.085 ;
        RECT 47.420 126.040 47.770 126.085 ;
        RECT 37.330 125.900 39.935 126.040 ;
        RECT 47.255 125.900 47.770 126.040 ;
        RECT 37.330 125.840 37.650 125.900 ;
        RECT 39.645 125.855 39.935 125.900 ;
        RECT 47.420 125.855 47.770 125.900 ;
        RECT 47.450 125.840 47.770 125.855 ;
        RECT 32.730 125.560 37.100 125.700 ;
        RECT 38.250 125.700 38.570 125.760 ;
        RECT 41.930 125.700 42.250 125.760 ;
        RECT 44.705 125.700 44.995 125.745 ;
        RECT 38.250 125.560 44.995 125.700 ;
        RECT 26.305 125.515 26.595 125.560 ;
        RECT 32.730 125.500 33.050 125.560 ;
        RECT 35.505 125.515 35.795 125.560 ;
        RECT 38.250 125.500 38.570 125.560 ;
        RECT 41.930 125.500 42.250 125.560 ;
        RECT 44.705 125.515 44.995 125.560 ;
        RECT 46.530 125.700 46.850 125.760 ;
        RECT 59.425 125.700 59.715 125.745 ;
        RECT 46.530 125.560 59.715 125.700 ;
        RECT 46.530 125.500 46.850 125.560 ;
        RECT 59.425 125.515 59.715 125.560 ;
        RECT 5.520 124.880 84.180 125.360 ;
        RECT 20.770 124.480 21.090 124.740 ;
        RECT 28.130 124.480 28.450 124.740 ;
        RECT 39.645 124.495 39.935 124.725 ;
        RECT 37.790 124.340 38.110 124.400 ;
        RECT 29.600 124.200 38.110 124.340 ;
        RECT 26.405 124.000 26.695 124.045 ;
        RECT 27.210 124.000 27.530 124.060 ;
        RECT 26.405 123.860 27.530 124.000 ;
        RECT 26.405 123.815 26.695 123.860 ;
        RECT 27.210 123.800 27.530 123.860 ;
        RECT 29.600 123.720 29.740 124.200 ;
        RECT 37.790 124.140 38.110 124.200 ;
        RECT 29.985 124.000 30.275 124.045 ;
        RECT 37.330 124.000 37.650 124.060 ;
        RECT 29.985 123.860 37.650 124.000 ;
        RECT 29.985 123.815 30.275 123.860 ;
        RECT 37.330 123.800 37.650 123.860 ;
        RECT 38.250 123.800 38.570 124.060 ;
        RECT 39.720 124.000 39.860 124.495 ;
        RECT 41.385 124.000 41.675 124.045 ;
        RECT 39.720 123.860 41.675 124.000 ;
        RECT 41.385 123.815 41.675 123.860 ;
        RECT 23.095 123.660 23.385 123.705 ;
        RECT 25.615 123.660 25.905 123.705 ;
        RECT 26.805 123.660 27.095 123.705 ;
        RECT 23.095 123.520 27.095 123.660 ;
        RECT 23.095 123.475 23.385 123.520 ;
        RECT 25.615 123.475 25.905 123.520 ;
        RECT 26.805 123.475 27.095 123.520 ;
        RECT 27.685 123.475 27.975 123.705 ;
        RECT 23.530 123.320 23.820 123.365 ;
        RECT 25.100 123.320 25.390 123.365 ;
        RECT 27.200 123.320 27.490 123.365 ;
        RECT 23.530 123.180 27.490 123.320 ;
        RECT 27.760 123.320 27.900 123.475 ;
        RECT 29.510 123.460 29.830 123.720 ;
        RECT 32.270 123.660 32.590 123.720 ;
        RECT 32.745 123.660 33.035 123.705 ;
        RECT 32.270 123.520 33.035 123.660 ;
        RECT 32.270 123.460 32.590 123.520 ;
        RECT 32.745 123.475 33.035 123.520 ;
        RECT 34.110 123.660 34.430 123.720 ;
        RECT 36.410 123.660 36.730 123.720 ;
        RECT 34.110 123.520 36.730 123.660 ;
        RECT 34.110 123.460 34.430 123.520 ;
        RECT 36.410 123.460 36.730 123.520 ;
        RECT 36.885 123.660 37.175 123.705 ;
        RECT 37.790 123.660 38.110 123.720 ;
        RECT 36.885 123.520 38.110 123.660 ;
        RECT 36.885 123.475 37.175 123.520 ;
        RECT 37.790 123.460 38.110 123.520 ;
        RECT 38.710 123.460 39.030 123.720 ;
        RECT 40.105 123.475 40.395 123.705 ;
        RECT 40.985 123.660 41.275 123.705 ;
        RECT 42.175 123.660 42.465 123.705 ;
        RECT 44.695 123.660 44.985 123.705 ;
        RECT 40.985 123.520 44.985 123.660 ;
        RECT 40.985 123.475 41.275 123.520 ;
        RECT 42.175 123.475 42.465 123.520 ;
        RECT 44.695 123.475 44.985 123.520 ;
        RECT 29.050 123.320 29.370 123.380 ;
        RECT 40.180 123.320 40.320 123.475 ;
        RECT 27.760 123.180 40.320 123.320 ;
        RECT 40.590 123.320 40.880 123.365 ;
        RECT 42.690 123.320 42.980 123.365 ;
        RECT 44.260 123.320 44.550 123.365 ;
        RECT 40.590 123.180 44.550 123.320 ;
        RECT 23.530 123.135 23.820 123.180 ;
        RECT 25.100 123.135 25.390 123.180 ;
        RECT 27.200 123.135 27.490 123.180 ;
        RECT 29.050 123.120 29.370 123.180 ;
        RECT 36.960 123.040 37.100 123.180 ;
        RECT 40.590 123.135 40.880 123.180 ;
        RECT 42.690 123.135 42.980 123.180 ;
        RECT 44.260 123.135 44.550 123.180 ;
        RECT 45.610 123.320 45.930 123.380 ;
        RECT 47.005 123.320 47.295 123.365 ;
        RECT 45.610 123.180 47.295 123.320 ;
        RECT 45.610 123.120 45.930 123.180 ;
        RECT 47.005 123.135 47.295 123.180 ;
        RECT 31.810 122.980 32.130 123.040 ;
        RECT 34.110 122.980 34.430 123.040 ;
        RECT 31.810 122.840 34.430 122.980 ;
        RECT 31.810 122.780 32.130 122.840 ;
        RECT 34.110 122.780 34.430 122.840 ;
        RECT 35.950 122.780 36.270 123.040 ;
        RECT 36.870 122.780 37.190 123.040 ;
        RECT 37.790 122.980 38.110 123.040 ;
        RECT 41.010 122.980 41.330 123.040 ;
        RECT 37.790 122.840 41.330 122.980 ;
        RECT 37.790 122.780 38.110 122.840 ;
        RECT 41.010 122.780 41.330 122.840 ;
        RECT 5.520 122.160 84.180 122.640 ;
        RECT 27.210 121.760 27.530 122.020 ;
        RECT 32.270 121.760 32.590 122.020 ;
        RECT 32.745 121.960 33.035 122.005 ;
        RECT 35.030 121.960 35.350 122.020 ;
        RECT 32.745 121.820 35.350 121.960 ;
        RECT 32.745 121.775 33.035 121.820 ;
        RECT 35.030 121.760 35.350 121.820 ;
        RECT 37.330 121.960 37.650 122.020 ;
        RECT 39.170 121.960 39.490 122.020 ;
        RECT 40.550 121.960 40.870 122.020 ;
        RECT 41.025 121.960 41.315 122.005 ;
        RECT 37.330 121.820 38.435 121.960 ;
        RECT 37.330 121.760 37.650 121.820 ;
        RECT 28.605 121.620 28.895 121.665 ;
        RECT 29.510 121.620 29.830 121.680 ;
        RECT 28.605 121.480 29.830 121.620 ;
        RECT 28.605 121.435 28.895 121.480 ;
        RECT 29.510 121.420 29.830 121.480 ;
        RECT 33.650 121.420 33.970 121.680 ;
        RECT 34.150 121.620 34.440 121.665 ;
        RECT 36.250 121.620 36.540 121.665 ;
        RECT 37.820 121.620 38.110 121.665 ;
        RECT 34.150 121.480 38.110 121.620 ;
        RECT 38.295 121.620 38.435 121.820 ;
        RECT 39.170 121.820 41.315 121.960 ;
        RECT 39.170 121.760 39.490 121.820 ;
        RECT 40.550 121.760 40.870 121.820 ;
        RECT 41.025 121.775 41.315 121.820 ;
        RECT 46.085 121.620 46.375 121.665 ;
        RECT 38.295 121.480 46.375 121.620 ;
        RECT 34.150 121.435 34.440 121.480 ;
        RECT 36.250 121.435 36.540 121.480 ;
        RECT 37.820 121.435 38.110 121.480 ;
        RECT 46.085 121.435 46.375 121.480 ;
        RECT 18.930 121.280 19.250 121.340 ;
        RECT 20.325 121.280 20.615 121.325 ;
        RECT 18.930 121.140 20.615 121.280 ;
        RECT 18.930 121.080 19.250 121.140 ;
        RECT 20.325 121.095 20.615 121.140 ;
        RECT 29.050 121.080 29.370 121.340 ;
        RECT 33.740 121.280 33.880 121.420 ;
        RECT 30.520 121.140 33.880 121.280 ;
        RECT 34.545 121.280 34.835 121.325 ;
        RECT 35.735 121.280 36.025 121.325 ;
        RECT 38.255 121.280 38.545 121.325 ;
        RECT 34.545 121.140 38.545 121.280 ;
        RECT 28.145 120.755 28.435 120.985 ;
        RECT 29.525 120.940 29.815 120.985 ;
        RECT 29.970 120.940 30.290 121.000 ;
        RECT 30.520 120.985 30.660 121.140 ;
        RECT 34.545 121.095 34.835 121.140 ;
        RECT 35.735 121.095 36.025 121.140 ;
        RECT 38.255 121.095 38.545 121.140 ;
        RECT 41.470 121.080 41.790 121.340 ;
        RECT 58.045 121.280 58.335 121.325 ;
        RECT 58.505 121.280 58.795 121.325 ;
        RECT 58.045 121.140 58.795 121.280 ;
        RECT 58.045 121.095 58.335 121.140 ;
        RECT 58.505 121.095 58.795 121.140 ;
        RECT 29.525 120.800 30.290 120.940 ;
        RECT 29.525 120.755 29.815 120.800 ;
        RECT 28.220 120.600 28.360 120.755 ;
        RECT 29.970 120.740 30.290 120.800 ;
        RECT 30.445 120.755 30.735 120.985 ;
        RECT 31.350 120.740 31.670 121.000 ;
        RECT 31.810 120.740 32.130 121.000 ;
        RECT 33.205 120.755 33.495 120.985 ;
        RECT 33.665 120.940 33.955 120.985 ;
        RECT 36.870 120.940 37.190 121.000 ;
        RECT 33.665 120.800 37.190 120.940 ;
        RECT 33.665 120.755 33.955 120.800 ;
        RECT 32.730 120.600 33.050 120.660 ;
        RECT 28.220 120.460 33.050 120.600 ;
        RECT 32.730 120.400 33.050 120.460 ;
        RECT 23.545 120.260 23.835 120.305 ;
        RECT 23.990 120.260 24.310 120.320 ;
        RECT 23.545 120.120 24.310 120.260 ;
        RECT 33.280 120.260 33.420 120.755 ;
        RECT 36.870 120.740 37.190 120.800 ;
        RECT 41.010 120.740 41.330 121.000 ;
        RECT 52.050 120.740 52.370 121.000 ;
        RECT 59.870 120.740 60.190 121.000 ;
        RECT 60.330 120.740 60.650 121.000 ;
        RECT 60.805 120.755 61.095 120.985 ;
        RECT 61.250 120.940 61.570 121.000 ;
        RECT 61.725 120.940 62.015 120.985 ;
        RECT 61.250 120.800 62.015 120.940 ;
        RECT 35.000 120.600 35.290 120.645 ;
        RECT 35.950 120.600 36.270 120.660 ;
        RECT 35.000 120.460 36.270 120.600 ;
        RECT 35.000 120.415 35.290 120.460 ;
        RECT 35.950 120.400 36.270 120.460 ;
        RECT 45.165 120.415 45.455 120.645 ;
        RECT 58.030 120.600 58.350 120.660 ;
        RECT 60.880 120.600 61.020 120.755 ;
        RECT 61.250 120.740 61.570 120.800 ;
        RECT 61.725 120.755 62.015 120.800 ;
        RECT 58.030 120.460 61.020 120.600 ;
        RECT 38.710 120.260 39.030 120.320 ;
        RECT 33.280 120.120 39.030 120.260 ;
        RECT 23.545 120.075 23.835 120.120 ;
        RECT 23.990 120.060 24.310 120.120 ;
        RECT 38.710 120.060 39.030 120.120 ;
        RECT 42.865 120.260 43.155 120.305 ;
        RECT 43.310 120.260 43.630 120.320 ;
        RECT 45.240 120.260 45.380 120.415 ;
        RECT 58.030 120.400 58.350 120.460 ;
        RECT 42.865 120.120 45.380 120.260 ;
        RECT 48.830 120.260 49.150 120.320 ;
        RECT 49.305 120.260 49.595 120.305 ;
        RECT 48.830 120.120 49.595 120.260 ;
        RECT 42.865 120.075 43.155 120.120 ;
        RECT 43.310 120.060 43.630 120.120 ;
        RECT 48.830 120.060 49.150 120.120 ;
        RECT 49.305 120.075 49.595 120.120 ;
        RECT 53.890 120.260 54.210 120.320 ;
        RECT 54.825 120.260 55.115 120.305 ;
        RECT 53.890 120.120 55.115 120.260 ;
        RECT 53.890 120.060 54.210 120.120 ;
        RECT 54.825 120.075 55.115 120.120 ;
        RECT 5.520 119.440 84.180 119.920 ;
        RECT 22.165 119.240 22.455 119.285 ;
        RECT 23.070 119.240 23.390 119.300 ;
        RECT 22.165 119.100 23.390 119.240 ;
        RECT 22.165 119.055 22.455 119.100 ;
        RECT 23.070 119.040 23.390 119.100 ;
        RECT 38.710 119.240 39.030 119.300 ;
        RECT 40.105 119.240 40.395 119.285 ;
        RECT 38.710 119.100 40.395 119.240 ;
        RECT 38.710 119.040 39.030 119.100 ;
        RECT 40.105 119.055 40.395 119.100 ;
        RECT 41.010 119.240 41.330 119.300 ;
        RECT 55.285 119.240 55.575 119.285 ;
        RECT 41.010 119.100 55.575 119.240 ;
        RECT 41.010 119.040 41.330 119.100 ;
        RECT 55.285 119.055 55.575 119.100 ;
        RECT 38.265 118.900 38.555 118.945 ;
        RECT 50.210 118.900 50.530 118.960 ;
        RECT 38.265 118.760 40.780 118.900 ;
        RECT 38.265 118.715 38.555 118.760 ;
        RECT 40.640 118.620 40.780 118.760 ;
        RECT 47.540 118.760 50.530 118.900 ;
        RECT 15.250 118.360 15.570 118.620 ;
        RECT 15.710 118.560 16.030 118.620 ;
        RECT 16.545 118.560 16.835 118.605 ;
        RECT 15.710 118.420 16.835 118.560 ;
        RECT 15.710 118.360 16.030 118.420 ;
        RECT 16.545 118.375 16.835 118.420 ;
        RECT 39.185 118.375 39.475 118.605 ;
        RECT 40.550 118.560 40.870 118.620 ;
        RECT 41.025 118.560 41.315 118.605 ;
        RECT 40.550 118.420 41.315 118.560 ;
        RECT 16.145 118.220 16.435 118.265 ;
        RECT 17.335 118.220 17.625 118.265 ;
        RECT 19.855 118.220 20.145 118.265 ;
        RECT 16.145 118.080 20.145 118.220 ;
        RECT 39.260 118.220 39.400 118.375 ;
        RECT 40.550 118.360 40.870 118.420 ;
        RECT 41.025 118.375 41.315 118.420 ;
        RECT 41.930 118.360 42.250 118.620 ;
        RECT 47.540 118.605 47.680 118.760 ;
        RECT 50.210 118.700 50.530 118.760 ;
        RECT 48.830 118.605 49.150 118.620 ;
        RECT 47.465 118.375 47.755 118.605 ;
        RECT 48.800 118.560 49.150 118.605 ;
        RECT 54.825 118.560 55.115 118.605 ;
        RECT 48.635 118.420 49.150 118.560 ;
        RECT 48.800 118.375 49.150 118.420 ;
        RECT 48.830 118.360 49.150 118.375 ;
        RECT 54.440 118.420 55.115 118.560 ;
        RECT 42.020 118.220 42.160 118.360 ;
        RECT 39.260 118.080 42.160 118.220 ;
        RECT 48.345 118.220 48.635 118.265 ;
        RECT 49.535 118.220 49.825 118.265 ;
        RECT 52.055 118.220 52.345 118.265 ;
        RECT 48.345 118.080 52.345 118.220 ;
        RECT 16.145 118.035 16.435 118.080 ;
        RECT 17.335 118.035 17.625 118.080 ;
        RECT 19.855 118.035 20.145 118.080 ;
        RECT 48.345 118.035 48.635 118.080 ;
        RECT 49.535 118.035 49.825 118.080 ;
        RECT 52.055 118.035 52.345 118.080 ;
        RECT 15.750 117.880 16.040 117.925 ;
        RECT 17.850 117.880 18.140 117.925 ;
        RECT 19.420 117.880 19.710 117.925 ;
        RECT 15.750 117.740 19.710 117.880 ;
        RECT 15.750 117.695 16.040 117.740 ;
        RECT 17.850 117.695 18.140 117.740 ;
        RECT 19.420 117.695 19.710 117.740 ;
        RECT 33.190 117.880 33.510 117.940 ;
        RECT 54.440 117.925 54.580 118.420 ;
        RECT 54.825 118.375 55.115 118.420 ;
        RECT 55.745 118.560 56.035 118.605 ;
        RECT 59.410 118.560 59.730 118.620 ;
        RECT 55.745 118.420 59.730 118.560 ;
        RECT 55.745 118.375 56.035 118.420 ;
        RECT 59.410 118.360 59.730 118.420 ;
        RECT 65.045 118.560 65.335 118.605 ;
        RECT 65.850 118.560 66.170 118.620 ;
        RECT 65.045 118.420 66.170 118.560 ;
        RECT 65.045 118.375 65.335 118.420 ;
        RECT 65.850 118.360 66.170 118.420 ;
        RECT 66.310 118.560 66.630 118.620 ;
        RECT 69.070 118.560 69.390 118.620 ;
        RECT 66.310 118.420 69.390 118.560 ;
        RECT 66.310 118.360 66.630 118.420 ;
        RECT 69.070 118.360 69.390 118.420 ;
        RECT 61.735 118.220 62.025 118.265 ;
        RECT 64.255 118.220 64.545 118.265 ;
        RECT 65.445 118.220 65.735 118.265 ;
        RECT 61.735 118.080 65.735 118.220 ;
        RECT 61.735 118.035 62.025 118.080 ;
        RECT 64.255 118.035 64.545 118.080 ;
        RECT 65.445 118.035 65.735 118.080 ;
        RECT 41.945 117.880 42.235 117.925 ;
        RECT 33.190 117.740 42.235 117.880 ;
        RECT 33.190 117.680 33.510 117.740 ;
        RECT 41.945 117.695 42.235 117.740 ;
        RECT 47.950 117.880 48.240 117.925 ;
        RECT 50.050 117.880 50.340 117.925 ;
        RECT 51.620 117.880 51.910 117.925 ;
        RECT 47.950 117.740 51.910 117.880 ;
        RECT 47.950 117.695 48.240 117.740 ;
        RECT 50.050 117.695 50.340 117.740 ;
        RECT 51.620 117.695 51.910 117.740 ;
        RECT 54.365 117.695 54.655 117.925 ;
        RECT 62.170 117.880 62.460 117.925 ;
        RECT 63.740 117.880 64.030 117.925 ;
        RECT 65.840 117.880 66.130 117.925 ;
        RECT 62.170 117.740 66.130 117.880 ;
        RECT 62.170 117.695 62.460 117.740 ;
        RECT 63.740 117.695 64.030 117.740 ;
        RECT 65.840 117.695 66.130 117.740 ;
        RECT 37.330 117.340 37.650 117.600 ;
        RECT 59.425 117.540 59.715 117.585 ;
        RECT 60.790 117.540 61.110 117.600 ;
        RECT 59.425 117.400 61.110 117.540 ;
        RECT 59.425 117.355 59.715 117.400 ;
        RECT 60.790 117.340 61.110 117.400 ;
        RECT 5.520 116.720 84.180 117.200 ;
        RECT 15.710 116.320 16.030 116.580 ;
        RECT 16.630 116.520 16.950 116.580 ;
        RECT 23.530 116.520 23.850 116.580 ;
        RECT 16.630 116.380 23.850 116.520 ;
        RECT 16.630 116.320 16.950 116.380 ;
        RECT 23.530 116.320 23.850 116.380 ;
        RECT 59.410 116.320 59.730 116.580 ;
        RECT 59.870 116.320 60.190 116.580 ;
        RECT 65.850 116.520 66.170 116.580 ;
        RECT 66.325 116.520 66.615 116.565 ;
        RECT 65.850 116.380 66.615 116.520 ;
        RECT 65.850 116.320 66.170 116.380 ;
        RECT 66.325 116.335 66.615 116.380 ;
        RECT 11.110 116.180 11.400 116.225 ;
        RECT 12.680 116.180 12.970 116.225 ;
        RECT 14.780 116.180 15.070 116.225 ;
        RECT 19.430 116.180 19.720 116.225 ;
        RECT 21.530 116.180 21.820 116.225 ;
        RECT 23.100 116.180 23.390 116.225 ;
        RECT 11.110 116.040 15.070 116.180 ;
        RECT 11.110 115.995 11.400 116.040 ;
        RECT 12.680 115.995 12.970 116.040 ;
        RECT 14.780 115.995 15.070 116.040 ;
        RECT 15.340 116.040 19.160 116.180 ;
        RECT 15.340 115.900 15.480 116.040 ;
        RECT 10.675 115.840 10.965 115.885 ;
        RECT 13.195 115.840 13.485 115.885 ;
        RECT 14.385 115.840 14.675 115.885 ;
        RECT 10.675 115.700 14.675 115.840 ;
        RECT 10.675 115.655 10.965 115.700 ;
        RECT 13.195 115.655 13.485 115.700 ;
        RECT 14.385 115.655 14.675 115.700 ;
        RECT 15.250 115.640 15.570 115.900 ;
        RECT 19.020 115.885 19.160 116.040 ;
        RECT 19.430 116.040 23.390 116.180 ;
        RECT 19.430 115.995 19.720 116.040 ;
        RECT 21.530 115.995 21.820 116.040 ;
        RECT 23.100 115.995 23.390 116.040 ;
        RECT 45.190 116.180 45.480 116.225 ;
        RECT 47.290 116.180 47.580 116.225 ;
        RECT 48.860 116.180 49.150 116.225 ;
        RECT 45.190 116.040 49.150 116.180 ;
        RECT 45.190 115.995 45.480 116.040 ;
        RECT 47.290 115.995 47.580 116.040 ;
        RECT 48.860 115.995 49.150 116.040 ;
        RECT 53.010 116.180 53.300 116.225 ;
        RECT 55.110 116.180 55.400 116.225 ;
        RECT 56.680 116.180 56.970 116.225 ;
        RECT 53.010 116.040 56.970 116.180 ;
        RECT 53.010 115.995 53.300 116.040 ;
        RECT 55.110 115.995 55.400 116.040 ;
        RECT 56.680 115.995 56.970 116.040 ;
        RECT 18.945 115.655 19.235 115.885 ;
        RECT 19.825 115.840 20.115 115.885 ;
        RECT 21.015 115.840 21.305 115.885 ;
        RECT 23.535 115.840 23.825 115.885 ;
        RECT 19.825 115.700 23.825 115.840 ;
        RECT 19.825 115.655 20.115 115.700 ;
        RECT 21.015 115.655 21.305 115.700 ;
        RECT 23.535 115.655 23.825 115.700 ;
        RECT 45.585 115.840 45.875 115.885 ;
        RECT 46.775 115.840 47.065 115.885 ;
        RECT 49.295 115.840 49.585 115.885 ;
        RECT 45.585 115.700 49.585 115.840 ;
        RECT 45.585 115.655 45.875 115.700 ;
        RECT 46.775 115.655 47.065 115.700 ;
        RECT 49.295 115.655 49.585 115.700 ;
        RECT 53.405 115.840 53.695 115.885 ;
        RECT 54.595 115.840 54.885 115.885 ;
        RECT 57.115 115.840 57.405 115.885 ;
        RECT 53.405 115.700 57.405 115.840 ;
        RECT 59.500 115.840 59.640 116.320 ;
        RECT 62.645 115.840 62.935 115.885 ;
        RECT 59.500 115.700 62.935 115.840 ;
        RECT 53.405 115.655 53.695 115.700 ;
        RECT 54.595 115.655 54.885 115.700 ;
        RECT 57.115 115.655 57.405 115.700 ;
        RECT 62.645 115.655 62.935 115.700 ;
        RECT 16.630 115.300 16.950 115.560 ;
        RECT 17.090 115.500 17.410 115.560 ;
        RECT 17.565 115.500 17.855 115.545 ;
        RECT 17.090 115.360 17.855 115.500 ;
        RECT 17.090 115.300 17.410 115.360 ;
        RECT 17.565 115.315 17.855 115.360 ;
        RECT 18.025 115.315 18.315 115.545 ;
        RECT 29.065 115.500 29.355 115.545 ;
        RECT 25.920 115.360 29.355 115.500 ;
        RECT 14.040 115.160 14.330 115.205 ;
        RECT 16.170 115.160 16.490 115.220 ;
        RECT 14.040 115.020 16.490 115.160 ;
        RECT 14.040 114.975 14.330 115.020 ;
        RECT 16.170 114.960 16.490 115.020 ;
        RECT 8.365 114.820 8.655 114.865 ;
        RECT 10.190 114.820 10.510 114.880 ;
        RECT 8.365 114.680 10.510 114.820 ;
        RECT 8.365 114.635 8.655 114.680 ;
        RECT 10.190 114.620 10.510 114.680 ;
        RECT 16.630 114.820 16.950 114.880 ;
        RECT 18.100 114.820 18.240 115.315 ;
        RECT 18.470 115.160 18.790 115.220 ;
        RECT 20.170 115.160 20.460 115.205 ;
        RECT 18.470 115.020 20.460 115.160 ;
        RECT 18.470 114.960 18.790 115.020 ;
        RECT 20.170 114.975 20.460 115.020 ;
        RECT 16.630 114.680 18.240 114.820 ;
        RECT 23.070 114.820 23.390 114.880 ;
        RECT 25.920 114.865 26.060 115.360 ;
        RECT 29.065 115.315 29.355 115.360 ;
        RECT 33.190 115.300 33.510 115.560 ;
        RECT 42.390 115.500 42.710 115.560 ;
        RECT 44.705 115.500 44.995 115.545 ;
        RECT 50.210 115.500 50.530 115.560 ;
        RECT 53.890 115.545 54.210 115.560 ;
        RECT 52.525 115.500 52.815 115.545 ;
        RECT 53.860 115.500 54.210 115.545 ;
        RECT 42.390 115.360 52.815 115.500 ;
        RECT 53.695 115.360 54.210 115.500 ;
        RECT 42.390 115.300 42.710 115.360 ;
        RECT 44.705 115.315 44.995 115.360 ;
        RECT 50.210 115.300 50.530 115.360 ;
        RECT 52.525 115.315 52.815 115.360 ;
        RECT 53.860 115.315 54.210 115.360 ;
        RECT 53.890 115.300 54.210 115.315 ;
        RECT 60.790 115.500 61.110 115.560 ;
        RECT 63.565 115.500 63.855 115.545 ;
        RECT 64.010 115.500 64.330 115.560 ;
        RECT 60.790 115.360 64.330 115.500 ;
        RECT 60.790 115.300 61.110 115.360 ;
        RECT 63.565 115.315 63.855 115.360 ;
        RECT 64.010 115.300 64.330 115.360 ;
        RECT 65.390 115.300 65.710 115.560 ;
        RECT 46.070 115.205 46.390 115.220 ;
        RECT 46.040 114.975 46.390 115.205 ;
        RECT 46.070 114.960 46.390 114.975 ;
        RECT 58.490 115.160 58.810 115.220 ;
        RECT 64.485 115.160 64.775 115.205 ;
        RECT 58.490 115.020 64.775 115.160 ;
        RECT 58.490 114.960 58.810 115.020 ;
        RECT 64.485 114.975 64.775 115.020 ;
        RECT 64.930 114.960 65.250 115.220 ;
        RECT 25.845 114.820 26.135 114.865 ;
        RECT 23.070 114.680 26.135 114.820 ;
        RECT 16.630 114.620 16.950 114.680 ;
        RECT 23.070 114.620 23.390 114.680 ;
        RECT 25.845 114.635 26.135 114.680 ;
        RECT 26.290 114.620 26.610 114.880 ;
        RECT 29.970 114.820 30.290 114.880 ;
        RECT 30.445 114.820 30.735 114.865 ;
        RECT 29.970 114.680 30.735 114.820 ;
        RECT 29.970 114.620 30.290 114.680 ;
        RECT 30.445 114.635 30.735 114.680 ;
        RECT 49.290 114.820 49.610 114.880 ;
        RECT 51.605 114.820 51.895 114.865 ;
        RECT 49.290 114.680 51.895 114.820 ;
        RECT 49.290 114.620 49.610 114.680 ;
        RECT 51.605 114.635 51.895 114.680 ;
        RECT 5.520 114.000 84.180 114.480 ;
        RECT 18.025 113.615 18.315 113.845 ;
        RECT 31.350 113.800 31.670 113.860 ;
        RECT 32.285 113.800 32.575 113.845 ;
        RECT 31.350 113.660 32.575 113.800 ;
        RECT 16.170 113.460 16.490 113.520 ;
        RECT 18.100 113.460 18.240 113.615 ;
        RECT 31.350 113.600 31.670 113.660 ;
        RECT 32.285 113.615 32.575 113.660 ;
        RECT 49.305 113.800 49.595 113.845 ;
        RECT 52.050 113.800 52.370 113.860 ;
        RECT 49.305 113.660 52.370 113.800 ;
        RECT 49.305 113.615 49.595 113.660 ;
        RECT 52.050 113.600 52.370 113.660 ;
        RECT 58.490 113.600 58.810 113.860 ;
        RECT 60.330 113.800 60.650 113.860 ;
        RECT 61.265 113.800 61.555 113.845 ;
        RECT 60.330 113.660 61.555 113.800 ;
        RECT 60.330 113.600 60.650 113.660 ;
        RECT 61.265 113.615 61.555 113.660 ;
        RECT 16.170 113.320 18.240 113.460 ;
        RECT 18.865 113.460 19.155 113.505 ;
        RECT 19.390 113.460 19.710 113.520 ;
        RECT 18.865 113.320 19.710 113.460 ;
        RECT 16.170 113.260 16.490 113.320 ;
        RECT 18.865 113.275 19.155 113.320 ;
        RECT 19.390 113.260 19.710 113.320 ;
        RECT 19.865 113.460 20.155 113.505 ;
        RECT 26.290 113.460 26.610 113.520 ;
        RECT 31.440 113.460 31.580 113.600 ;
        RECT 19.865 113.320 26.610 113.460 ;
        RECT 19.865 113.275 20.155 113.320 ;
        RECT 26.290 113.260 26.610 113.320 ;
        RECT 29.600 113.320 31.580 113.460 ;
        RECT 4.210 113.120 4.530 113.180 ;
        RECT 7.445 113.120 7.735 113.165 ;
        RECT 4.210 112.980 7.735 113.120 ;
        RECT 4.210 112.920 4.530 112.980 ;
        RECT 7.445 112.935 7.735 112.980 ;
        RECT 17.090 112.920 17.410 113.180 ;
        RECT 17.565 113.120 17.855 113.165 ;
        RECT 20.325 113.120 20.615 113.165 ;
        RECT 17.565 112.980 20.615 113.120 ;
        RECT 17.565 112.935 17.855 112.980 ;
        RECT 20.325 112.935 20.615 112.980 ;
        RECT 23.990 112.920 24.310 113.180 ;
        RECT 29.600 113.165 29.740 113.320 ;
        RECT 24.925 112.935 25.215 113.165 ;
        RECT 29.525 112.935 29.815 113.165 ;
        RECT 17.180 112.780 17.320 112.920 ;
        RECT 19.390 112.780 19.710 112.840 ;
        RECT 17.180 112.640 19.710 112.780 ;
        RECT 19.390 112.580 19.710 112.640 ;
        RECT 23.545 112.780 23.835 112.825 ;
        RECT 24.465 112.780 24.755 112.825 ;
        RECT 23.545 112.640 24.755 112.780 ;
        RECT 23.545 112.595 23.835 112.640 ;
        RECT 24.465 112.595 24.755 112.640 ;
        RECT 8.365 112.440 8.655 112.485 ;
        RECT 8.810 112.440 9.130 112.500 ;
        RECT 8.365 112.300 9.130 112.440 ;
        RECT 8.365 112.255 8.655 112.300 ;
        RECT 8.810 112.240 9.130 112.300 ;
        RECT 16.185 112.440 16.475 112.485 ;
        RECT 18.470 112.440 18.790 112.500 ;
        RECT 16.185 112.300 18.790 112.440 ;
        RECT 16.185 112.255 16.475 112.300 ;
        RECT 18.470 112.240 18.790 112.300 ;
        RECT 23.070 112.440 23.390 112.500 ;
        RECT 25.000 112.440 25.140 112.935 ;
        RECT 29.050 112.580 29.370 112.840 ;
        RECT 23.070 112.300 25.140 112.440 ;
        RECT 23.070 112.240 23.390 112.300 ;
        RECT 29.600 112.160 29.740 112.935 ;
        RECT 29.970 112.920 30.290 113.180 ;
        RECT 32.285 112.935 32.575 113.165 ;
        RECT 32.730 113.120 33.050 113.180 ;
        RECT 33.205 113.120 33.495 113.165 ;
        RECT 34.110 113.120 34.430 113.180 ;
        RECT 32.730 112.980 34.430 113.120 ;
        RECT 30.445 112.595 30.735 112.825 ;
        RECT 32.360 112.780 32.500 112.935 ;
        RECT 32.730 112.920 33.050 112.980 ;
        RECT 33.205 112.935 33.495 112.980 ;
        RECT 34.110 112.920 34.430 112.980 ;
        RECT 36.410 113.120 36.730 113.180 ;
        RECT 37.330 113.120 37.650 113.180 ;
        RECT 36.410 112.980 37.650 113.120 ;
        RECT 36.410 112.920 36.730 112.980 ;
        RECT 37.330 112.920 37.650 112.980 ;
        RECT 38.265 112.935 38.555 113.165 ;
        RECT 33.650 112.780 33.970 112.840 ;
        RECT 32.360 112.640 33.970 112.780 ;
        RECT 30.520 112.440 30.660 112.595 ;
        RECT 33.650 112.580 33.970 112.640 ;
        RECT 35.030 112.440 35.350 112.500 ;
        RECT 30.520 112.300 35.350 112.440 ;
        RECT 35.030 112.240 35.350 112.300 ;
        RECT 37.330 112.440 37.650 112.500 ;
        RECT 38.340 112.440 38.480 112.935 ;
        RECT 42.390 112.920 42.710 113.180 ;
        RECT 43.770 113.165 44.090 113.180 ;
        RECT 43.740 112.935 44.090 113.165 ;
        RECT 43.770 112.920 44.090 112.935 ;
        RECT 58.030 112.920 58.350 113.180 ;
        RECT 58.965 113.120 59.255 113.165 ;
        RECT 60.420 113.120 60.560 113.600 ;
        RECT 58.965 112.980 60.560 113.120 ;
        RECT 58.965 112.935 59.255 112.980 ;
        RECT 41.930 112.580 42.250 112.840 ;
        RECT 43.285 112.780 43.575 112.825 ;
        RECT 44.475 112.780 44.765 112.825 ;
        RECT 46.995 112.780 47.285 112.825 ;
        RECT 43.285 112.640 47.285 112.780 ;
        RECT 43.285 112.595 43.575 112.640 ;
        RECT 44.475 112.595 44.765 112.640 ;
        RECT 46.995 112.595 47.285 112.640 ;
        RECT 38.725 112.440 39.015 112.485 ;
        RECT 37.330 112.300 39.015 112.440 ;
        RECT 37.330 112.240 37.650 112.300 ;
        RECT 38.725 112.255 39.015 112.300 ;
        RECT 42.890 112.440 43.180 112.485 ;
        RECT 44.990 112.440 45.280 112.485 ;
        RECT 46.560 112.440 46.850 112.485 ;
        RECT 42.890 112.300 46.850 112.440 ;
        RECT 60.420 112.440 60.560 112.980 ;
        RECT 60.790 112.920 61.110 113.180 ;
        RECT 61.725 113.120 62.015 113.165 ;
        RECT 62.170 113.120 62.490 113.180 ;
        RECT 61.725 112.980 62.490 113.120 ;
        RECT 61.725 112.935 62.015 112.980 ;
        RECT 62.170 112.920 62.490 112.980 ;
        RECT 80.570 113.120 80.890 113.180 ;
        RECT 81.045 113.120 81.335 113.165 ;
        RECT 80.570 112.980 81.335 113.120 ;
        RECT 80.570 112.920 80.890 112.980 ;
        RECT 81.045 112.935 81.335 112.980 ;
        RECT 64.010 112.780 64.330 112.840 ;
        RECT 64.485 112.780 64.775 112.825 ;
        RECT 64.010 112.640 64.775 112.780 ;
        RECT 64.010 112.580 64.330 112.640 ;
        RECT 64.485 112.595 64.775 112.640 ;
        RECT 65.865 112.440 66.155 112.485 ;
        RECT 60.420 112.300 66.155 112.440 ;
        RECT 42.890 112.255 43.180 112.300 ;
        RECT 44.990 112.255 45.280 112.300 ;
        RECT 46.560 112.255 46.850 112.300 ;
        RECT 65.865 112.255 66.155 112.300 ;
        RECT 81.950 112.240 82.270 112.500 ;
        RECT 18.945 112.100 19.235 112.145 ;
        RECT 23.990 112.100 24.310 112.160 ;
        RECT 18.945 111.960 24.310 112.100 ;
        RECT 18.945 111.915 19.235 111.960 ;
        RECT 23.990 111.900 24.310 111.960 ;
        RECT 28.130 111.900 28.450 112.160 ;
        RECT 29.510 111.900 29.830 112.160 ;
        RECT 35.950 112.100 36.270 112.160 ;
        RECT 36.885 112.100 37.175 112.145 ;
        RECT 35.950 111.960 37.175 112.100 ;
        RECT 35.950 111.900 36.270 111.960 ;
        RECT 36.885 111.915 37.175 111.960 ;
        RECT 37.790 111.900 38.110 112.160 ;
        RECT 66.785 112.100 67.075 112.145 ;
        RECT 71.370 112.100 71.690 112.160 ;
        RECT 66.785 111.960 71.690 112.100 ;
        RECT 66.785 111.915 67.075 111.960 ;
        RECT 71.370 111.900 71.690 111.960 ;
        RECT 5.520 111.280 84.180 111.760 ;
        RECT 49.305 111.080 49.595 111.125 ;
        RECT 49.750 111.080 50.070 111.140 ;
        RECT 49.305 110.940 50.070 111.080 ;
        RECT 49.305 110.895 49.595 110.940 ;
        RECT 49.750 110.880 50.070 110.940 ;
        RECT 80.570 110.880 80.890 111.140 ;
        RECT 27.250 110.740 27.540 110.785 ;
        RECT 29.350 110.740 29.640 110.785 ;
        RECT 30.920 110.740 31.210 110.785 ;
        RECT 27.250 110.600 31.210 110.740 ;
        RECT 27.250 110.555 27.540 110.600 ;
        RECT 29.350 110.555 29.640 110.600 ;
        RECT 30.920 110.555 31.210 110.600 ;
        RECT 37.370 110.740 37.660 110.785 ;
        RECT 39.470 110.740 39.760 110.785 ;
        RECT 41.040 110.740 41.330 110.785 ;
        RECT 37.370 110.600 41.330 110.740 ;
        RECT 37.370 110.555 37.660 110.600 ;
        RECT 39.470 110.555 39.760 110.600 ;
        RECT 41.040 110.555 41.330 110.600 ;
        RECT 41.930 110.740 42.250 110.800 ;
        RECT 43.785 110.740 44.075 110.785 ;
        RECT 41.930 110.600 44.075 110.740 ;
        RECT 41.930 110.540 42.250 110.600 ;
        RECT 43.785 110.555 44.075 110.600 ;
        RECT 51.170 110.740 51.460 110.785 ;
        RECT 53.270 110.740 53.560 110.785 ;
        RECT 54.840 110.740 55.130 110.785 ;
        RECT 51.170 110.600 55.130 110.740 ;
        RECT 51.170 110.555 51.460 110.600 ;
        RECT 53.270 110.555 53.560 110.600 ;
        RECT 54.840 110.555 55.130 110.600 ;
        RECT 62.170 110.540 62.490 110.800 ;
        RECT 64.930 110.740 65.220 110.785 ;
        RECT 66.500 110.740 66.790 110.785 ;
        RECT 68.600 110.740 68.890 110.785 ;
        RECT 64.930 110.600 68.890 110.740 ;
        RECT 64.930 110.555 65.220 110.600 ;
        RECT 66.500 110.555 66.790 110.600 ;
        RECT 68.600 110.555 68.890 110.600 ;
        RECT 27.645 110.400 27.935 110.445 ;
        RECT 28.835 110.400 29.125 110.445 ;
        RECT 31.355 110.400 31.645 110.445 ;
        RECT 27.645 110.260 31.645 110.400 ;
        RECT 27.645 110.215 27.935 110.260 ;
        RECT 28.835 110.215 29.125 110.260 ;
        RECT 31.355 110.215 31.645 110.260 ;
        RECT 36.870 110.200 37.190 110.460 ;
        RECT 37.765 110.400 38.055 110.445 ;
        RECT 38.955 110.400 39.245 110.445 ;
        RECT 41.475 110.400 41.765 110.445 ;
        RECT 37.765 110.260 41.765 110.400 ;
        RECT 37.765 110.215 38.055 110.260 ;
        RECT 38.955 110.215 39.245 110.260 ;
        RECT 41.475 110.215 41.765 110.260 ;
        RECT 4.210 110.060 4.530 110.120 ;
        RECT 6.985 110.060 7.275 110.105 ;
        RECT 4.210 109.920 7.275 110.060 ;
        RECT 4.210 109.860 4.530 109.920 ;
        RECT 6.985 109.875 7.275 109.920 ;
        RECT 8.365 110.060 8.655 110.105 ;
        RECT 9.270 110.060 9.590 110.120 ;
        RECT 13.870 110.060 14.190 110.120 ;
        RECT 14.345 110.060 14.635 110.105 ;
        RECT 8.365 109.920 12.720 110.060 ;
        RECT 8.365 109.875 8.655 109.920 ;
        RECT 9.270 109.860 9.590 109.920 ;
        RECT 0.530 109.720 0.850 109.780 ;
        RECT 12.580 109.720 12.720 109.920 ;
        RECT 13.870 109.920 14.635 110.060 ;
        RECT 13.870 109.860 14.190 109.920 ;
        RECT 14.345 109.875 14.635 109.920 ;
        RECT 15.250 110.060 15.570 110.120 ;
        RECT 23.530 110.060 23.850 110.120 ;
        RECT 26.765 110.060 27.055 110.105 ;
        RECT 15.250 109.920 27.055 110.060 ;
        RECT 15.250 109.860 15.570 109.920 ;
        RECT 23.530 109.860 23.850 109.920 ;
        RECT 26.765 109.875 27.055 109.920 ;
        RECT 27.760 109.920 34.800 110.060 ;
        RECT 18.930 109.720 19.250 109.780 ;
        RECT 27.760 109.720 27.900 109.920 ;
        RECT 0.530 109.580 12.260 109.720 ;
        RECT 12.580 109.580 27.900 109.720 ;
        RECT 28.100 109.720 28.390 109.765 ;
        RECT 34.125 109.720 34.415 109.765 ;
        RECT 28.100 109.580 34.415 109.720 ;
        RECT 0.530 109.520 0.850 109.580 ;
        RECT 11.570 109.180 11.890 109.440 ;
        RECT 12.120 109.380 12.260 109.580 ;
        RECT 18.930 109.520 19.250 109.580 ;
        RECT 28.100 109.535 28.390 109.580 ;
        RECT 34.125 109.535 34.415 109.580 ;
        RECT 29.050 109.380 29.370 109.440 ;
        RECT 12.120 109.240 29.370 109.380 ;
        RECT 29.050 109.180 29.370 109.240 ;
        RECT 32.730 109.380 33.050 109.440 ;
        RECT 33.650 109.380 33.970 109.440 ;
        RECT 32.730 109.240 33.970 109.380 ;
        RECT 34.660 109.380 34.800 109.920 ;
        RECT 35.030 109.860 35.350 110.120 ;
        RECT 35.950 109.860 36.270 110.120 ;
        RECT 36.410 110.060 36.730 110.120 ;
        RECT 42.020 110.060 42.160 110.540 ;
        RECT 50.210 110.400 50.530 110.460 ;
        RECT 50.685 110.400 50.975 110.445 ;
        RECT 50.210 110.260 50.975 110.400 ;
        RECT 50.210 110.200 50.530 110.260 ;
        RECT 50.685 110.215 50.975 110.260 ;
        RECT 51.565 110.400 51.855 110.445 ;
        RECT 52.755 110.400 53.045 110.445 ;
        RECT 55.275 110.400 55.565 110.445 ;
        RECT 51.565 110.260 55.565 110.400 ;
        RECT 51.565 110.215 51.855 110.260 ;
        RECT 52.755 110.215 53.045 110.260 ;
        RECT 55.275 110.215 55.565 110.260 ;
        RECT 64.495 110.400 64.785 110.445 ;
        RECT 67.015 110.400 67.305 110.445 ;
        RECT 68.205 110.400 68.495 110.445 ;
        RECT 64.495 110.260 68.495 110.400 ;
        RECT 64.495 110.215 64.785 110.260 ;
        RECT 67.015 110.215 67.305 110.260 ;
        RECT 68.205 110.215 68.495 110.260 ;
        RECT 36.410 109.920 36.910 110.060 ;
        RECT 37.880 109.920 42.160 110.060 ;
        RECT 36.410 109.860 36.730 109.920 ;
        RECT 36.870 109.720 37.190 109.780 ;
        RECT 37.880 109.720 38.020 109.920 ;
        RECT 47.465 109.875 47.755 110.105 ;
        RECT 56.650 110.060 56.970 110.120 ;
        RECT 58.045 110.060 58.335 110.105 ;
        RECT 56.650 109.920 58.335 110.060 ;
        RECT 38.250 109.765 38.570 109.780 ;
        RECT 36.870 109.580 38.020 109.720 ;
        RECT 36.870 109.520 37.190 109.580 ;
        RECT 38.220 109.535 38.570 109.765 ;
        RECT 38.250 109.520 38.570 109.535 ;
        RECT 47.540 109.380 47.680 109.875 ;
        RECT 56.650 109.860 56.970 109.920 ;
        RECT 58.045 109.875 58.335 109.920 ;
        RECT 58.965 109.875 59.255 110.105 ;
        RECT 61.725 110.060 62.015 110.105 ;
        RECT 62.630 110.060 62.950 110.120 ;
        RECT 64.930 110.060 65.250 110.120 ;
        RECT 61.725 109.920 65.250 110.060 ;
        RECT 61.725 109.875 62.015 109.920 ;
        RECT 49.290 109.520 49.610 109.780 ;
        RECT 52.020 109.720 52.310 109.765 ;
        RECT 58.505 109.720 58.795 109.765 ;
        RECT 52.020 109.580 58.795 109.720 ;
        RECT 59.040 109.720 59.180 109.875 ;
        RECT 62.630 109.860 62.950 109.920 ;
        RECT 64.930 109.860 65.250 109.920 ;
        RECT 69.070 110.060 69.390 110.120 ;
        RECT 71.830 110.060 72.150 110.120 ;
        RECT 69.070 109.920 72.150 110.060 ;
        RECT 69.070 109.860 69.390 109.920 ;
        RECT 71.830 109.860 72.150 109.920 ;
        RECT 79.650 109.860 79.970 110.120 ;
        RECT 80.570 110.060 80.890 110.120 ;
        RECT 81.045 110.060 81.335 110.105 ;
        RECT 80.570 109.920 81.335 110.060 ;
        RECT 80.570 109.860 80.890 109.920 ;
        RECT 81.045 109.875 81.335 109.920 ;
        RECT 63.090 109.720 63.410 109.780 ;
        RECT 59.040 109.580 63.410 109.720 ;
        RECT 52.020 109.535 52.310 109.580 ;
        RECT 58.505 109.535 58.795 109.580 ;
        RECT 63.090 109.520 63.410 109.580 ;
        RECT 66.770 109.720 67.090 109.780 ;
        RECT 67.750 109.720 68.040 109.765 ;
        RECT 66.770 109.580 68.040 109.720 ;
        RECT 66.770 109.520 67.090 109.580 ;
        RECT 67.750 109.535 68.040 109.580 ;
        RECT 48.370 109.380 48.690 109.440 ;
        RECT 34.660 109.240 48.690 109.380 ;
        RECT 32.730 109.180 33.050 109.240 ;
        RECT 33.650 109.180 33.970 109.240 ;
        RECT 48.370 109.180 48.690 109.240 ;
        RECT 50.225 109.380 50.515 109.425 ;
        RECT 57.110 109.380 57.430 109.440 ;
        RECT 50.225 109.240 57.430 109.380 ;
        RECT 50.225 109.195 50.515 109.240 ;
        RECT 57.110 109.180 57.430 109.240 ;
        RECT 57.585 109.380 57.875 109.425 ;
        RECT 58.950 109.380 59.270 109.440 ;
        RECT 60.790 109.380 61.110 109.440 ;
        RECT 57.585 109.240 61.110 109.380 ;
        RECT 57.585 109.195 57.875 109.240 ;
        RECT 58.950 109.180 59.270 109.240 ;
        RECT 60.790 109.180 61.110 109.240 ;
        RECT 61.250 109.380 61.570 109.440 ;
        RECT 66.310 109.380 66.630 109.440 ;
        RECT 61.250 109.240 66.630 109.380 ;
        RECT 61.250 109.180 61.570 109.240 ;
        RECT 66.310 109.180 66.630 109.240 ;
        RECT 81.950 109.180 82.270 109.440 ;
        RECT 5.520 108.560 84.180 109.040 ;
        RECT 13.425 108.360 13.715 108.405 ;
        RECT 14.330 108.360 14.650 108.420 ;
        RECT 13.425 108.220 14.650 108.360 ;
        RECT 13.425 108.175 13.715 108.220 ;
        RECT 14.330 108.160 14.650 108.220 ;
        RECT 15.250 108.160 15.570 108.420 ;
        RECT 30.445 108.360 30.735 108.405 ;
        RECT 35.030 108.360 35.350 108.420 ;
        RECT 30.445 108.220 32.960 108.360 ;
        RECT 30.445 108.175 30.735 108.220 ;
        RECT 15.340 108.020 15.480 108.160 ;
        RECT 13.960 107.880 15.480 108.020 ;
        RECT 24.880 108.020 25.170 108.065 ;
        RECT 28.130 108.020 28.450 108.080 ;
        RECT 24.880 107.880 28.450 108.020 ;
        RECT 13.960 107.740 14.100 107.880 ;
        RECT 24.880 107.835 25.170 107.880 ;
        RECT 28.130 107.820 28.450 107.880 ;
        RECT 8.365 107.680 8.655 107.725 ;
        RECT 8.810 107.680 9.130 107.740 ;
        RECT 8.365 107.540 9.130 107.680 ;
        RECT 8.365 107.495 8.655 107.540 ;
        RECT 8.810 107.480 9.130 107.540 ;
        RECT 10.190 107.480 10.510 107.740 ;
        RECT 13.870 107.480 14.190 107.740 ;
        RECT 15.250 107.725 15.570 107.740 ;
        RECT 15.220 107.495 15.570 107.725 ;
        RECT 15.250 107.480 15.570 107.495 ;
        RECT 19.390 107.680 19.710 107.740 ;
        RECT 21.245 107.680 21.535 107.725 ;
        RECT 19.390 107.540 21.535 107.680 ;
        RECT 19.390 107.480 19.710 107.540 ;
        RECT 21.245 107.495 21.535 107.540 ;
        RECT 22.165 107.680 22.455 107.725 ;
        RECT 23.070 107.680 23.390 107.740 ;
        RECT 22.165 107.540 23.390 107.680 ;
        RECT 22.165 107.495 22.455 107.540 ;
        RECT 23.070 107.480 23.390 107.540 ;
        RECT 23.530 107.480 23.850 107.740 ;
        RECT 28.590 107.680 28.910 107.740 ;
        RECT 32.820 107.725 32.960 108.220 ;
        RECT 35.030 108.220 36.180 108.360 ;
        RECT 35.030 108.160 35.350 108.220 ;
        RECT 33.650 108.020 33.970 108.080 ;
        RECT 35.505 108.020 35.795 108.065 ;
        RECT 33.650 107.880 35.795 108.020 ;
        RECT 36.040 108.020 36.180 108.220 ;
        RECT 38.250 108.160 38.570 108.420 ;
        RECT 56.650 108.160 56.970 108.420 ;
        RECT 57.110 108.360 57.430 108.420 ;
        RECT 59.425 108.360 59.715 108.405 ;
        RECT 57.110 108.220 59.715 108.360 ;
        RECT 57.110 108.160 57.430 108.220 ;
        RECT 59.425 108.175 59.715 108.220 ;
        RECT 60.805 108.175 61.095 108.405 ;
        RECT 62.185 108.360 62.475 108.405 ;
        RECT 62.630 108.360 62.950 108.420 ;
        RECT 62.185 108.220 62.950 108.360 ;
        RECT 62.185 108.175 62.475 108.220 ;
        RECT 39.185 108.020 39.475 108.065 ;
        RECT 36.040 107.880 39.475 108.020 ;
        RECT 33.650 107.820 33.970 107.880 ;
        RECT 35.505 107.835 35.795 107.880 ;
        RECT 39.185 107.835 39.475 107.880 ;
        RECT 31.825 107.680 32.115 107.725 ;
        RECT 28.590 107.540 32.115 107.680 ;
        RECT 28.590 107.480 28.910 107.540 ;
        RECT 31.825 107.495 32.115 107.540 ;
        RECT 32.745 107.680 33.035 107.725 ;
        RECT 33.190 107.680 33.510 107.740 ;
        RECT 32.745 107.540 33.510 107.680 ;
        RECT 32.745 107.495 33.035 107.540 ;
        RECT 33.190 107.480 33.510 107.540 ;
        RECT 34.570 107.680 34.890 107.740 ;
        RECT 36.410 107.680 36.730 107.740 ;
        RECT 34.570 107.540 36.730 107.680 ;
        RECT 34.570 107.480 34.890 107.540 ;
        RECT 36.410 107.480 36.730 107.540 ;
        RECT 36.885 107.680 37.175 107.725 ;
        RECT 37.330 107.680 37.650 107.740 ;
        RECT 36.885 107.540 37.650 107.680 ;
        RECT 36.885 107.495 37.175 107.540 ;
        RECT 37.330 107.480 37.650 107.540 ;
        RECT 38.725 107.495 39.015 107.725 ;
        RECT 9.730 107.140 10.050 107.400 ;
        RECT 14.765 107.340 15.055 107.385 ;
        RECT 15.955 107.340 16.245 107.385 ;
        RECT 18.475 107.340 18.765 107.385 ;
        RECT 14.765 107.200 18.765 107.340 ;
        RECT 14.765 107.155 15.055 107.200 ;
        RECT 15.955 107.155 16.245 107.200 ;
        RECT 18.475 107.155 18.765 107.200 ;
        RECT 24.425 107.340 24.715 107.385 ;
        RECT 25.615 107.340 25.905 107.385 ;
        RECT 28.135 107.340 28.425 107.385 ;
        RECT 24.425 107.200 28.425 107.340 ;
        RECT 24.425 107.155 24.715 107.200 ;
        RECT 25.615 107.155 25.905 107.200 ;
        RECT 28.135 107.155 28.425 107.200 ;
        RECT 37.790 107.340 38.110 107.400 ;
        RECT 38.265 107.340 38.555 107.385 ;
        RECT 37.790 107.200 38.555 107.340 ;
        RECT 37.790 107.140 38.110 107.200 ;
        RECT 38.265 107.155 38.555 107.200 ;
        RECT 8.825 107.000 9.115 107.045 ;
        RECT 14.370 107.000 14.660 107.045 ;
        RECT 16.470 107.000 16.760 107.045 ;
        RECT 18.040 107.000 18.330 107.045 ;
        RECT 8.825 106.860 13.870 107.000 ;
        RECT 8.825 106.815 9.115 106.860 ;
        RECT 9.285 106.660 9.575 106.705 ;
        RECT 10.650 106.660 10.970 106.720 ;
        RECT 9.285 106.520 10.970 106.660 ;
        RECT 13.730 106.660 13.870 106.860 ;
        RECT 14.370 106.860 18.330 107.000 ;
        RECT 14.370 106.815 14.660 106.860 ;
        RECT 16.470 106.815 16.760 106.860 ;
        RECT 18.040 106.815 18.330 106.860 ;
        RECT 24.030 107.000 24.320 107.045 ;
        RECT 26.130 107.000 26.420 107.045 ;
        RECT 27.700 107.000 27.990 107.045 ;
        RECT 24.030 106.860 27.990 107.000 ;
        RECT 24.030 106.815 24.320 106.860 ;
        RECT 26.130 106.815 26.420 106.860 ;
        RECT 27.700 106.815 27.990 106.860 ;
        RECT 33.665 107.000 33.955 107.045 ;
        RECT 38.800 107.000 38.940 107.495 ;
        RECT 48.370 107.480 48.690 107.740 ;
        RECT 49.290 107.480 49.610 107.740 ;
        RECT 49.750 107.480 50.070 107.740 ;
        RECT 55.730 107.480 56.050 107.740 ;
        RECT 59.500 107.680 59.640 108.175 ;
        RECT 60.880 108.020 61.020 108.175 ;
        RECT 62.630 108.160 62.950 108.220 ;
        RECT 63.090 108.020 63.410 108.080 ;
        RECT 65.390 108.020 65.710 108.080 ;
        RECT 65.865 108.020 66.155 108.065 ;
        RECT 60.880 107.880 66.155 108.020 ;
        RECT 63.090 107.820 63.410 107.880 ;
        RECT 65.390 107.820 65.710 107.880 ;
        RECT 65.865 107.835 66.155 107.880 ;
        RECT 61.710 107.680 62.030 107.740 ;
        RECT 59.500 107.540 62.030 107.680 ;
        RECT 61.710 107.480 62.030 107.540 ;
        RECT 67.230 107.680 67.550 107.740 ;
        RECT 67.705 107.680 67.995 107.725 ;
        RECT 67.230 107.540 67.995 107.680 ;
        RECT 67.230 107.480 67.550 107.540 ;
        RECT 67.705 107.495 67.995 107.540 ;
        RECT 71.830 107.480 72.150 107.740 ;
        RECT 73.210 107.725 73.530 107.740 ;
        RECT 73.180 107.495 73.530 107.725 ;
        RECT 73.210 107.480 73.530 107.495 ;
        RECT 48.830 107.340 49.150 107.400 ;
        RECT 49.840 107.340 49.980 107.480 ;
        RECT 48.830 107.200 49.980 107.340 ;
        RECT 54.365 107.340 54.655 107.385 ;
        RECT 57.585 107.340 57.875 107.385 ;
        RECT 54.365 107.200 57.875 107.340 ;
        RECT 48.830 107.140 49.150 107.200 ;
        RECT 54.365 107.155 54.655 107.200 ;
        RECT 57.585 107.155 57.875 107.200 ;
        RECT 33.665 106.860 38.940 107.000 ;
        RECT 51.605 107.000 51.895 107.045 ;
        RECT 54.825 107.000 55.115 107.045 ;
        RECT 56.190 107.000 56.510 107.060 ;
        RECT 51.605 106.860 56.510 107.000 ;
        RECT 57.660 107.000 57.800 107.155 ;
        RECT 58.950 107.140 59.270 107.400 ;
        RECT 59.870 107.385 60.190 107.400 ;
        RECT 59.870 107.155 60.300 107.385 ;
        RECT 64.945 107.155 65.235 107.385 ;
        RECT 66.310 107.340 66.630 107.400 ;
        RECT 66.785 107.340 67.075 107.385 ;
        RECT 66.310 107.200 67.075 107.340 ;
        RECT 59.870 107.140 60.190 107.155 ;
        RECT 60.790 107.000 61.110 107.060 ;
        RECT 57.660 106.860 61.110 107.000 ;
        RECT 33.665 106.815 33.955 106.860 ;
        RECT 51.605 106.815 51.895 106.860 ;
        RECT 54.825 106.815 55.115 106.860 ;
        RECT 56.190 106.800 56.510 106.860 ;
        RECT 60.790 106.800 61.110 106.860 ;
        RECT 62.630 107.000 62.950 107.060 ;
        RECT 64.470 107.000 64.790 107.060 ;
        RECT 65.020 107.000 65.160 107.155 ;
        RECT 66.310 107.140 66.630 107.200 ;
        RECT 66.785 107.155 67.075 107.200 ;
        RECT 72.725 107.340 73.015 107.385 ;
        RECT 73.915 107.340 74.205 107.385 ;
        RECT 76.435 107.340 76.725 107.385 ;
        RECT 79.650 107.340 79.970 107.400 ;
        RECT 81.965 107.340 82.255 107.385 ;
        RECT 72.725 107.200 76.725 107.340 ;
        RECT 72.725 107.155 73.015 107.200 ;
        RECT 73.915 107.155 74.205 107.200 ;
        RECT 76.435 107.155 76.725 107.200 ;
        RECT 78.820 107.200 82.255 107.340 ;
        RECT 67.245 107.000 67.535 107.045 ;
        RECT 70.910 107.000 71.230 107.060 ;
        RECT 78.820 107.045 78.960 107.200 ;
        RECT 79.650 107.140 79.970 107.200 ;
        RECT 81.965 107.155 82.255 107.200 ;
        RECT 62.630 106.860 65.160 107.000 ;
        RECT 66.400 106.860 71.230 107.000 ;
        RECT 62.630 106.800 62.950 106.860 ;
        RECT 64.470 106.800 64.790 106.860 ;
        RECT 19.850 106.660 20.170 106.720 ;
        RECT 13.730 106.520 20.170 106.660 ;
        RECT 9.285 106.475 9.575 106.520 ;
        RECT 10.650 106.460 10.970 106.520 ;
        RECT 19.850 106.460 20.170 106.520 ;
        RECT 20.310 106.660 20.630 106.720 ;
        RECT 20.785 106.660 21.075 106.705 ;
        RECT 20.310 106.520 21.075 106.660 ;
        RECT 20.310 106.460 20.630 106.520 ;
        RECT 20.785 106.475 21.075 106.520 ;
        RECT 21.245 106.660 21.535 106.705 ;
        RECT 32.270 106.660 32.590 106.720 ;
        RECT 21.245 106.520 32.590 106.660 ;
        RECT 21.245 106.475 21.535 106.520 ;
        RECT 32.270 106.460 32.590 106.520 ;
        RECT 32.730 106.460 33.050 106.720 ;
        RECT 36.425 106.660 36.715 106.705 ;
        RECT 36.870 106.660 37.190 106.720 ;
        RECT 37.345 106.660 37.635 106.705 ;
        RECT 36.425 106.520 37.635 106.660 ;
        RECT 36.425 106.475 36.715 106.520 ;
        RECT 36.870 106.460 37.190 106.520 ;
        RECT 37.345 106.475 37.635 106.520 ;
        RECT 58.030 106.660 58.350 106.720 ;
        RECT 66.400 106.660 66.540 106.860 ;
        RECT 67.245 106.815 67.535 106.860 ;
        RECT 70.910 106.800 71.230 106.860 ;
        RECT 72.330 107.000 72.620 107.045 ;
        RECT 74.430 107.000 74.720 107.045 ;
        RECT 76.000 107.000 76.290 107.045 ;
        RECT 72.330 106.860 76.290 107.000 ;
        RECT 72.330 106.815 72.620 106.860 ;
        RECT 74.430 106.815 74.720 106.860 ;
        RECT 76.000 106.815 76.290 106.860 ;
        RECT 78.745 106.815 79.035 107.045 ;
        RECT 58.030 106.520 66.540 106.660 ;
        RECT 58.030 106.460 58.350 106.520 ;
        RECT 66.770 106.460 67.090 106.720 ;
        RECT 79.190 106.460 79.510 106.720 ;
        RECT 5.520 105.840 84.180 106.320 ;
        RECT 13.410 105.640 13.730 105.700 ;
        RECT 13.885 105.640 14.175 105.685 ;
        RECT 13.410 105.500 14.175 105.640 ;
        RECT 13.410 105.440 13.730 105.500 ;
        RECT 13.885 105.455 14.175 105.500 ;
        RECT 15.250 105.440 15.570 105.700 ;
        RECT 16.185 105.640 16.475 105.685 ;
        RECT 19.390 105.640 19.710 105.700 ;
        RECT 16.185 105.500 19.710 105.640 ;
        RECT 16.185 105.455 16.475 105.500 ;
        RECT 7.470 105.300 7.760 105.345 ;
        RECT 9.570 105.300 9.860 105.345 ;
        RECT 11.140 105.300 11.430 105.345 ;
        RECT 7.470 105.160 11.430 105.300 ;
        RECT 7.470 105.115 7.760 105.160 ;
        RECT 9.570 105.115 9.860 105.160 ;
        RECT 11.140 105.115 11.430 105.160 ;
        RECT 14.805 105.300 15.095 105.345 ;
        RECT 16.260 105.300 16.400 105.455 ;
        RECT 19.390 105.440 19.710 105.500 ;
        RECT 19.850 105.640 20.170 105.700 ;
        RECT 23.085 105.640 23.375 105.685 ;
        RECT 19.850 105.500 23.375 105.640 ;
        RECT 19.850 105.440 20.170 105.500 ;
        RECT 23.085 105.455 23.375 105.500 ;
        RECT 24.005 105.455 24.295 105.685 ;
        RECT 28.590 105.640 28.910 105.700 ;
        RECT 29.065 105.640 29.355 105.685 ;
        RECT 28.590 105.500 29.355 105.640 ;
        RECT 18.470 105.300 18.790 105.360 ;
        RECT 20.310 105.300 20.630 105.360 ;
        RECT 24.080 105.300 24.220 105.455 ;
        RECT 28.590 105.440 28.910 105.500 ;
        RECT 29.065 105.455 29.355 105.500 ;
        RECT 31.365 105.640 31.655 105.685 ;
        RECT 34.570 105.640 34.890 105.700 ;
        RECT 31.365 105.500 34.890 105.640 ;
        RECT 31.365 105.455 31.655 105.500 ;
        RECT 34.570 105.440 34.890 105.500 ;
        RECT 42.865 105.455 43.155 105.685 ;
        RECT 14.805 105.160 16.400 105.300 ;
        RECT 17.640 105.160 24.220 105.300 ;
        RECT 14.805 105.115 15.095 105.160 ;
        RECT 7.865 104.960 8.155 105.005 ;
        RECT 9.055 104.960 9.345 105.005 ;
        RECT 11.575 104.960 11.865 105.005 ;
        RECT 7.865 104.820 11.865 104.960 ;
        RECT 7.865 104.775 8.155 104.820 ;
        RECT 9.055 104.775 9.345 104.820 ;
        RECT 11.575 104.775 11.865 104.820 ;
        RECT 15.710 104.760 16.030 105.020 ;
        RECT 6.985 104.620 7.275 104.665 ;
        RECT 13.870 104.620 14.190 104.680 ;
        RECT 6.985 104.480 14.190 104.620 ;
        RECT 6.985 104.435 7.275 104.480 ;
        RECT 13.870 104.420 14.190 104.480 ;
        RECT 14.345 104.620 14.635 104.665 ;
        RECT 14.790 104.620 15.110 104.680 ;
        RECT 16.630 104.620 16.950 104.680 ;
        RECT 14.345 104.480 16.950 104.620 ;
        RECT 14.345 104.435 14.635 104.480 ;
        RECT 14.790 104.420 15.110 104.480 ;
        RECT 16.630 104.420 16.950 104.480 ;
        RECT 17.105 104.630 17.395 104.665 ;
        RECT 17.640 104.630 17.780 105.160 ;
        RECT 18.470 105.100 18.790 105.160 ;
        RECT 20.310 105.100 20.630 105.160 ;
        RECT 28.680 104.960 28.820 105.440 ;
        RECT 31.810 105.300 32.130 105.360 ;
        RECT 32.285 105.300 32.575 105.345 ;
        RECT 31.810 105.160 32.575 105.300 ;
        RECT 31.810 105.100 32.130 105.160 ;
        RECT 32.285 105.115 32.575 105.160 ;
        RECT 32.730 105.300 33.050 105.360 ;
        RECT 42.940 105.300 43.080 105.455 ;
        RECT 51.130 105.440 51.450 105.700 ;
        RECT 55.730 105.640 56.050 105.700 ;
        RECT 57.570 105.640 57.890 105.700 ;
        RECT 58.965 105.640 59.255 105.685 ;
        RECT 55.730 105.500 59.255 105.640 ;
        RECT 55.730 105.440 56.050 105.500 ;
        RECT 57.570 105.440 57.890 105.500 ;
        RECT 58.965 105.455 59.255 105.500 ;
        RECT 61.250 105.640 61.570 105.700 ;
        RECT 62.185 105.640 62.475 105.685 ;
        RECT 61.250 105.500 62.475 105.640 ;
        RECT 49.290 105.300 49.610 105.360 ;
        RECT 32.730 105.160 49.610 105.300 ;
        RECT 32.730 105.100 33.050 105.160 ;
        RECT 49.290 105.100 49.610 105.160 ;
        RECT 18.100 104.820 25.140 104.960 ;
        RECT 18.100 104.680 18.240 104.820 ;
        RECT 17.105 104.490 17.780 104.630 ;
        RECT 17.105 104.435 17.395 104.490 ;
        RECT 18.010 104.420 18.330 104.680 ;
        RECT 20.785 104.620 21.075 104.665 ;
        RECT 22.625 104.620 22.915 104.665 ;
        RECT 18.560 104.480 21.075 104.620 ;
        RECT 7.430 104.280 7.750 104.340 ;
        RECT 8.210 104.280 8.500 104.325 ;
        RECT 7.430 104.140 8.500 104.280 ;
        RECT 7.430 104.080 7.750 104.140 ;
        RECT 8.210 104.095 8.500 104.140 ;
        RECT 8.810 104.280 9.130 104.340 ;
        RECT 18.560 104.280 18.700 104.480 ;
        RECT 20.785 104.435 21.075 104.480 ;
        RECT 21.320 104.480 22.915 104.620 ;
        RECT 8.810 104.140 18.700 104.280 ;
        RECT 8.810 104.080 9.130 104.140 ;
        RECT 18.560 103.940 18.700 104.140 ;
        RECT 18.930 104.280 19.250 104.340 ;
        RECT 21.320 104.280 21.460 104.480 ;
        RECT 22.625 104.435 22.915 104.480 ;
        RECT 23.070 104.620 23.390 104.680 ;
        RECT 25.000 104.665 25.140 104.820 ;
        RECT 27.760 104.820 28.820 104.960 ;
        RECT 29.050 104.960 29.370 105.020 ;
        RECT 59.040 104.960 59.180 105.455 ;
        RECT 61.250 105.440 61.570 105.500 ;
        RECT 62.185 105.455 62.475 105.500 ;
        RECT 64.470 105.440 64.790 105.700 ;
        RECT 65.390 105.640 65.710 105.700 ;
        RECT 67.230 105.640 67.550 105.700 ;
        RECT 65.390 105.500 67.550 105.640 ;
        RECT 65.390 105.440 65.710 105.500 ;
        RECT 67.230 105.440 67.550 105.500 ;
        RECT 73.210 105.640 73.530 105.700 ;
        RECT 74.145 105.640 74.435 105.685 ;
        RECT 73.210 105.500 74.435 105.640 ;
        RECT 73.210 105.440 73.530 105.500 ;
        RECT 74.145 105.455 74.435 105.500 ;
        RECT 80.570 105.440 80.890 105.700 ;
        RECT 60.790 105.300 61.110 105.360 ;
        RECT 64.010 105.300 64.330 105.360 ;
        RECT 66.325 105.300 66.615 105.345 ;
        RECT 67.690 105.300 68.010 105.360 ;
        RECT 60.790 105.160 65.160 105.300 ;
        RECT 60.790 105.100 61.110 105.160 ;
        RECT 64.010 105.100 64.330 105.160 ;
        RECT 65.020 105.005 65.160 105.160 ;
        RECT 66.325 105.160 70.680 105.300 ;
        RECT 66.325 105.115 66.615 105.160 ;
        RECT 67.690 105.100 68.010 105.160 ;
        RECT 29.050 104.820 44.920 104.960 ;
        RECT 59.040 104.820 64.700 104.960 ;
        RECT 27.760 104.665 27.900 104.820 ;
        RECT 29.050 104.760 29.370 104.820 ;
        RECT 24.005 104.620 24.295 104.665 ;
        RECT 23.070 104.480 24.295 104.620 ;
        RECT 23.070 104.420 23.390 104.480 ;
        RECT 24.005 104.435 24.295 104.480 ;
        RECT 24.925 104.435 25.215 104.665 ;
        RECT 27.685 104.435 27.975 104.665 ;
        RECT 28.605 104.620 28.895 104.665 ;
        RECT 29.510 104.620 29.830 104.680 ;
        RECT 28.605 104.480 29.830 104.620 ;
        RECT 28.605 104.435 28.895 104.480 ;
        RECT 29.510 104.420 29.830 104.480 ;
        RECT 30.445 104.435 30.735 104.665 ;
        RECT 31.825 104.620 32.115 104.665 ;
        RECT 34.110 104.620 34.430 104.680 ;
        RECT 31.825 104.480 34.430 104.620 ;
        RECT 31.825 104.435 32.115 104.480 ;
        RECT 18.930 104.140 21.460 104.280 ;
        RECT 21.835 104.280 22.125 104.325 ;
        RECT 23.530 104.280 23.850 104.340 ;
        RECT 30.520 104.280 30.660 104.435 ;
        RECT 34.110 104.420 34.430 104.480 ;
        RECT 35.045 104.435 35.335 104.665 ;
        RECT 30.890 104.280 31.210 104.340 ;
        RECT 35.120 104.280 35.260 104.435 ;
        RECT 36.410 104.420 36.730 104.680 ;
        RECT 36.885 104.620 37.175 104.665 ;
        RECT 37.330 104.620 37.650 104.680 ;
        RECT 36.885 104.480 37.650 104.620 ;
        RECT 36.885 104.435 37.175 104.480 ;
        RECT 37.330 104.420 37.650 104.480 ;
        RECT 37.790 104.420 38.110 104.680 ;
        RECT 44.780 104.665 44.920 104.820 ;
        RECT 44.705 104.435 44.995 104.665 ;
        RECT 58.505 104.620 58.795 104.665 ;
        RECT 58.950 104.620 59.270 104.680 ;
        RECT 60.790 104.620 61.110 104.680 ;
        RECT 64.560 104.665 64.700 104.820 ;
        RECT 64.945 104.775 65.235 105.005 ;
        RECT 65.480 104.820 67.920 104.960 ;
        RECT 58.505 104.480 64.240 104.620 ;
        RECT 58.505 104.435 58.795 104.480 ;
        RECT 58.950 104.420 59.270 104.480 ;
        RECT 60.790 104.420 61.110 104.480 ;
        RECT 39.170 104.280 39.490 104.340 ;
        RECT 21.835 104.140 23.850 104.280 ;
        RECT 18.930 104.080 19.250 104.140 ;
        RECT 21.835 104.095 22.125 104.140 ;
        RECT 23.530 104.080 23.850 104.140 ;
        RECT 28.220 104.140 30.200 104.280 ;
        RECT 30.520 104.140 39.490 104.280 ;
        RECT 28.220 103.940 28.360 104.140 ;
        RECT 18.560 103.800 28.360 103.940 ;
        RECT 28.590 103.740 28.910 104.000 ;
        RECT 30.060 103.940 30.200 104.140 ;
        RECT 30.890 104.080 31.210 104.140 ;
        RECT 39.170 104.080 39.490 104.140 ;
        RECT 41.930 104.080 42.250 104.340 ;
        RECT 48.830 104.280 49.150 104.340 ;
        RECT 64.100 104.280 64.240 104.480 ;
        RECT 64.485 104.435 64.775 104.665 ;
        RECT 65.480 104.620 65.620 104.820 ;
        RECT 67.780 104.665 67.920 104.820 ;
        RECT 70.540 104.665 70.680 105.160 ;
        RECT 76.890 104.760 77.210 105.020 ;
        RECT 66.785 104.620 67.075 104.665 ;
        RECT 65.020 104.480 65.620 104.620 ;
        RECT 65.940 104.480 67.075 104.620 ;
        RECT 65.020 104.280 65.160 104.480 ;
        RECT 42.480 104.140 49.150 104.280 ;
        RECT 42.480 103.940 42.620 104.140 ;
        RECT 48.830 104.080 49.150 104.140 ;
        RECT 61.340 104.140 63.780 104.280 ;
        RECT 64.100 104.140 65.160 104.280 ;
        RECT 61.340 104.000 61.480 104.140 ;
        RECT 30.060 103.800 42.620 103.940 ;
        RECT 42.850 103.985 43.170 104.000 ;
        RECT 42.850 103.755 43.235 103.985 ;
        RECT 42.850 103.740 43.170 103.755 ;
        RECT 43.770 103.740 44.090 104.000 ;
        RECT 61.250 103.740 61.570 104.000 ;
        RECT 62.170 103.740 62.490 104.000 ;
        RECT 63.640 103.940 63.780 104.140 ;
        RECT 65.940 103.940 66.080 104.480 ;
        RECT 66.785 104.435 67.075 104.480 ;
        RECT 67.705 104.435 67.995 104.665 ;
        RECT 70.465 104.435 70.755 104.665 ;
        RECT 70.910 104.620 71.230 104.680 ;
        RECT 75.985 104.620 76.275 104.665 ;
        RECT 79.190 104.620 79.510 104.680 ;
        RECT 70.910 104.480 71.425 104.620 ;
        RECT 75.985 104.480 79.510 104.620 ;
        RECT 70.910 104.420 71.230 104.480 ;
        RECT 75.985 104.435 76.275 104.480 ;
        RECT 79.190 104.420 79.510 104.480 ;
        RECT 79.650 104.420 79.970 104.680 ;
        RECT 63.640 103.800 66.080 103.940 ;
        RECT 69.070 103.940 69.390 104.000 ;
        RECT 72.305 103.940 72.595 103.985 ;
        RECT 69.070 103.800 72.595 103.940 ;
        RECT 69.070 103.740 69.390 103.800 ;
        RECT 72.305 103.755 72.595 103.800 ;
        RECT 75.050 103.940 75.370 104.000 ;
        RECT 76.445 103.940 76.735 103.985 ;
        RECT 75.050 103.800 76.735 103.940 ;
        RECT 75.050 103.740 75.370 103.800 ;
        RECT 76.445 103.755 76.735 103.800 ;
        RECT 5.520 103.120 84.180 103.600 ;
        RECT 7.430 102.720 7.750 102.980 ;
        RECT 15.710 102.920 16.030 102.980 ;
        RECT 17.105 102.920 17.395 102.965 ;
        RECT 15.710 102.780 17.395 102.920 ;
        RECT 15.710 102.720 16.030 102.780 ;
        RECT 17.105 102.735 17.395 102.780 ;
        RECT 30.890 102.720 31.210 102.980 ;
        RECT 31.810 102.920 32.130 102.980 ;
        RECT 32.285 102.920 32.575 102.965 ;
        RECT 31.810 102.780 32.575 102.920 ;
        RECT 31.810 102.720 32.130 102.780 ;
        RECT 32.285 102.735 32.575 102.780 ;
        RECT 34.110 102.920 34.430 102.980 ;
        RECT 35.045 102.920 35.335 102.965 ;
        RECT 37.330 102.920 37.650 102.980 ;
        RECT 49.290 102.965 49.610 102.980 ;
        RECT 42.865 102.920 43.155 102.965 ;
        RECT 34.110 102.780 35.335 102.920 ;
        RECT 34.110 102.720 34.430 102.780 ;
        RECT 35.045 102.735 35.335 102.780 ;
        RECT 35.580 102.780 43.155 102.920 ;
        RECT 8.810 102.380 9.130 102.640 ;
        RECT 9.270 102.380 9.590 102.640 ;
        RECT 9.975 102.580 10.265 102.625 ;
        RECT 11.570 102.580 11.890 102.640 ;
        RECT 14.330 102.580 14.650 102.640 ;
        RECT 17.550 102.580 17.870 102.640 ;
        RECT 28.590 102.580 28.910 102.640 ;
        RECT 9.975 102.440 11.890 102.580 ;
        RECT 9.975 102.395 10.265 102.440 ;
        RECT 11.570 102.380 11.890 102.440 ;
        RECT 13.960 102.440 14.650 102.580 ;
        RECT 8.365 102.055 8.655 102.285 ;
        RECT 8.440 101.900 8.580 102.055 ;
        RECT 10.650 102.040 10.970 102.300 ;
        RECT 12.505 102.240 12.795 102.285 ;
        RECT 13.410 102.240 13.730 102.300 ;
        RECT 13.960 102.285 14.100 102.440 ;
        RECT 14.330 102.380 14.650 102.440 ;
        RECT 14.880 102.440 18.700 102.580 ;
        RECT 14.880 102.285 15.020 102.440 ;
        RECT 17.550 102.380 17.870 102.440 ;
        RECT 18.560 102.300 18.700 102.440 ;
        RECT 28.590 102.440 33.420 102.580 ;
        RECT 28.590 102.380 28.910 102.440 ;
        RECT 12.505 102.100 13.730 102.240 ;
        RECT 12.505 102.055 12.795 102.100 ;
        RECT 13.410 102.040 13.730 102.100 ;
        RECT 13.885 102.055 14.175 102.285 ;
        RECT 14.805 102.055 15.095 102.285 ;
        RECT 15.250 102.040 15.570 102.300 ;
        RECT 18.470 102.040 18.790 102.300 ;
        RECT 18.930 102.240 19.250 102.300 ;
        RECT 24.005 102.240 24.295 102.285 ;
        RECT 18.930 102.100 24.295 102.240 ;
        RECT 18.930 102.040 19.250 102.100 ;
        RECT 24.005 102.055 24.295 102.100 ;
        RECT 25.340 102.240 25.630 102.285 ;
        RECT 25.340 102.100 29.740 102.240 ;
        RECT 25.340 102.055 25.630 102.100 ;
        RECT 9.730 101.900 10.050 101.960 ;
        RECT 14.345 101.900 14.635 101.945 ;
        RECT 15.710 101.900 16.030 101.960 ;
        RECT 17.105 101.900 17.395 101.945 ;
        RECT 8.440 101.760 12.260 101.900 ;
        RECT 9.730 101.700 10.050 101.760 ;
        RECT 6.510 101.560 6.830 101.620 ;
        RECT 11.585 101.560 11.875 101.605 ;
        RECT 6.510 101.420 11.875 101.560 ;
        RECT 12.120 101.560 12.260 101.760 ;
        RECT 14.345 101.760 17.395 101.900 ;
        RECT 14.345 101.715 14.635 101.760 ;
        RECT 15.710 101.700 16.030 101.760 ;
        RECT 17.105 101.715 17.395 101.760 ;
        RECT 18.010 101.900 18.330 101.960 ;
        RECT 23.085 101.900 23.375 101.945 ;
        RECT 18.010 101.760 23.375 101.900 ;
        RECT 18.010 101.700 18.330 101.760 ;
        RECT 23.085 101.715 23.375 101.760 ;
        RECT 24.885 101.900 25.175 101.945 ;
        RECT 26.075 101.900 26.365 101.945 ;
        RECT 28.595 101.900 28.885 101.945 ;
        RECT 24.885 101.760 28.885 101.900 ;
        RECT 29.600 101.900 29.740 102.100 ;
        RECT 31.810 102.040 32.130 102.300 ;
        RECT 33.280 102.285 33.420 102.440 ;
        RECT 33.205 102.055 33.495 102.285 ;
        RECT 34.585 102.240 34.875 102.285 ;
        RECT 35.030 102.240 35.350 102.300 ;
        RECT 35.580 102.285 35.720 102.780 ;
        RECT 37.330 102.720 37.650 102.780 ;
        RECT 42.865 102.735 43.155 102.780 ;
        RECT 49.290 102.735 49.675 102.965 ;
        RECT 56.190 102.920 56.510 102.980 ;
        RECT 59.410 102.920 59.730 102.980 ;
        RECT 68.150 102.920 68.470 102.980 ;
        RECT 70.925 102.920 71.215 102.965 ;
        RECT 76.890 102.920 77.210 102.980 ;
        RECT 56.190 102.780 69.760 102.920 ;
        RECT 49.290 102.720 49.610 102.735 ;
        RECT 56.190 102.720 56.510 102.780 ;
        RECT 59.410 102.720 59.730 102.780 ;
        RECT 68.150 102.720 68.470 102.780 ;
        RECT 48.370 102.380 48.690 102.640 ;
        RECT 58.950 102.580 59.270 102.640 ;
        RECT 59.870 102.580 60.190 102.640 ;
        RECT 58.950 102.440 69.300 102.580 ;
        RECT 58.950 102.380 59.270 102.440 ;
        RECT 59.870 102.380 60.190 102.440 ;
        RECT 69.160 102.300 69.300 102.440 ;
        RECT 34.585 102.100 35.350 102.240 ;
        RECT 34.585 102.055 34.875 102.100 ;
        RECT 35.030 102.040 35.350 102.100 ;
        RECT 35.505 102.055 35.795 102.285 ;
        RECT 37.300 102.240 37.590 102.285 ;
        RECT 38.710 102.240 39.030 102.300 ;
        RECT 37.300 102.100 39.030 102.240 ;
        RECT 37.300 102.055 37.590 102.100 ;
        RECT 38.710 102.040 39.030 102.100 ;
        RECT 57.570 102.040 57.890 102.300 ;
        RECT 61.250 102.240 61.570 102.300 ;
        RECT 65.405 102.240 65.695 102.285 ;
        RECT 61.250 102.100 65.695 102.240 ;
        RECT 61.250 102.040 61.570 102.100 ;
        RECT 65.405 102.055 65.695 102.100 ;
        RECT 66.325 102.240 66.615 102.285 ;
        RECT 67.230 102.240 67.550 102.300 ;
        RECT 66.325 102.100 67.550 102.240 ;
        RECT 66.325 102.055 66.615 102.100 ;
        RECT 67.230 102.040 67.550 102.100 ;
        RECT 67.705 102.055 67.995 102.285 ;
        RECT 34.125 101.900 34.415 101.945 ;
        RECT 29.600 101.760 34.415 101.900 ;
        RECT 24.885 101.715 25.175 101.760 ;
        RECT 26.075 101.715 26.365 101.760 ;
        RECT 28.595 101.715 28.885 101.760 ;
        RECT 34.125 101.715 34.415 101.760 ;
        RECT 35.950 101.700 36.270 101.960 ;
        RECT 36.845 101.900 37.135 101.945 ;
        RECT 38.035 101.900 38.325 101.945 ;
        RECT 40.555 101.900 40.845 101.945 ;
        RECT 36.845 101.760 40.845 101.900 ;
        RECT 36.845 101.715 37.135 101.760 ;
        RECT 38.035 101.715 38.325 101.760 ;
        RECT 40.555 101.715 40.845 101.760 ;
        RECT 46.070 101.900 46.390 101.960 ;
        RECT 47.005 101.900 47.295 101.945 ;
        RECT 46.070 101.760 47.295 101.900 ;
        RECT 46.070 101.700 46.390 101.760 ;
        RECT 47.005 101.715 47.295 101.760 ;
        RECT 47.450 101.900 47.770 101.960 ;
        RECT 50.685 101.900 50.975 101.945 ;
        RECT 47.450 101.760 50.975 101.900 ;
        RECT 47.450 101.700 47.770 101.760 ;
        RECT 50.685 101.715 50.975 101.760 ;
        RECT 58.965 101.900 59.255 101.945 ;
        RECT 61.340 101.900 61.480 102.040 ;
        RECT 58.965 101.760 61.480 101.900 ;
        RECT 65.850 101.900 66.170 101.960 ;
        RECT 67.780 101.900 67.920 102.055 ;
        RECT 68.610 102.040 68.930 102.300 ;
        RECT 69.070 102.040 69.390 102.300 ;
        RECT 69.620 102.285 69.760 102.780 ;
        RECT 70.925 102.780 77.210 102.920 ;
        RECT 70.925 102.735 71.215 102.780 ;
        RECT 76.890 102.720 77.210 102.780 ;
        RECT 69.545 102.055 69.835 102.285 ;
        RECT 72.765 102.055 73.055 102.285 ;
        RECT 65.850 101.760 67.920 101.900 ;
        RECT 58.965 101.715 59.255 101.760 ;
        RECT 65.850 101.700 66.170 101.760 ;
        RECT 16.185 101.560 16.475 101.605 ;
        RECT 16.630 101.560 16.950 101.620 ;
        RECT 24.490 101.560 24.780 101.605 ;
        RECT 26.590 101.560 26.880 101.605 ;
        RECT 28.160 101.560 28.450 101.605 ;
        RECT 12.120 101.420 21.000 101.560 ;
        RECT 6.510 101.360 6.830 101.420 ;
        RECT 11.585 101.375 11.875 101.420 ;
        RECT 16.185 101.375 16.475 101.420 ;
        RECT 16.630 101.360 16.950 101.420 ;
        RECT 18.010 101.020 18.330 101.280 ;
        RECT 18.470 101.220 18.790 101.280 ;
        RECT 20.325 101.220 20.615 101.265 ;
        RECT 18.470 101.080 20.615 101.220 ;
        RECT 20.860 101.220 21.000 101.420 ;
        RECT 24.490 101.420 28.450 101.560 ;
        RECT 24.490 101.375 24.780 101.420 ;
        RECT 26.590 101.375 26.880 101.420 ;
        RECT 28.160 101.375 28.450 101.420 ;
        RECT 36.450 101.560 36.740 101.605 ;
        RECT 38.550 101.560 38.840 101.605 ;
        RECT 40.120 101.560 40.410 101.605 ;
        RECT 36.450 101.420 40.410 101.560 ;
        RECT 36.450 101.375 36.740 101.420 ;
        RECT 38.550 101.375 38.840 101.420 ;
        RECT 40.120 101.375 40.410 101.420 ;
        RECT 50.225 101.560 50.515 101.605 ;
        RECT 72.290 101.560 72.610 101.620 ;
        RECT 72.840 101.560 72.980 102.055 ;
        RECT 79.650 101.900 79.970 101.960 ;
        RECT 81.045 101.900 81.335 101.945 ;
        RECT 79.650 101.760 81.335 101.900 ;
        RECT 79.650 101.700 79.970 101.760 ;
        RECT 81.045 101.715 81.335 101.760 ;
        RECT 50.225 101.420 72.980 101.560 ;
        RECT 50.225 101.375 50.515 101.420 ;
        RECT 72.290 101.360 72.610 101.420 ;
        RECT 41.930 101.220 42.250 101.280 ;
        RECT 20.860 101.080 42.250 101.220 ;
        RECT 18.470 101.020 18.790 101.080 ;
        RECT 20.325 101.035 20.615 101.080 ;
        RECT 41.930 101.020 42.250 101.080 ;
        RECT 44.230 101.020 44.550 101.280 ;
        RECT 48.830 101.220 49.150 101.280 ;
        RECT 49.305 101.220 49.595 101.265 ;
        RECT 48.830 101.080 49.595 101.220 ;
        RECT 48.830 101.020 49.150 101.080 ;
        RECT 49.305 101.035 49.595 101.080 ;
        RECT 53.890 101.020 54.210 101.280 ;
        RECT 57.570 101.220 57.890 101.280 ;
        RECT 58.045 101.220 58.335 101.265 ;
        RECT 57.570 101.080 58.335 101.220 ;
        RECT 57.570 101.020 57.890 101.080 ;
        RECT 58.045 101.035 58.335 101.080 ;
        RECT 58.505 101.220 58.795 101.265 ;
        RECT 59.870 101.220 60.190 101.280 ;
        RECT 58.505 101.080 60.190 101.220 ;
        RECT 58.505 101.035 58.795 101.080 ;
        RECT 59.870 101.020 60.190 101.080 ;
        RECT 65.850 101.220 66.170 101.280 ;
        RECT 66.785 101.220 67.075 101.265 ;
        RECT 65.850 101.080 67.075 101.220 ;
        RECT 65.850 101.020 66.170 101.080 ;
        RECT 66.785 101.035 67.075 101.080 ;
        RECT 67.230 101.220 67.550 101.280 ;
        RECT 69.070 101.220 69.390 101.280 ;
        RECT 71.845 101.220 72.135 101.265 ;
        RECT 67.230 101.080 72.135 101.220 ;
        RECT 67.230 101.020 67.550 101.080 ;
        RECT 69.070 101.020 69.390 101.080 ;
        RECT 71.845 101.035 72.135 101.080 ;
        RECT 76.430 101.220 76.750 101.280 ;
        RECT 78.285 101.220 78.575 101.265 ;
        RECT 76.430 101.080 78.575 101.220 ;
        RECT 76.430 101.020 76.750 101.080 ;
        RECT 78.285 101.035 78.575 101.080 ;
        RECT 5.520 100.400 84.180 100.880 ;
        RECT 7.905 100.200 8.195 100.245 ;
        RECT 13.870 100.200 14.190 100.260 ;
        RECT 14.790 100.200 15.110 100.260 ;
        RECT 25.845 100.200 26.135 100.245 ;
        RECT 7.905 100.060 15.110 100.200 ;
        RECT 7.905 100.015 8.195 100.060 ;
        RECT 13.870 100.000 14.190 100.060 ;
        RECT 14.790 100.000 15.110 100.060 ;
        RECT 16.260 100.060 26.135 100.200 ;
        RECT 16.260 99.920 16.400 100.060 ;
        RECT 25.845 100.015 26.135 100.060 ;
        RECT 30.905 100.200 31.195 100.245 ;
        RECT 31.810 100.200 32.130 100.260 ;
        RECT 30.905 100.060 32.130 100.200 ;
        RECT 30.905 100.015 31.195 100.060 ;
        RECT 31.810 100.000 32.130 100.060 ;
        RECT 32.285 100.200 32.575 100.245 ;
        RECT 35.490 100.200 35.810 100.260 ;
        RECT 32.285 100.060 35.810 100.200 ;
        RECT 32.285 100.015 32.575 100.060 ;
        RECT 35.490 100.000 35.810 100.060 ;
        RECT 38.710 100.000 39.030 100.260 ;
        RECT 42.850 100.200 43.170 100.260 ;
        RECT 43.325 100.200 43.615 100.245 ;
        RECT 42.850 100.060 43.615 100.200 ;
        RECT 42.850 100.000 43.170 100.060 ;
        RECT 43.325 100.015 43.615 100.060 ;
        RECT 45.625 100.200 45.915 100.245 ;
        RECT 47.450 100.200 47.770 100.260 ;
        RECT 45.625 100.060 47.770 100.200 ;
        RECT 45.625 100.015 45.915 100.060 ;
        RECT 47.450 100.000 47.770 100.060 ;
        RECT 79.650 100.000 79.970 100.260 ;
        RECT 16.170 99.860 16.490 99.920 ;
        RECT 10.740 99.720 16.490 99.860 ;
        RECT 4.210 99.180 4.530 99.240 ;
        RECT 7.445 99.180 7.735 99.225 ;
        RECT 4.210 99.040 7.735 99.180 ;
        RECT 4.210 98.980 4.530 99.040 ;
        RECT 7.445 98.995 7.735 99.040 ;
        RECT 9.745 99.180 10.035 99.225 ;
        RECT 10.190 99.180 10.510 99.240 ;
        RECT 10.740 99.225 10.880 99.720 ;
        RECT 16.170 99.660 16.490 99.720 ;
        RECT 19.430 99.860 19.720 99.905 ;
        RECT 21.530 99.860 21.820 99.905 ;
        RECT 23.100 99.860 23.390 99.905 ;
        RECT 37.345 99.860 37.635 99.905 ;
        RECT 19.430 99.720 23.390 99.860 ;
        RECT 19.430 99.675 19.720 99.720 ;
        RECT 21.530 99.675 21.820 99.720 ;
        RECT 23.100 99.675 23.390 99.720 ;
        RECT 33.740 99.720 37.635 99.860 ;
        RECT 15.710 99.320 16.030 99.580 ;
        RECT 18.930 99.320 19.250 99.580 ;
        RECT 19.825 99.520 20.115 99.565 ;
        RECT 21.015 99.520 21.305 99.565 ;
        RECT 23.535 99.520 23.825 99.565 ;
        RECT 33.740 99.520 33.880 99.720 ;
        RECT 37.345 99.675 37.635 99.720 ;
        RECT 48.370 99.860 48.660 99.905 ;
        RECT 49.940 99.860 50.230 99.905 ;
        RECT 52.040 99.860 52.330 99.905 ;
        RECT 48.370 99.720 52.330 99.860 ;
        RECT 48.370 99.675 48.660 99.720 ;
        RECT 49.940 99.675 50.230 99.720 ;
        RECT 52.040 99.675 52.330 99.720 ;
        RECT 58.045 99.860 58.335 99.905 ;
        RECT 60.330 99.860 60.650 99.920 ;
        RECT 69.530 99.860 69.850 99.920 ;
        RECT 58.045 99.720 60.650 99.860 ;
        RECT 58.045 99.675 58.335 99.720 ;
        RECT 60.330 99.660 60.650 99.720 ;
        RECT 66.400 99.720 69.850 99.860 ;
        RECT 36.870 99.520 37.190 99.580 ;
        RECT 19.825 99.380 23.825 99.520 ;
        RECT 19.825 99.335 20.115 99.380 ;
        RECT 21.015 99.335 21.305 99.380 ;
        RECT 23.535 99.335 23.825 99.380 ;
        RECT 31.440 99.380 33.880 99.520 ;
        RECT 9.745 99.040 10.510 99.180 ;
        RECT 9.745 98.995 10.035 99.040 ;
        RECT 10.190 98.980 10.510 99.040 ;
        RECT 10.665 98.995 10.955 99.225 ;
        RECT 11.570 98.980 11.890 99.240 ;
        RECT 16.185 99.180 16.475 99.225 ;
        RECT 18.470 99.180 18.790 99.240 ;
        RECT 31.440 99.225 31.580 99.380 ;
        RECT 16.185 99.040 18.790 99.180 ;
        RECT 16.185 98.995 16.475 99.040 ;
        RECT 18.470 98.980 18.790 99.040 ;
        RECT 30.445 98.995 30.735 99.225 ;
        RECT 31.365 98.995 31.655 99.225 ;
        RECT 10.280 98.840 10.420 98.980 ;
        RECT 15.710 98.840 16.030 98.900 ;
        RECT 20.170 98.840 20.460 98.885 ;
        RECT 10.280 98.700 16.030 98.840 ;
        RECT 15.710 98.640 16.030 98.700 ;
        RECT 18.100 98.700 20.460 98.840 ;
        RECT 30.520 98.840 30.660 98.995 ;
        RECT 33.190 98.980 33.510 99.240 ;
        RECT 33.740 99.225 33.880 99.380 ;
        RECT 34.660 99.380 37.190 99.520 ;
        RECT 33.665 99.180 33.955 99.225 ;
        RECT 34.110 99.180 34.430 99.240 ;
        RECT 34.660 99.225 34.800 99.380 ;
        RECT 36.870 99.320 37.190 99.380 ;
        RECT 47.935 99.520 48.225 99.565 ;
        RECT 50.455 99.520 50.745 99.565 ;
        RECT 51.645 99.520 51.935 99.565 ;
        RECT 47.935 99.380 51.935 99.520 ;
        RECT 47.935 99.335 48.225 99.380 ;
        RECT 50.455 99.335 50.745 99.380 ;
        RECT 51.645 99.335 51.935 99.380 ;
        RECT 53.890 99.520 54.210 99.580 ;
        RECT 55.285 99.520 55.575 99.565 ;
        RECT 53.890 99.380 55.575 99.520 ;
        RECT 53.890 99.320 54.210 99.380 ;
        RECT 55.285 99.335 55.575 99.380 ;
        RECT 56.205 99.520 56.495 99.565 ;
        RECT 65.405 99.520 65.695 99.565 ;
        RECT 56.205 99.380 65.695 99.520 ;
        RECT 56.205 99.335 56.495 99.380 ;
        RECT 65.405 99.335 65.695 99.380 ;
        RECT 33.665 99.040 34.430 99.180 ;
        RECT 33.665 98.995 33.955 99.040 ;
        RECT 34.110 98.980 34.430 99.040 ;
        RECT 34.585 98.995 34.875 99.225 ;
        RECT 35.030 98.980 35.350 99.240 ;
        RECT 35.505 98.995 35.795 99.225 ;
        RECT 36.425 99.180 36.715 99.225 ;
        RECT 37.330 99.180 37.650 99.240 ;
        RECT 36.425 99.040 37.650 99.180 ;
        RECT 36.425 98.995 36.715 99.040 ;
        RECT 35.580 98.840 35.720 98.995 ;
        RECT 37.330 98.980 37.650 99.040 ;
        RECT 37.790 98.980 38.110 99.240 ;
        RECT 43.785 99.180 44.075 99.225 ;
        RECT 49.290 99.180 49.610 99.240 ;
        RECT 52.525 99.180 52.815 99.225 ;
        RECT 43.785 99.040 48.140 99.180 ;
        RECT 43.785 98.995 44.075 99.040 ;
        RECT 48.000 98.900 48.140 99.040 ;
        RECT 49.290 99.040 52.815 99.180 ;
        RECT 49.290 98.980 49.610 99.040 ;
        RECT 52.525 98.995 52.815 99.040 ;
        RECT 57.110 98.980 57.430 99.240 ;
        RECT 58.950 98.980 59.270 99.240 ;
        RECT 59.410 99.180 59.730 99.240 ;
        RECT 66.400 99.225 66.540 99.720 ;
        RECT 69.530 99.660 69.850 99.720 ;
        RECT 73.250 99.860 73.540 99.905 ;
        RECT 75.350 99.860 75.640 99.905 ;
        RECT 76.920 99.860 77.210 99.905 ;
        RECT 73.250 99.720 77.210 99.860 ;
        RECT 73.250 99.675 73.540 99.720 ;
        RECT 75.350 99.675 75.640 99.720 ;
        RECT 76.920 99.675 77.210 99.720 ;
        RECT 66.785 99.520 67.075 99.565 ;
        RECT 67.230 99.520 67.550 99.580 ;
        RECT 69.070 99.520 69.390 99.580 ;
        RECT 66.785 99.380 67.550 99.520 ;
        RECT 66.785 99.335 67.075 99.380 ;
        RECT 67.230 99.320 67.550 99.380 ;
        RECT 67.780 99.380 69.390 99.520 ;
        RECT 67.780 99.225 67.920 99.380 ;
        RECT 69.070 99.320 69.390 99.380 ;
        RECT 73.645 99.520 73.935 99.565 ;
        RECT 74.835 99.520 75.125 99.565 ;
        RECT 77.355 99.520 77.645 99.565 ;
        RECT 73.645 99.380 77.645 99.520 ;
        RECT 73.645 99.335 73.935 99.380 ;
        RECT 74.835 99.335 75.125 99.380 ;
        RECT 77.355 99.335 77.645 99.380 ;
        RECT 59.885 99.180 60.175 99.225 ;
        RECT 59.410 99.040 60.175 99.180 ;
        RECT 59.410 98.980 59.730 99.040 ;
        RECT 59.885 98.995 60.175 99.040 ;
        RECT 64.945 98.995 65.235 99.225 ;
        RECT 65.865 98.995 66.155 99.225 ;
        RECT 66.325 98.995 66.615 99.225 ;
        RECT 67.705 98.995 67.995 99.225 ;
        RECT 68.165 98.995 68.455 99.225 ;
        RECT 30.520 98.700 35.720 98.840 ;
        RECT 10.650 98.300 10.970 98.560 ;
        RECT 14.330 98.300 14.650 98.560 ;
        RECT 18.100 98.545 18.240 98.700 ;
        RECT 20.170 98.655 20.460 98.700 ;
        RECT 33.740 98.560 33.880 98.700 ;
        RECT 47.910 98.640 48.230 98.900 ;
        RECT 51.300 98.840 51.590 98.885 ;
        RECT 54.825 98.840 55.115 98.885 ;
        RECT 59.040 98.840 59.180 98.980 ;
        RECT 51.300 98.700 53.200 98.840 ;
        RECT 51.300 98.655 51.590 98.700 ;
        RECT 18.025 98.315 18.315 98.545 ;
        RECT 33.650 98.300 33.970 98.560 ;
        RECT 53.060 98.545 53.200 98.700 ;
        RECT 54.825 98.700 59.180 98.840 ;
        RECT 54.825 98.655 55.115 98.700 ;
        RECT 52.985 98.315 53.275 98.545 ;
        RECT 58.490 98.500 58.810 98.560 ;
        RECT 59.425 98.500 59.715 98.545 ;
        RECT 58.490 98.360 59.715 98.500 ;
        RECT 65.020 98.500 65.160 98.995 ;
        RECT 65.940 98.840 66.080 98.995 ;
        RECT 66.770 98.840 67.090 98.900 ;
        RECT 68.240 98.840 68.380 98.995 ;
        RECT 72.750 98.980 73.070 99.240 ;
        RECT 65.940 98.700 68.380 98.840 ;
        RECT 74.100 98.840 74.390 98.885 ;
        RECT 74.590 98.840 74.910 98.900 ;
        RECT 74.100 98.700 74.910 98.840 ;
        RECT 66.770 98.640 67.090 98.700 ;
        RECT 74.100 98.655 74.390 98.700 ;
        RECT 74.590 98.640 74.910 98.700 ;
        RECT 67.230 98.500 67.550 98.560 ;
        RECT 65.020 98.360 67.550 98.500 ;
        RECT 58.490 98.300 58.810 98.360 ;
        RECT 59.425 98.315 59.715 98.360 ;
        RECT 67.230 98.300 67.550 98.360 ;
        RECT 69.085 98.500 69.375 98.545 ;
        RECT 77.350 98.500 77.670 98.560 ;
        RECT 69.085 98.360 77.670 98.500 ;
        RECT 69.085 98.315 69.375 98.360 ;
        RECT 77.350 98.300 77.670 98.360 ;
        RECT 5.520 97.680 84.180 98.160 ;
        RECT 15.710 97.280 16.030 97.540 ;
        RECT 16.170 97.280 16.490 97.540 ;
        RECT 33.190 97.480 33.510 97.540 ;
        RECT 35.045 97.480 35.335 97.525 ;
        RECT 33.190 97.340 35.335 97.480 ;
        RECT 33.190 97.280 33.510 97.340 ;
        RECT 35.045 97.295 35.335 97.340 ;
        RECT 36.885 97.480 37.175 97.525 ;
        RECT 46.070 97.480 46.390 97.540 ;
        RECT 36.885 97.340 46.390 97.480 ;
        RECT 36.885 97.295 37.175 97.340 ;
        RECT 46.070 97.280 46.390 97.340 ;
        RECT 56.665 97.480 56.955 97.525 ;
        RECT 57.110 97.480 57.430 97.540 ;
        RECT 56.665 97.340 57.430 97.480 ;
        RECT 56.665 97.295 56.955 97.340 ;
        RECT 57.110 97.280 57.430 97.340 ;
        RECT 57.585 97.295 57.875 97.525 ;
        RECT 58.030 97.480 58.350 97.540 ;
        RECT 59.870 97.480 60.190 97.540 ;
        RECT 58.030 97.340 60.190 97.480 ;
        RECT 8.320 97.140 8.610 97.185 ;
        RECT 18.485 97.140 18.775 97.185 ;
        RECT 8.320 97.000 18.775 97.140 ;
        RECT 8.320 96.955 8.610 97.000 ;
        RECT 18.485 96.955 18.775 97.000 ;
        RECT 35.950 97.140 36.270 97.200 ;
        RECT 41.010 97.140 41.330 97.200 ;
        RECT 35.950 97.000 41.330 97.140 ;
        RECT 35.950 96.940 36.270 97.000 ;
        RECT 6.970 96.600 7.290 96.860 ;
        RECT 14.330 96.800 14.650 96.860 ;
        RECT 18.025 96.800 18.315 96.845 ;
        RECT 14.330 96.660 18.315 96.800 ;
        RECT 14.330 96.600 14.650 96.660 ;
        RECT 18.025 96.615 18.315 96.660 ;
        RECT 18.945 96.615 19.235 96.845 ;
        RECT 37.345 96.800 37.635 96.845 ;
        RECT 38.250 96.800 38.570 96.860 ;
        RECT 39.260 96.845 39.400 97.000 ;
        RECT 41.010 96.940 41.330 97.000 ;
        RECT 48.830 97.140 49.150 97.200 ;
        RECT 49.305 97.140 49.595 97.185 ;
        RECT 48.830 97.000 49.595 97.140 ;
        RECT 48.830 96.940 49.150 97.000 ;
        RECT 49.305 96.955 49.595 97.000 ;
        RECT 51.100 97.140 51.390 97.185 ;
        RECT 57.660 97.140 57.800 97.295 ;
        RECT 58.030 97.280 58.350 97.340 ;
        RECT 59.870 97.280 60.190 97.340 ;
        RECT 66.770 97.280 67.090 97.540 ;
        RECT 68.610 97.480 68.930 97.540 ;
        RECT 69.545 97.480 69.835 97.525 ;
        RECT 68.610 97.340 69.835 97.480 ;
        RECT 68.610 97.280 68.930 97.340 ;
        RECT 69.545 97.295 69.835 97.340 ;
        RECT 74.590 97.280 74.910 97.540 ;
        RECT 76.430 97.280 76.750 97.540 ;
        RECT 72.765 97.140 73.055 97.185 ;
        RECT 51.100 97.000 57.800 97.140 ;
        RECT 68.700 97.000 73.055 97.140 ;
        RECT 51.100 96.955 51.390 97.000 ;
        RECT 40.550 96.845 40.870 96.860 ;
        RECT 37.345 96.660 38.570 96.800 ;
        RECT 37.345 96.615 37.635 96.660 ;
        RECT 7.865 96.460 8.155 96.505 ;
        RECT 9.055 96.460 9.345 96.505 ;
        RECT 11.575 96.460 11.865 96.505 ;
        RECT 15.140 96.460 15.430 96.505 ;
        RECT 7.865 96.320 11.865 96.460 ;
        RECT 7.865 96.275 8.155 96.320 ;
        RECT 9.055 96.275 9.345 96.320 ;
        RECT 11.575 96.275 11.865 96.320 ;
        RECT 13.960 96.320 15.430 96.460 ;
        RECT 7.470 96.120 7.760 96.165 ;
        RECT 9.570 96.120 9.860 96.165 ;
        RECT 11.140 96.120 11.430 96.165 ;
        RECT 7.470 95.980 11.430 96.120 ;
        RECT 7.470 95.935 7.760 95.980 ;
        RECT 9.570 95.935 9.860 95.980 ;
        RECT 11.140 95.935 11.430 95.980 ;
        RECT 13.960 95.840 14.100 96.320 ;
        RECT 15.140 96.275 15.430 96.320 ;
        RECT 17.550 96.260 17.870 96.520 ;
        RECT 18.470 96.460 18.790 96.520 ;
        RECT 19.020 96.460 19.160 96.615 ;
        RECT 38.250 96.600 38.570 96.660 ;
        RECT 39.185 96.615 39.475 96.845 ;
        RECT 40.520 96.615 40.870 96.845 ;
        RECT 40.550 96.600 40.870 96.615 ;
        RECT 48.370 96.600 48.690 96.860 ;
        RECT 58.490 96.800 58.810 96.860 ;
        RECT 59.425 96.800 59.715 96.845 ;
        RECT 58.490 96.660 59.715 96.800 ;
        RECT 58.490 96.600 58.810 96.660 ;
        RECT 59.425 96.615 59.715 96.660 ;
        RECT 61.250 96.800 61.570 96.860 ;
        RECT 64.485 96.800 64.775 96.845 ;
        RECT 61.250 96.660 64.775 96.800 ;
        RECT 61.250 96.600 61.570 96.660 ;
        RECT 64.485 96.615 64.775 96.660 ;
        RECT 65.865 96.800 66.155 96.845 ;
        RECT 66.310 96.800 66.630 96.860 ;
        RECT 65.865 96.660 66.630 96.800 ;
        RECT 65.865 96.615 66.155 96.660 ;
        RECT 66.310 96.600 66.630 96.660 ;
        RECT 67.690 96.600 68.010 96.860 ;
        RECT 68.150 96.800 68.470 96.860 ;
        RECT 68.700 96.845 68.840 97.000 ;
        RECT 72.765 96.955 73.055 97.000 ;
        RECT 68.625 96.800 68.915 96.845 ;
        RECT 71.385 96.800 71.675 96.845 ;
        RECT 68.150 96.660 68.915 96.800 ;
        RECT 68.150 96.600 68.470 96.660 ;
        RECT 68.625 96.615 68.915 96.660 ;
        RECT 69.160 96.660 71.675 96.800 ;
        RECT 18.470 96.320 19.160 96.460 ;
        RECT 18.470 96.260 18.790 96.320 ;
        RECT 37.805 96.275 38.095 96.505 ;
        RECT 40.065 96.460 40.355 96.505 ;
        RECT 41.255 96.460 41.545 96.505 ;
        RECT 43.775 96.460 44.065 96.505 ;
        RECT 49.765 96.460 50.055 96.505 ;
        RECT 40.065 96.320 44.065 96.460 ;
        RECT 40.065 96.275 40.355 96.320 ;
        RECT 41.255 96.275 41.545 96.320 ;
        RECT 43.775 96.275 44.065 96.320 ;
        RECT 49.380 96.320 50.055 96.460 ;
        RECT 37.880 96.120 38.020 96.275 ;
        RECT 49.380 96.180 49.520 96.320 ;
        RECT 49.765 96.275 50.055 96.320 ;
        RECT 50.645 96.460 50.935 96.505 ;
        RECT 51.835 96.460 52.125 96.505 ;
        RECT 54.355 96.460 54.645 96.505 ;
        RECT 50.645 96.320 54.645 96.460 ;
        RECT 50.645 96.275 50.935 96.320 ;
        RECT 51.835 96.275 52.125 96.320 ;
        RECT 54.355 96.275 54.645 96.320 ;
        RECT 60.330 96.460 60.650 96.520 ;
        RECT 62.630 96.460 62.950 96.520 ;
        RECT 60.330 96.320 62.950 96.460 ;
        RECT 60.330 96.260 60.650 96.320 ;
        RECT 62.630 96.260 62.950 96.320 ;
        RECT 65.405 96.460 65.695 96.505 ;
        RECT 66.770 96.460 67.090 96.520 ;
        RECT 67.780 96.460 67.920 96.600 ;
        RECT 65.405 96.320 67.920 96.460 ;
        RECT 65.405 96.275 65.695 96.320 ;
        RECT 66.770 96.260 67.090 96.320 ;
        RECT 39.170 96.120 39.490 96.180 ;
        RECT 37.880 95.980 39.490 96.120 ;
        RECT 39.170 95.920 39.490 95.980 ;
        RECT 39.670 96.120 39.960 96.165 ;
        RECT 41.770 96.120 42.060 96.165 ;
        RECT 43.340 96.120 43.630 96.165 ;
        RECT 39.670 95.980 43.630 96.120 ;
        RECT 39.670 95.935 39.960 95.980 ;
        RECT 41.770 95.935 42.060 95.980 ;
        RECT 43.340 95.935 43.630 95.980 ;
        RECT 43.860 95.980 48.600 96.120 ;
        RECT 13.870 95.580 14.190 95.840 ;
        RECT 14.330 95.580 14.650 95.840 ;
        RECT 26.290 95.780 26.610 95.840 ;
        RECT 43.860 95.780 44.000 95.980 ;
        RECT 26.290 95.640 44.000 95.780 ;
        RECT 26.290 95.580 26.610 95.640 ;
        RECT 47.910 95.580 48.230 95.840 ;
        RECT 48.460 95.780 48.600 95.980 ;
        RECT 49.290 95.920 49.610 96.180 ;
        RECT 50.250 96.120 50.540 96.165 ;
        RECT 52.350 96.120 52.640 96.165 ;
        RECT 53.920 96.120 54.210 96.165 ;
        RECT 50.250 95.980 54.210 96.120 ;
        RECT 50.250 95.935 50.540 95.980 ;
        RECT 52.350 95.935 52.640 95.980 ;
        RECT 53.920 95.935 54.210 95.980 ;
        RECT 64.930 95.920 65.250 96.180 ;
        RECT 67.690 95.920 68.010 96.180 ;
        RECT 68.610 96.120 68.930 96.180 ;
        RECT 69.160 96.120 69.300 96.660 ;
        RECT 71.385 96.615 71.675 96.660 ;
        RECT 71.830 96.600 72.150 96.860 ;
        RECT 70.450 96.460 70.770 96.520 ;
        RECT 70.925 96.460 71.215 96.505 ;
        RECT 70.450 96.320 71.215 96.460 ;
        RECT 70.450 96.260 70.770 96.320 ;
        RECT 70.925 96.275 71.215 96.320 ;
        RECT 76.890 96.260 77.210 96.520 ;
        RECT 77.350 96.260 77.670 96.520 ;
        RECT 68.610 95.980 69.300 96.120 ;
        RECT 69.530 96.120 69.850 96.180 ;
        RECT 73.670 96.120 73.990 96.180 ;
        RECT 69.530 95.980 73.990 96.120 ;
        RECT 68.610 95.920 68.930 95.980 ;
        RECT 69.530 95.920 69.850 95.980 ;
        RECT 73.670 95.920 73.990 95.980 ;
        RECT 69.990 95.780 70.310 95.840 ;
        RECT 48.460 95.640 70.310 95.780 ;
        RECT 69.990 95.580 70.310 95.640 ;
        RECT 71.370 95.580 71.690 95.840 ;
        RECT 5.520 94.960 84.180 95.440 ;
        RECT 10.650 94.760 10.970 94.820 ;
        RECT 11.125 94.760 11.415 94.805 ;
        RECT 10.650 94.620 11.415 94.760 ;
        RECT 10.650 94.560 10.970 94.620 ;
        RECT 11.125 94.575 11.415 94.620 ;
        RECT 11.570 94.560 11.890 94.820 ;
        RECT 29.970 94.760 30.290 94.820 ;
        RECT 33.665 94.760 33.955 94.805 ;
        RECT 29.970 94.620 33.955 94.760 ;
        RECT 29.970 94.560 30.290 94.620 ;
        RECT 33.665 94.575 33.955 94.620 ;
        RECT 40.105 94.760 40.395 94.805 ;
        RECT 40.550 94.760 40.870 94.820 ;
        RECT 40.105 94.620 40.870 94.760 ;
        RECT 40.105 94.575 40.395 94.620 ;
        RECT 40.550 94.560 40.870 94.620 ;
        RECT 60.345 94.760 60.635 94.805 ;
        RECT 61.250 94.760 61.570 94.820 ;
        RECT 60.345 94.620 61.570 94.760 ;
        RECT 60.345 94.575 60.635 94.620 ;
        RECT 61.250 94.560 61.570 94.620 ;
        RECT 66.770 94.560 67.090 94.820 ;
        RECT 67.230 94.760 67.550 94.820 ;
        RECT 68.165 94.760 68.455 94.805 ;
        RECT 70.450 94.760 70.770 94.820 ;
        RECT 67.230 94.620 68.455 94.760 ;
        RECT 67.230 94.560 67.550 94.620 ;
        RECT 68.165 94.575 68.455 94.620 ;
        RECT 69.620 94.620 70.770 94.760 ;
        RECT 26.790 94.420 27.080 94.465 ;
        RECT 28.890 94.420 29.180 94.465 ;
        RECT 30.460 94.420 30.750 94.465 ;
        RECT 26.790 94.280 30.750 94.420 ;
        RECT 26.790 94.235 27.080 94.280 ;
        RECT 28.890 94.235 29.180 94.280 ;
        RECT 30.460 94.235 30.750 94.280 ;
        RECT 33.205 94.420 33.495 94.465 ;
        RECT 42.850 94.420 43.170 94.480 ;
        RECT 66.310 94.420 66.630 94.480 ;
        RECT 69.620 94.420 69.760 94.620 ;
        RECT 70.450 94.560 70.770 94.620 ;
        RECT 75.065 94.760 75.355 94.805 ;
        RECT 76.890 94.760 77.210 94.820 ;
        RECT 75.065 94.620 77.210 94.760 ;
        RECT 75.065 94.575 75.355 94.620 ;
        RECT 76.890 94.560 77.210 94.620 ;
        RECT 33.205 94.280 36.640 94.420 ;
        RECT 33.205 94.235 33.495 94.280 ;
        RECT 12.045 94.080 12.335 94.125 ;
        RECT 12.505 94.080 12.795 94.125 ;
        RECT 12.045 93.940 12.795 94.080 ;
        RECT 12.045 93.895 12.335 93.940 ;
        RECT 12.505 93.895 12.795 93.940 ;
        RECT 18.930 94.080 19.250 94.140 ;
        RECT 36.500 94.125 36.640 94.280 ;
        RECT 42.850 94.280 46.760 94.420 ;
        RECT 42.850 94.220 43.170 94.280 ;
        RECT 26.305 94.080 26.595 94.125 ;
        RECT 18.930 93.940 26.595 94.080 ;
        RECT 18.930 93.880 19.250 93.940 ;
        RECT 26.305 93.895 26.595 93.940 ;
        RECT 27.185 94.080 27.475 94.125 ;
        RECT 28.375 94.080 28.665 94.125 ;
        RECT 30.895 94.080 31.185 94.125 ;
        RECT 27.185 93.940 31.185 94.080 ;
        RECT 27.185 93.895 27.475 93.940 ;
        RECT 28.375 93.895 28.665 93.940 ;
        RECT 30.895 93.895 31.185 93.940 ;
        RECT 36.425 94.080 36.715 94.125 ;
        RECT 37.330 94.080 37.650 94.140 ;
        RECT 36.425 93.940 37.650 94.080 ;
        RECT 36.425 93.895 36.715 93.940 ;
        RECT 37.330 93.880 37.650 93.940 ;
        RECT 43.310 93.880 43.630 94.140 ;
        RECT 10.665 93.555 10.955 93.785 ;
        RECT 13.870 93.740 14.190 93.800 ;
        RECT 15.265 93.740 15.555 93.785 ;
        RECT 13.870 93.600 15.555 93.740 ;
        RECT 10.740 93.400 10.880 93.555 ;
        RECT 13.870 93.540 14.190 93.600 ;
        RECT 15.265 93.555 15.555 93.600 ;
        RECT 42.405 93.740 42.695 93.785 ;
        RECT 44.230 93.740 44.550 93.800 ;
        RECT 46.620 93.785 46.760 94.280 ;
        RECT 66.310 94.280 69.760 94.420 ;
        RECT 69.990 94.420 70.310 94.480 ;
        RECT 69.990 94.280 72.980 94.420 ;
        RECT 66.310 94.220 66.630 94.280 ;
        RECT 69.990 94.220 70.310 94.280 ;
        RECT 47.910 94.080 48.230 94.140 ;
        RECT 50.670 94.080 50.990 94.140 ;
        RECT 47.910 93.940 50.990 94.080 ;
        RECT 47.910 93.880 48.230 93.940 ;
        RECT 50.670 93.880 50.990 93.940 ;
        RECT 57.570 94.080 57.890 94.140 ;
        RECT 57.570 93.940 61.940 94.080 ;
        RECT 57.570 93.880 57.890 93.940 ;
        RECT 61.800 93.800 61.940 93.940 ;
        RECT 72.290 93.880 72.610 94.140 ;
        RECT 72.840 94.125 72.980 94.280 ;
        RECT 72.765 93.895 73.055 94.125 ;
        RECT 42.405 93.600 44.550 93.740 ;
        RECT 42.405 93.555 42.695 93.600 ;
        RECT 44.230 93.540 44.550 93.600 ;
        RECT 46.545 93.555 46.835 93.785 ;
        RECT 53.890 93.540 54.210 93.800 ;
        RECT 57.125 93.740 57.415 93.785 ;
        RECT 60.330 93.740 60.650 93.800 ;
        RECT 57.125 93.600 60.650 93.740 ;
        RECT 57.125 93.555 57.415 93.600 ;
        RECT 60.330 93.540 60.650 93.600 ;
        RECT 61.710 93.540 62.030 93.800 ;
        RECT 62.630 93.540 62.950 93.800 ;
        RECT 64.930 93.740 65.250 93.800 ;
        RECT 66.325 93.740 66.615 93.785 ;
        RECT 64.930 93.600 66.615 93.740 ;
        RECT 64.930 93.540 65.250 93.600 ;
        RECT 66.325 93.555 66.615 93.600 ;
        RECT 66.770 93.540 67.090 93.800 ;
        RECT 14.790 93.400 15.110 93.460 ;
        RECT 17.550 93.400 17.870 93.460 ;
        RECT 27.670 93.445 27.990 93.460 ;
        RECT 10.740 93.260 17.870 93.400 ;
        RECT 14.790 93.200 15.110 93.260 ;
        RECT 17.550 93.200 17.870 93.260 ;
        RECT 27.640 93.215 27.990 93.445 ;
        RECT 41.945 93.400 42.235 93.445 ;
        RECT 47.005 93.400 47.295 93.445 ;
        RECT 47.450 93.400 47.770 93.460 ;
        RECT 41.945 93.260 44.920 93.400 ;
        RECT 41.945 93.215 42.235 93.260 ;
        RECT 27.670 93.200 27.990 93.215 ;
        RECT 44.780 93.105 44.920 93.260 ;
        RECT 47.005 93.260 47.770 93.400 ;
        RECT 47.005 93.215 47.295 93.260 ;
        RECT 47.450 93.200 47.770 93.260 ;
        RECT 60.790 93.400 61.110 93.460 ;
        RECT 61.265 93.400 61.555 93.445 ;
        RECT 64.470 93.400 64.790 93.460 ;
        RECT 60.790 93.260 61.555 93.400 ;
        RECT 60.790 93.200 61.110 93.260 ;
        RECT 61.265 93.215 61.555 93.260 ;
        RECT 61.800 93.260 64.790 93.400 ;
        RECT 44.705 92.875 44.995 93.105 ;
        RECT 59.410 92.860 59.730 93.120 ;
        RECT 60.265 93.060 60.555 93.105 ;
        RECT 61.800 93.060 61.940 93.260 ;
        RECT 64.470 93.200 64.790 93.260 ;
        RECT 60.265 92.920 61.940 93.060 ;
        RECT 62.170 93.060 62.490 93.120 ;
        RECT 68.610 93.060 68.930 93.120 ;
        RECT 62.170 92.920 68.930 93.060 ;
        RECT 60.265 92.875 60.555 92.920 ;
        RECT 62.170 92.860 62.490 92.920 ;
        RECT 68.610 92.860 68.930 92.920 ;
        RECT 73.210 92.860 73.530 93.120 ;
        RECT 5.520 92.240 84.180 92.720 ;
        RECT 14.805 92.040 15.095 92.085 ;
        RECT 15.250 92.040 15.570 92.100 ;
        RECT 18.470 92.040 18.790 92.100 ;
        RECT 14.805 91.900 18.790 92.040 ;
        RECT 14.805 91.855 15.095 91.900 ;
        RECT 15.250 91.840 15.570 91.900 ;
        RECT 18.470 91.840 18.790 91.900 ;
        RECT 25.385 92.040 25.675 92.085 ;
        RECT 26.290 92.040 26.610 92.100 ;
        RECT 25.385 91.900 26.610 92.040 ;
        RECT 25.385 91.855 25.675 91.900 ;
        RECT 26.290 91.840 26.610 91.900 ;
        RECT 27.225 92.040 27.515 92.085 ;
        RECT 27.670 92.040 27.990 92.100 ;
        RECT 37.330 92.085 37.650 92.100 ;
        RECT 27.225 91.900 27.990 92.040 ;
        RECT 27.225 91.855 27.515 91.900 ;
        RECT 27.670 91.840 27.990 91.900 ;
        RECT 29.065 92.040 29.355 92.085 ;
        RECT 32.285 92.040 32.575 92.085 ;
        RECT 29.065 91.900 32.575 92.040 ;
        RECT 29.065 91.855 29.355 91.900 ;
        RECT 32.285 91.855 32.575 91.900 ;
        RECT 37.330 91.855 37.715 92.085 ;
        RECT 47.465 92.040 47.755 92.085 ;
        RECT 53.890 92.040 54.210 92.100 ;
        RECT 47.465 91.900 54.210 92.040 ;
        RECT 47.465 91.855 47.755 91.900 ;
        RECT 37.330 91.840 37.650 91.855 ;
        RECT 10.650 91.700 10.970 91.760 ;
        RECT 29.525 91.700 29.815 91.745 ;
        RECT 29.970 91.700 30.290 91.760 ;
        RECT 10.650 91.560 13.180 91.700 ;
        RECT 10.650 91.500 10.970 91.560 ;
        RECT 13.040 91.405 13.180 91.560 ;
        RECT 29.525 91.560 30.290 91.700 ;
        RECT 29.525 91.515 29.815 91.560 ;
        RECT 29.970 91.500 30.290 91.560 ;
        RECT 36.410 91.500 36.730 91.760 ;
        RECT 10.205 91.360 10.495 91.405 ;
        RECT 10.205 91.220 12.720 91.360 ;
        RECT 10.205 91.175 10.495 91.220 ;
        RECT 10.665 90.835 10.955 91.065 ;
        RECT 10.740 90.680 10.880 90.835 ;
        RECT 11.110 90.820 11.430 91.080 ;
        RECT 12.580 91.020 12.720 91.220 ;
        RECT 12.965 91.175 13.255 91.405 ;
        RECT 13.885 91.360 14.175 91.405 ;
        RECT 14.790 91.360 15.110 91.420 ;
        RECT 13.885 91.220 15.110 91.360 ;
        RECT 13.885 91.175 14.175 91.220 ;
        RECT 14.790 91.160 15.110 91.220 ;
        RECT 18.485 91.360 18.775 91.405 ;
        RECT 18.930 91.360 19.250 91.420 ;
        RECT 19.850 91.405 20.170 91.420 ;
        RECT 18.485 91.220 19.250 91.360 ;
        RECT 18.485 91.175 18.775 91.220 ;
        RECT 18.930 91.160 19.250 91.220 ;
        RECT 19.820 91.175 20.170 91.405 ;
        RECT 19.850 91.160 20.170 91.175 ;
        RECT 34.110 91.160 34.430 91.420 ;
        RECT 34.585 91.360 34.875 91.405 ;
        RECT 47.540 91.360 47.680 91.855 ;
        RECT 53.890 91.840 54.210 91.900 ;
        RECT 57.585 91.855 57.875 92.085 ;
        RECT 68.165 92.040 68.455 92.085 ;
        RECT 73.210 92.040 73.530 92.100 ;
        RECT 68.165 91.900 73.530 92.040 ;
        RECT 68.165 91.855 68.455 91.900 ;
        RECT 53.140 91.700 53.430 91.745 ;
        RECT 57.660 91.700 57.800 91.855 ;
        RECT 73.210 91.840 73.530 91.900 ;
        RECT 74.605 92.040 74.895 92.085 ;
        RECT 75.050 92.040 75.370 92.100 ;
        RECT 74.605 91.900 75.370 92.040 ;
        RECT 74.605 91.855 74.895 91.900 ;
        RECT 75.050 91.840 75.370 91.900 ;
        RECT 53.140 91.560 57.800 91.700 ;
        RECT 53.140 91.515 53.430 91.560 ;
        RECT 58.950 91.500 59.270 91.760 ;
        RECT 59.425 91.700 59.715 91.745 ;
        RECT 61.265 91.700 61.555 91.745 ;
        RECT 59.425 91.560 61.555 91.700 ;
        RECT 59.425 91.515 59.715 91.560 ;
        RECT 61.265 91.515 61.555 91.560 ;
        RECT 63.180 91.560 73.440 91.700 ;
        RECT 34.585 91.220 47.680 91.360 ;
        RECT 48.460 91.220 55.040 91.360 ;
        RECT 34.585 91.175 34.875 91.220 ;
        RECT 13.410 91.020 13.730 91.080 ;
        RECT 17.550 91.020 17.870 91.080 ;
        RECT 12.580 90.880 17.870 91.020 ;
        RECT 13.410 90.820 13.730 90.880 ;
        RECT 17.550 90.820 17.870 90.880 ;
        RECT 19.365 91.020 19.655 91.065 ;
        RECT 20.555 91.020 20.845 91.065 ;
        RECT 23.075 91.020 23.365 91.065 ;
        RECT 19.365 90.880 23.365 91.020 ;
        RECT 19.365 90.835 19.655 90.880 ;
        RECT 20.555 90.835 20.845 90.880 ;
        RECT 23.075 90.835 23.365 90.880 ;
        RECT 30.430 90.820 30.750 91.080 ;
        RECT 35.505 91.020 35.795 91.065 ;
        RECT 47.910 91.020 48.230 91.080 ;
        RECT 35.505 90.880 48.230 91.020 ;
        RECT 35.505 90.835 35.795 90.880 ;
        RECT 47.910 90.820 48.230 90.880 ;
        RECT 14.790 90.680 15.110 90.740 ;
        RECT 17.090 90.680 17.410 90.740 ;
        RECT 18.970 90.680 19.260 90.725 ;
        RECT 21.070 90.680 21.360 90.725 ;
        RECT 22.640 90.680 22.930 90.725 ;
        RECT 48.460 90.680 48.600 91.220 ;
        RECT 49.775 91.020 50.065 91.065 ;
        RECT 52.295 91.020 52.585 91.065 ;
        RECT 53.485 91.020 53.775 91.065 ;
        RECT 49.775 90.880 53.775 91.020 ;
        RECT 49.775 90.835 50.065 90.880 ;
        RECT 52.295 90.835 52.585 90.880 ;
        RECT 53.485 90.835 53.775 90.880 ;
        RECT 54.365 90.835 54.655 91.065 ;
        RECT 10.740 90.540 18.700 90.680 ;
        RECT 14.790 90.480 15.110 90.540 ;
        RECT 17.090 90.480 17.410 90.540 ;
        RECT 8.350 90.140 8.670 90.400 ;
        RECT 13.870 90.140 14.190 90.400 ;
        RECT 18.560 90.340 18.700 90.540 ;
        RECT 18.970 90.540 22.930 90.680 ;
        RECT 18.970 90.495 19.260 90.540 ;
        RECT 21.070 90.495 21.360 90.540 ;
        RECT 22.640 90.495 22.930 90.540 ;
        RECT 23.620 90.540 48.600 90.680 ;
        RECT 50.210 90.680 50.500 90.725 ;
        RECT 51.780 90.680 52.070 90.725 ;
        RECT 53.880 90.680 54.170 90.725 ;
        RECT 50.210 90.540 54.170 90.680 ;
        RECT 23.620 90.340 23.760 90.540 ;
        RECT 50.210 90.495 50.500 90.540 ;
        RECT 51.780 90.495 52.070 90.540 ;
        RECT 53.880 90.495 54.170 90.540 ;
        RECT 18.560 90.200 23.760 90.340 ;
        RECT 37.330 90.140 37.650 90.400 ;
        RECT 38.265 90.340 38.555 90.385 ;
        RECT 40.550 90.340 40.870 90.400 ;
        RECT 38.265 90.200 40.870 90.340 ;
        RECT 38.265 90.155 38.555 90.200 ;
        RECT 40.550 90.140 40.870 90.200 ;
        RECT 49.290 90.340 49.610 90.400 ;
        RECT 54.440 90.340 54.580 90.835 ;
        RECT 54.900 90.680 55.040 91.220 ;
        RECT 58.505 91.175 58.795 91.405 ;
        RECT 58.580 91.020 58.720 91.175 ;
        RECT 60.330 91.160 60.650 91.420 ;
        RECT 62.170 91.160 62.490 91.420 ;
        RECT 62.630 91.160 62.950 91.420 ;
        RECT 61.250 91.020 61.570 91.080 ;
        RECT 58.580 90.880 61.570 91.020 ;
        RECT 61.250 90.820 61.570 90.880 ;
        RECT 63.180 90.680 63.320 91.560 ;
        RECT 63.565 91.175 63.855 91.405 ;
        RECT 63.640 91.020 63.780 91.175 ;
        RECT 64.010 91.160 64.330 91.420 ;
        RECT 64.930 91.360 65.250 91.420 ;
        RECT 66.325 91.360 66.615 91.405 ;
        RECT 64.930 91.220 66.615 91.360 ;
        RECT 64.930 91.160 65.250 91.220 ;
        RECT 66.325 91.175 66.615 91.220 ;
        RECT 68.610 91.160 68.930 91.420 ;
        RECT 69.545 91.360 69.835 91.405 ;
        RECT 69.990 91.360 70.310 91.420 ;
        RECT 69.545 91.220 70.310 91.360 ;
        RECT 69.545 91.175 69.835 91.220 ;
        RECT 69.990 91.160 70.310 91.220 ;
        RECT 70.465 91.360 70.755 91.405 ;
        RECT 71.845 91.360 72.135 91.405 ;
        RECT 70.465 91.220 72.135 91.360 ;
        RECT 70.465 91.175 70.755 91.220 ;
        RECT 71.845 91.175 72.135 91.220 ;
        RECT 72.290 91.360 72.610 91.420 ;
        RECT 73.300 91.405 73.440 91.560 ;
        RECT 72.765 91.360 73.055 91.405 ;
        RECT 72.290 91.220 73.055 91.360 ;
        RECT 72.290 91.160 72.610 91.220 ;
        RECT 72.765 91.175 73.055 91.220 ;
        RECT 73.225 91.175 73.515 91.405 ;
        RECT 73.685 91.175 73.975 91.405 ;
        RECT 65.390 91.020 65.710 91.080 ;
        RECT 63.640 90.880 65.710 91.020 ;
        RECT 65.390 90.820 65.710 90.880 ;
        RECT 66.785 90.835 67.075 91.065 ;
        RECT 69.070 91.020 69.390 91.080 ;
        RECT 71.370 91.020 71.690 91.080 ;
        RECT 73.760 91.020 73.900 91.175 ;
        RECT 69.070 90.880 73.900 91.020 ;
        RECT 54.900 90.540 63.320 90.680 ;
        RECT 66.860 90.680 67.000 90.835 ;
        RECT 69.070 90.820 69.390 90.880 ;
        RECT 71.370 90.820 71.690 90.880 ;
        RECT 69.990 90.680 70.310 90.740 ;
        RECT 66.860 90.540 70.310 90.680 ;
        RECT 69.990 90.480 70.310 90.540 ;
        RECT 49.290 90.200 54.580 90.340 ;
        RECT 59.410 90.340 59.730 90.400 ;
        RECT 61.710 90.340 62.030 90.400 ;
        RECT 64.010 90.340 64.330 90.400 ;
        RECT 59.410 90.200 64.330 90.340 ;
        RECT 49.290 90.140 49.610 90.200 ;
        RECT 59.410 90.140 59.730 90.200 ;
        RECT 61.710 90.140 62.030 90.200 ;
        RECT 64.010 90.140 64.330 90.200 ;
        RECT 67.245 90.340 67.535 90.385 ;
        RECT 70.910 90.340 71.230 90.400 ;
        RECT 67.245 90.200 71.230 90.340 ;
        RECT 67.245 90.155 67.535 90.200 ;
        RECT 70.910 90.140 71.230 90.200 ;
        RECT 5.520 89.520 84.180 90.000 ;
        RECT 13.885 89.320 14.175 89.365 ;
        RECT 14.790 89.320 15.110 89.380 ;
        RECT 13.885 89.180 15.110 89.320 ;
        RECT 13.885 89.135 14.175 89.180 ;
        RECT 14.790 89.120 15.110 89.180 ;
        RECT 16.630 89.120 16.950 89.380 ;
        RECT 17.565 89.320 17.855 89.365 ;
        RECT 18.010 89.320 18.330 89.380 ;
        RECT 17.565 89.180 18.330 89.320 ;
        RECT 17.565 89.135 17.855 89.180 ;
        RECT 18.010 89.120 18.330 89.180 ;
        RECT 19.405 89.320 19.695 89.365 ;
        RECT 19.850 89.320 20.170 89.380 ;
        RECT 19.405 89.180 20.170 89.320 ;
        RECT 19.405 89.135 19.695 89.180 ;
        RECT 19.850 89.120 20.170 89.180 ;
        RECT 41.025 89.320 41.315 89.365 ;
        RECT 41.470 89.320 41.790 89.380 ;
        RECT 41.025 89.180 41.790 89.320 ;
        RECT 41.025 89.135 41.315 89.180 ;
        RECT 41.470 89.120 41.790 89.180 ;
        RECT 64.485 89.135 64.775 89.365 ;
        RECT 64.930 89.320 65.250 89.380 ;
        RECT 65.405 89.320 65.695 89.365 ;
        RECT 64.930 89.180 65.695 89.320 ;
        RECT 7.470 88.980 7.760 89.025 ;
        RECT 9.570 88.980 9.860 89.025 ;
        RECT 11.140 88.980 11.430 89.025 ;
        RECT 7.470 88.840 11.430 88.980 ;
        RECT 7.470 88.795 7.760 88.840 ;
        RECT 9.570 88.795 9.860 88.840 ;
        RECT 11.140 88.795 11.430 88.840 ;
        RECT 6.970 88.440 7.290 88.700 ;
        RECT 7.865 88.640 8.155 88.685 ;
        RECT 9.055 88.640 9.345 88.685 ;
        RECT 11.575 88.640 11.865 88.685 ;
        RECT 15.250 88.640 15.570 88.700 ;
        RECT 7.865 88.500 11.865 88.640 ;
        RECT 7.865 88.455 8.155 88.500 ;
        RECT 9.055 88.455 9.345 88.500 ;
        RECT 11.575 88.455 11.865 88.500 ;
        RECT 14.420 88.500 15.570 88.640 ;
        RECT 18.100 88.640 18.240 89.120 ;
        RECT 22.165 88.640 22.455 88.685 ;
        RECT 18.100 88.500 22.455 88.640 ;
        RECT 7.060 88.300 7.200 88.440 ;
        RECT 13.870 88.300 14.190 88.360 ;
        RECT 7.060 88.160 14.190 88.300 ;
        RECT 13.870 88.100 14.190 88.160 ;
        RECT 8.350 88.005 8.670 88.020 ;
        RECT 8.320 87.960 8.670 88.005 ;
        RECT 8.155 87.820 8.670 87.960 ;
        RECT 8.320 87.775 8.670 87.820 ;
        RECT 8.350 87.760 8.670 87.775 ;
        RECT 11.110 87.960 11.430 88.020 ;
        RECT 14.420 87.960 14.560 88.500 ;
        RECT 15.250 88.440 15.570 88.500 ;
        RECT 22.165 88.455 22.455 88.500 ;
        RECT 30.890 88.640 31.210 88.700 ;
        RECT 33.205 88.640 33.495 88.685 ;
        RECT 34.110 88.640 34.430 88.700 ;
        RECT 60.790 88.640 61.110 88.700 ;
        RECT 64.560 88.640 64.700 89.135 ;
        RECT 64.930 89.120 65.250 89.180 ;
        RECT 65.405 89.135 65.695 89.180 ;
        RECT 30.890 88.500 34.430 88.640 ;
        RECT 30.890 88.440 31.210 88.500 ;
        RECT 33.205 88.455 33.495 88.500 ;
        RECT 34.110 88.440 34.430 88.500 ;
        RECT 60.420 88.500 64.700 88.640 ;
        RECT 17.550 88.300 17.870 88.360 ;
        RECT 19.850 88.300 20.170 88.360 ;
        RECT 21.705 88.300 21.995 88.345 ;
        RECT 17.550 88.160 21.995 88.300 ;
        RECT 17.550 88.100 17.870 88.160 ;
        RECT 19.850 88.100 20.170 88.160 ;
        RECT 21.705 88.115 21.995 88.160 ;
        RECT 40.105 88.115 40.395 88.345 ;
        RECT 40.550 88.300 40.870 88.360 ;
        RECT 60.420 88.345 60.560 88.500 ;
        RECT 60.790 88.440 61.110 88.500 ;
        RECT 72.290 88.440 72.610 88.700 ;
        RECT 41.025 88.300 41.315 88.345 ;
        RECT 40.550 88.160 41.315 88.300 ;
        RECT 11.110 87.820 14.560 87.960 ;
        RECT 15.250 87.960 15.570 88.020 ;
        RECT 15.725 87.960 16.015 88.005 ;
        RECT 15.250 87.820 16.015 87.960 ;
        RECT 11.110 87.760 11.430 87.820 ;
        RECT 15.250 87.760 15.570 87.820 ;
        RECT 15.725 87.775 16.015 87.820 ;
        RECT 21.245 87.960 21.535 88.005 ;
        RECT 26.290 87.960 26.610 88.020 ;
        RECT 21.245 87.820 26.610 87.960 ;
        RECT 21.245 87.775 21.535 87.820 ;
        RECT 26.290 87.760 26.610 87.820 ;
        RECT 38.725 87.960 39.015 88.005 ;
        RECT 39.170 87.960 39.490 88.020 ;
        RECT 38.725 87.820 39.490 87.960 ;
        RECT 40.180 87.960 40.320 88.115 ;
        RECT 40.550 88.100 40.870 88.160 ;
        RECT 41.025 88.115 41.315 88.160 ;
        RECT 60.345 88.115 60.635 88.345 ;
        RECT 61.265 88.300 61.555 88.345 ;
        RECT 64.930 88.300 65.250 88.360 ;
        RECT 61.265 88.160 65.250 88.300 ;
        RECT 61.265 88.115 61.555 88.160 ;
        RECT 64.640 88.100 65.250 88.160 ;
        RECT 70.910 88.100 71.230 88.360 ;
        RECT 71.370 88.100 71.690 88.360 ;
        RECT 73.685 88.300 73.975 88.345 ;
        RECT 74.130 88.300 74.450 88.360 ;
        RECT 73.685 88.160 74.450 88.300 ;
        RECT 73.685 88.115 73.975 88.160 ;
        RECT 74.130 88.100 74.450 88.160 ;
        RECT 81.950 88.100 82.270 88.360 ;
        RECT 44.690 87.960 45.010 88.020 ;
        RECT 40.180 87.820 45.010 87.960 ;
        RECT 38.725 87.775 39.015 87.820 ;
        RECT 39.170 87.760 39.490 87.820 ;
        RECT 44.690 87.760 45.010 87.820 ;
        RECT 59.410 87.760 59.730 88.020 ;
        RECT 62.630 87.960 62.950 88.020 ;
        RECT 63.565 87.960 63.855 88.005 ;
        RECT 64.640 87.990 65.005 88.100 ;
        RECT 62.630 87.820 63.855 87.960 ;
        RECT 64.715 87.945 65.005 87.990 ;
        RECT 62.630 87.760 62.950 87.820 ;
        RECT 63.565 87.775 63.855 87.820 ;
        RECT 14.330 87.620 14.650 87.680 ;
        RECT 16.725 87.620 17.015 87.665 ;
        RECT 14.330 87.480 17.015 87.620 ;
        RECT 14.330 87.420 14.650 87.480 ;
        RECT 16.725 87.435 17.015 87.480 ;
        RECT 33.650 87.620 33.970 87.680 ;
        RECT 35.965 87.620 36.255 87.665 ;
        RECT 33.650 87.480 36.255 87.620 ;
        RECT 33.650 87.420 33.970 87.480 ;
        RECT 35.965 87.435 36.255 87.480 ;
        RECT 41.930 87.420 42.250 87.680 ;
        RECT 62.170 87.620 62.490 87.680 ;
        RECT 69.990 87.620 70.310 87.680 ;
        RECT 73.225 87.620 73.515 87.665 ;
        RECT 62.170 87.480 73.515 87.620 ;
        RECT 62.170 87.420 62.490 87.480 ;
        RECT 69.990 87.420 70.310 87.480 ;
        RECT 73.225 87.435 73.515 87.480 ;
        RECT 79.190 87.420 79.510 87.680 ;
        RECT 5.520 86.800 84.180 87.280 ;
        RECT 9.285 86.600 9.575 86.645 ;
        RECT 10.650 86.600 10.970 86.660 ;
        RECT 16.630 86.600 16.950 86.660 ;
        RECT 9.285 86.460 10.970 86.600 ;
        RECT 9.285 86.415 9.575 86.460 ;
        RECT 10.650 86.400 10.970 86.460 ;
        RECT 11.200 86.460 16.950 86.600 ;
        RECT 11.200 86.260 11.340 86.460 ;
        RECT 16.630 86.400 16.950 86.460 ;
        RECT 18.470 86.600 18.790 86.660 ;
        RECT 18.470 86.460 19.160 86.600 ;
        RECT 18.470 86.400 18.790 86.460 ;
        RECT 13.870 86.260 14.190 86.320 ;
        RECT 19.020 86.305 19.160 86.460 ;
        RECT 30.890 86.400 31.210 86.660 ;
        RECT 31.825 86.415 32.115 86.645 ;
        RECT 10.280 86.120 11.340 86.260 ;
        RECT 11.660 86.120 18.700 86.260 ;
        RECT 10.280 84.945 10.420 86.120 ;
        RECT 11.110 85.720 11.430 85.980 ;
        RECT 11.660 85.965 11.800 86.120 ;
        RECT 13.870 86.060 14.190 86.120 ;
        RECT 11.585 85.735 11.875 85.965 ;
        RECT 12.920 85.920 13.210 85.965 ;
        RECT 14.330 85.920 14.650 85.980 ;
        RECT 12.920 85.780 14.650 85.920 ;
        RECT 18.560 85.920 18.700 86.120 ;
        RECT 18.945 86.075 19.235 86.305 ;
        RECT 19.390 86.260 19.710 86.320 ;
        RECT 19.945 86.260 20.235 86.305 ;
        RECT 19.390 86.120 20.235 86.260 ;
        RECT 19.390 86.060 19.710 86.120 ;
        RECT 19.945 86.075 20.235 86.120 ;
        RECT 25.340 86.260 25.630 86.305 ;
        RECT 31.900 86.260 32.040 86.415 ;
        RECT 33.650 86.400 33.970 86.660 ;
        RECT 35.030 86.600 35.350 86.660 ;
        RECT 37.805 86.600 38.095 86.645 ;
        RECT 35.030 86.460 38.095 86.600 ;
        RECT 35.030 86.400 35.350 86.460 ;
        RECT 37.805 86.415 38.095 86.460 ;
        RECT 41.470 86.400 41.790 86.660 ;
        RECT 44.230 86.600 44.550 86.660 ;
        RECT 42.020 86.460 44.550 86.600 ;
        RECT 42.020 86.260 42.160 86.460 ;
        RECT 44.230 86.400 44.550 86.460 ;
        RECT 44.690 86.400 45.010 86.660 ;
        RECT 56.205 86.600 56.495 86.645 ;
        RECT 60.790 86.600 61.110 86.660 ;
        RECT 56.205 86.460 61.110 86.600 ;
        RECT 56.205 86.415 56.495 86.460 ;
        RECT 60.790 86.400 61.110 86.460 ;
        RECT 64.470 86.400 64.790 86.660 ;
        RECT 66.325 86.600 66.615 86.645 ;
        RECT 66.770 86.600 67.090 86.660 ;
        RECT 66.325 86.460 67.090 86.600 ;
        RECT 66.325 86.415 66.615 86.460 ;
        RECT 66.770 86.400 67.090 86.460 ;
        RECT 79.650 86.600 79.970 86.660 ;
        RECT 80.585 86.600 80.875 86.645 ;
        RECT 81.950 86.600 82.270 86.660 ;
        RECT 79.650 86.460 82.270 86.600 ;
        RECT 79.650 86.400 79.970 86.460 ;
        RECT 80.585 86.415 80.875 86.460 ;
        RECT 81.950 86.400 82.270 86.460 ;
        RECT 25.340 86.120 32.040 86.260 ;
        RECT 39.260 86.120 42.160 86.260 ;
        RECT 42.405 86.260 42.695 86.305 ;
        RECT 48.830 86.260 49.150 86.320 ;
        RECT 42.405 86.120 49.150 86.260 ;
        RECT 25.340 86.075 25.630 86.120 ;
        RECT 36.410 85.920 36.730 85.980 ;
        RECT 39.260 85.965 39.400 86.120 ;
        RECT 42.405 86.075 42.695 86.120 ;
        RECT 48.830 86.060 49.150 86.120 ;
        RECT 59.425 86.260 59.715 86.305 ;
        RECT 61.710 86.260 62.030 86.320 ;
        RECT 59.425 86.120 65.620 86.260 ;
        RECT 59.425 86.075 59.715 86.120 ;
        RECT 61.710 86.060 62.030 86.120 ;
        RECT 39.185 85.920 39.475 85.965 ;
        RECT 18.560 85.780 19.160 85.920 ;
        RECT 12.920 85.735 13.210 85.780 ;
        RECT 14.330 85.720 14.650 85.780 ;
        RECT 19.020 85.640 19.160 85.780 ;
        RECT 36.410 85.780 39.475 85.920 ;
        RECT 36.410 85.720 36.730 85.780 ;
        RECT 39.185 85.735 39.475 85.780 ;
        RECT 39.645 85.735 39.935 85.965 ;
        RECT 10.665 85.395 10.955 85.625 ;
        RECT 12.465 85.580 12.755 85.625 ;
        RECT 13.655 85.580 13.945 85.625 ;
        RECT 16.175 85.580 16.465 85.625 ;
        RECT 12.465 85.440 16.465 85.580 ;
        RECT 12.465 85.395 12.755 85.440 ;
        RECT 13.655 85.395 13.945 85.440 ;
        RECT 16.175 85.395 16.465 85.440 ;
        RECT 18.930 85.580 19.250 85.640 ;
        RECT 24.005 85.580 24.295 85.625 ;
        RECT 18.930 85.440 24.295 85.580 ;
        RECT 10.205 84.715 10.495 84.945 ;
        RECT 10.740 84.900 10.880 85.395 ;
        RECT 18.930 85.380 19.250 85.440 ;
        RECT 24.005 85.395 24.295 85.440 ;
        RECT 24.885 85.580 25.175 85.625 ;
        RECT 26.075 85.580 26.365 85.625 ;
        RECT 28.595 85.580 28.885 85.625 ;
        RECT 24.885 85.440 28.885 85.580 ;
        RECT 24.885 85.395 25.175 85.440 ;
        RECT 26.075 85.395 26.365 85.440 ;
        RECT 28.595 85.395 28.885 85.440 ;
        RECT 29.050 85.580 29.370 85.640 ;
        RECT 34.125 85.580 34.415 85.625 ;
        RECT 29.050 85.440 34.415 85.580 ;
        RECT 29.050 85.380 29.370 85.440 ;
        RECT 34.125 85.395 34.415 85.440 ;
        RECT 35.045 85.395 35.335 85.625 ;
        RECT 39.720 85.580 39.860 85.735 ;
        RECT 40.090 85.720 40.410 85.980 ;
        RECT 41.025 85.920 41.315 85.965 ;
        RECT 41.930 85.920 42.250 85.980 ;
        RECT 41.025 85.780 42.250 85.920 ;
        RECT 41.025 85.735 41.315 85.780 ;
        RECT 41.930 85.720 42.250 85.780 ;
        RECT 44.230 85.720 44.550 85.980 ;
        RECT 50.640 85.920 50.930 85.965 ;
        RECT 57.585 85.920 57.875 85.965 ;
        RECT 50.640 85.780 57.875 85.920 ;
        RECT 50.640 85.735 50.930 85.780 ;
        RECT 57.585 85.735 57.875 85.780 ;
        RECT 58.490 85.720 58.810 85.980 ;
        RECT 58.950 85.720 59.270 85.980 ;
        RECT 60.015 85.920 60.305 85.965 ;
        RECT 59.500 85.780 60.305 85.920 ;
        RECT 47.005 85.580 47.295 85.625 ;
        RECT 39.720 85.440 47.295 85.580 ;
        RECT 12.070 85.240 12.360 85.285 ;
        RECT 14.170 85.240 14.460 85.285 ;
        RECT 15.740 85.240 16.030 85.285 ;
        RECT 12.070 85.100 16.030 85.240 ;
        RECT 12.070 85.055 12.360 85.100 ;
        RECT 14.170 85.055 14.460 85.100 ;
        RECT 15.740 85.055 16.030 85.100 ;
        RECT 16.630 85.240 16.950 85.300 ;
        RECT 24.490 85.240 24.780 85.285 ;
        RECT 26.590 85.240 26.880 85.285 ;
        RECT 28.160 85.240 28.450 85.285 ;
        RECT 16.630 85.100 20.080 85.240 ;
        RECT 16.630 85.040 16.950 85.100 ;
        RECT 15.250 84.900 15.570 84.960 ;
        RECT 18.470 84.900 18.790 84.960 ;
        RECT 19.940 84.945 20.080 85.100 ;
        RECT 24.490 85.100 28.450 85.240 ;
        RECT 35.120 85.240 35.260 85.395 ;
        RECT 41.470 85.240 41.790 85.300 ;
        RECT 35.120 85.100 41.790 85.240 ;
        RECT 24.490 85.055 24.780 85.100 ;
        RECT 26.590 85.055 26.880 85.100 ;
        RECT 28.160 85.055 28.450 85.100 ;
        RECT 41.470 85.040 41.790 85.100 ;
        RECT 42.480 84.960 42.620 85.440 ;
        RECT 47.005 85.395 47.295 85.440 ;
        RECT 49.290 85.380 49.610 85.640 ;
        RECT 50.185 85.580 50.475 85.625 ;
        RECT 51.375 85.580 51.665 85.625 ;
        RECT 53.895 85.580 54.185 85.625 ;
        RECT 50.185 85.440 54.185 85.580 ;
        RECT 50.185 85.395 50.475 85.440 ;
        RECT 51.375 85.395 51.665 85.440 ;
        RECT 53.895 85.395 54.185 85.440 ;
        RECT 58.030 85.580 58.350 85.640 ;
        RECT 59.500 85.580 59.640 85.780 ;
        RECT 60.015 85.735 60.305 85.780 ;
        RECT 60.790 85.920 61.110 85.980 ;
        RECT 62.185 85.920 62.475 85.965 ;
        RECT 62.630 85.920 62.950 85.980 ;
        RECT 60.790 85.780 62.950 85.920 ;
        RECT 60.790 85.720 61.110 85.780 ;
        RECT 62.185 85.735 62.475 85.780 ;
        RECT 62.630 85.720 62.950 85.780 ;
        RECT 64.930 85.720 65.250 85.980 ;
        RECT 65.480 85.965 65.620 86.120 ;
        RECT 65.405 85.735 65.695 85.965 ;
        RECT 66.860 85.920 67.000 86.400 ;
        RECT 70.910 86.260 71.230 86.320 ;
        RECT 72.290 86.260 72.610 86.320 ;
        RECT 70.910 86.120 72.610 86.260 ;
        RECT 70.910 86.060 71.230 86.120 ;
        RECT 72.290 86.060 72.610 86.120 ;
        RECT 70.005 85.920 70.295 85.965 ;
        RECT 66.860 85.780 70.295 85.920 ;
        RECT 70.005 85.735 70.295 85.780 ;
        RECT 71.370 85.720 71.690 85.980 ;
        RECT 71.830 85.720 72.150 85.980 ;
        RECT 72.750 85.920 73.070 85.980 ;
        RECT 75.050 85.965 75.370 85.980 ;
        RECT 73.685 85.920 73.975 85.965 ;
        RECT 72.750 85.780 73.975 85.920 ;
        RECT 72.750 85.720 73.070 85.780 ;
        RECT 73.685 85.735 73.975 85.780 ;
        RECT 75.020 85.735 75.370 85.965 ;
        RECT 75.050 85.720 75.370 85.735 ;
        RECT 81.030 85.720 81.350 85.980 ;
        RECT 58.030 85.440 59.640 85.580 ;
        RECT 58.030 85.380 58.350 85.440 ;
        RECT 45.610 85.040 45.930 85.300 ;
        RECT 49.790 85.240 50.080 85.285 ;
        RECT 51.890 85.240 52.180 85.285 ;
        RECT 53.460 85.240 53.750 85.285 ;
        RECT 49.790 85.100 53.750 85.240 ;
        RECT 49.790 85.055 50.080 85.100 ;
        RECT 51.890 85.055 52.180 85.100 ;
        RECT 53.460 85.055 53.750 85.100 ;
        RECT 64.025 85.240 64.315 85.285 ;
        RECT 65.020 85.240 65.160 85.720 ;
        RECT 66.310 85.580 66.630 85.640 ;
        RECT 67.230 85.580 67.550 85.640 ;
        RECT 66.310 85.440 67.550 85.580 ;
        RECT 66.310 85.380 66.630 85.440 ;
        RECT 67.230 85.380 67.550 85.440 ;
        RECT 74.565 85.580 74.855 85.625 ;
        RECT 75.755 85.580 76.045 85.625 ;
        RECT 78.275 85.580 78.565 85.625 ;
        RECT 74.565 85.440 78.565 85.580 ;
        RECT 74.565 85.395 74.855 85.440 ;
        RECT 75.755 85.395 76.045 85.440 ;
        RECT 78.275 85.395 78.565 85.440 ;
        RECT 64.025 85.100 65.160 85.240 ;
        RECT 74.170 85.240 74.460 85.285 ;
        RECT 76.270 85.240 76.560 85.285 ;
        RECT 77.840 85.240 78.130 85.285 ;
        RECT 74.170 85.100 78.130 85.240 ;
        RECT 64.025 85.055 64.315 85.100 ;
        RECT 74.170 85.055 74.460 85.100 ;
        RECT 76.270 85.055 76.560 85.100 ;
        RECT 77.840 85.055 78.130 85.100 ;
        RECT 81.950 85.040 82.270 85.300 ;
        RECT 10.740 84.760 18.790 84.900 ;
        RECT 15.250 84.700 15.570 84.760 ;
        RECT 18.470 84.700 18.790 84.760 ;
        RECT 19.865 84.715 20.155 84.945 ;
        RECT 20.785 84.900 21.075 84.945 ;
        RECT 23.070 84.900 23.390 84.960 ;
        RECT 20.785 84.760 23.390 84.900 ;
        RECT 20.785 84.715 21.075 84.760 ;
        RECT 23.070 84.700 23.390 84.760 ;
        RECT 42.390 84.700 42.710 84.960 ;
        RECT 57.110 84.900 57.430 84.960 ;
        RECT 60.790 84.900 61.110 84.960 ;
        RECT 57.110 84.760 61.110 84.900 ;
        RECT 57.110 84.700 57.430 84.760 ;
        RECT 60.790 84.700 61.110 84.760 ;
        RECT 66.310 84.900 66.630 84.960 ;
        RECT 67.690 84.900 68.010 84.960 ;
        RECT 66.310 84.760 68.010 84.900 ;
        RECT 66.310 84.700 66.630 84.760 ;
        RECT 67.690 84.700 68.010 84.760 ;
        RECT 72.765 84.900 73.055 84.945 ;
        RECT 76.890 84.900 77.210 84.960 ;
        RECT 72.765 84.760 77.210 84.900 ;
        RECT 72.765 84.715 73.055 84.760 ;
        RECT 76.890 84.700 77.210 84.760 ;
        RECT 5.520 84.080 84.180 84.560 ;
        RECT 14.330 83.680 14.650 83.940 ;
        RECT 17.565 83.880 17.855 83.925 ;
        RECT 19.390 83.880 19.710 83.940 ;
        RECT 17.565 83.740 19.710 83.880 ;
        RECT 17.565 83.695 17.855 83.740 ;
        RECT 19.390 83.680 19.710 83.740 ;
        RECT 37.330 83.880 37.650 83.940 ;
        RECT 37.805 83.880 38.095 83.925 ;
        RECT 42.390 83.880 42.710 83.940 ;
        RECT 37.330 83.740 42.710 83.880 ;
        RECT 37.330 83.680 37.650 83.740 ;
        RECT 37.805 83.695 38.095 83.740 ;
        RECT 42.390 83.680 42.710 83.740 ;
        RECT 59.885 83.880 60.175 83.925 ;
        RECT 60.330 83.880 60.650 83.940 ;
        RECT 61.710 83.880 62.030 83.940 ;
        RECT 65.405 83.880 65.695 83.925 ;
        RECT 67.690 83.880 68.010 83.940 ;
        RECT 75.050 83.880 75.370 83.940 ;
        RECT 75.525 83.880 75.815 83.925 ;
        RECT 59.885 83.740 65.695 83.880 ;
        RECT 59.885 83.695 60.175 83.740 ;
        RECT 60.330 83.680 60.650 83.740 ;
        RECT 61.710 83.680 62.030 83.740 ;
        RECT 65.405 83.695 65.695 83.740 ;
        RECT 66.040 83.740 72.980 83.880 ;
        RECT 15.710 83.340 16.030 83.600 ;
        RECT 20.350 83.540 20.640 83.585 ;
        RECT 22.450 83.540 22.740 83.585 ;
        RECT 24.020 83.540 24.310 83.585 ;
        RECT 20.350 83.400 24.310 83.540 ;
        RECT 20.350 83.355 20.640 83.400 ;
        RECT 22.450 83.355 22.740 83.400 ;
        RECT 24.020 83.355 24.310 83.400 ;
        RECT 35.965 83.540 36.255 83.585 ;
        RECT 36.410 83.540 36.730 83.600 ;
        RECT 35.965 83.400 36.730 83.540 ;
        RECT 35.965 83.355 36.255 83.400 ;
        RECT 36.410 83.340 36.730 83.400 ;
        RECT 40.550 83.340 40.870 83.600 ;
        RECT 41.470 83.540 41.790 83.600 ;
        RECT 43.310 83.540 43.630 83.600 ;
        RECT 41.470 83.400 43.630 83.540 ;
        RECT 41.470 83.340 41.790 83.400 ;
        RECT 43.310 83.340 43.630 83.400 ;
        RECT 49.790 83.540 50.080 83.585 ;
        RECT 51.890 83.540 52.180 83.585 ;
        RECT 53.460 83.540 53.750 83.585 ;
        RECT 49.790 83.400 53.750 83.540 ;
        RECT 49.790 83.355 50.080 83.400 ;
        RECT 51.890 83.355 52.180 83.400 ;
        RECT 53.460 83.355 53.750 83.400 ;
        RECT 56.205 83.540 56.495 83.585 ;
        RECT 66.040 83.540 66.180 83.740 ;
        RECT 67.690 83.680 68.010 83.740 ;
        RECT 69.990 83.540 70.310 83.600 ;
        RECT 56.205 83.400 58.260 83.540 ;
        RECT 56.205 83.355 56.495 83.400 ;
        RECT 13.885 83.200 14.175 83.245 ;
        RECT 15.800 83.200 15.940 83.340 ;
        RECT 17.550 83.200 17.870 83.260 ;
        RECT 13.885 83.060 15.480 83.200 ;
        RECT 15.800 83.060 17.870 83.200 ;
        RECT 13.885 83.015 14.175 83.060 ;
        RECT 15.340 82.905 15.480 83.060 ;
        RECT 15.265 82.675 15.555 82.905 ;
        RECT 15.710 82.660 16.030 82.920 ;
        RECT 17.180 82.905 17.320 83.060 ;
        RECT 17.550 83.000 17.870 83.060 ;
        RECT 18.930 83.200 19.250 83.260 ;
        RECT 19.865 83.200 20.155 83.245 ;
        RECT 18.930 83.060 20.155 83.200 ;
        RECT 18.930 83.000 19.250 83.060 ;
        RECT 19.865 83.015 20.155 83.060 ;
        RECT 20.745 83.200 21.035 83.245 ;
        RECT 21.935 83.200 22.225 83.245 ;
        RECT 24.455 83.200 24.745 83.245 ;
        RECT 20.745 83.060 24.745 83.200 ;
        RECT 20.745 83.015 21.035 83.060 ;
        RECT 21.935 83.015 22.225 83.060 ;
        RECT 24.455 83.015 24.745 83.060 ;
        RECT 47.910 83.000 48.230 83.260 ;
        RECT 49.290 83.000 49.610 83.260 ;
        RECT 50.185 83.200 50.475 83.245 ;
        RECT 51.375 83.200 51.665 83.245 ;
        RECT 53.895 83.200 54.185 83.245 ;
        RECT 56.665 83.200 56.955 83.245 ;
        RECT 50.185 83.060 54.185 83.200 ;
        RECT 50.185 83.015 50.475 83.060 ;
        RECT 51.375 83.015 51.665 83.060 ;
        RECT 53.895 83.015 54.185 83.060 ;
        RECT 54.440 83.060 56.955 83.200 ;
        RECT 17.105 82.675 17.395 82.905 ;
        RECT 35.505 82.675 35.795 82.905 ;
        RECT 50.640 82.860 50.930 82.905 ;
        RECT 54.440 82.860 54.580 83.060 ;
        RECT 56.665 83.015 56.955 83.060 ;
        RECT 50.640 82.720 54.580 82.860 ;
        RECT 50.640 82.675 50.930 82.720 ;
        RECT 12.045 82.520 12.335 82.565 ;
        RECT 12.965 82.520 13.255 82.565 ;
        RECT 14.330 82.520 14.650 82.580 ;
        RECT 12.045 82.380 12.720 82.520 ;
        RECT 12.045 82.335 12.335 82.380 ;
        RECT 12.580 82.240 12.720 82.380 ;
        RECT 12.965 82.380 14.650 82.520 ;
        RECT 12.965 82.335 13.255 82.380 ;
        RECT 14.330 82.320 14.650 82.380 ;
        RECT 20.310 82.520 20.630 82.580 ;
        RECT 21.090 82.520 21.380 82.565 ;
        RECT 20.310 82.380 21.380 82.520 ;
        RECT 35.580 82.520 35.720 82.675 ;
        RECT 57.570 82.660 57.890 82.920 ;
        RECT 58.120 82.905 58.260 83.400 ;
        RECT 65.480 83.400 66.180 83.540 ;
        RECT 66.400 83.400 70.310 83.540 ;
        RECT 65.480 83.260 65.620 83.400 ;
        RECT 61.800 83.060 62.860 83.200 ;
        RECT 58.045 82.860 58.335 82.905 ;
        RECT 58.490 82.860 58.810 82.920 ;
        RECT 58.045 82.720 58.810 82.860 ;
        RECT 58.045 82.675 58.335 82.720 ;
        RECT 58.490 82.660 58.810 82.720 ;
        RECT 58.965 82.675 59.255 82.905 ;
        RECT 59.425 82.860 59.715 82.905 ;
        RECT 59.870 82.860 60.190 82.920 ;
        RECT 59.425 82.720 60.190 82.860 ;
        RECT 59.425 82.675 59.715 82.720 ;
        RECT 37.790 82.520 38.110 82.580 ;
        RECT 35.580 82.380 38.110 82.520 ;
        RECT 20.310 82.320 20.630 82.380 ;
        RECT 21.090 82.335 21.380 82.380 ;
        RECT 37.790 82.320 38.110 82.380 ;
        RECT 42.390 82.520 42.710 82.580 ;
        RECT 45.150 82.520 45.470 82.580 ;
        RECT 42.390 82.380 45.470 82.520 ;
        RECT 42.390 82.320 42.710 82.380 ;
        RECT 45.150 82.320 45.470 82.380 ;
        RECT 12.490 82.180 12.810 82.240 ;
        RECT 14.790 82.180 15.110 82.240 ;
        RECT 12.490 82.040 15.110 82.180 ;
        RECT 12.490 81.980 12.810 82.040 ;
        RECT 14.790 81.980 15.110 82.040 ;
        RECT 26.750 81.980 27.070 82.240 ;
        RECT 32.270 81.980 32.590 82.240 ;
        RECT 38.710 81.980 39.030 82.240 ;
        RECT 40.105 82.180 40.395 82.225 ;
        RECT 41.470 82.180 41.790 82.240 ;
        RECT 40.105 82.040 41.790 82.180 ;
        RECT 40.105 81.995 40.395 82.040 ;
        RECT 41.470 81.980 41.790 82.040 ;
        RECT 44.690 81.980 45.010 82.240 ;
        RECT 46.530 81.980 46.850 82.240 ;
        RECT 47.005 82.180 47.295 82.225 ;
        RECT 49.750 82.180 50.070 82.240 ;
        RECT 47.005 82.040 50.070 82.180 ;
        RECT 47.005 81.995 47.295 82.040 ;
        RECT 49.750 81.980 50.070 82.040 ;
        RECT 58.030 82.180 58.350 82.240 ;
        RECT 59.040 82.180 59.180 82.675 ;
        RECT 59.870 82.660 60.190 82.720 ;
        RECT 60.790 82.660 61.110 82.920 ;
        RECT 61.800 82.905 61.940 83.060 ;
        RECT 62.720 82.920 62.860 83.060 ;
        RECT 65.390 83.000 65.710 83.260 ;
        RECT 66.400 83.245 66.540 83.400 ;
        RECT 69.990 83.340 70.310 83.400 ;
        RECT 66.325 83.015 66.615 83.245 ;
        RECT 69.070 83.200 69.390 83.260 ;
        RECT 69.545 83.200 69.835 83.245 ;
        RECT 72.305 83.200 72.595 83.245 ;
        RECT 69.070 83.060 72.595 83.200 ;
        RECT 69.070 83.000 69.390 83.060 ;
        RECT 69.545 83.015 69.835 83.060 ;
        RECT 72.305 83.015 72.595 83.060 ;
        RECT 61.725 82.675 62.015 82.905 ;
        RECT 62.185 82.675 62.475 82.905 ;
        RECT 62.630 82.860 62.950 82.920 ;
        RECT 63.105 82.860 63.395 82.905 ;
        RECT 62.630 82.720 63.395 82.860 ;
        RECT 58.030 82.040 59.180 82.180 ;
        RECT 60.880 82.180 61.020 82.660 ;
        RECT 62.260 82.180 62.400 82.675 ;
        RECT 62.630 82.660 62.950 82.720 ;
        RECT 63.105 82.675 63.395 82.720 ;
        RECT 64.930 82.660 65.250 82.920 ;
        RECT 66.770 82.860 67.090 82.920 ;
        RECT 67.705 82.860 67.995 82.905 ;
        RECT 66.770 82.720 67.995 82.860 ;
        RECT 66.770 82.660 67.090 82.720 ;
        RECT 67.705 82.675 67.995 82.720 ;
        RECT 70.465 82.675 70.755 82.905 ;
        RECT 71.385 82.675 71.675 82.905 ;
        RECT 71.845 82.860 72.135 82.905 ;
        RECT 72.840 82.860 72.980 83.740 ;
        RECT 75.050 83.740 75.815 83.880 ;
        RECT 75.050 83.680 75.370 83.740 ;
        RECT 75.525 83.695 75.815 83.740 ;
        RECT 80.585 83.880 80.875 83.925 ;
        RECT 81.030 83.880 81.350 83.940 ;
        RECT 80.585 83.740 81.350 83.880 ;
        RECT 80.585 83.695 80.875 83.740 ;
        RECT 81.030 83.680 81.350 83.740 ;
        RECT 74.145 83.200 74.435 83.245 ;
        RECT 78.285 83.200 78.575 83.245 ;
        RECT 74.145 83.060 78.575 83.200 ;
        RECT 74.145 83.015 74.435 83.060 ;
        RECT 78.285 83.015 78.575 83.060 ;
        RECT 71.845 82.720 72.980 82.860 ;
        RECT 73.225 82.860 73.515 82.905 ;
        RECT 73.670 82.860 73.990 82.920 ;
        RECT 73.225 82.720 73.990 82.860 ;
        RECT 71.845 82.675 72.135 82.720 ;
        RECT 73.225 82.675 73.515 82.720 ;
        RECT 68.610 82.320 68.930 82.580 ;
        RECT 69.530 82.520 69.850 82.580 ;
        RECT 70.540 82.520 70.680 82.675 ;
        RECT 69.530 82.380 70.680 82.520 ;
        RECT 69.530 82.320 69.850 82.380 ;
        RECT 60.880 82.040 62.400 82.180 ;
        RECT 58.030 81.980 58.350 82.040 ;
        RECT 62.630 81.980 62.950 82.240 ;
        RECT 66.325 82.180 66.615 82.225 ;
        RECT 68.150 82.180 68.470 82.240 ;
        RECT 71.460 82.180 71.600 82.675 ;
        RECT 73.670 82.660 73.990 82.720 ;
        RECT 77.365 82.860 77.655 82.905 ;
        RECT 79.190 82.860 79.510 82.920 ;
        RECT 77.365 82.720 79.510 82.860 ;
        RECT 77.365 82.675 77.655 82.720 ;
        RECT 79.190 82.660 79.510 82.720 ;
        RECT 79.650 82.660 79.970 82.920 ;
        RECT 76.890 82.520 77.210 82.580 ;
        RECT 77.825 82.520 78.115 82.565 ;
        RECT 76.890 82.380 78.115 82.520 ;
        RECT 76.890 82.320 77.210 82.380 ;
        RECT 77.825 82.335 78.115 82.380 ;
        RECT 66.325 82.040 71.600 82.180 ;
        RECT 66.325 81.995 66.615 82.040 ;
        RECT 68.150 81.980 68.470 82.040 ;
        RECT 5.520 81.360 84.180 81.840 ;
        RECT 20.310 80.960 20.630 81.220 ;
        RECT 37.790 81.160 38.110 81.220 ;
        RECT 38.725 81.160 39.015 81.205 ;
        RECT 37.790 81.020 39.015 81.160 ;
        RECT 37.790 80.960 38.110 81.020 ;
        RECT 38.725 80.975 39.015 81.020 ;
        RECT 39.185 81.160 39.475 81.205 ;
        RECT 40.090 81.160 40.410 81.220 ;
        RECT 39.185 81.020 40.410 81.160 ;
        RECT 39.185 80.975 39.475 81.020 ;
        RECT 40.090 80.960 40.410 81.020 ;
        RECT 48.830 81.160 49.150 81.220 ;
        RECT 49.305 81.160 49.595 81.205 ;
        RECT 48.830 81.020 49.595 81.160 ;
        RECT 48.830 80.960 49.150 81.020 ;
        RECT 49.305 80.975 49.595 81.020 ;
        RECT 19.850 80.820 20.170 80.880 ;
        RECT 22.625 80.820 22.915 80.865 ;
        RECT 34.570 80.820 34.890 80.880 ;
        RECT 41.010 80.820 41.330 80.880 ;
        RECT 19.850 80.680 22.915 80.820 ;
        RECT 19.850 80.620 20.170 80.680 ;
        RECT 22.625 80.635 22.915 80.680 ;
        RECT 31.900 80.680 41.330 80.820 ;
        RECT 22.165 80.480 22.455 80.525 ;
        RECT 23.530 80.480 23.850 80.540 ;
        RECT 26.750 80.480 27.070 80.540 ;
        RECT 31.900 80.525 32.040 80.680 ;
        RECT 34.570 80.620 34.890 80.680 ;
        RECT 41.010 80.620 41.330 80.680 ;
        RECT 41.470 80.620 41.790 80.880 ;
        RECT 43.740 80.820 44.030 80.865 ;
        RECT 44.690 80.820 45.010 80.880 ;
        RECT 43.740 80.680 45.010 80.820 ;
        RECT 43.740 80.635 44.030 80.680 ;
        RECT 44.690 80.620 45.010 80.680 ;
        RECT 33.190 80.525 33.510 80.540 ;
        RECT 22.165 80.340 27.070 80.480 ;
        RECT 22.165 80.295 22.455 80.340 ;
        RECT 23.530 80.280 23.850 80.340 ;
        RECT 26.750 80.280 27.070 80.340 ;
        RECT 31.825 80.295 32.115 80.525 ;
        RECT 33.160 80.295 33.510 80.525 ;
        RECT 33.190 80.280 33.510 80.295 ;
        RECT 39.170 80.480 39.490 80.540 ;
        RECT 40.105 80.480 40.395 80.525 ;
        RECT 39.170 80.340 40.395 80.480 ;
        RECT 49.380 80.480 49.520 80.975 ;
        RECT 49.750 80.960 50.070 81.220 ;
        RECT 58.950 81.160 59.270 81.220 ;
        RECT 60.345 81.160 60.635 81.205 ;
        RECT 61.250 81.160 61.570 81.220 ;
        RECT 62.630 81.160 62.950 81.220 ;
        RECT 58.950 81.020 62.950 81.160 ;
        RECT 58.950 80.960 59.270 81.020 ;
        RECT 60.345 80.975 60.635 81.020 ;
        RECT 61.250 80.960 61.570 81.020 ;
        RECT 62.630 80.960 62.950 81.020 ;
        RECT 63.550 81.160 63.870 81.220 ;
        RECT 66.310 81.160 66.630 81.220 ;
        RECT 68.035 81.160 68.325 81.205 ;
        RECT 63.550 81.020 68.325 81.160 ;
        RECT 63.550 80.960 63.870 81.020 ;
        RECT 66.310 80.960 66.630 81.020 ;
        RECT 68.035 80.975 68.325 81.020 ;
        RECT 64.025 80.820 64.315 80.865 ;
        RECT 64.930 80.820 65.250 80.880 ;
        RECT 58.625 80.680 65.250 80.820 ;
        RECT 58.625 80.540 58.765 80.680 ;
        RECT 64.025 80.635 64.315 80.680 ;
        RECT 64.930 80.620 65.250 80.680 ;
        RECT 69.070 80.620 69.390 80.880 ;
        RECT 52.525 80.480 52.815 80.525 ;
        RECT 49.380 80.340 52.815 80.480 ;
        RECT 39.170 80.280 39.490 80.340 ;
        RECT 40.105 80.295 40.395 80.340 ;
        RECT 52.525 80.295 52.815 80.340 ;
        RECT 58.490 80.280 58.810 80.540 ;
        RECT 71.370 80.480 71.690 80.540 ;
        RECT 59.040 80.340 71.690 80.480 ;
        RECT 23.070 79.940 23.390 80.200 ;
        RECT 32.705 80.140 32.995 80.185 ;
        RECT 33.895 80.140 34.185 80.185 ;
        RECT 36.415 80.140 36.705 80.185 ;
        RECT 32.705 80.000 36.705 80.140 ;
        RECT 32.705 79.955 32.995 80.000 ;
        RECT 33.895 79.955 34.185 80.000 ;
        RECT 36.415 79.955 36.705 80.000 ;
        RECT 38.710 80.140 39.030 80.200 ;
        RECT 40.565 80.140 40.855 80.185 ;
        RECT 38.710 80.000 40.855 80.140 ;
        RECT 38.710 79.940 39.030 80.000 ;
        RECT 40.565 79.955 40.855 80.000 ;
        RECT 41.010 80.140 41.330 80.200 ;
        RECT 42.405 80.140 42.695 80.185 ;
        RECT 41.010 80.000 42.695 80.140 ;
        RECT 41.010 79.940 41.330 80.000 ;
        RECT 42.405 79.955 42.695 80.000 ;
        RECT 43.285 80.140 43.575 80.185 ;
        RECT 44.475 80.140 44.765 80.185 ;
        RECT 46.995 80.140 47.285 80.185 ;
        RECT 43.285 80.000 47.285 80.140 ;
        RECT 43.285 79.955 43.575 80.000 ;
        RECT 44.475 79.955 44.765 80.000 ;
        RECT 46.995 79.955 47.285 80.000 ;
        RECT 32.310 79.800 32.600 79.845 ;
        RECT 34.410 79.800 34.700 79.845 ;
        RECT 35.980 79.800 36.270 79.845 ;
        RECT 42.890 79.800 43.180 79.845 ;
        RECT 44.990 79.800 45.280 79.845 ;
        RECT 46.560 79.800 46.850 79.845 ;
        RECT 32.310 79.660 36.270 79.800 ;
        RECT 32.310 79.615 32.600 79.660 ;
        RECT 34.410 79.615 34.700 79.660 ;
        RECT 35.980 79.615 36.270 79.660 ;
        RECT 36.500 79.660 42.115 79.800 ;
        RECT 26.750 79.460 27.070 79.520 ;
        RECT 36.500 79.460 36.640 79.660 ;
        RECT 26.750 79.320 36.640 79.460 ;
        RECT 26.750 79.260 27.070 79.320 ;
        RECT 41.470 79.260 41.790 79.520 ;
        RECT 41.975 79.460 42.115 79.660 ;
        RECT 42.890 79.660 46.850 79.800 ;
        RECT 42.890 79.615 43.180 79.660 ;
        RECT 44.990 79.615 45.280 79.660 ;
        RECT 46.560 79.615 46.850 79.660 ;
        RECT 59.040 79.460 59.180 80.340 ;
        RECT 71.370 80.280 71.690 80.340 ;
        RECT 77.825 80.480 78.115 80.525 ;
        RECT 80.570 80.480 80.890 80.540 ;
        RECT 81.965 80.480 82.255 80.525 ;
        RECT 77.825 80.340 82.255 80.480 ;
        RECT 77.825 80.295 78.115 80.340 ;
        RECT 80.570 80.280 80.890 80.340 ;
        RECT 81.965 80.295 82.255 80.340 ;
        RECT 64.470 80.140 64.790 80.200 ;
        RECT 61.340 80.000 64.790 80.140 ;
        RECT 61.340 79.845 61.480 80.000 ;
        RECT 64.470 79.940 64.790 80.000 ;
        RECT 61.265 79.615 61.555 79.845 ;
        RECT 62.170 79.600 62.490 79.860 ;
        RECT 66.770 79.800 67.090 79.860 ;
        RECT 64.640 79.660 67.090 79.800 ;
        RECT 41.975 79.320 59.180 79.460 ;
        RECT 60.330 79.260 60.650 79.520 ;
        RECT 61.725 79.460 62.015 79.505 ;
        RECT 64.640 79.460 64.780 79.660 ;
        RECT 66.770 79.600 67.090 79.660 ;
        RECT 61.725 79.320 64.780 79.460 ;
        RECT 64.930 79.460 65.250 79.520 ;
        RECT 67.245 79.460 67.535 79.505 ;
        RECT 64.930 79.320 67.535 79.460 ;
        RECT 61.725 79.275 62.015 79.320 ;
        RECT 64.930 79.260 65.250 79.320 ;
        RECT 67.245 79.275 67.535 79.320 ;
        RECT 68.150 79.260 68.470 79.520 ;
        RECT 78.730 79.260 79.050 79.520 ;
        RECT 79.190 79.260 79.510 79.520 ;
        RECT 5.520 78.640 84.180 79.120 ;
        RECT 14.790 78.440 15.110 78.500 ;
        RECT 15.725 78.440 16.015 78.485 ;
        RECT 16.630 78.440 16.950 78.500 ;
        RECT 11.200 78.300 16.950 78.440 ;
        RECT 11.200 77.805 11.340 78.300 ;
        RECT 14.790 78.240 15.110 78.300 ;
        RECT 15.725 78.255 16.015 78.300 ;
        RECT 16.630 78.240 16.950 78.300 ;
        RECT 33.190 78.440 33.510 78.500 ;
        RECT 34.585 78.440 34.875 78.485 ;
        RECT 33.190 78.300 34.875 78.440 ;
        RECT 33.190 78.240 33.510 78.300 ;
        RECT 34.585 78.255 34.875 78.300 ;
        RECT 41.470 78.440 41.790 78.500 ;
        RECT 44.705 78.440 44.995 78.485 ;
        RECT 41.470 78.300 44.995 78.440 ;
        RECT 41.470 78.240 41.790 78.300 ;
        RECT 44.705 78.255 44.995 78.300 ;
        RECT 45.150 78.440 45.470 78.500 ;
        RECT 45.625 78.440 45.915 78.485 ;
        RECT 45.150 78.300 45.915 78.440 ;
        RECT 45.150 78.240 45.470 78.300 ;
        RECT 45.625 78.255 45.915 78.300 ;
        RECT 46.530 78.440 46.850 78.500 ;
        RECT 47.005 78.440 47.295 78.485 ;
        RECT 46.530 78.300 47.295 78.440 ;
        RECT 46.530 78.240 46.850 78.300 ;
        RECT 47.005 78.255 47.295 78.300 ;
        RECT 60.330 78.440 60.650 78.500 ;
        RECT 61.265 78.440 61.555 78.485 ;
        RECT 60.330 78.300 61.555 78.440 ;
        RECT 60.330 78.240 60.650 78.300 ;
        RECT 61.265 78.255 61.555 78.300 ;
        RECT 69.545 78.440 69.835 78.485 ;
        RECT 78.270 78.440 78.590 78.500 ;
        RECT 69.545 78.300 78.590 78.440 ;
        RECT 69.545 78.255 69.835 78.300 ;
        RECT 78.270 78.240 78.590 78.300 ;
        RECT 80.570 78.240 80.890 78.500 ;
        RECT 81.950 78.240 82.270 78.500 ;
        RECT 14.330 78.100 14.650 78.160 ;
        RECT 18.025 78.100 18.315 78.145 ;
        RECT 27.670 78.100 27.990 78.160 ;
        RECT 65.850 78.100 66.170 78.160 ;
        RECT 69.070 78.100 69.390 78.160 ;
        RECT 11.660 77.960 16.860 78.100 ;
        RECT 11.125 77.575 11.415 77.805 ;
        RECT 11.660 77.465 11.800 77.960 ;
        RECT 14.330 77.900 14.650 77.960 ;
        RECT 12.045 77.760 12.335 77.805 ;
        RECT 15.710 77.760 16.030 77.820 ;
        RECT 12.045 77.620 16.030 77.760 ;
        RECT 12.045 77.575 12.335 77.620 ;
        RECT 10.205 77.235 10.495 77.465 ;
        RECT 11.585 77.235 11.875 77.465 ;
        RECT 10.280 77.080 10.420 77.235 ;
        RECT 12.490 77.220 12.810 77.480 ;
        RECT 13.040 77.465 13.180 77.620 ;
        RECT 15.710 77.560 16.030 77.620 ;
        RECT 12.965 77.235 13.255 77.465 ;
        RECT 13.885 77.420 14.175 77.465 ;
        RECT 14.790 77.420 15.110 77.480 ;
        RECT 16.720 77.465 16.860 77.960 ;
        RECT 18.025 77.960 23.300 78.100 ;
        RECT 18.025 77.915 18.315 77.960 ;
        RECT 23.160 77.805 23.300 77.960 ;
        RECT 27.670 77.960 62.170 78.100 ;
        RECT 27.670 77.900 27.990 77.960 ;
        RECT 23.085 77.575 23.375 77.805 ;
        RECT 30.430 77.760 30.750 77.820 ;
        RECT 31.365 77.760 31.655 77.805 ;
        RECT 30.430 77.620 31.655 77.760 ;
        RECT 30.430 77.560 30.750 77.620 ;
        RECT 31.365 77.575 31.655 77.620 ;
        RECT 13.885 77.280 15.110 77.420 ;
        RECT 13.885 77.235 14.175 77.280 ;
        RECT 13.040 77.080 13.180 77.235 ;
        RECT 14.790 77.220 15.110 77.280 ;
        RECT 15.265 77.235 15.555 77.465 ;
        RECT 16.645 77.235 16.935 77.465 ;
        RECT 19.850 77.420 20.170 77.480 ;
        RECT 22.165 77.420 22.455 77.465 ;
        RECT 19.850 77.280 22.455 77.420 ;
        RECT 31.440 77.420 31.580 77.575 ;
        RECT 32.270 77.560 32.590 77.820 ;
        RECT 38.250 77.760 38.570 77.820 ;
        RECT 39.645 77.760 39.935 77.805 ;
        RECT 38.250 77.620 39.935 77.760 ;
        RECT 38.250 77.560 38.570 77.620 ;
        RECT 39.645 77.575 39.935 77.620 ;
        RECT 40.550 77.560 40.870 77.820 ;
        RECT 49.765 77.760 50.055 77.805 ;
        RECT 50.670 77.760 50.990 77.820 ;
        RECT 49.765 77.620 50.990 77.760 ;
        RECT 62.030 77.760 62.170 77.960 ;
        RECT 65.850 77.960 69.390 78.100 ;
        RECT 65.850 77.900 66.170 77.960 ;
        RECT 69.070 77.900 69.390 77.960 ;
        RECT 74.170 78.100 74.460 78.145 ;
        RECT 76.270 78.100 76.560 78.145 ;
        RECT 77.840 78.100 78.130 78.145 ;
        RECT 74.170 77.960 78.130 78.100 ;
        RECT 74.170 77.915 74.460 77.960 ;
        RECT 76.270 77.915 76.560 77.960 ;
        RECT 77.840 77.915 78.130 77.960 ;
        RECT 72.750 77.760 73.070 77.820 ;
        RECT 73.685 77.760 73.975 77.805 ;
        RECT 62.030 77.620 72.060 77.760 ;
        RECT 49.765 77.575 50.055 77.620 ;
        RECT 50.670 77.560 50.990 77.620 ;
        RECT 34.110 77.420 34.430 77.480 ;
        RECT 31.440 77.280 34.430 77.420 ;
        RECT 10.280 76.940 13.180 77.080 ;
        RECT 13.410 76.880 13.730 77.140 ;
        RECT 9.285 76.740 9.575 76.785 ;
        RECT 10.650 76.740 10.970 76.800 ;
        RECT 9.285 76.600 10.970 76.740 ;
        RECT 9.285 76.555 9.575 76.600 ;
        RECT 10.650 76.540 10.970 76.600 ;
        RECT 12.950 76.740 13.270 76.800 ;
        RECT 15.340 76.740 15.480 77.235 ;
        RECT 15.710 77.080 16.030 77.140 ;
        RECT 16.720 77.080 16.860 77.235 ;
        RECT 19.850 77.220 20.170 77.280 ;
        RECT 22.165 77.235 22.455 77.280 ;
        RECT 34.110 77.220 34.430 77.280 ;
        RECT 49.305 77.420 49.595 77.465 ;
        RECT 50.210 77.420 50.530 77.480 ;
        RECT 56.665 77.420 56.955 77.465 ;
        RECT 49.305 77.280 56.955 77.420 ;
        RECT 49.305 77.235 49.595 77.280 ;
        RECT 50.210 77.220 50.530 77.280 ;
        RECT 56.665 77.235 56.955 77.280 ;
        RECT 59.885 77.420 60.175 77.465 ;
        RECT 63.090 77.420 63.410 77.480 ;
        RECT 59.885 77.280 63.410 77.420 ;
        RECT 59.885 77.235 60.175 77.280 ;
        RECT 63.090 77.220 63.410 77.280 ;
        RECT 65.850 77.220 66.170 77.480 ;
        RECT 66.785 77.235 67.075 77.465 ;
        RECT 67.245 77.235 67.535 77.465 ;
        RECT 15.710 76.940 16.860 77.080 ;
        RECT 44.230 77.080 44.550 77.140 ;
        RECT 46.545 77.080 46.835 77.125 ;
        RECT 44.230 76.940 46.835 77.080 ;
        RECT 15.710 76.880 16.030 76.940 ;
        RECT 44.230 76.880 44.550 76.940 ;
        RECT 46.545 76.895 46.835 76.940 ;
        RECT 58.490 77.080 58.810 77.140 ;
        RECT 61.250 77.125 61.570 77.140 ;
        RECT 60.345 77.080 60.635 77.125 ;
        RECT 58.490 76.940 60.635 77.080 ;
        RECT 58.490 76.880 58.810 76.940 ;
        RECT 60.345 76.895 60.635 76.940 ;
        RECT 61.250 76.895 61.635 77.125 ;
        RECT 61.250 76.880 61.570 76.895 ;
        RECT 12.950 76.600 15.480 76.740 ;
        RECT 20.325 76.740 20.615 76.785 ;
        RECT 21.230 76.740 21.550 76.800 ;
        RECT 20.325 76.600 21.550 76.740 ;
        RECT 12.950 76.540 13.270 76.600 ;
        RECT 20.325 76.555 20.615 76.600 ;
        RECT 21.230 76.540 21.550 76.600 ;
        RECT 22.625 76.740 22.915 76.785 ;
        RECT 27.670 76.740 27.990 76.800 ;
        RECT 22.625 76.600 27.990 76.740 ;
        RECT 22.625 76.555 22.915 76.600 ;
        RECT 27.670 76.540 27.990 76.600 ;
        RECT 32.745 76.740 33.035 76.785 ;
        RECT 35.030 76.740 35.350 76.800 ;
        RECT 32.745 76.600 35.350 76.740 ;
        RECT 32.745 76.555 33.035 76.600 ;
        RECT 35.030 76.540 35.350 76.600 ;
        RECT 36.870 76.540 37.190 76.800 ;
        RECT 43.770 76.540 44.090 76.800 ;
        RECT 45.545 76.740 45.835 76.785 ;
        RECT 47.450 76.740 47.770 76.800 ;
        RECT 45.545 76.600 47.770 76.740 ;
        RECT 45.545 76.555 45.835 76.600 ;
        RECT 47.450 76.540 47.770 76.600 ;
        RECT 48.845 76.740 49.135 76.785 ;
        RECT 51.590 76.740 51.910 76.800 ;
        RECT 48.845 76.600 51.910 76.740 ;
        RECT 48.845 76.555 49.135 76.600 ;
        RECT 51.590 76.540 51.910 76.600 ;
        RECT 62.170 76.740 62.490 76.800 ;
        RECT 66.860 76.740 67.000 77.235 ;
        RECT 67.320 77.080 67.460 77.235 ;
        RECT 67.690 77.220 68.010 77.480 ;
        RECT 68.150 77.420 68.470 77.480 ;
        RECT 68.625 77.420 68.915 77.465 ;
        RECT 68.150 77.280 68.915 77.420 ;
        RECT 68.150 77.220 68.470 77.280 ;
        RECT 68.625 77.235 68.915 77.280 ;
        RECT 70.450 77.220 70.770 77.480 ;
        RECT 70.910 77.420 71.230 77.480 ;
        RECT 71.920 77.465 72.060 77.620 ;
        RECT 72.750 77.620 73.975 77.760 ;
        RECT 72.750 77.560 73.070 77.620 ;
        RECT 73.685 77.575 73.975 77.620 ;
        RECT 74.565 77.760 74.855 77.805 ;
        RECT 75.755 77.760 76.045 77.805 ;
        RECT 78.275 77.760 78.565 77.805 ;
        RECT 74.565 77.620 78.565 77.760 ;
        RECT 74.565 77.575 74.855 77.620 ;
        RECT 75.755 77.575 76.045 77.620 ;
        RECT 78.275 77.575 78.565 77.620 ;
        RECT 71.385 77.420 71.675 77.465 ;
        RECT 70.910 77.280 71.675 77.420 ;
        RECT 70.910 77.220 71.230 77.280 ;
        RECT 71.385 77.235 71.675 77.280 ;
        RECT 71.845 77.235 72.135 77.465 ;
        RECT 72.290 77.220 72.610 77.480 ;
        RECT 78.730 77.420 79.050 77.480 ;
        RECT 81.045 77.420 81.335 77.465 ;
        RECT 78.730 77.280 81.335 77.420 ;
        RECT 78.730 77.220 79.050 77.280 ;
        RECT 81.045 77.235 81.335 77.280 ;
        RECT 73.670 77.080 73.990 77.140 ;
        RECT 67.320 76.940 73.990 77.080 ;
        RECT 71.460 76.800 71.600 76.940 ;
        RECT 73.670 76.880 73.990 76.940 ;
        RECT 75.020 77.080 75.310 77.125 ;
        RECT 75.510 77.080 75.830 77.140 ;
        RECT 75.020 76.940 75.830 77.080 ;
        RECT 75.020 76.895 75.310 76.940 ;
        RECT 75.510 76.880 75.830 76.940 ;
        RECT 62.170 76.600 67.000 76.740 ;
        RECT 62.170 76.540 62.490 76.600 ;
        RECT 71.370 76.540 71.690 76.800 ;
        RECT 73.225 76.740 73.515 76.785 ;
        RECT 77.810 76.740 78.130 76.800 ;
        RECT 73.225 76.600 78.130 76.740 ;
        RECT 73.225 76.555 73.515 76.600 ;
        RECT 77.810 76.540 78.130 76.600 ;
        RECT 5.520 75.920 84.180 76.400 ;
        RECT 14.790 75.520 15.110 75.780 ;
        RECT 27.670 75.520 27.990 75.780 ;
        RECT 38.250 75.720 38.570 75.780 ;
        RECT 38.725 75.720 39.015 75.765 ;
        RECT 38.250 75.580 39.015 75.720 ;
        RECT 38.250 75.520 38.570 75.580 ;
        RECT 38.725 75.535 39.015 75.580 ;
        RECT 39.645 75.720 39.935 75.765 ;
        RECT 40.550 75.720 40.870 75.780 ;
        RECT 39.645 75.580 40.870 75.720 ;
        RECT 39.645 75.535 39.935 75.580 ;
        RECT 40.550 75.520 40.870 75.580 ;
        RECT 49.765 75.720 50.055 75.765 ;
        RECT 50.210 75.720 50.530 75.780 ;
        RECT 62.630 75.720 62.950 75.780 ;
        RECT 65.390 75.720 65.710 75.780 ;
        RECT 70.005 75.720 70.295 75.765 ;
        RECT 70.450 75.720 70.770 75.780 ;
        RECT 49.765 75.580 50.530 75.720 ;
        RECT 49.765 75.535 50.055 75.580 ;
        RECT 50.210 75.520 50.530 75.580 ;
        RECT 58.580 75.580 67.920 75.720 ;
        RECT 13.870 75.380 14.190 75.440 ;
        RECT 7.980 75.240 14.190 75.380 ;
        RECT 14.880 75.380 15.020 75.520 ;
        RECT 34.570 75.380 34.890 75.440 ;
        RECT 14.880 75.240 18.700 75.380 ;
        RECT 7.980 75.085 8.120 75.240 ;
        RECT 13.870 75.180 14.190 75.240 ;
        RECT 9.270 75.085 9.590 75.100 ;
        RECT 7.905 74.855 8.195 75.085 ;
        RECT 9.240 74.855 9.590 75.085 ;
        RECT 9.270 74.840 9.590 74.855 ;
        RECT 15.710 75.040 16.030 75.100 ;
        RECT 18.560 75.085 18.700 75.240 ;
        RECT 20.860 75.240 34.890 75.380 ;
        RECT 20.860 75.085 21.000 75.240 ;
        RECT 17.105 75.040 17.395 75.085 ;
        RECT 15.710 74.900 17.395 75.040 ;
        RECT 15.710 74.840 16.030 74.900 ;
        RECT 17.105 74.855 17.395 74.900 ;
        RECT 18.485 74.855 18.775 75.085 ;
        RECT 20.785 74.855 21.075 75.085 ;
        RECT 21.230 75.040 21.550 75.100 ;
        RECT 31.900 75.085 32.040 75.240 ;
        RECT 34.570 75.180 34.890 75.240 ;
        RECT 44.230 75.380 44.550 75.440 ;
        RECT 47.910 75.380 48.230 75.440 ;
        RECT 44.230 75.240 48.230 75.380 ;
        RECT 44.230 75.180 44.550 75.240 ;
        RECT 47.910 75.180 48.230 75.240 ;
        RECT 55.440 75.380 55.730 75.425 ;
        RECT 57.585 75.380 57.875 75.425 ;
        RECT 55.440 75.240 57.875 75.380 ;
        RECT 55.440 75.195 55.730 75.240 ;
        RECT 57.585 75.195 57.875 75.240 ;
        RECT 33.190 75.085 33.510 75.100 ;
        RECT 22.065 75.040 22.355 75.085 ;
        RECT 21.230 74.900 22.355 75.040 ;
        RECT 21.230 74.840 21.550 74.900 ;
        RECT 22.065 74.855 22.355 74.900 ;
        RECT 31.825 74.855 32.115 75.085 ;
        RECT 33.160 74.855 33.510 75.085 ;
        RECT 33.190 74.840 33.510 74.855 ;
        RECT 45.150 75.085 45.470 75.100 ;
        RECT 45.150 74.855 45.500 75.085 ;
        RECT 56.190 75.040 56.510 75.100 ;
        RECT 58.580 75.085 58.720 75.580 ;
        RECT 62.630 75.520 62.950 75.580 ;
        RECT 65.390 75.520 65.710 75.580 ;
        RECT 62.170 75.380 62.490 75.440 ;
        RECT 65.850 75.380 66.170 75.440 ;
        RECT 67.245 75.380 67.535 75.425 ;
        RECT 61.800 75.240 62.490 75.380 ;
        RECT 56.665 75.040 56.955 75.085 ;
        RECT 56.190 74.900 56.955 75.040 ;
        RECT 45.150 74.840 45.470 74.855 ;
        RECT 56.190 74.840 56.510 74.900 ;
        RECT 56.665 74.855 56.955 74.900 ;
        RECT 58.505 74.855 58.795 75.085 ;
        RECT 58.965 75.040 59.255 75.085 ;
        RECT 59.410 75.040 59.730 75.100 ;
        RECT 61.800 75.085 61.940 75.240 ;
        RECT 62.170 75.180 62.490 75.240 ;
        RECT 62.720 75.240 67.535 75.380 ;
        RECT 67.780 75.380 67.920 75.580 ;
        RECT 70.005 75.580 70.770 75.720 ;
        RECT 70.005 75.535 70.295 75.580 ;
        RECT 70.450 75.520 70.770 75.580 ;
        RECT 75.510 75.520 75.830 75.780 ;
        RECT 77.365 75.720 77.655 75.765 ;
        RECT 79.190 75.720 79.510 75.780 ;
        RECT 77.365 75.580 79.510 75.720 ;
        RECT 77.365 75.535 77.655 75.580 ;
        RECT 79.190 75.520 79.510 75.580 ;
        RECT 68.165 75.380 68.455 75.425 ;
        RECT 67.780 75.240 68.455 75.380 ;
        RECT 58.965 74.900 59.730 75.040 ;
        RECT 58.965 74.855 59.255 74.900 ;
        RECT 59.410 74.840 59.730 74.900 ;
        RECT 59.885 74.855 60.175 75.085 ;
        RECT 61.725 74.855 62.015 75.085 ;
        RECT 62.720 75.040 62.860 75.240 ;
        RECT 65.850 75.180 66.170 75.240 ;
        RECT 67.245 75.195 67.535 75.240 ;
        RECT 68.165 75.195 68.455 75.240 ;
        RECT 77.810 75.180 78.130 75.440 ;
        RECT 62.260 74.900 62.860 75.040 ;
        RECT 8.785 74.700 9.075 74.745 ;
        RECT 9.975 74.700 10.265 74.745 ;
        RECT 12.495 74.700 12.785 74.745 ;
        RECT 8.785 74.560 12.785 74.700 ;
        RECT 8.785 74.515 9.075 74.560 ;
        RECT 9.975 74.515 10.265 74.560 ;
        RECT 12.495 74.515 12.785 74.560 ;
        RECT 21.665 74.700 21.955 74.745 ;
        RECT 22.855 74.700 23.145 74.745 ;
        RECT 25.375 74.700 25.665 74.745 ;
        RECT 21.665 74.560 25.665 74.700 ;
        RECT 21.665 74.515 21.955 74.560 ;
        RECT 22.855 74.515 23.145 74.560 ;
        RECT 25.375 74.515 25.665 74.560 ;
        RECT 32.705 74.700 32.995 74.745 ;
        RECT 33.895 74.700 34.185 74.745 ;
        RECT 36.415 74.700 36.705 74.745 ;
        RECT 32.705 74.560 36.705 74.700 ;
        RECT 32.705 74.515 32.995 74.560 ;
        RECT 33.895 74.515 34.185 74.560 ;
        RECT 36.415 74.515 36.705 74.560 ;
        RECT 41.955 74.700 42.245 74.745 ;
        RECT 44.475 74.700 44.765 74.745 ;
        RECT 45.665 74.700 45.955 74.745 ;
        RECT 41.955 74.560 45.955 74.700 ;
        RECT 41.955 74.515 42.245 74.560 ;
        RECT 44.475 74.515 44.765 74.560 ;
        RECT 45.665 74.515 45.955 74.560 ;
        RECT 46.545 74.515 46.835 74.745 ;
        RECT 52.075 74.700 52.365 74.745 ;
        RECT 54.595 74.700 54.885 74.745 ;
        RECT 55.785 74.700 56.075 74.745 ;
        RECT 52.075 74.560 56.075 74.700 ;
        RECT 59.960 74.700 60.100 74.855 ;
        RECT 62.260 74.745 62.400 74.900 ;
        RECT 63.090 74.840 63.410 75.100 ;
        RECT 64.010 75.040 64.330 75.100 ;
        RECT 64.945 75.040 65.235 75.085 ;
        RECT 64.010 74.900 65.235 75.040 ;
        RECT 64.010 74.840 64.330 74.900 ;
        RECT 64.945 74.855 65.235 74.900 ;
        RECT 60.805 74.700 61.095 74.745 ;
        RECT 59.960 74.560 61.095 74.700 ;
        RECT 52.075 74.515 52.365 74.560 ;
        RECT 54.595 74.515 54.885 74.560 ;
        RECT 55.785 74.515 56.075 74.560 ;
        RECT 60.805 74.515 61.095 74.560 ;
        RECT 62.185 74.515 62.475 74.745 ;
        RECT 62.630 74.700 62.950 74.760 ;
        RECT 63.550 74.700 63.870 74.760 ;
        RECT 62.630 74.560 63.870 74.700 ;
        RECT 65.020 74.700 65.160 74.855 ;
        RECT 66.310 74.840 66.630 75.100 ;
        RECT 67.705 74.855 67.995 75.085 ;
        RECT 69.085 75.040 69.375 75.085 ;
        RECT 70.450 75.040 70.770 75.100 ;
        RECT 69.085 74.900 70.770 75.040 ;
        RECT 69.085 74.855 69.375 74.900 ;
        RECT 67.780 74.700 67.920 74.855 ;
        RECT 70.450 74.840 70.770 74.900 ;
        RECT 79.665 75.040 79.955 75.085 ;
        RECT 80.570 75.040 80.890 75.100 ;
        RECT 79.665 74.900 80.890 75.040 ;
        RECT 79.665 74.855 79.955 74.900 ;
        RECT 80.570 74.840 80.890 74.900 ;
        RECT 71.830 74.700 72.150 74.760 ;
        RECT 65.020 74.560 72.150 74.700 ;
        RECT 8.390 74.360 8.680 74.405 ;
        RECT 10.490 74.360 10.780 74.405 ;
        RECT 12.060 74.360 12.350 74.405 ;
        RECT 8.390 74.220 12.350 74.360 ;
        RECT 8.390 74.175 8.680 74.220 ;
        RECT 10.490 74.175 10.780 74.220 ;
        RECT 12.060 74.175 12.350 74.220 ;
        RECT 17.090 74.360 17.410 74.420 ;
        RECT 19.865 74.360 20.155 74.405 ;
        RECT 17.090 74.220 20.155 74.360 ;
        RECT 17.090 74.160 17.410 74.220 ;
        RECT 19.865 74.175 20.155 74.220 ;
        RECT 21.270 74.360 21.560 74.405 ;
        RECT 23.370 74.360 23.660 74.405 ;
        RECT 24.940 74.360 25.230 74.405 ;
        RECT 21.270 74.220 25.230 74.360 ;
        RECT 21.270 74.175 21.560 74.220 ;
        RECT 23.370 74.175 23.660 74.220 ;
        RECT 24.940 74.175 25.230 74.220 ;
        RECT 32.310 74.360 32.600 74.405 ;
        RECT 34.410 74.360 34.700 74.405 ;
        RECT 35.980 74.360 36.270 74.405 ;
        RECT 32.310 74.220 36.270 74.360 ;
        RECT 32.310 74.175 32.600 74.220 ;
        RECT 34.410 74.175 34.700 74.220 ;
        RECT 35.980 74.175 36.270 74.220 ;
        RECT 42.390 74.360 42.680 74.405 ;
        RECT 43.960 74.360 44.250 74.405 ;
        RECT 46.060 74.360 46.350 74.405 ;
        RECT 42.390 74.220 46.350 74.360 ;
        RECT 42.390 74.175 42.680 74.220 ;
        RECT 43.960 74.175 44.250 74.220 ;
        RECT 46.060 74.175 46.350 74.220 ;
        RECT 17.550 73.820 17.870 74.080 ;
        RECT 44.690 74.020 45.010 74.080 ;
        RECT 46.620 74.020 46.760 74.515 ;
        RECT 62.630 74.500 62.950 74.560 ;
        RECT 63.550 74.500 63.870 74.560 ;
        RECT 71.830 74.500 72.150 74.560 ;
        RECT 78.270 74.500 78.590 74.760 ;
        RECT 52.510 74.360 52.800 74.405 ;
        RECT 54.080 74.360 54.370 74.405 ;
        RECT 56.180 74.360 56.470 74.405 ;
        RECT 52.510 74.220 56.470 74.360 ;
        RECT 52.510 74.175 52.800 74.220 ;
        RECT 54.080 74.175 54.370 74.220 ;
        RECT 56.180 74.175 56.470 74.220 ;
        RECT 59.410 74.160 59.730 74.420 ;
        RECT 66.310 74.360 66.630 74.420 ;
        RECT 67.690 74.360 68.010 74.420 ;
        RECT 66.310 74.220 68.010 74.360 ;
        RECT 66.310 74.160 66.630 74.220 ;
        RECT 67.690 74.160 68.010 74.220 ;
        RECT 44.690 73.880 46.760 74.020 ;
        RECT 80.585 74.020 80.875 74.065 ;
        RECT 81.030 74.020 81.350 74.080 ;
        RECT 80.585 73.880 81.350 74.020 ;
        RECT 44.690 73.820 45.010 73.880 ;
        RECT 80.585 73.835 80.875 73.880 ;
        RECT 81.030 73.820 81.350 73.880 ;
        RECT 5.520 73.200 84.180 73.680 ;
        RECT 8.825 73.000 9.115 73.045 ;
        RECT 9.270 73.000 9.590 73.060 ;
        RECT 8.825 72.860 9.590 73.000 ;
        RECT 8.825 72.815 9.115 72.860 ;
        RECT 9.270 72.800 9.590 72.860 ;
        RECT 13.425 73.000 13.715 73.045 ;
        RECT 14.790 73.000 15.110 73.060 ;
        RECT 13.425 72.860 15.110 73.000 ;
        RECT 13.425 72.815 13.715 72.860 ;
        RECT 14.790 72.800 15.110 72.860 ;
        RECT 15.710 72.800 16.030 73.060 ;
        RECT 33.190 73.000 33.510 73.060 ;
        RECT 34.585 73.000 34.875 73.045 ;
        RECT 44.230 73.000 44.550 73.060 ;
        RECT 33.190 72.860 34.875 73.000 ;
        RECT 33.190 72.800 33.510 72.860 ;
        RECT 34.585 72.815 34.875 72.860 ;
        RECT 37.420 72.860 44.550 73.000 ;
        RECT 11.585 72.660 11.875 72.705 ;
        RECT 15.800 72.660 15.940 72.800 ;
        RECT 11.585 72.520 15.940 72.660 ;
        RECT 21.730 72.660 22.020 72.705 ;
        RECT 23.830 72.660 24.120 72.705 ;
        RECT 25.400 72.660 25.690 72.705 ;
        RECT 21.730 72.520 25.690 72.660 ;
        RECT 11.585 72.475 11.875 72.520 ;
        RECT 21.730 72.475 22.020 72.520 ;
        RECT 23.830 72.475 24.120 72.520 ;
        RECT 25.400 72.475 25.690 72.520 ;
        RECT 34.110 72.660 34.430 72.720 ;
        RECT 37.420 72.660 37.560 72.860 ;
        RECT 44.230 72.800 44.550 72.860 ;
        RECT 44.705 73.000 44.995 73.045 ;
        RECT 45.150 73.000 45.470 73.060 ;
        RECT 44.705 72.860 45.470 73.000 ;
        RECT 44.705 72.815 44.995 72.860 ;
        RECT 45.150 72.800 45.470 72.860 ;
        RECT 49.305 73.000 49.595 73.045 ;
        RECT 64.930 73.000 65.250 73.060 ;
        RECT 65.405 73.000 65.695 73.045 ;
        RECT 68.610 73.000 68.930 73.060 ;
        RECT 49.305 72.860 56.880 73.000 ;
        RECT 49.305 72.815 49.595 72.860 ;
        RECT 49.380 72.660 49.520 72.815 ;
        RECT 34.110 72.520 37.560 72.660 ;
        RECT 34.110 72.460 34.430 72.520 ;
        RECT 10.190 72.320 10.510 72.380 ;
        RECT 13.410 72.320 13.730 72.380 ;
        RECT 9.820 72.180 13.730 72.320 ;
        RECT 9.820 72.025 9.960 72.180 ;
        RECT 10.190 72.120 10.510 72.180 ;
        RECT 13.410 72.120 13.730 72.180 ;
        RECT 22.125 72.320 22.415 72.365 ;
        RECT 23.315 72.320 23.605 72.365 ;
        RECT 25.835 72.320 26.125 72.365 ;
        RECT 22.125 72.180 26.125 72.320 ;
        RECT 22.125 72.135 22.415 72.180 ;
        RECT 23.315 72.135 23.605 72.180 ;
        RECT 25.835 72.135 26.125 72.180 ;
        RECT 36.870 72.120 37.190 72.380 ;
        RECT 37.420 72.365 37.560 72.520 ;
        RECT 41.100 72.520 49.520 72.660 ;
        RECT 52.050 72.660 52.340 72.705 ;
        RECT 53.620 72.660 53.910 72.705 ;
        RECT 55.720 72.660 56.010 72.705 ;
        RECT 52.050 72.520 56.010 72.660 ;
        RECT 41.100 72.365 41.240 72.520 ;
        RECT 52.050 72.475 52.340 72.520 ;
        RECT 53.620 72.475 53.910 72.520 ;
        RECT 55.720 72.475 56.010 72.520 ;
        RECT 37.345 72.135 37.635 72.365 ;
        RECT 41.025 72.135 41.315 72.365 ;
        RECT 41.485 72.135 41.775 72.365 ;
        RECT 43.770 72.320 44.090 72.380 ;
        RECT 47.005 72.320 47.295 72.365 ;
        RECT 43.770 72.180 47.295 72.320 ;
        RECT 9.745 71.795 10.035 72.025 ;
        RECT 10.650 71.780 10.970 72.040 ;
        RECT 14.790 71.980 15.110 72.040 ;
        RECT 15.265 71.980 15.555 72.025 ;
        RECT 14.790 71.840 15.555 71.980 ;
        RECT 14.790 71.780 15.110 71.840 ;
        RECT 15.265 71.795 15.555 71.840 ;
        RECT 17.105 71.980 17.395 72.025 ;
        RECT 17.550 71.980 17.870 72.040 ;
        RECT 17.105 71.840 17.870 71.980 ;
        RECT 17.105 71.795 17.395 71.840 ;
        RECT 17.550 71.780 17.870 71.840 ;
        RECT 21.245 71.980 21.535 72.025 ;
        RECT 33.665 71.980 33.955 72.025 ;
        RECT 34.570 71.980 34.890 72.040 ;
        RECT 21.245 71.840 34.890 71.980 ;
        RECT 21.245 71.795 21.535 71.840 ;
        RECT 33.665 71.795 33.955 71.840 ;
        RECT 34.570 71.780 34.890 71.840 ;
        RECT 39.630 71.980 39.950 72.040 ;
        RECT 41.560 71.980 41.700 72.135 ;
        RECT 43.770 72.120 44.090 72.180 ;
        RECT 47.005 72.135 47.295 72.180 ;
        RECT 47.910 72.120 48.230 72.380 ;
        RECT 56.740 72.365 56.880 72.860 ;
        RECT 64.930 72.860 68.930 73.000 ;
        RECT 64.930 72.800 65.250 72.860 ;
        RECT 65.405 72.815 65.695 72.860 ;
        RECT 68.610 72.800 68.930 72.860 ;
        RECT 80.570 72.800 80.890 73.060 ;
        RECT 59.410 72.660 59.730 72.720 ;
        RECT 74.170 72.660 74.460 72.705 ;
        RECT 76.270 72.660 76.560 72.705 ;
        RECT 77.840 72.660 78.130 72.705 ;
        RECT 59.410 72.520 63.320 72.660 ;
        RECT 59.410 72.460 59.730 72.520 ;
        RECT 51.615 72.320 51.905 72.365 ;
        RECT 54.135 72.320 54.425 72.365 ;
        RECT 55.325 72.320 55.615 72.365 ;
        RECT 51.615 72.180 55.615 72.320 ;
        RECT 51.615 72.135 51.905 72.180 ;
        RECT 54.135 72.135 54.425 72.180 ;
        RECT 55.325 72.135 55.615 72.180 ;
        RECT 56.665 72.135 56.955 72.365 ;
        RECT 59.885 72.320 60.175 72.365 ;
        RECT 59.885 72.180 61.940 72.320 ;
        RECT 59.885 72.135 60.175 72.180 ;
        RECT 39.630 71.840 41.700 71.980 ;
        RECT 44.690 71.980 45.010 72.040 ;
        RECT 49.290 71.980 49.610 72.040 ;
        RECT 56.190 71.980 56.510 72.040 ;
        RECT 44.690 71.840 56.510 71.980 ;
        RECT 39.630 71.780 39.950 71.840 ;
        RECT 44.690 71.780 45.010 71.840 ;
        RECT 49.290 71.780 49.610 71.840 ;
        RECT 56.190 71.780 56.510 71.840 ;
        RECT 58.030 71.980 58.350 72.040 ;
        RECT 61.250 71.980 61.570 72.040 ;
        RECT 61.800 72.025 61.940 72.180 ;
        RECT 62.630 72.120 62.950 72.380 ;
        RECT 63.180 72.025 63.320 72.520 ;
        RECT 74.170 72.520 78.130 72.660 ;
        RECT 74.170 72.475 74.460 72.520 ;
        RECT 76.270 72.475 76.560 72.520 ;
        RECT 77.840 72.475 78.130 72.520 ;
        RECT 63.550 72.320 63.870 72.380 ;
        RECT 65.390 72.320 65.710 72.380 ;
        RECT 63.550 72.180 65.710 72.320 ;
        RECT 63.550 72.120 63.870 72.180 ;
        RECT 65.390 72.120 65.710 72.180 ;
        RECT 69.070 72.320 69.390 72.380 ;
        RECT 70.910 72.320 71.230 72.380 ;
        RECT 69.070 72.180 71.230 72.320 ;
        RECT 69.070 72.120 69.390 72.180 ;
        RECT 70.910 72.120 71.230 72.180 ;
        RECT 72.750 72.320 73.070 72.380 ;
        RECT 73.670 72.320 73.990 72.380 ;
        RECT 72.750 72.180 73.990 72.320 ;
        RECT 72.750 72.120 73.070 72.180 ;
        RECT 73.670 72.120 73.990 72.180 ;
        RECT 74.565 72.320 74.855 72.365 ;
        RECT 75.755 72.320 76.045 72.365 ;
        RECT 78.275 72.320 78.565 72.365 ;
        RECT 74.565 72.180 78.565 72.320 ;
        RECT 74.565 72.135 74.855 72.180 ;
        RECT 75.755 72.135 76.045 72.180 ;
        RECT 78.275 72.135 78.565 72.180 ;
        RECT 58.030 71.840 61.570 71.980 ;
        RECT 58.030 71.780 58.350 71.840 ;
        RECT 61.250 71.780 61.570 71.840 ;
        RECT 61.725 71.795 62.015 72.025 ;
        RECT 63.105 71.795 63.395 72.025 ;
        RECT 64.470 71.780 64.790 72.040 ;
        RECT 65.480 71.980 65.620 72.120 ;
        RECT 65.865 71.980 66.155 72.025 ;
        RECT 65.480 71.840 66.155 71.980 ;
        RECT 65.865 71.795 66.155 71.840 ;
        RECT 66.770 71.780 67.090 72.040 ;
        RECT 67.230 71.980 67.550 72.040 ;
        RECT 67.705 71.980 67.995 72.025 ;
        RECT 80.110 71.980 80.430 72.040 ;
        RECT 67.230 71.840 80.430 71.980 ;
        RECT 67.230 71.780 67.550 71.840 ;
        RECT 67.705 71.795 67.995 71.840 ;
        RECT 80.110 71.780 80.430 71.840 ;
        RECT 81.030 71.780 81.350 72.040 ;
        RECT 12.950 71.640 13.270 71.700 ;
        RECT 13.425 71.640 13.715 71.685 ;
        RECT 12.950 71.500 13.715 71.640 ;
        RECT 12.950 71.440 13.270 71.500 ;
        RECT 13.425 71.455 13.715 71.500 ;
        RECT 20.310 71.640 20.630 71.700 ;
        RECT 22.470 71.640 22.760 71.685 ;
        RECT 29.970 71.640 30.290 71.700 ;
        RECT 54.980 71.640 55.270 71.685 ;
        RECT 60.345 71.640 60.635 71.685 ;
        RECT 20.310 71.500 22.760 71.640 ;
        RECT 20.310 71.440 20.630 71.500 ;
        RECT 22.470 71.455 22.760 71.500 ;
        RECT 28.220 71.500 48.370 71.640 ;
        RECT 14.330 71.100 14.650 71.360 ;
        RECT 18.010 71.100 18.330 71.360 ;
        RECT 28.220 71.345 28.360 71.500 ;
        RECT 29.970 71.440 30.290 71.500 ;
        RECT 28.145 71.115 28.435 71.345 ;
        RECT 36.425 71.300 36.715 71.345 ;
        RECT 38.725 71.300 39.015 71.345 ;
        RECT 36.425 71.160 39.015 71.300 ;
        RECT 36.425 71.115 36.715 71.160 ;
        RECT 38.725 71.115 39.015 71.160 ;
        RECT 40.550 71.100 40.870 71.360 ;
        RECT 46.530 71.100 46.850 71.360 ;
        RECT 48.230 71.300 48.370 71.500 ;
        RECT 54.980 71.500 60.635 71.640 ;
        RECT 54.980 71.455 55.270 71.500 ;
        RECT 60.345 71.455 60.635 71.500 ;
        RECT 62.630 71.640 62.950 71.700 ;
        RECT 65.390 71.640 65.710 71.700 ;
        RECT 73.210 71.640 73.530 71.700 ;
        RECT 75.050 71.685 75.370 71.700 ;
        RECT 62.630 71.500 65.710 71.640 ;
        RECT 62.630 71.440 62.950 71.500 ;
        RECT 65.390 71.440 65.710 71.500 ;
        RECT 66.400 71.500 73.530 71.640 ;
        RECT 66.400 71.360 66.540 71.500 ;
        RECT 73.210 71.440 73.530 71.500 ;
        RECT 75.020 71.455 75.370 71.685 ;
        RECT 75.050 71.440 75.370 71.455 ;
        RECT 65.850 71.300 66.170 71.360 ;
        RECT 48.230 71.160 66.170 71.300 ;
        RECT 65.850 71.100 66.170 71.160 ;
        RECT 66.310 71.100 66.630 71.360 ;
        RECT 67.690 71.300 68.010 71.360 ;
        RECT 68.625 71.300 68.915 71.345 ;
        RECT 74.130 71.300 74.450 71.360 ;
        RECT 67.690 71.160 74.450 71.300 ;
        RECT 67.690 71.100 68.010 71.160 ;
        RECT 68.625 71.115 68.915 71.160 ;
        RECT 74.130 71.100 74.450 71.160 ;
        RECT 81.950 71.100 82.270 71.360 ;
        RECT 5.520 70.480 84.180 70.960 ;
        RECT 9.745 70.280 10.035 70.325 ;
        RECT 14.790 70.280 15.110 70.340 ;
        RECT 18.485 70.280 18.775 70.325 ;
        RECT 19.850 70.280 20.170 70.340 ;
        RECT 9.745 70.140 20.170 70.280 ;
        RECT 9.745 70.095 10.035 70.140 ;
        RECT 14.790 70.080 15.110 70.140 ;
        RECT 18.485 70.095 18.775 70.140 ;
        RECT 19.850 70.080 20.170 70.140 ;
        RECT 20.310 70.080 20.630 70.340 ;
        RECT 51.130 70.280 51.450 70.340 ;
        RECT 32.820 70.140 51.450 70.280 ;
        RECT 13.870 69.940 14.190 70.000 ;
        RECT 18.930 69.940 19.250 70.000 ;
        RECT 24.465 69.940 24.755 69.985 ;
        RECT 13.870 69.800 24.755 69.940 ;
        RECT 13.870 69.740 14.190 69.800 ;
        RECT 18.930 69.740 19.250 69.800 ;
        RECT 24.465 69.755 24.755 69.800 ;
        RECT 31.810 69.940 32.130 70.000 ;
        RECT 32.820 69.985 32.960 70.140 ;
        RECT 51.130 70.080 51.450 70.140 ;
        RECT 59.410 70.280 59.730 70.340 ;
        RECT 60.805 70.280 61.095 70.325 ;
        RECT 59.410 70.140 61.095 70.280 ;
        RECT 59.410 70.080 59.730 70.140 ;
        RECT 60.805 70.095 61.095 70.140 ;
        RECT 62.170 70.080 62.490 70.340 ;
        RECT 62.630 70.080 62.950 70.340 ;
        RECT 63.090 70.080 63.410 70.340 ;
        RECT 65.850 70.280 66.170 70.340 ;
        RECT 65.850 70.140 66.540 70.280 ;
        RECT 65.850 70.080 66.170 70.140 ;
        RECT 32.745 69.940 33.035 69.985 ;
        RECT 31.810 69.800 33.035 69.940 ;
        RECT 31.810 69.740 32.130 69.800 ;
        RECT 32.745 69.755 33.035 69.800 ;
        RECT 33.190 69.940 33.510 70.000 ;
        RECT 34.570 69.940 34.890 70.000 ;
        RECT 36.425 69.940 36.715 69.985 ;
        RECT 33.190 69.800 36.715 69.940 ;
        RECT 33.190 69.740 33.510 69.800 ;
        RECT 34.570 69.740 34.890 69.800 ;
        RECT 36.425 69.755 36.715 69.800 ;
        RECT 45.610 69.940 45.930 70.000 ;
        RECT 58.490 69.940 58.810 70.000 ;
        RECT 62.260 69.940 62.400 70.080 ;
        RECT 45.610 69.800 55.500 69.940 ;
        RECT 9.285 69.415 9.575 69.645 ;
        RECT 9.360 68.920 9.500 69.415 ;
        RECT 13.410 69.400 13.730 69.660 ;
        RECT 14.790 69.600 15.110 69.660 ;
        RECT 13.960 69.460 15.110 69.600 ;
        RECT 10.190 69.060 10.510 69.320 ;
        RECT 13.960 69.305 14.100 69.460 ;
        RECT 14.790 69.400 15.110 69.460 ;
        RECT 20.785 69.600 21.075 69.645 ;
        RECT 31.900 69.600 32.040 69.740 ;
        RECT 20.785 69.460 32.040 69.600 ;
        RECT 36.500 69.600 36.640 69.755 ;
        RECT 45.610 69.740 45.930 69.800 ;
        RECT 40.565 69.600 40.855 69.645 ;
        RECT 36.500 69.460 40.855 69.600 ;
        RECT 20.785 69.415 21.075 69.460 ;
        RECT 40.565 69.415 40.855 69.460 ;
        RECT 41.900 69.600 42.190 69.645 ;
        RECT 41.900 69.460 48.140 69.600 ;
        RECT 41.900 69.415 42.190 69.460 ;
        RECT 13.885 69.075 14.175 69.305 ;
        RECT 14.330 69.060 14.650 69.320 ;
        RECT 17.090 69.060 17.410 69.320 ;
        RECT 18.025 69.260 18.315 69.305 ;
        RECT 29.970 69.260 30.290 69.320 ;
        RECT 18.025 69.120 30.290 69.260 ;
        RECT 18.025 69.075 18.315 69.120 ;
        RECT 29.970 69.060 30.290 69.120 ;
        RECT 41.445 69.260 41.735 69.305 ;
        RECT 42.635 69.260 42.925 69.305 ;
        RECT 45.155 69.260 45.445 69.305 ;
        RECT 41.445 69.120 45.445 69.260 ;
        RECT 41.445 69.075 41.735 69.120 ;
        RECT 42.635 69.075 42.925 69.120 ;
        RECT 45.155 69.075 45.445 69.120 ;
        RECT 45.610 69.260 45.930 69.320 ;
        RECT 45.610 69.120 47.680 69.260 ;
        RECT 45.610 69.060 45.930 69.120 ;
        RECT 12.950 68.920 13.270 68.980 ;
        RECT 47.540 68.965 47.680 69.120 ;
        RECT 48.000 68.965 48.140 69.460 ;
        RECT 49.750 69.400 50.070 69.660 ;
        RECT 55.360 69.645 55.500 69.800 ;
        RECT 58.490 69.800 62.400 69.940 ;
        RECT 58.490 69.740 58.810 69.800 ;
        RECT 50.225 69.600 50.515 69.645 ;
        RECT 52.065 69.600 52.355 69.645 ;
        RECT 50.225 69.460 52.355 69.600 ;
        RECT 50.225 69.415 50.515 69.460 ;
        RECT 52.065 69.415 52.355 69.460 ;
        RECT 55.285 69.415 55.575 69.645 ;
        RECT 56.190 69.600 56.510 69.660 ;
        RECT 58.045 69.600 58.335 69.645 ;
        RECT 56.190 69.460 58.335 69.600 ;
        RECT 56.190 69.400 56.510 69.460 ;
        RECT 58.045 69.415 58.335 69.460 ;
        RECT 60.790 69.400 61.110 69.660 ;
        RECT 61.800 69.645 61.940 69.800 ;
        RECT 61.725 69.415 62.015 69.645 ;
        RECT 62.170 69.400 62.490 69.660 ;
        RECT 63.180 69.645 63.320 70.080 ;
        RECT 64.530 69.800 65.160 69.940 ;
        RECT 64.530 69.645 64.670 69.800 ;
        RECT 63.105 69.600 63.395 69.645 ;
        RECT 62.720 69.460 63.395 69.600 ;
        RECT 50.685 69.075 50.975 69.305 ;
        RECT 41.050 68.920 41.340 68.965 ;
        RECT 43.150 68.920 43.440 68.965 ;
        RECT 44.720 68.920 45.010 68.965 ;
        RECT 9.360 68.780 13.870 68.920 ;
        RECT 12.950 68.720 13.270 68.780 ;
        RECT 7.430 68.380 7.750 68.640 ;
        RECT 11.110 68.580 11.430 68.640 ;
        RECT 11.585 68.580 11.875 68.625 ;
        RECT 11.110 68.440 11.875 68.580 ;
        RECT 13.730 68.580 13.870 68.780 ;
        RECT 41.050 68.780 45.010 68.920 ;
        RECT 41.050 68.735 41.340 68.780 ;
        RECT 43.150 68.735 43.440 68.780 ;
        RECT 44.720 68.735 45.010 68.780 ;
        RECT 47.465 68.735 47.755 68.965 ;
        RECT 47.925 68.735 48.215 68.965 ;
        RECT 48.370 68.920 48.690 68.980 ;
        RECT 50.760 68.920 50.900 69.075 ;
        RECT 62.720 68.980 62.860 69.460 ;
        RECT 63.105 69.415 63.395 69.460 ;
        RECT 63.595 69.415 63.885 69.645 ;
        RECT 64.455 69.415 64.745 69.645 ;
        RECT 48.370 68.780 50.900 68.920 ;
        RECT 48.370 68.720 48.690 68.780 ;
        RECT 62.630 68.720 62.950 68.980 ;
        RECT 63.645 68.920 63.785 69.415 ;
        RECT 65.020 69.260 65.160 69.800 ;
        RECT 65.850 69.400 66.170 69.660 ;
        RECT 66.400 69.615 66.540 70.140 ;
        RECT 68.625 70.095 68.915 70.325 ;
        RECT 69.070 70.280 69.390 70.340 ;
        RECT 72.290 70.280 72.610 70.340 ;
        RECT 69.070 70.140 72.610 70.280 ;
        RECT 66.785 69.940 67.075 69.985 ;
        RECT 68.150 69.940 68.470 70.000 ;
        RECT 66.785 69.800 68.470 69.940 ;
        RECT 68.700 69.940 68.840 70.095 ;
        RECT 69.070 70.080 69.390 70.140 ;
        RECT 72.290 70.080 72.610 70.140 ;
        RECT 75.050 70.080 75.370 70.340 ;
        RECT 77.365 69.940 77.655 69.985 ;
        RECT 68.700 69.800 77.655 69.940 ;
        RECT 66.785 69.755 67.075 69.800 ;
        RECT 68.150 69.740 68.470 69.800 ;
        RECT 77.365 69.755 77.655 69.800 ;
        RECT 66.400 69.600 67.000 69.615 ;
        RECT 67.245 69.600 67.535 69.645 ;
        RECT 66.400 69.475 67.535 69.600 ;
        RECT 66.860 69.460 67.535 69.475 ;
        RECT 67.245 69.415 67.535 69.460 ;
        RECT 67.705 69.415 67.995 69.645 ;
        RECT 69.085 69.600 69.375 69.645 ;
        RECT 69.530 69.600 69.850 69.660 ;
        RECT 69.085 69.460 69.850 69.600 ;
        RECT 69.085 69.415 69.375 69.460 ;
        RECT 66.310 69.260 66.630 69.320 ;
        RECT 65.020 69.120 66.630 69.260 ;
        RECT 67.780 69.260 67.920 69.415 ;
        RECT 69.530 69.400 69.850 69.460 ;
        RECT 69.990 69.400 70.310 69.660 ;
        RECT 70.465 69.415 70.755 69.645 ;
        RECT 70.925 69.600 71.215 69.645 ;
        RECT 71.370 69.600 71.690 69.660 ;
        RECT 70.925 69.460 71.690 69.600 ;
        RECT 70.925 69.415 71.215 69.460 ;
        RECT 68.150 69.260 68.470 69.320 ;
        RECT 67.780 69.120 68.470 69.260 ;
        RECT 70.540 69.260 70.680 69.415 ;
        RECT 71.370 69.400 71.690 69.460 ;
        RECT 76.905 69.600 77.195 69.645 ;
        RECT 79.205 69.600 79.495 69.645 ;
        RECT 76.905 69.460 79.495 69.600 ;
        RECT 76.905 69.415 77.195 69.460 ;
        RECT 79.205 69.415 79.495 69.460 ;
        RECT 80.570 69.600 80.890 69.660 ;
        RECT 81.965 69.600 82.255 69.645 ;
        RECT 80.570 69.460 82.255 69.600 ;
        RECT 80.570 69.400 80.890 69.460 ;
        RECT 81.965 69.415 82.255 69.460 ;
        RECT 71.830 69.260 72.150 69.320 ;
        RECT 70.540 69.120 72.150 69.260 ;
        RECT 66.310 69.060 66.630 69.120 ;
        RECT 68.150 69.060 68.470 69.120 ;
        RECT 71.830 69.060 72.150 69.120 ;
        RECT 77.825 69.075 78.115 69.305 ;
        RECT 72.305 68.920 72.595 68.965 ;
        RECT 77.900 68.920 78.040 69.075 ;
        RECT 63.645 68.780 65.160 68.920 ;
        RECT 58.950 68.580 59.270 68.640 ;
        RECT 13.730 68.440 59.270 68.580 ;
        RECT 11.110 68.380 11.430 68.440 ;
        RECT 11.585 68.395 11.875 68.440 ;
        RECT 58.950 68.380 59.270 68.440 ;
        RECT 64.470 68.380 64.790 68.640 ;
        RECT 65.020 68.580 65.160 68.780 ;
        RECT 72.305 68.780 78.040 68.920 ;
        RECT 72.305 68.735 72.595 68.780 ;
        RECT 67.690 68.580 68.010 68.640 ;
        RECT 65.020 68.440 68.010 68.580 ;
        RECT 67.690 68.380 68.010 68.440 ;
        RECT 5.520 67.760 84.180 68.240 ;
        RECT 11.570 67.560 11.890 67.620 ;
        RECT 12.950 67.560 13.270 67.620 ;
        RECT 13.885 67.560 14.175 67.605 ;
        RECT 11.570 67.420 14.175 67.560 ;
        RECT 11.570 67.360 11.890 67.420 ;
        RECT 12.950 67.360 13.270 67.420 ;
        RECT 13.885 67.375 14.175 67.420 ;
        RECT 65.850 67.360 66.170 67.620 ;
        RECT 67.690 67.360 68.010 67.620 ;
        RECT 68.625 67.560 68.915 67.605 ;
        RECT 69.990 67.560 70.310 67.620 ;
        RECT 68.625 67.420 70.310 67.560 ;
        RECT 68.625 67.375 68.915 67.420 ;
        RECT 69.990 67.360 70.310 67.420 ;
        RECT 7.470 67.220 7.760 67.265 ;
        RECT 9.570 67.220 9.860 67.265 ;
        RECT 11.140 67.220 11.430 67.265 ;
        RECT 7.470 67.080 11.430 67.220 ;
        RECT 7.470 67.035 7.760 67.080 ;
        RECT 9.570 67.035 9.860 67.080 ;
        RECT 11.140 67.035 11.430 67.080 ;
        RECT 13.410 67.220 13.730 67.280 ;
        RECT 17.090 67.220 17.410 67.280 ;
        RECT 13.410 67.080 17.410 67.220 ;
        RECT 13.410 67.020 13.730 67.080 ;
        RECT 17.090 67.020 17.410 67.080 ;
        RECT 19.430 67.220 19.720 67.265 ;
        RECT 21.530 67.220 21.820 67.265 ;
        RECT 23.100 67.220 23.390 67.265 ;
        RECT 19.430 67.080 23.390 67.220 ;
        RECT 19.430 67.035 19.720 67.080 ;
        RECT 21.530 67.035 21.820 67.080 ;
        RECT 23.100 67.035 23.390 67.080 ;
        RECT 33.230 67.220 33.520 67.265 ;
        RECT 35.330 67.220 35.620 67.265 ;
        RECT 36.900 67.220 37.190 67.265 ;
        RECT 33.230 67.080 37.190 67.220 ;
        RECT 33.230 67.035 33.520 67.080 ;
        RECT 35.330 67.035 35.620 67.080 ;
        RECT 36.900 67.035 37.190 67.080 ;
        RECT 39.645 67.220 39.935 67.265 ;
        RECT 64.470 67.220 64.790 67.280 ;
        RECT 66.310 67.220 66.630 67.280 ;
        RECT 67.780 67.220 67.920 67.360 ;
        RECT 39.645 67.080 47.680 67.220 ;
        RECT 39.645 67.035 39.935 67.080 ;
        RECT 47.540 66.940 47.680 67.080 ;
        RECT 64.470 67.080 67.920 67.220 ;
        RECT 69.070 67.220 69.390 67.280 ;
        RECT 71.370 67.220 71.690 67.280 ;
        RECT 69.070 67.080 71.690 67.220 ;
        RECT 64.470 67.020 64.790 67.080 ;
        RECT 66.310 67.020 66.630 67.080 ;
        RECT 69.070 67.020 69.390 67.080 ;
        RECT 71.370 67.020 71.690 67.080 ;
        RECT 7.865 66.880 8.155 66.925 ;
        RECT 9.055 66.880 9.345 66.925 ;
        RECT 11.575 66.880 11.865 66.925 ;
        RECT 7.865 66.740 11.865 66.880 ;
        RECT 7.865 66.695 8.155 66.740 ;
        RECT 9.055 66.695 9.345 66.740 ;
        RECT 11.575 66.695 11.865 66.740 ;
        RECT 18.930 66.680 19.250 66.940 ;
        RECT 19.825 66.880 20.115 66.925 ;
        RECT 21.015 66.880 21.305 66.925 ;
        RECT 23.535 66.880 23.825 66.925 ;
        RECT 19.825 66.740 23.825 66.880 ;
        RECT 19.825 66.695 20.115 66.740 ;
        RECT 21.015 66.695 21.305 66.740 ;
        RECT 23.535 66.695 23.825 66.740 ;
        RECT 31.825 66.880 32.115 66.925 ;
        RECT 33.625 66.880 33.915 66.925 ;
        RECT 34.815 66.880 35.105 66.925 ;
        RECT 37.335 66.880 37.625 66.925 ;
        RECT 31.825 66.740 32.500 66.880 ;
        RECT 31.825 66.695 32.115 66.740 ;
        RECT 6.985 66.540 7.275 66.585 ;
        RECT 13.870 66.540 14.190 66.600 ;
        RECT 6.985 66.400 14.190 66.540 ;
        RECT 6.985 66.355 7.275 66.400 ;
        RECT 13.870 66.340 14.190 66.400 ;
        RECT 7.430 66.200 7.750 66.260 ;
        RECT 8.210 66.200 8.500 66.245 ;
        RECT 7.430 66.060 8.500 66.200 ;
        RECT 7.430 66.000 7.750 66.060 ;
        RECT 8.210 66.015 8.500 66.060 ;
        RECT 20.280 66.200 20.570 66.245 ;
        RECT 21.230 66.200 21.550 66.260 ;
        RECT 20.280 66.060 21.550 66.200 ;
        RECT 32.360 66.200 32.500 66.740 ;
        RECT 33.625 66.740 37.625 66.880 ;
        RECT 33.625 66.695 33.915 66.740 ;
        RECT 34.815 66.695 35.105 66.740 ;
        RECT 37.335 66.695 37.625 66.740 ;
        RECT 43.325 66.880 43.615 66.925 ;
        RECT 44.230 66.880 44.550 66.940 ;
        RECT 43.325 66.740 44.550 66.880 ;
        RECT 43.325 66.695 43.615 66.740 ;
        RECT 44.230 66.680 44.550 66.740 ;
        RECT 47.450 66.680 47.770 66.940 ;
        RECT 56.190 66.880 56.510 66.940 ;
        RECT 56.665 66.880 56.955 66.925 ;
        RECT 56.190 66.740 56.955 66.880 ;
        RECT 56.190 66.680 56.510 66.740 ;
        RECT 56.665 66.695 56.955 66.740 ;
        RECT 60.330 66.880 60.650 66.940 ;
        RECT 61.725 66.880 62.015 66.925 ;
        RECT 60.330 66.740 67.000 66.880 ;
        RECT 60.330 66.680 60.650 66.740 ;
        RECT 61.725 66.695 62.015 66.740 ;
        RECT 32.745 66.540 33.035 66.585 ;
        RECT 33.190 66.540 33.510 66.600 ;
        RECT 41.010 66.540 41.330 66.600 ;
        RECT 32.745 66.400 33.510 66.540 ;
        RECT 32.745 66.355 33.035 66.400 ;
        RECT 33.190 66.340 33.510 66.400 ;
        RECT 33.740 66.400 41.330 66.540 ;
        RECT 33.740 66.200 33.880 66.400 ;
        RECT 41.010 66.340 41.330 66.400 ;
        RECT 51.130 66.540 51.450 66.600 ;
        RECT 52.985 66.540 53.275 66.585 ;
        RECT 57.570 66.540 57.890 66.600 ;
        RECT 51.130 66.400 57.890 66.540 ;
        RECT 51.130 66.340 51.450 66.400 ;
        RECT 52.985 66.355 53.275 66.400 ;
        RECT 57.570 66.340 57.890 66.400 ;
        RECT 58.045 66.355 58.335 66.585 ;
        RECT 32.360 66.060 33.880 66.200 ;
        RECT 34.080 66.200 34.370 66.245 ;
        RECT 49.290 66.200 49.610 66.260 ;
        RECT 58.120 66.200 58.260 66.355 ;
        RECT 62.630 66.340 62.950 66.600 ;
        RECT 63.090 66.540 63.410 66.600 ;
        RECT 64.485 66.540 64.775 66.585 ;
        RECT 63.090 66.400 64.775 66.540 ;
        RECT 63.090 66.340 63.410 66.400 ;
        RECT 64.485 66.355 64.775 66.400 ;
        RECT 64.945 66.355 65.235 66.585 ;
        RECT 34.080 66.060 40.320 66.200 ;
        RECT 20.280 66.015 20.570 66.060 ;
        RECT 21.230 66.000 21.550 66.060 ;
        RECT 34.080 66.015 34.370 66.060 ;
        RECT 25.845 65.860 26.135 65.905 ;
        RECT 26.290 65.860 26.610 65.920 ;
        RECT 25.845 65.720 26.610 65.860 ;
        RECT 25.845 65.675 26.135 65.720 ;
        RECT 26.290 65.660 26.610 65.720 ;
        RECT 28.590 65.660 28.910 65.920 ;
        RECT 30.430 65.660 30.750 65.920 ;
        RECT 30.890 65.660 31.210 65.920 ;
        RECT 40.180 65.905 40.320 66.060 ;
        RECT 49.290 66.060 58.260 66.200 ;
        RECT 58.950 66.200 59.270 66.260 ;
        RECT 63.550 66.200 63.870 66.260 ;
        RECT 65.020 66.200 65.160 66.355 ;
        RECT 65.390 66.340 65.710 66.600 ;
        RECT 66.860 66.585 67.000 66.740 ;
        RECT 67.230 66.680 67.550 66.940 ;
        RECT 72.290 66.880 72.610 66.940 ;
        RECT 72.290 66.740 73.440 66.880 ;
        RECT 72.290 66.680 72.610 66.740 ;
        RECT 66.325 66.355 66.615 66.585 ;
        RECT 66.785 66.355 67.075 66.585 ;
        RECT 58.950 66.060 62.170 66.200 ;
        RECT 49.290 66.000 49.610 66.060 ;
        RECT 58.950 66.000 59.270 66.060 ;
        RECT 40.105 65.675 40.395 65.905 ;
        RECT 41.930 65.660 42.250 65.920 ;
        RECT 42.405 65.860 42.695 65.905 ;
        RECT 44.705 65.860 44.995 65.905 ;
        RECT 42.405 65.720 44.995 65.860 ;
        RECT 42.405 65.675 42.695 65.720 ;
        RECT 44.705 65.675 44.995 65.720 ;
        RECT 59.410 65.860 59.730 65.920 ;
        RECT 61.265 65.860 61.555 65.905 ;
        RECT 59.410 65.720 61.555 65.860 ;
        RECT 62.030 65.860 62.170 66.060 ;
        RECT 63.550 66.060 65.160 66.200 ;
        RECT 65.850 66.200 66.170 66.260 ;
        RECT 66.400 66.200 66.540 66.355 ;
        RECT 67.320 66.200 67.460 66.680 ;
        RECT 71.370 66.340 71.690 66.600 ;
        RECT 73.300 66.585 73.440 66.740 ;
        RECT 73.225 66.355 73.515 66.585 ;
        RECT 78.745 66.540 79.035 66.585 ;
        RECT 79.650 66.540 79.970 66.600 ;
        RECT 78.745 66.400 79.970 66.540 ;
        RECT 78.745 66.355 79.035 66.400 ;
        RECT 79.650 66.340 79.970 66.400 ;
        RECT 81.950 66.340 82.270 66.600 ;
        RECT 65.850 66.060 67.460 66.200 ;
        RECT 70.910 66.200 71.230 66.260 ;
        RECT 71.830 66.200 72.150 66.260 ;
        RECT 72.305 66.200 72.595 66.245 ;
        RECT 70.910 66.060 72.595 66.200 ;
        RECT 63.550 66.000 63.870 66.060 ;
        RECT 65.850 66.000 66.170 66.060 ;
        RECT 70.910 66.000 71.230 66.060 ;
        RECT 71.830 66.000 72.150 66.060 ;
        RECT 72.305 66.015 72.595 66.060 ;
        RECT 72.765 66.200 73.055 66.245 ;
        RECT 75.050 66.200 75.370 66.260 ;
        RECT 72.765 66.060 75.370 66.200 ;
        RECT 72.765 66.015 73.055 66.060 ;
        RECT 72.840 65.860 72.980 66.015 ;
        RECT 75.050 66.000 75.370 66.060 ;
        RECT 62.030 65.720 72.980 65.860 ;
        RECT 74.145 65.860 74.435 65.905 ;
        RECT 76.890 65.860 77.210 65.920 ;
        RECT 74.145 65.720 77.210 65.860 ;
        RECT 59.410 65.660 59.730 65.720 ;
        RECT 61.265 65.675 61.555 65.720 ;
        RECT 74.145 65.675 74.435 65.720 ;
        RECT 76.890 65.660 77.210 65.720 ;
        RECT 77.810 65.660 78.130 65.920 ;
        RECT 79.190 65.660 79.510 65.920 ;
        RECT 5.520 65.040 84.180 65.520 ;
        RECT 6.510 64.840 6.830 64.900 ;
        RECT 7.445 64.840 7.735 64.885 ;
        RECT 6.510 64.700 7.735 64.840 ;
        RECT 6.510 64.640 6.830 64.700 ;
        RECT 7.445 64.655 7.735 64.700 ;
        RECT 8.440 64.700 15.940 64.840 ;
        RECT 8.440 64.205 8.580 64.700 ;
        RECT 13.870 64.500 14.190 64.560 ;
        RECT 9.820 64.360 14.190 64.500 ;
        RECT 9.820 64.205 9.960 64.360 ;
        RECT 13.870 64.300 14.190 64.360 ;
        RECT 11.110 64.205 11.430 64.220 ;
        RECT 8.365 63.975 8.655 64.205 ;
        RECT 9.745 63.975 10.035 64.205 ;
        RECT 11.080 64.160 11.430 64.205 ;
        RECT 10.915 64.020 11.430 64.160 ;
        RECT 15.800 64.160 15.940 64.700 ;
        RECT 16.645 64.655 16.935 64.885 ;
        RECT 19.405 64.840 19.695 64.885 ;
        RECT 19.850 64.840 20.170 64.900 ;
        RECT 19.405 64.700 20.170 64.840 ;
        RECT 19.405 64.655 19.695 64.700 ;
        RECT 16.720 64.500 16.860 64.655 ;
        RECT 19.850 64.640 20.170 64.700 ;
        RECT 21.230 64.640 21.550 64.900 ;
        RECT 30.430 64.840 30.750 64.900 ;
        RECT 32.285 64.840 32.575 64.885 ;
        RECT 30.430 64.700 32.575 64.840 ;
        RECT 30.430 64.640 30.750 64.700 ;
        RECT 32.285 64.655 32.575 64.700 ;
        RECT 35.490 64.840 35.810 64.900 ;
        RECT 40.550 64.840 40.870 64.900 ;
        RECT 35.490 64.700 40.870 64.840 ;
        RECT 35.490 64.640 35.810 64.700 ;
        RECT 40.550 64.640 40.870 64.700 ;
        RECT 45.165 64.840 45.455 64.885 ;
        RECT 46.530 64.840 46.850 64.900 ;
        RECT 45.165 64.700 46.850 64.840 ;
        RECT 45.165 64.655 45.455 64.700 ;
        RECT 46.530 64.640 46.850 64.700 ;
        RECT 47.465 64.840 47.755 64.885 ;
        RECT 49.290 64.840 49.610 64.900 ;
        RECT 47.465 64.700 49.610 64.840 ;
        RECT 47.465 64.655 47.755 64.700 ;
        RECT 49.290 64.640 49.610 64.700 ;
        RECT 57.585 64.655 57.875 64.885 ;
        RECT 17.090 64.500 17.410 64.560 ;
        RECT 54.980 64.500 55.270 64.545 ;
        RECT 57.660 64.500 57.800 64.655 ;
        RECT 59.410 64.640 59.730 64.900 ;
        RECT 66.785 64.655 67.075 64.885 ;
        RECT 70.465 64.840 70.755 64.885 ;
        RECT 78.730 64.840 79.050 64.900 ;
        RECT 70.465 64.700 79.050 64.840 ;
        RECT 70.465 64.655 70.755 64.700 ;
        RECT 16.720 64.360 51.820 64.500 ;
        RECT 17.090 64.300 17.410 64.360 ;
        RECT 15.800 64.020 23.300 64.160 ;
        RECT 11.080 63.975 11.430 64.020 ;
        RECT 11.110 63.960 11.430 63.975 ;
        RECT 10.625 63.820 10.915 63.865 ;
        RECT 11.815 63.820 12.105 63.865 ;
        RECT 14.335 63.820 14.625 63.865 ;
        RECT 10.625 63.680 14.625 63.820 ;
        RECT 10.625 63.635 10.915 63.680 ;
        RECT 11.815 63.635 12.105 63.680 ;
        RECT 14.335 63.635 14.625 63.680 ;
        RECT 18.010 63.620 18.330 63.880 ;
        RECT 18.945 63.820 19.235 63.865 ;
        RECT 20.310 63.820 20.630 63.880 ;
        RECT 18.945 63.680 20.630 63.820 ;
        RECT 23.160 63.820 23.300 64.020 ;
        RECT 35.490 63.960 35.810 64.220 ;
        RECT 35.950 63.960 36.270 64.220 ;
        RECT 36.425 64.160 36.715 64.205 ;
        RECT 36.870 64.160 37.190 64.220 ;
        RECT 36.425 64.020 37.190 64.160 ;
        RECT 36.425 63.975 36.715 64.020 ;
        RECT 36.870 63.960 37.190 64.020 ;
        RECT 37.345 63.975 37.635 64.205 ;
        RECT 37.805 64.160 38.095 64.205 ;
        RECT 41.470 64.160 41.790 64.220 ;
        RECT 37.805 64.020 41.790 64.160 ;
        RECT 37.805 63.975 38.095 64.020 ;
        RECT 23.530 63.820 23.850 63.880 ;
        RECT 37.420 63.820 37.560 63.975 ;
        RECT 41.470 63.960 41.790 64.020 ;
        RECT 47.005 64.160 47.295 64.205 ;
        RECT 51.130 64.160 51.450 64.220 ;
        RECT 47.005 64.020 51.450 64.160 ;
        RECT 51.680 64.160 51.820 64.360 ;
        RECT 54.980 64.360 57.800 64.500 ;
        RECT 58.120 64.360 66.540 64.500 ;
        RECT 54.980 64.315 55.270 64.360 ;
        RECT 58.120 64.160 58.260 64.360 ;
        RECT 51.680 64.020 58.260 64.160 ;
        RECT 59.885 64.160 60.175 64.205 ;
        RECT 60.790 64.160 61.110 64.220 ;
        RECT 63.090 64.160 63.410 64.220 ;
        RECT 59.885 64.020 63.410 64.160 ;
        RECT 47.005 63.975 47.295 64.020 ;
        RECT 51.130 63.960 51.450 64.020 ;
        RECT 59.885 63.975 60.175 64.020 ;
        RECT 60.790 63.960 61.110 64.020 ;
        RECT 63.090 63.960 63.410 64.020 ;
        RECT 64.470 64.160 64.790 64.220 ;
        RECT 64.945 64.160 65.235 64.205 ;
        RECT 64.470 64.020 65.235 64.160 ;
        RECT 64.470 63.960 64.790 64.020 ;
        RECT 64.945 63.975 65.235 64.020 ;
        RECT 65.850 63.960 66.170 64.220 ;
        RECT 23.160 63.680 37.560 63.820 ;
        RECT 18.945 63.635 19.235 63.680 ;
        RECT 20.310 63.620 20.630 63.680 ;
        RECT 23.530 63.620 23.850 63.680 ;
        RECT 40.550 63.620 40.870 63.880 ;
        RECT 43.310 63.620 43.630 63.880 ;
        RECT 47.925 63.635 48.215 63.865 ;
        RECT 51.615 63.820 51.905 63.865 ;
        RECT 54.135 63.820 54.425 63.865 ;
        RECT 55.325 63.820 55.615 63.865 ;
        RECT 51.615 63.680 55.615 63.820 ;
        RECT 51.615 63.635 51.905 63.680 ;
        RECT 54.135 63.635 54.425 63.680 ;
        RECT 55.325 63.635 55.615 63.680 ;
        RECT 56.205 63.820 56.495 63.865 ;
        RECT 56.650 63.820 56.970 63.880 ;
        RECT 56.205 63.680 56.970 63.820 ;
        RECT 56.205 63.635 56.495 63.680 ;
        RECT 10.230 63.480 10.520 63.525 ;
        RECT 12.330 63.480 12.620 63.525 ;
        RECT 13.900 63.480 14.190 63.525 ;
        RECT 10.230 63.340 14.190 63.480 ;
        RECT 10.230 63.295 10.520 63.340 ;
        RECT 12.330 63.295 12.620 63.340 ;
        RECT 13.900 63.295 14.190 63.340 ;
        RECT 38.725 63.480 39.015 63.525 ;
        RECT 45.150 63.480 45.470 63.540 ;
        RECT 38.725 63.340 45.470 63.480 ;
        RECT 38.725 63.295 39.015 63.340 ;
        RECT 45.150 63.280 45.470 63.340 ;
        RECT 11.570 63.140 11.890 63.200 ;
        RECT 13.410 63.140 13.730 63.200 ;
        RECT 11.570 63.000 13.730 63.140 ;
        RECT 11.570 62.940 11.890 63.000 ;
        RECT 13.410 62.940 13.730 63.000 ;
        RECT 39.630 63.140 39.950 63.200 ;
        RECT 48.000 63.140 48.140 63.635 ;
        RECT 56.650 63.620 56.970 63.680 ;
        RECT 60.345 63.820 60.635 63.865 ;
        RECT 61.710 63.820 62.030 63.880 ;
        RECT 60.345 63.680 62.030 63.820 ;
        RECT 66.400 63.820 66.540 64.360 ;
        RECT 66.860 64.160 67.000 64.655 ;
        RECT 78.730 64.640 79.050 64.700 ;
        RECT 80.570 64.840 80.890 64.900 ;
        RECT 81.045 64.840 81.335 64.885 ;
        RECT 81.950 64.840 82.270 64.900 ;
        RECT 80.570 64.700 82.270 64.840 ;
        RECT 80.570 64.640 80.890 64.700 ;
        RECT 81.045 64.655 81.335 64.700 ;
        RECT 81.950 64.640 82.270 64.700 ;
        RECT 69.530 64.500 69.850 64.560 ;
        RECT 68.240 64.360 69.850 64.500 ;
        RECT 68.240 64.205 68.380 64.360 ;
        RECT 69.530 64.300 69.850 64.360 ;
        RECT 71.830 64.300 72.150 64.560 ;
        RECT 75.480 64.500 75.770 64.545 ;
        RECT 75.970 64.500 76.290 64.560 ;
        RECT 75.480 64.360 76.290 64.500 ;
        RECT 75.480 64.315 75.770 64.360 ;
        RECT 75.970 64.300 76.290 64.360 ;
        RECT 67.245 64.160 67.535 64.205 ;
        RECT 66.860 64.020 67.535 64.160 ;
        RECT 67.245 63.975 67.535 64.020 ;
        RECT 68.165 63.975 68.455 64.205 ;
        RECT 68.610 63.960 68.930 64.220 ;
        RECT 69.070 63.960 69.390 64.220 ;
        RECT 70.910 63.960 71.230 64.220 ;
        RECT 72.305 63.975 72.595 64.205 ;
        RECT 72.380 63.820 72.520 63.975 ;
        RECT 72.750 63.960 73.070 64.220 ;
        RECT 73.670 64.160 73.990 64.220 ;
        RECT 74.145 64.160 74.435 64.205 ;
        RECT 73.670 64.020 74.435 64.160 ;
        RECT 73.670 63.960 73.990 64.020 ;
        RECT 74.145 63.975 74.435 64.020 ;
        RECT 74.590 63.960 74.910 64.220 ;
        RECT 82.410 63.960 82.730 64.220 ;
        RECT 74.680 63.820 74.820 63.960 ;
        RECT 66.400 63.680 74.820 63.820 ;
        RECT 75.025 63.820 75.315 63.865 ;
        RECT 76.215 63.820 76.505 63.865 ;
        RECT 78.735 63.820 79.025 63.865 ;
        RECT 75.025 63.680 79.025 63.820 ;
        RECT 60.345 63.635 60.635 63.680 ;
        RECT 61.710 63.620 62.030 63.680 ;
        RECT 75.025 63.635 75.315 63.680 ;
        RECT 76.215 63.635 76.505 63.680 ;
        RECT 78.735 63.635 79.025 63.680 ;
        RECT 52.050 63.480 52.340 63.525 ;
        RECT 53.620 63.480 53.910 63.525 ;
        RECT 55.720 63.480 56.010 63.525 ;
        RECT 52.050 63.340 56.010 63.480 ;
        RECT 52.050 63.295 52.340 63.340 ;
        RECT 53.620 63.295 53.910 63.340 ;
        RECT 55.720 63.295 56.010 63.340 ;
        RECT 64.010 63.480 64.330 63.540 ;
        RECT 68.610 63.480 68.930 63.540 ;
        RECT 64.010 63.340 68.930 63.480 ;
        RECT 64.010 63.280 64.330 63.340 ;
        RECT 68.610 63.280 68.930 63.340 ;
        RECT 69.530 63.480 69.850 63.540 ;
        RECT 72.750 63.480 73.070 63.540 ;
        RECT 69.530 63.340 73.070 63.480 ;
        RECT 69.530 63.280 69.850 63.340 ;
        RECT 72.750 63.280 73.070 63.340 ;
        RECT 74.630 63.480 74.920 63.525 ;
        RECT 76.730 63.480 77.020 63.525 ;
        RECT 78.300 63.480 78.590 63.525 ;
        RECT 74.630 63.340 78.590 63.480 ;
        RECT 74.630 63.295 74.920 63.340 ;
        RECT 76.730 63.295 77.020 63.340 ;
        RECT 78.300 63.295 78.590 63.340 ;
        RECT 80.110 63.480 80.430 63.540 ;
        RECT 81.505 63.480 81.795 63.525 ;
        RECT 80.110 63.340 81.795 63.480 ;
        RECT 80.110 63.280 80.430 63.340 ;
        RECT 81.505 63.295 81.795 63.340 ;
        RECT 50.670 63.140 50.990 63.200 ;
        RECT 52.510 63.140 52.830 63.200 ;
        RECT 39.630 63.000 52.830 63.140 ;
        RECT 39.630 62.940 39.950 63.000 ;
        RECT 50.670 62.940 50.990 63.000 ;
        RECT 52.510 62.940 52.830 63.000 ;
        RECT 64.930 62.940 65.250 63.200 ;
        RECT 73.685 63.140 73.975 63.185 ;
        RECT 77.810 63.140 78.130 63.200 ;
        RECT 73.685 63.000 78.130 63.140 ;
        RECT 73.685 62.955 73.975 63.000 ;
        RECT 77.810 62.940 78.130 63.000 ;
        RECT 5.520 62.320 84.180 62.800 ;
        RECT 20.310 62.120 20.630 62.180 ;
        RECT 26.290 62.120 26.610 62.180 ;
        RECT 32.730 62.120 33.050 62.180 ;
        RECT 20.310 61.980 33.050 62.120 ;
        RECT 20.310 61.920 20.630 61.980 ;
        RECT 26.290 61.920 26.610 61.980 ;
        RECT 32.730 61.920 33.050 61.980 ;
        RECT 33.665 62.120 33.955 62.165 ;
        RECT 35.490 62.120 35.810 62.180 ;
        RECT 33.665 61.980 35.810 62.120 ;
        RECT 33.665 61.935 33.955 61.980 ;
        RECT 35.490 61.920 35.810 61.980 ;
        RECT 41.470 62.120 41.790 62.180 ;
        RECT 42.390 62.120 42.710 62.180 ;
        RECT 41.470 61.980 42.710 62.120 ;
        RECT 41.470 61.920 41.790 61.980 ;
        RECT 42.390 61.920 42.710 61.980 ;
        RECT 51.590 61.920 51.910 62.180 ;
        RECT 69.545 62.120 69.835 62.165 ;
        RECT 70.910 62.120 71.230 62.180 ;
        RECT 69.545 61.980 71.230 62.120 ;
        RECT 69.545 61.935 69.835 61.980 ;
        RECT 70.910 61.920 71.230 61.980 ;
        RECT 75.970 61.920 76.290 62.180 ;
        RECT 26.750 61.780 27.070 61.840 ;
        RECT 10.280 61.640 27.070 61.780 ;
        RECT 8.350 60.900 8.670 61.160 ;
        RECT 10.280 61.145 10.420 61.640 ;
        RECT 26.750 61.580 27.070 61.640 ;
        RECT 27.250 61.780 27.540 61.825 ;
        RECT 29.350 61.780 29.640 61.825 ;
        RECT 30.920 61.780 31.210 61.825 ;
        RECT 27.250 61.640 31.210 61.780 ;
        RECT 27.250 61.595 27.540 61.640 ;
        RECT 29.350 61.595 29.640 61.640 ;
        RECT 30.920 61.595 31.210 61.640 ;
        RECT 45.190 61.780 45.480 61.825 ;
        RECT 47.290 61.780 47.580 61.825 ;
        RECT 48.860 61.780 49.150 61.825 ;
        RECT 45.190 61.640 49.150 61.780 ;
        RECT 45.190 61.595 45.480 61.640 ;
        RECT 47.290 61.595 47.580 61.640 ;
        RECT 48.860 61.595 49.150 61.640 ;
        RECT 19.390 61.440 19.710 61.500 ;
        RECT 27.645 61.440 27.935 61.485 ;
        RECT 28.835 61.440 29.125 61.485 ;
        RECT 31.355 61.440 31.645 61.485 ;
        RECT 19.390 61.300 20.540 61.440 ;
        RECT 19.390 61.240 19.710 61.300 ;
        RECT 10.205 60.915 10.495 61.145 ;
        RECT 13.425 61.100 13.715 61.145 ;
        RECT 14.790 61.100 15.110 61.160 ;
        RECT 20.400 61.145 20.540 61.300 ;
        RECT 27.645 61.300 31.645 61.440 ;
        RECT 27.645 61.255 27.935 61.300 ;
        RECT 28.835 61.255 29.125 61.300 ;
        RECT 31.355 61.255 31.645 61.300 ;
        RECT 40.105 61.440 40.395 61.485 ;
        RECT 41.010 61.440 41.330 61.500 ;
        RECT 40.105 61.300 41.330 61.440 ;
        RECT 40.105 61.255 40.395 61.300 ;
        RECT 41.010 61.240 41.330 61.300 ;
        RECT 44.690 61.240 45.010 61.500 ;
        RECT 45.585 61.440 45.875 61.485 ;
        RECT 46.775 61.440 47.065 61.485 ;
        RECT 49.295 61.440 49.585 61.485 ;
        RECT 45.585 61.300 49.585 61.440 ;
        RECT 51.680 61.440 51.820 61.920 ;
        RECT 81.950 61.580 82.270 61.840 ;
        RECT 54.825 61.440 55.115 61.485 ;
        RECT 51.680 61.300 55.115 61.440 ;
        RECT 45.585 61.255 45.875 61.300 ;
        RECT 46.775 61.255 47.065 61.300 ;
        RECT 49.295 61.255 49.585 61.300 ;
        RECT 54.825 61.255 55.115 61.300 ;
        RECT 59.425 61.440 59.715 61.485 ;
        RECT 59.870 61.440 60.190 61.500 ;
        RECT 62.630 61.440 62.950 61.500 ;
        RECT 65.850 61.440 66.170 61.500 ;
        RECT 59.425 61.300 60.190 61.440 ;
        RECT 59.425 61.255 59.715 61.300 ;
        RECT 59.870 61.240 60.190 61.300 ;
        RECT 60.880 61.300 66.170 61.440 ;
        RECT 13.425 60.960 15.110 61.100 ;
        RECT 13.425 60.915 13.715 60.960 ;
        RECT 14.790 60.900 15.110 60.960 ;
        RECT 20.325 60.915 20.615 61.145 ;
        RECT 20.785 60.915 21.075 61.145 ;
        RECT 21.245 60.915 21.535 61.145 ;
        RECT 19.390 60.760 19.710 60.820 ;
        RECT 20.860 60.760 21.000 60.915 ;
        RECT 19.390 60.620 21.000 60.760 ;
        RECT 19.390 60.560 19.710 60.620 ;
        RECT 4.210 60.420 4.530 60.480 ;
        RECT 7.445 60.420 7.735 60.465 ;
        RECT 4.210 60.280 7.735 60.420 ;
        RECT 4.210 60.220 4.530 60.280 ;
        RECT 7.445 60.235 7.735 60.280 ;
        RECT 9.270 60.220 9.590 60.480 ;
        RECT 12.505 60.420 12.795 60.465 ;
        RECT 15.250 60.420 15.570 60.480 ;
        RECT 12.505 60.280 15.570 60.420 ;
        RECT 12.505 60.235 12.795 60.280 ;
        RECT 15.250 60.220 15.570 60.280 ;
        RECT 18.010 60.420 18.330 60.480 ;
        RECT 18.945 60.420 19.235 60.465 ;
        RECT 18.010 60.280 19.235 60.420 ;
        RECT 18.010 60.220 18.330 60.280 ;
        RECT 18.945 60.235 19.235 60.280 ;
        RECT 20.310 60.420 20.630 60.480 ;
        RECT 21.320 60.420 21.460 60.915 ;
        RECT 22.150 60.900 22.470 61.160 ;
        RECT 23.530 60.900 23.850 61.160 ;
        RECT 26.765 61.100 27.055 61.145 ;
        RECT 33.190 61.100 33.510 61.160 ;
        RECT 26.765 60.960 33.510 61.100 ;
        RECT 26.765 60.915 27.055 60.960 ;
        RECT 33.190 60.900 33.510 60.960 ;
        RECT 38.725 61.100 39.015 61.145 ;
        RECT 40.550 61.100 40.870 61.160 ;
        RECT 38.725 60.960 40.870 61.100 ;
        RECT 38.725 60.915 39.015 60.960 ;
        RECT 40.550 60.900 40.870 60.960 ;
        RECT 43.325 61.100 43.615 61.145 ;
        RECT 43.770 61.100 44.090 61.160 ;
        RECT 43.325 60.960 44.090 61.100 ;
        RECT 43.325 60.915 43.615 60.960 ;
        RECT 43.770 60.900 44.090 60.960 ;
        RECT 50.210 61.100 50.530 61.160 ;
        RECT 55.745 61.100 56.035 61.145 ;
        RECT 50.210 60.960 56.035 61.100 ;
        RECT 50.210 60.900 50.530 60.960 ;
        RECT 55.745 60.915 56.035 60.960 ;
        RECT 58.030 61.100 58.350 61.160 ;
        RECT 60.330 61.100 60.650 61.160 ;
        RECT 60.880 61.145 61.020 61.300 ;
        RECT 62.630 61.240 62.950 61.300 ;
        RECT 65.850 61.240 66.170 61.300 ;
        RECT 66.325 61.440 66.615 61.485 ;
        RECT 69.070 61.440 69.390 61.500 ;
        RECT 73.670 61.440 73.990 61.500 ;
        RECT 66.325 61.300 73.990 61.440 ;
        RECT 66.325 61.255 66.615 61.300 ;
        RECT 69.070 61.240 69.390 61.300 ;
        RECT 73.670 61.240 73.990 61.300 ;
        RECT 77.810 61.440 78.130 61.500 ;
        RECT 78.285 61.440 78.575 61.485 ;
        RECT 77.810 61.300 78.575 61.440 ;
        RECT 77.810 61.240 78.130 61.300 ;
        RECT 78.285 61.255 78.575 61.300 ;
        RECT 78.730 61.240 79.050 61.500 ;
        RECT 58.030 60.960 60.650 61.100 ;
        RECT 58.030 60.900 58.350 60.960 ;
        RECT 60.330 60.900 60.650 60.960 ;
        RECT 60.805 60.915 61.095 61.145 ;
        RECT 64.930 61.100 65.250 61.160 ;
        RECT 67.705 61.100 67.995 61.145 ;
        RECT 64.930 60.960 67.995 61.100 ;
        RECT 64.930 60.900 65.250 60.960 ;
        RECT 67.705 60.915 67.995 60.960 ;
        RECT 68.625 61.100 68.915 61.145 ;
        RECT 69.990 61.100 70.310 61.160 ;
        RECT 71.830 61.100 72.150 61.160 ;
        RECT 68.625 60.960 72.150 61.100 ;
        RECT 68.625 60.915 68.915 60.960 ;
        RECT 69.990 60.900 70.310 60.960 ;
        RECT 71.830 60.900 72.150 60.960 ;
        RECT 72.765 61.100 73.055 61.145 ;
        RECT 80.110 61.100 80.430 61.160 ;
        RECT 72.765 60.960 80.430 61.100 ;
        RECT 72.765 60.915 73.055 60.960 ;
        RECT 80.110 60.900 80.430 60.960 ;
        RECT 81.045 61.100 81.335 61.145 ;
        RECT 81.490 61.100 81.810 61.160 ;
        RECT 81.045 60.960 81.810 61.100 ;
        RECT 81.045 60.915 81.335 60.960 ;
        RECT 81.490 60.900 81.810 60.960 ;
        RECT 22.625 60.575 22.915 60.805 ;
        RECT 28.100 60.760 28.390 60.805 ;
        RECT 28.590 60.760 28.910 60.820 ;
        RECT 28.100 60.620 28.910 60.760 ;
        RECT 28.100 60.575 28.390 60.620 ;
        RECT 20.310 60.280 21.460 60.420 ;
        RECT 21.690 60.420 22.010 60.480 ;
        RECT 22.700 60.420 22.840 60.575 ;
        RECT 28.590 60.560 28.910 60.620 ;
        RECT 46.040 60.760 46.330 60.805 ;
        RECT 47.450 60.760 47.770 60.820 ;
        RECT 46.040 60.620 47.770 60.760 ;
        RECT 46.040 60.575 46.330 60.620 ;
        RECT 47.450 60.560 47.770 60.620 ;
        RECT 57.570 60.760 57.890 60.820 ;
        RECT 59.870 60.760 60.190 60.820 ;
        RECT 62.185 60.760 62.475 60.805 ;
        RECT 57.570 60.620 62.475 60.760 ;
        RECT 57.570 60.560 57.890 60.620 ;
        RECT 59.870 60.560 60.190 60.620 ;
        RECT 62.185 60.575 62.475 60.620 ;
        RECT 77.825 60.760 78.115 60.805 ;
        RECT 79.190 60.760 79.510 60.820 ;
        RECT 77.825 60.620 79.510 60.760 ;
        RECT 77.825 60.575 78.115 60.620 ;
        RECT 79.190 60.560 79.510 60.620 ;
        RECT 21.690 60.280 22.840 60.420 ;
        RECT 23.990 60.420 24.310 60.480 ;
        RECT 24.465 60.420 24.755 60.465 ;
        RECT 23.990 60.280 24.755 60.420 ;
        RECT 20.310 60.220 20.630 60.280 ;
        RECT 21.690 60.220 22.010 60.280 ;
        RECT 23.990 60.220 24.310 60.280 ;
        RECT 24.465 60.235 24.755 60.280 ;
        RECT 36.870 60.220 37.190 60.480 ;
        RECT 39.170 60.220 39.490 60.480 ;
        RECT 41.470 60.420 41.790 60.480 ;
        RECT 42.865 60.420 43.155 60.465 ;
        RECT 44.690 60.420 45.010 60.480 ;
        RECT 41.470 60.280 45.010 60.420 ;
        RECT 41.470 60.220 41.790 60.280 ;
        RECT 42.865 60.235 43.155 60.280 ;
        RECT 44.690 60.220 45.010 60.280 ;
        RECT 52.050 60.220 52.370 60.480 ;
        RECT 58.950 60.220 59.270 60.480 ;
        RECT 59.410 60.220 59.730 60.480 ;
        RECT 75.525 60.420 75.815 60.465 ;
        RECT 77.350 60.420 77.670 60.480 ;
        RECT 75.525 60.280 77.670 60.420 ;
        RECT 75.525 60.235 75.815 60.280 ;
        RECT 77.350 60.220 77.670 60.280 ;
        RECT 5.520 59.600 84.180 60.080 ;
        RECT 18.930 59.400 19.250 59.460 ;
        RECT 21.690 59.400 22.010 59.460 ;
        RECT 8.440 59.260 22.010 59.400 ;
        RECT 8.440 59.105 8.580 59.260 ;
        RECT 18.930 59.200 19.250 59.260 ;
        RECT 21.690 59.200 22.010 59.260 ;
        RECT 23.530 59.400 23.850 59.460 ;
        RECT 30.905 59.400 31.195 59.445 ;
        RECT 23.530 59.260 31.195 59.400 ;
        RECT 23.530 59.200 23.850 59.260 ;
        RECT 30.905 59.215 31.195 59.260 ;
        RECT 41.485 59.400 41.775 59.445 ;
        RECT 43.310 59.400 43.630 59.460 ;
        RECT 41.485 59.260 43.630 59.400 ;
        RECT 41.485 59.215 41.775 59.260 ;
        RECT 43.310 59.200 43.630 59.260 ;
        RECT 45.150 59.200 45.470 59.460 ;
        RECT 47.450 59.200 47.770 59.460 ;
        RECT 49.765 59.400 50.055 59.445 ;
        RECT 50.210 59.400 50.530 59.460 ;
        RECT 49.765 59.260 50.530 59.400 ;
        RECT 49.765 59.215 50.055 59.260 ;
        RECT 50.210 59.200 50.530 59.260 ;
        RECT 57.585 59.215 57.875 59.445 ;
        RECT 58.950 59.400 59.270 59.460 ;
        RECT 58.950 59.260 60.560 59.400 ;
        RECT 8.365 58.875 8.655 59.105 ;
        RECT 9.285 59.060 9.575 59.105 ;
        RECT 14.330 59.060 14.650 59.120 ;
        RECT 24.450 59.060 24.770 59.120 ;
        RECT 27.670 59.060 27.990 59.120 ;
        RECT 9.285 58.920 14.650 59.060 ;
        RECT 9.285 58.875 9.575 58.920 ;
        RECT 14.330 58.860 14.650 58.920 ;
        RECT 16.720 58.920 24.220 59.060 ;
        RECT 13.870 58.720 14.190 58.780 ;
        RECT 16.720 58.765 16.860 58.920 ;
        RECT 18.010 58.765 18.330 58.780 ;
        RECT 24.080 58.765 24.220 58.920 ;
        RECT 24.450 58.920 27.990 59.060 ;
        RECT 24.450 58.860 24.770 58.920 ;
        RECT 27.670 58.860 27.990 58.920 ;
        RECT 35.920 59.060 36.210 59.105 ;
        RECT 36.870 59.060 37.190 59.120 ;
        RECT 35.920 58.920 37.190 59.060 ;
        RECT 35.920 58.875 36.210 58.920 ;
        RECT 36.870 58.860 37.190 58.920 ;
        RECT 45.625 59.060 45.915 59.105 ;
        RECT 52.050 59.060 52.370 59.120 ;
        RECT 45.625 58.920 52.370 59.060 ;
        RECT 45.625 58.875 45.915 58.920 ;
        RECT 52.050 58.860 52.370 58.920 ;
        RECT 55.440 59.060 55.730 59.105 ;
        RECT 57.660 59.060 57.800 59.215 ;
        RECT 58.950 59.200 59.270 59.260 ;
        RECT 55.440 58.920 57.800 59.060 ;
        RECT 55.440 58.875 55.730 58.920 ;
        RECT 59.410 58.860 59.730 59.120 ;
        RECT 25.370 58.765 25.690 58.780 ;
        RECT 16.645 58.720 16.935 58.765 ;
        RECT 17.980 58.720 18.330 58.765 ;
        RECT 13.870 58.580 16.935 58.720 ;
        RECT 17.815 58.580 18.330 58.720 ;
        RECT 13.870 58.520 14.190 58.580 ;
        RECT 16.645 58.535 16.935 58.580 ;
        RECT 17.980 58.535 18.330 58.580 ;
        RECT 24.005 58.535 24.295 58.765 ;
        RECT 25.340 58.535 25.690 58.765 ;
        RECT 18.010 58.520 18.330 58.535 ;
        RECT 25.370 58.520 25.690 58.535 ;
        RECT 33.190 58.720 33.510 58.780 ;
        RECT 34.585 58.720 34.875 58.765 ;
        RECT 33.190 58.580 34.875 58.720 ;
        RECT 33.190 58.520 33.510 58.580 ;
        RECT 34.585 58.535 34.875 58.580 ;
        RECT 56.650 58.520 56.970 58.780 ;
        RECT 58.030 58.720 58.350 58.780 ;
        RECT 58.505 58.720 58.795 58.765 ;
        RECT 58.030 58.580 58.795 58.720 ;
        RECT 58.030 58.520 58.350 58.580 ;
        RECT 58.505 58.535 58.795 58.580 ;
        RECT 58.950 58.520 59.270 58.780 ;
        RECT 60.420 58.765 60.560 59.260 ;
        RECT 63.090 59.200 63.410 59.460 ;
        RECT 71.370 59.400 71.690 59.460 ;
        RECT 73.685 59.400 73.975 59.445 ;
        RECT 71.370 59.260 73.975 59.400 ;
        RECT 71.370 59.200 71.690 59.260 ;
        RECT 73.685 59.215 73.975 59.260 ;
        RECT 77.350 59.200 77.670 59.460 ;
        RECT 79.650 59.200 79.970 59.460 ;
        RECT 63.180 59.060 63.320 59.200 ;
        RECT 66.770 59.060 67.090 59.120 ;
        RECT 61.800 58.920 67.090 59.060 ;
        RECT 60.345 58.535 60.635 58.765 ;
        RECT 60.790 58.520 61.110 58.780 ;
        RECT 61.800 58.765 61.940 58.920 ;
        RECT 66.770 58.860 67.090 58.920 ;
        RECT 61.725 58.535 62.015 58.765 ;
        RECT 63.105 58.720 63.395 58.765 ;
        RECT 69.070 58.720 69.390 58.780 ;
        RECT 63.105 58.580 69.390 58.720 ;
        RECT 63.105 58.535 63.395 58.580 ;
        RECT 14.790 58.180 15.110 58.440 ;
        RECT 16.170 58.180 16.490 58.440 ;
        RECT 17.525 58.380 17.815 58.425 ;
        RECT 18.715 58.380 19.005 58.425 ;
        RECT 21.235 58.380 21.525 58.425 ;
        RECT 17.525 58.240 21.525 58.380 ;
        RECT 17.525 58.195 17.815 58.240 ;
        RECT 18.715 58.195 19.005 58.240 ;
        RECT 21.235 58.195 21.525 58.240 ;
        RECT 24.885 58.380 25.175 58.425 ;
        RECT 26.075 58.380 26.365 58.425 ;
        RECT 28.595 58.380 28.885 58.425 ;
        RECT 24.885 58.240 28.885 58.380 ;
        RECT 24.885 58.195 25.175 58.240 ;
        RECT 26.075 58.195 26.365 58.240 ;
        RECT 28.595 58.195 28.885 58.240 ;
        RECT 35.465 58.380 35.755 58.425 ;
        RECT 36.655 58.380 36.945 58.425 ;
        RECT 39.175 58.380 39.465 58.425 ;
        RECT 35.465 58.240 39.465 58.380 ;
        RECT 35.465 58.195 35.755 58.240 ;
        RECT 36.655 58.195 36.945 58.240 ;
        RECT 39.175 58.195 39.465 58.240 ;
        RECT 44.690 58.380 45.010 58.440 ;
        RECT 47.910 58.380 48.230 58.440 ;
        RECT 44.690 58.240 48.230 58.380 ;
        RECT 44.690 58.180 45.010 58.240 ;
        RECT 47.910 58.180 48.230 58.240 ;
        RECT 52.075 58.380 52.365 58.425 ;
        RECT 54.595 58.380 54.885 58.425 ;
        RECT 55.785 58.380 56.075 58.425 ;
        RECT 52.075 58.240 56.075 58.380 ;
        RECT 56.740 58.380 56.880 58.520 ;
        RECT 63.180 58.380 63.320 58.535 ;
        RECT 69.070 58.520 69.390 58.580 ;
        RECT 69.990 58.720 70.310 58.780 ;
        RECT 73.210 58.720 73.530 58.780 ;
        RECT 69.990 58.580 73.530 58.720 ;
        RECT 69.990 58.520 70.310 58.580 ;
        RECT 73.210 58.520 73.530 58.580 ;
        RECT 74.145 58.535 74.435 58.765 ;
        RECT 56.740 58.240 63.320 58.380 ;
        RECT 65.850 58.380 66.170 58.440 ;
        RECT 74.220 58.380 74.360 58.535 ;
        RECT 80.570 58.520 80.890 58.780 ;
        RECT 81.030 58.520 81.350 58.780 ;
        RECT 65.850 58.240 74.360 58.380 ;
        RECT 52.075 58.195 52.365 58.240 ;
        RECT 54.595 58.195 54.885 58.240 ;
        RECT 55.785 58.195 56.075 58.240 ;
        RECT 65.850 58.180 66.170 58.240 ;
        RECT 77.810 58.180 78.130 58.440 ;
        RECT 78.285 58.195 78.575 58.425 ;
        RECT 8.350 58.040 8.670 58.100 ;
        RECT 17.130 58.040 17.420 58.085 ;
        RECT 19.230 58.040 19.520 58.085 ;
        RECT 20.800 58.040 21.090 58.085 ;
        RECT 8.350 57.900 13.870 58.040 ;
        RECT 8.350 57.840 8.670 57.900 ;
        RECT 10.205 57.700 10.495 57.745 ;
        RECT 10.650 57.700 10.970 57.760 ;
        RECT 10.205 57.560 10.970 57.700 ;
        RECT 13.730 57.700 13.870 57.900 ;
        RECT 17.130 57.900 21.090 58.040 ;
        RECT 17.130 57.855 17.420 57.900 ;
        RECT 19.230 57.855 19.520 57.900 ;
        RECT 20.800 57.855 21.090 57.900 ;
        RECT 24.490 58.040 24.780 58.085 ;
        RECT 26.590 58.040 26.880 58.085 ;
        RECT 28.160 58.040 28.450 58.085 ;
        RECT 24.490 57.900 28.450 58.040 ;
        RECT 24.490 57.855 24.780 57.900 ;
        RECT 26.590 57.855 26.880 57.900 ;
        RECT 28.160 57.855 28.450 57.900 ;
        RECT 35.070 58.040 35.360 58.085 ;
        RECT 37.170 58.040 37.460 58.085 ;
        RECT 38.740 58.040 39.030 58.085 ;
        RECT 35.070 57.900 39.030 58.040 ;
        RECT 35.070 57.855 35.360 57.900 ;
        RECT 37.170 57.855 37.460 57.900 ;
        RECT 38.740 57.855 39.030 57.900 ;
        RECT 52.510 58.040 52.800 58.085 ;
        RECT 54.080 58.040 54.370 58.085 ;
        RECT 56.180 58.040 56.470 58.085 ;
        RECT 52.510 57.900 56.470 58.040 ;
        RECT 52.510 57.855 52.800 57.900 ;
        RECT 54.080 57.855 54.370 57.900 ;
        RECT 56.180 57.855 56.470 57.900 ;
        RECT 69.530 58.040 69.850 58.100 ;
        RECT 78.360 58.040 78.500 58.195 ;
        RECT 69.530 57.900 78.500 58.040 ;
        RECT 69.530 57.840 69.850 57.900 ;
        RECT 81.950 57.840 82.270 58.100 ;
        RECT 19.850 57.700 20.170 57.760 ;
        RECT 23.545 57.700 23.835 57.745 ;
        RECT 27.670 57.700 27.990 57.760 ;
        RECT 13.730 57.560 27.990 57.700 ;
        RECT 10.205 57.515 10.495 57.560 ;
        RECT 10.650 57.500 10.970 57.560 ;
        RECT 19.850 57.500 20.170 57.560 ;
        RECT 23.545 57.515 23.835 57.560 ;
        RECT 27.670 57.500 27.990 57.560 ;
        RECT 61.265 57.700 61.555 57.745 ;
        RECT 62.170 57.700 62.490 57.760 ;
        RECT 61.265 57.560 62.490 57.700 ;
        RECT 61.265 57.515 61.555 57.560 ;
        RECT 62.170 57.500 62.490 57.560 ;
        RECT 65.850 57.700 66.170 57.760 ;
        RECT 72.750 57.700 73.070 57.760 ;
        RECT 65.850 57.560 73.070 57.700 ;
        RECT 65.850 57.500 66.170 57.560 ;
        RECT 72.750 57.500 73.070 57.560 ;
        RECT 75.510 57.500 75.830 57.760 ;
        RECT 5.520 56.880 84.180 57.360 ;
        RECT 5.590 56.680 5.910 56.740 ;
        RECT 7.445 56.680 7.735 56.725 ;
        RECT 5.590 56.540 7.735 56.680 ;
        RECT 5.590 56.480 5.910 56.540 ;
        RECT 7.445 56.495 7.735 56.540 ;
        RECT 14.790 56.680 15.110 56.740 ;
        RECT 18.470 56.680 18.790 56.740 ;
        RECT 14.790 56.540 18.790 56.680 ;
        RECT 14.790 56.480 15.110 56.540 ;
        RECT 18.470 56.480 18.790 56.540 ;
        RECT 20.310 56.680 20.630 56.740 ;
        RECT 20.785 56.680 21.075 56.725 ;
        RECT 20.310 56.540 21.075 56.680 ;
        RECT 20.310 56.480 20.630 56.540 ;
        RECT 20.785 56.495 21.075 56.540 ;
        RECT 24.925 56.680 25.215 56.725 ;
        RECT 25.370 56.680 25.690 56.740 ;
        RECT 24.925 56.540 25.690 56.680 ;
        RECT 24.925 56.495 25.215 56.540 ;
        RECT 25.370 56.480 25.690 56.540 ;
        RECT 34.585 56.680 34.875 56.725 ;
        RECT 35.030 56.680 35.350 56.740 ;
        RECT 34.585 56.540 35.350 56.680 ;
        RECT 34.585 56.495 34.875 56.540 ;
        RECT 35.030 56.480 35.350 56.540 ;
        RECT 41.930 56.680 42.250 56.740 ;
        RECT 42.865 56.680 43.155 56.725 ;
        RECT 41.930 56.540 43.155 56.680 ;
        RECT 41.930 56.480 42.250 56.540 ;
        RECT 42.865 56.495 43.155 56.540 ;
        RECT 48.385 56.680 48.675 56.725 ;
        RECT 49.750 56.680 50.070 56.740 ;
        RECT 48.385 56.540 50.070 56.680 ;
        RECT 48.385 56.495 48.675 56.540 ;
        RECT 49.750 56.480 50.070 56.540 ;
        RECT 58.950 56.680 59.270 56.740 ;
        RECT 64.470 56.680 64.790 56.740 ;
        RECT 58.950 56.540 64.790 56.680 ;
        RECT 58.950 56.480 59.270 56.540 ;
        RECT 64.470 56.480 64.790 56.540 ;
        RECT 64.930 56.680 65.250 56.740 ;
        RECT 69.070 56.680 69.390 56.740 ;
        RECT 64.930 56.540 69.390 56.680 ;
        RECT 64.930 56.480 65.250 56.540 ;
        RECT 69.070 56.480 69.390 56.540 ;
        RECT 69.530 56.480 69.850 56.740 ;
        RECT 73.225 56.680 73.515 56.725 ;
        RECT 77.810 56.680 78.130 56.740 ;
        RECT 73.225 56.540 78.130 56.680 ;
        RECT 73.225 56.495 73.515 56.540 ;
        RECT 77.810 56.480 78.130 56.540 ;
        RECT 80.110 56.680 80.430 56.740 ;
        RECT 81.045 56.680 81.335 56.725 ;
        RECT 80.110 56.540 81.335 56.680 ;
        RECT 80.110 56.480 80.430 56.540 ;
        RECT 81.045 56.495 81.335 56.540 ;
        RECT 9.310 56.340 9.600 56.385 ;
        RECT 11.410 56.340 11.700 56.385 ;
        RECT 12.980 56.340 13.270 56.385 ;
        RECT 9.310 56.200 13.270 56.340 ;
        RECT 9.310 56.155 9.600 56.200 ;
        RECT 11.410 56.155 11.700 56.200 ;
        RECT 12.980 56.155 13.270 56.200 ;
        RECT 14.330 56.340 14.650 56.400 ;
        RECT 15.725 56.340 16.015 56.385 ;
        RECT 17.090 56.340 17.410 56.400 ;
        RECT 23.070 56.340 23.390 56.400 ;
        RECT 14.330 56.200 17.410 56.340 ;
        RECT 14.330 56.140 14.650 56.200 ;
        RECT 15.725 56.155 16.015 56.200 ;
        RECT 17.090 56.140 17.410 56.200 ;
        RECT 22.140 56.200 23.390 56.340 ;
        RECT 9.705 56.000 9.995 56.045 ;
        RECT 10.895 56.000 11.185 56.045 ;
        RECT 13.415 56.000 13.705 56.045 ;
        RECT 9.705 55.860 13.705 56.000 ;
        RECT 9.705 55.815 9.995 55.860 ;
        RECT 10.895 55.815 11.185 55.860 ;
        RECT 13.415 55.815 13.705 55.860 ;
        RECT 8.365 55.475 8.655 55.705 ;
        RECT 8.440 55.320 8.580 55.475 ;
        RECT 8.810 55.460 9.130 55.720 ;
        RECT 14.330 55.660 14.650 55.720 ;
        RECT 9.820 55.520 14.650 55.660 ;
        RECT 9.820 55.320 9.960 55.520 ;
        RECT 14.330 55.460 14.650 55.520 ;
        RECT 18.930 55.460 19.250 55.720 ;
        RECT 19.850 55.460 20.170 55.720 ;
        RECT 21.705 55.660 21.995 55.705 ;
        RECT 22.140 55.660 22.280 56.200 ;
        RECT 23.070 56.140 23.390 56.200 ;
        RECT 27.710 56.340 28.000 56.385 ;
        RECT 29.810 56.340 30.100 56.385 ;
        RECT 31.380 56.340 31.670 56.385 ;
        RECT 27.710 56.200 31.670 56.340 ;
        RECT 27.710 56.155 28.000 56.200 ;
        RECT 29.810 56.155 30.100 56.200 ;
        RECT 31.380 56.155 31.670 56.200 ;
        RECT 32.730 56.340 33.050 56.400 ;
        RECT 57.570 56.340 57.890 56.400 ;
        RECT 65.390 56.340 65.710 56.400 ;
        RECT 74.630 56.340 74.920 56.385 ;
        RECT 76.730 56.340 77.020 56.385 ;
        RECT 78.300 56.340 78.590 56.385 ;
        RECT 32.730 56.200 60.560 56.340 ;
        RECT 32.730 56.140 33.050 56.200 ;
        RECT 57.570 56.140 57.890 56.200 ;
        RECT 23.990 56.000 24.310 56.060 ;
        RECT 22.700 55.860 24.310 56.000 ;
        RECT 22.700 55.705 22.840 55.860 ;
        RECT 23.990 55.800 24.310 55.860 ;
        RECT 28.105 56.000 28.395 56.045 ;
        RECT 29.295 56.000 29.585 56.045 ;
        RECT 31.815 56.000 32.105 56.045 ;
        RECT 28.105 55.860 32.105 56.000 ;
        RECT 28.105 55.815 28.395 55.860 ;
        RECT 29.295 55.815 29.585 55.860 ;
        RECT 31.815 55.815 32.105 55.860 ;
        RECT 37.805 56.000 38.095 56.045 ;
        RECT 39.630 56.000 39.950 56.060 ;
        RECT 37.805 55.860 39.950 56.000 ;
        RECT 37.805 55.815 38.095 55.860 ;
        RECT 39.630 55.800 39.950 55.860 ;
        RECT 40.565 56.000 40.855 56.045 ;
        RECT 50.210 56.000 50.530 56.060 ;
        RECT 50.685 56.000 50.975 56.045 ;
        RECT 40.565 55.860 49.980 56.000 ;
        RECT 40.565 55.815 40.855 55.860 ;
        RECT 20.355 55.520 22.280 55.660 ;
        RECT 10.190 55.365 10.510 55.380 ;
        RECT 8.440 55.180 9.960 55.320 ;
        RECT 10.160 55.135 10.510 55.365 ;
        RECT 10.190 55.120 10.510 55.135 ;
        RECT 11.110 55.320 11.430 55.380 ;
        RECT 15.250 55.320 15.570 55.380 ;
        RECT 20.355 55.320 20.495 55.520 ;
        RECT 21.705 55.475 21.995 55.520 ;
        RECT 22.625 55.475 22.915 55.705 ;
        RECT 23.085 55.475 23.375 55.705 ;
        RECT 23.545 55.660 23.835 55.705 ;
        RECT 24.450 55.660 24.770 55.720 ;
        RECT 23.545 55.520 24.770 55.660 ;
        RECT 23.545 55.475 23.835 55.520 ;
        RECT 11.110 55.180 20.495 55.320 ;
        RECT 21.230 55.320 21.550 55.380 ;
        RECT 23.160 55.320 23.300 55.475 ;
        RECT 24.450 55.460 24.770 55.520 ;
        RECT 27.225 55.660 27.515 55.705 ;
        RECT 33.190 55.660 33.510 55.720 ;
        RECT 27.225 55.520 33.510 55.660 ;
        RECT 27.225 55.475 27.515 55.520 ;
        RECT 33.190 55.460 33.510 55.520 ;
        RECT 41.025 55.660 41.315 55.705 ;
        RECT 43.310 55.660 43.630 55.720 ;
        RECT 41.025 55.520 43.630 55.660 ;
        RECT 49.840 55.660 49.980 55.860 ;
        RECT 50.210 55.860 50.975 56.000 ;
        RECT 50.210 55.800 50.530 55.860 ;
        RECT 50.685 55.815 50.975 55.860 ;
        RECT 51.605 56.000 51.895 56.045 ;
        RECT 52.510 56.000 52.830 56.060 ;
        RECT 59.870 56.000 60.190 56.060 ;
        RECT 51.605 55.860 52.830 56.000 ;
        RECT 51.605 55.815 51.895 55.860 ;
        RECT 52.510 55.800 52.830 55.860 ;
        RECT 59.500 55.860 60.190 56.000 ;
        RECT 60.420 56.000 60.560 56.200 ;
        RECT 61.340 56.200 65.710 56.340 ;
        RECT 61.340 56.000 61.480 56.200 ;
        RECT 65.390 56.140 65.710 56.200 ;
        RECT 65.940 56.200 70.680 56.340 ;
        RECT 60.420 55.860 61.480 56.000 ;
        RECT 61.725 56.000 62.015 56.045 ;
        RECT 65.940 56.000 66.080 56.200 ;
        RECT 61.725 55.860 66.080 56.000 ;
        RECT 66.310 56.000 66.630 56.060 ;
        RECT 67.245 56.000 67.535 56.045 ;
        RECT 66.310 55.860 67.535 56.000 ;
        RECT 56.650 55.660 56.970 55.720 ;
        RECT 49.840 55.520 56.970 55.660 ;
        RECT 41.025 55.475 41.315 55.520 ;
        RECT 43.310 55.460 43.630 55.520 ;
        RECT 56.650 55.460 56.970 55.520 ;
        RECT 58.950 55.460 59.270 55.720 ;
        RECT 59.500 55.705 59.640 55.860 ;
        RECT 59.870 55.800 60.190 55.860 ;
        RECT 61.725 55.815 62.015 55.860 ;
        RECT 66.310 55.800 66.630 55.860 ;
        RECT 67.245 55.815 67.535 55.860 ;
        RECT 67.690 55.800 68.010 56.060 ;
        RECT 59.425 55.475 59.715 55.705 ;
        RECT 60.790 55.460 61.110 55.720 ;
        RECT 61.250 55.460 61.570 55.720 ;
        RECT 62.185 55.660 62.475 55.705 ;
        RECT 62.630 55.660 62.950 55.720 ;
        RECT 62.185 55.520 62.950 55.660 ;
        RECT 62.185 55.475 62.475 55.520 ;
        RECT 21.230 55.180 23.300 55.320 ;
        RECT 28.560 55.320 28.850 55.365 ;
        RECT 31.350 55.320 31.670 55.380 ;
        RECT 28.560 55.180 31.670 55.320 ;
        RECT 11.110 55.120 11.430 55.180 ;
        RECT 15.250 55.120 15.570 55.180 ;
        RECT 21.230 55.120 21.550 55.180 ;
        RECT 28.560 55.135 28.850 55.180 ;
        RECT 31.350 55.120 31.670 55.180 ;
        RECT 36.885 55.320 37.175 55.365 ;
        RECT 47.450 55.320 47.770 55.380 ;
        RECT 36.885 55.180 47.770 55.320 ;
        RECT 36.885 55.135 37.175 55.180 ;
        RECT 47.450 55.120 47.770 55.180 ;
        RECT 59.870 55.120 60.190 55.380 ;
        RECT 11.570 54.980 11.890 55.040 ;
        RECT 13.410 54.980 13.730 55.040 ;
        RECT 11.570 54.840 13.730 54.980 ;
        RECT 11.570 54.780 11.890 54.840 ;
        RECT 13.410 54.780 13.730 54.840 ;
        RECT 20.770 54.980 21.090 55.040 ;
        RECT 23.530 54.980 23.850 55.040 ;
        RECT 20.770 54.840 23.850 54.980 ;
        RECT 20.770 54.780 21.090 54.840 ;
        RECT 23.530 54.780 23.850 54.840 ;
        RECT 34.125 54.980 34.415 55.025 ;
        RECT 36.410 54.980 36.730 55.040 ;
        RECT 34.125 54.840 36.730 54.980 ;
        RECT 34.125 54.795 34.415 54.840 ;
        RECT 36.410 54.780 36.730 54.840 ;
        RECT 50.225 54.980 50.515 55.025 ;
        RECT 52.510 54.980 52.830 55.040 ;
        RECT 50.225 54.840 52.830 54.980 ;
        RECT 50.225 54.795 50.515 54.840 ;
        RECT 52.510 54.780 52.830 54.840 ;
        RECT 58.045 54.980 58.335 55.025 ;
        RECT 58.490 54.980 58.810 55.040 ;
        RECT 58.045 54.840 58.810 54.980 ;
        RECT 58.045 54.795 58.335 54.840 ;
        RECT 58.490 54.780 58.810 54.840 ;
        RECT 61.250 54.980 61.570 55.040 ;
        RECT 62.260 54.980 62.400 55.475 ;
        RECT 62.630 55.460 62.950 55.520 ;
        RECT 63.090 55.460 63.410 55.720 ;
        RECT 63.550 55.460 63.870 55.720 ;
        RECT 64.025 55.475 64.315 55.705 ;
        RECT 63.180 55.320 63.320 55.460 ;
        RECT 64.100 55.320 64.240 55.475 ;
        RECT 64.470 55.460 64.790 55.720 ;
        RECT 64.930 55.460 65.250 55.720 ;
        RECT 65.850 55.460 66.170 55.720 ;
        RECT 66.785 55.660 67.075 55.705 ;
        RECT 68.150 55.660 68.470 55.720 ;
        RECT 66.785 55.520 68.470 55.660 ;
        RECT 66.785 55.475 67.075 55.520 ;
        RECT 68.150 55.460 68.470 55.520 ;
        RECT 68.610 55.460 68.930 55.720 ;
        RECT 70.540 55.705 70.680 56.200 ;
        RECT 74.630 56.200 78.590 56.340 ;
        RECT 74.630 56.155 74.920 56.200 ;
        RECT 76.730 56.155 77.020 56.200 ;
        RECT 78.300 56.155 78.590 56.200 ;
        RECT 73.670 56.000 73.990 56.060 ;
        RECT 74.145 56.000 74.435 56.045 ;
        RECT 73.670 55.860 74.435 56.000 ;
        RECT 73.670 55.800 73.990 55.860 ;
        RECT 74.145 55.815 74.435 55.860 ;
        RECT 75.025 56.000 75.315 56.045 ;
        RECT 76.215 56.000 76.505 56.045 ;
        RECT 78.735 56.000 79.025 56.045 ;
        RECT 75.025 55.860 79.025 56.000 ;
        RECT 75.025 55.815 75.315 55.860 ;
        RECT 76.215 55.815 76.505 55.860 ;
        RECT 78.735 55.815 79.025 55.860 ;
        RECT 70.465 55.475 70.755 55.705 ;
        RECT 70.910 55.660 71.230 55.720 ;
        RECT 71.385 55.660 71.675 55.705 ;
        RECT 70.910 55.520 71.675 55.660 ;
        RECT 70.910 55.460 71.230 55.520 ;
        RECT 71.385 55.475 71.675 55.520 ;
        RECT 72.290 55.460 72.610 55.720 ;
        RECT 75.510 55.705 75.830 55.720 ;
        RECT 75.480 55.660 75.830 55.705 ;
        RECT 75.315 55.520 75.830 55.660 ;
        RECT 81.120 55.660 81.260 56.495 ;
        RECT 81.490 56.480 81.810 56.740 ;
        RECT 82.425 55.660 82.715 55.705 ;
        RECT 81.120 55.520 82.715 55.660 ;
        RECT 75.480 55.475 75.830 55.520 ;
        RECT 82.425 55.475 82.715 55.520 ;
        RECT 75.510 55.460 75.830 55.475 ;
        RECT 63.180 55.180 64.240 55.320 ;
        RECT 65.390 55.320 65.710 55.380 ;
        RECT 71.845 55.320 72.135 55.365 ;
        RECT 65.390 55.180 72.135 55.320 ;
        RECT 65.390 55.120 65.710 55.180 ;
        RECT 71.845 55.135 72.135 55.180 ;
        RECT 61.250 54.840 62.400 54.980 ;
        RECT 62.645 54.980 62.935 55.025 ;
        RECT 63.090 54.980 63.410 55.040 ;
        RECT 62.645 54.840 63.410 54.980 ;
        RECT 61.250 54.780 61.570 54.840 ;
        RECT 62.645 54.795 62.935 54.840 ;
        RECT 63.090 54.780 63.410 54.840 ;
        RECT 63.550 54.980 63.870 55.040 ;
        RECT 68.150 54.980 68.470 55.040 ;
        RECT 63.550 54.840 68.470 54.980 ;
        RECT 63.550 54.780 63.870 54.840 ;
        RECT 68.150 54.780 68.470 54.840 ;
        RECT 5.520 54.160 84.180 54.640 ;
        RECT 8.365 53.960 8.655 54.005 ;
        RECT 10.190 53.960 10.510 54.020 ;
        RECT 8.365 53.820 10.510 53.960 ;
        RECT 8.365 53.775 8.655 53.820 ;
        RECT 10.190 53.760 10.510 53.820 ;
        RECT 13.870 53.960 14.190 54.020 ;
        RECT 18.485 53.960 18.775 54.005 ;
        RECT 29.050 53.960 29.370 54.020 ;
        RECT 13.870 53.820 18.240 53.960 ;
        RECT 13.870 53.760 14.190 53.820 ;
        RECT 12.950 53.620 13.270 53.680 ;
        RECT 10.280 53.480 13.270 53.620 ;
        RECT 18.100 53.620 18.240 53.820 ;
        RECT 18.485 53.820 29.370 53.960 ;
        RECT 18.485 53.775 18.775 53.820 ;
        RECT 29.050 53.760 29.370 53.820 ;
        RECT 31.350 53.960 31.670 54.020 ;
        RECT 31.825 53.960 32.115 54.005 ;
        RECT 31.350 53.820 32.115 53.960 ;
        RECT 31.350 53.760 31.670 53.820 ;
        RECT 31.825 53.775 32.115 53.820 ;
        RECT 39.170 53.960 39.490 54.020 ;
        RECT 39.645 53.960 39.935 54.005 ;
        RECT 39.170 53.820 39.935 53.960 ;
        RECT 39.170 53.760 39.490 53.820 ;
        RECT 39.645 53.775 39.935 53.820 ;
        RECT 60.790 53.760 61.110 54.020 ;
        RECT 64.470 53.960 64.790 54.020 ;
        RECT 61.800 53.820 62.400 53.960 ;
        RECT 19.390 53.620 19.710 53.680 ;
        RECT 21.230 53.620 21.550 53.680 ;
        RECT 18.100 53.480 21.550 53.620 ;
        RECT 10.280 53.325 10.420 53.480 ;
        RECT 12.950 53.420 13.270 53.480 ;
        RECT 19.390 53.420 19.710 53.480 ;
        RECT 9.745 53.095 10.035 53.325 ;
        RECT 10.205 53.095 10.495 53.325 ;
        RECT 9.820 52.600 9.960 53.095 ;
        RECT 10.650 53.080 10.970 53.340 ;
        RECT 11.110 53.280 11.430 53.340 ;
        RECT 11.585 53.280 11.875 53.325 ;
        RECT 11.110 53.140 11.875 53.280 ;
        RECT 11.110 53.080 11.430 53.140 ;
        RECT 11.585 53.095 11.875 53.140 ;
        RECT 12.030 53.280 12.350 53.340 ;
        RECT 12.030 53.230 12.720 53.280 ;
        RECT 13.425 53.230 13.715 53.325 ;
        RECT 12.030 53.140 13.715 53.230 ;
        RECT 12.030 53.080 12.350 53.140 ;
        RECT 12.580 53.095 13.715 53.140 ;
        RECT 12.580 53.090 13.640 53.095 ;
        RECT 13.855 53.080 14.175 53.340 ;
        RECT 14.450 53.310 14.740 53.355 ;
        RECT 14.450 53.170 15.020 53.310 ;
        RECT 14.450 53.125 14.740 53.170 ;
        RECT 14.880 52.660 15.020 53.170 ;
        RECT 15.250 53.080 15.570 53.340 ;
        RECT 15.725 53.095 16.015 53.325 ;
        RECT 16.185 53.280 16.475 53.325 ;
        RECT 16.630 53.280 16.950 53.340 ;
        RECT 16.185 53.140 16.950 53.280 ;
        RECT 16.185 53.095 16.475 53.140 ;
        RECT 9.820 52.460 12.720 52.600 ;
        RECT 12.580 52.320 12.720 52.460 ;
        RECT 14.790 52.400 15.110 52.660 ;
        RECT 15.800 52.600 15.940 53.095 ;
        RECT 16.630 53.080 16.950 53.140 ;
        RECT 17.090 53.080 17.410 53.340 ;
        RECT 17.550 53.080 17.870 53.340 ;
        RECT 18.470 53.280 18.790 53.340 ;
        RECT 20.400 53.325 20.540 53.480 ;
        RECT 21.230 53.420 21.550 53.480 ;
        RECT 22.165 53.620 22.455 53.665 ;
        RECT 23.850 53.620 24.140 53.665 ;
        RECT 22.165 53.480 24.140 53.620 ;
        RECT 22.165 53.435 22.455 53.480 ;
        RECT 23.850 53.435 24.140 53.480 ;
        RECT 27.670 53.620 27.990 53.680 ;
        RECT 47.450 53.620 47.770 53.680 ;
        RECT 61.800 53.665 61.940 53.820 ;
        RECT 27.670 53.480 41.240 53.620 ;
        RECT 27.670 53.420 27.990 53.480 ;
        RECT 18.945 53.280 19.235 53.325 ;
        RECT 18.470 53.140 19.235 53.280 ;
        RECT 18.470 53.080 18.790 53.140 ;
        RECT 18.945 53.095 19.235 53.140 ;
        RECT 19.865 53.095 20.155 53.325 ;
        RECT 20.325 53.095 20.615 53.325 ;
        RECT 17.090 52.600 17.410 52.660 ;
        RECT 15.800 52.460 17.410 52.600 ;
        RECT 17.090 52.400 17.410 52.460 ;
        RECT 12.030 52.060 12.350 52.320 ;
        RECT 12.490 52.260 12.810 52.320 ;
        RECT 16.170 52.260 16.490 52.320 ;
        RECT 12.490 52.120 16.490 52.260 ;
        RECT 19.940 52.260 20.080 53.095 ;
        RECT 20.770 53.080 21.090 53.340 ;
        RECT 22.625 53.280 22.915 53.325 ;
        RECT 23.070 53.280 23.390 53.340 ;
        RECT 22.625 53.140 23.390 53.280 ;
        RECT 22.625 53.095 22.915 53.140 ;
        RECT 23.070 53.080 23.390 53.140 ;
        RECT 33.665 53.280 33.955 53.325 ;
        RECT 35.965 53.280 36.255 53.325 ;
        RECT 33.665 53.140 36.255 53.280 ;
        RECT 33.665 53.095 33.955 53.140 ;
        RECT 35.965 53.095 36.255 53.140 ;
        RECT 36.410 53.280 36.730 53.340 ;
        RECT 38.725 53.280 39.015 53.325 ;
        RECT 36.410 53.140 39.015 53.280 ;
        RECT 36.410 53.080 36.730 53.140 ;
        RECT 38.725 53.095 39.015 53.140 ;
        RECT 40.550 53.080 40.870 53.340 ;
        RECT 41.100 53.325 41.240 53.480 ;
        RECT 47.450 53.480 57.800 53.620 ;
        RECT 47.450 53.420 47.770 53.480 ;
        RECT 41.025 53.095 41.315 53.325 ;
        RECT 41.945 53.095 42.235 53.325 ;
        RECT 23.505 52.940 23.795 52.985 ;
        RECT 24.695 52.940 24.985 52.985 ;
        RECT 27.215 52.940 27.505 52.985 ;
        RECT 23.505 52.800 27.505 52.940 ;
        RECT 23.505 52.755 23.795 52.800 ;
        RECT 24.695 52.755 24.985 52.800 ;
        RECT 27.215 52.755 27.505 52.800 ;
        RECT 34.110 52.740 34.430 53.000 ;
        RECT 35.045 52.940 35.335 52.985 ;
        RECT 41.470 52.940 41.790 53.000 ;
        RECT 35.045 52.800 41.790 52.940 ;
        RECT 42.020 52.940 42.160 53.095 ;
        RECT 42.390 53.080 42.710 53.340 ;
        RECT 57.660 53.325 57.800 53.480 ;
        RECT 61.725 53.435 62.015 53.665 ;
        RECT 46.545 53.280 46.835 53.325 ;
        RECT 48.845 53.280 49.135 53.325 ;
        RECT 46.545 53.140 49.135 53.280 ;
        RECT 46.545 53.095 46.835 53.140 ;
        RECT 48.845 53.095 49.135 53.140 ;
        RECT 57.585 53.095 57.875 53.325 ;
        RECT 61.250 53.080 61.570 53.340 ;
        RECT 62.260 53.280 62.400 53.820 ;
        RECT 62.720 53.820 64.790 53.960 ;
        RECT 62.720 53.665 62.860 53.820 ;
        RECT 64.470 53.760 64.790 53.820 ;
        RECT 69.990 53.760 70.310 54.020 ;
        RECT 62.645 53.435 62.935 53.665 ;
        RECT 63.105 53.620 63.395 53.665 ;
        RECT 63.550 53.620 63.870 53.680 ;
        RECT 66.310 53.620 66.630 53.680 ;
        RECT 69.070 53.620 69.390 53.680 ;
        RECT 71.830 53.620 72.150 53.680 ;
        RECT 63.105 53.480 63.870 53.620 ;
        RECT 63.105 53.435 63.395 53.480 ;
        RECT 63.550 53.420 63.870 53.480 ;
        RECT 64.560 53.480 66.630 53.620 ;
        RECT 64.010 53.280 64.330 53.340 ;
        RECT 64.560 53.325 64.700 53.480 ;
        RECT 66.310 53.420 66.630 53.480 ;
        RECT 67.320 53.480 72.150 53.620 ;
        RECT 62.260 53.140 64.330 53.280 ;
        RECT 64.010 53.080 64.330 53.140 ;
        RECT 64.485 53.095 64.775 53.325 ;
        RECT 64.930 53.280 65.250 53.340 ;
        RECT 65.865 53.280 66.155 53.325 ;
        RECT 64.930 53.140 66.155 53.280 ;
        RECT 64.930 53.080 65.250 53.140 ;
        RECT 65.865 53.095 66.155 53.140 ;
        RECT 45.610 52.940 45.930 53.000 ;
        RECT 42.020 52.800 45.930 52.940 ;
        RECT 35.045 52.755 35.335 52.800 ;
        RECT 41.470 52.740 41.790 52.800 ;
        RECT 45.610 52.740 45.930 52.800 ;
        RECT 46.990 52.740 47.310 53.000 ;
        RECT 47.910 52.740 48.230 53.000 ;
        RECT 51.130 52.940 51.450 53.000 ;
        RECT 51.605 52.940 51.895 52.985 ;
        RECT 51.130 52.800 51.895 52.940 ;
        RECT 51.130 52.740 51.450 52.800 ;
        RECT 51.605 52.755 51.895 52.800 ;
        RECT 52.510 52.940 52.830 53.000 ;
        RECT 55.745 52.940 56.035 52.985 ;
        RECT 52.510 52.800 56.035 52.940 ;
        RECT 52.510 52.740 52.830 52.800 ;
        RECT 55.745 52.755 56.035 52.800 ;
        RECT 58.030 52.940 58.350 53.000 ;
        RECT 58.030 52.800 62.170 52.940 ;
        RECT 58.030 52.740 58.350 52.800 ;
        RECT 23.110 52.600 23.400 52.645 ;
        RECT 25.210 52.600 25.500 52.645 ;
        RECT 26.780 52.600 27.070 52.645 ;
        RECT 23.110 52.460 27.070 52.600 ;
        RECT 23.110 52.415 23.400 52.460 ;
        RECT 25.210 52.415 25.500 52.460 ;
        RECT 26.780 52.415 27.070 52.460 ;
        RECT 59.870 52.600 60.190 52.660 ;
        RECT 61.265 52.600 61.555 52.645 ;
        RECT 59.870 52.460 61.555 52.600 ;
        RECT 62.030 52.600 62.170 52.800 ;
        RECT 63.090 52.740 63.410 53.000 ;
        RECT 66.325 52.940 66.615 52.985 ;
        RECT 67.320 52.940 67.460 53.480 ;
        RECT 69.070 53.420 69.390 53.480 ;
        RECT 71.830 53.420 72.150 53.480 ;
        RECT 67.705 53.095 67.995 53.325 ;
        RECT 68.165 53.280 68.455 53.325 ;
        RECT 68.610 53.280 68.930 53.340 ;
        RECT 69.545 53.280 69.835 53.325 ;
        RECT 68.165 53.140 68.930 53.280 ;
        RECT 68.165 53.095 68.455 53.140 ;
        RECT 66.325 52.800 67.460 52.940 ;
        RECT 66.325 52.755 66.615 52.800 ;
        RECT 67.780 52.600 67.920 53.095 ;
        RECT 68.610 53.080 68.930 53.140 ;
        RECT 69.160 53.140 69.835 53.280 ;
        RECT 69.160 52.645 69.300 53.140 ;
        RECT 69.545 53.095 69.835 53.140 ;
        RECT 72.765 53.280 73.055 53.325 ;
        RECT 73.210 53.280 73.530 53.340 ;
        RECT 74.130 53.325 74.450 53.340 ;
        RECT 72.765 53.140 73.530 53.280 ;
        RECT 72.765 53.095 73.055 53.140 ;
        RECT 73.210 53.080 73.530 53.140 ;
        RECT 74.100 53.095 74.450 53.325 ;
        RECT 74.130 53.080 74.450 53.095 ;
        RECT 75.970 53.280 76.290 53.340 ;
        RECT 81.045 53.280 81.335 53.325 ;
        RECT 75.970 53.140 81.335 53.280 ;
        RECT 75.970 53.080 76.290 53.140 ;
        RECT 81.045 53.095 81.335 53.140 ;
        RECT 71.845 52.940 72.135 52.985 ;
        RECT 72.290 52.940 72.610 53.000 ;
        RECT 71.845 52.800 72.610 52.940 ;
        RECT 71.845 52.755 72.135 52.800 ;
        RECT 72.290 52.740 72.610 52.800 ;
        RECT 73.645 52.940 73.935 52.985 ;
        RECT 74.835 52.940 75.125 52.985 ;
        RECT 77.355 52.940 77.645 52.985 ;
        RECT 73.645 52.800 77.645 52.940 ;
        RECT 73.645 52.755 73.935 52.800 ;
        RECT 74.835 52.755 75.125 52.800 ;
        RECT 77.355 52.755 77.645 52.800 ;
        RECT 62.030 52.460 67.920 52.600 ;
        RECT 59.870 52.400 60.190 52.460 ;
        RECT 61.265 52.415 61.555 52.460 ;
        RECT 69.085 52.415 69.375 52.645 ;
        RECT 73.250 52.600 73.540 52.645 ;
        RECT 75.350 52.600 75.640 52.645 ;
        RECT 76.920 52.600 77.210 52.645 ;
        RECT 73.250 52.460 77.210 52.600 ;
        RECT 73.250 52.415 73.540 52.460 ;
        RECT 75.350 52.415 75.640 52.460 ;
        RECT 76.920 52.415 77.210 52.460 ;
        RECT 23.530 52.260 23.850 52.320 ;
        RECT 19.940 52.120 23.850 52.260 ;
        RECT 12.490 52.060 12.810 52.120 ;
        RECT 16.170 52.060 16.490 52.120 ;
        RECT 23.530 52.060 23.850 52.120 ;
        RECT 27.210 52.260 27.530 52.320 ;
        RECT 29.525 52.260 29.815 52.305 ;
        RECT 27.210 52.120 29.815 52.260 ;
        RECT 27.210 52.060 27.530 52.120 ;
        RECT 29.525 52.075 29.815 52.120 ;
        RECT 44.690 52.060 45.010 52.320 ;
        RECT 52.970 52.060 53.290 52.320 ;
        RECT 62.170 52.260 62.490 52.320 ;
        RECT 64.025 52.260 64.315 52.305 ;
        RECT 67.690 52.260 68.010 52.320 ;
        RECT 62.170 52.120 68.010 52.260 ;
        RECT 62.170 52.060 62.490 52.120 ;
        RECT 64.025 52.075 64.315 52.120 ;
        RECT 67.690 52.060 68.010 52.120 ;
        RECT 70.925 52.260 71.215 52.305 ;
        RECT 77.350 52.260 77.670 52.320 ;
        RECT 70.925 52.120 77.670 52.260 ;
        RECT 70.925 52.075 71.215 52.120 ;
        RECT 77.350 52.060 77.670 52.120 ;
        RECT 79.650 52.060 79.970 52.320 ;
        RECT 81.950 52.060 82.270 52.320 ;
        RECT 5.520 51.440 84.180 51.920 ;
        RECT 8.825 51.240 9.115 51.285 ;
        RECT 14.790 51.240 15.110 51.300 ;
        RECT 26.765 51.240 27.055 51.285 ;
        RECT 34.110 51.240 34.430 51.300 ;
        RECT 8.825 51.100 15.110 51.240 ;
        RECT 8.825 51.055 9.115 51.100 ;
        RECT 14.790 51.040 15.110 51.100 ;
        RECT 24.080 51.100 26.520 51.240 ;
        RECT 9.770 50.900 10.060 50.945 ;
        RECT 11.870 50.900 12.160 50.945 ;
        RECT 13.440 50.900 13.730 50.945 ;
        RECT 9.770 50.760 13.730 50.900 ;
        RECT 9.770 50.715 10.060 50.760 ;
        RECT 11.870 50.715 12.160 50.760 ;
        RECT 13.440 50.715 13.730 50.760 ;
        RECT 8.810 50.560 9.130 50.620 ;
        RECT 9.285 50.560 9.575 50.605 ;
        RECT 8.810 50.420 9.575 50.560 ;
        RECT 8.810 50.360 9.130 50.420 ;
        RECT 9.285 50.375 9.575 50.420 ;
        RECT 10.165 50.560 10.455 50.605 ;
        RECT 11.355 50.560 11.645 50.605 ;
        RECT 13.875 50.560 14.165 50.605 ;
        RECT 10.165 50.420 14.165 50.560 ;
        RECT 10.165 50.375 10.455 50.420 ;
        RECT 11.355 50.375 11.645 50.420 ;
        RECT 13.875 50.375 14.165 50.420 ;
        RECT 9.360 50.220 9.500 50.375 ;
        RECT 17.550 50.220 17.870 50.280 ;
        RECT 24.080 50.265 24.220 51.100 ;
        RECT 26.380 50.560 26.520 51.100 ;
        RECT 26.765 51.100 34.430 51.240 ;
        RECT 26.765 51.055 27.055 51.100 ;
        RECT 34.110 51.040 34.430 51.100 ;
        RECT 41.025 51.240 41.315 51.285 ;
        RECT 46.990 51.240 47.310 51.300 ;
        RECT 41.025 51.100 47.310 51.240 ;
        RECT 41.025 51.055 41.315 51.100 ;
        RECT 46.990 51.040 47.310 51.100 ;
        RECT 47.450 51.240 47.770 51.300 ;
        RECT 47.450 51.100 50.440 51.240 ;
        RECT 47.450 51.040 47.770 51.100 ;
        RECT 46.110 50.900 46.400 50.945 ;
        RECT 48.210 50.900 48.500 50.945 ;
        RECT 49.780 50.900 50.070 50.945 ;
        RECT 46.110 50.760 50.070 50.900 ;
        RECT 50.300 50.900 50.440 51.100 ;
        RECT 52.510 51.040 52.830 51.300 ;
        RECT 56.650 51.240 56.970 51.300 ;
        RECT 60.345 51.240 60.635 51.285 ;
        RECT 74.130 51.240 74.450 51.300 ;
        RECT 74.605 51.240 74.895 51.285 ;
        RECT 56.650 51.100 73.900 51.240 ;
        RECT 56.650 51.040 56.970 51.100 ;
        RECT 60.345 51.055 60.635 51.100 ;
        RECT 52.985 50.900 53.275 50.945 ;
        RECT 50.300 50.760 53.275 50.900 ;
        RECT 46.110 50.715 46.400 50.760 ;
        RECT 48.210 50.715 48.500 50.760 ;
        RECT 49.780 50.715 50.070 50.760 ;
        RECT 52.985 50.715 53.275 50.760 ;
        RECT 55.730 50.900 56.020 50.945 ;
        RECT 57.300 50.900 57.590 50.945 ;
        RECT 59.400 50.900 59.690 50.945 ;
        RECT 55.730 50.760 59.690 50.900 ;
        RECT 55.730 50.715 56.020 50.760 ;
        RECT 57.300 50.715 57.590 50.760 ;
        RECT 59.400 50.715 59.690 50.760 ;
        RECT 63.090 50.900 63.380 50.945 ;
        RECT 64.660 50.900 64.950 50.945 ;
        RECT 66.760 50.900 67.050 50.945 ;
        RECT 63.090 50.760 67.050 50.900 ;
        RECT 63.090 50.715 63.380 50.760 ;
        RECT 64.660 50.715 64.950 50.760 ;
        RECT 66.760 50.715 67.050 50.760 ;
        RECT 68.150 50.700 68.470 50.960 ;
        RECT 73.210 50.700 73.530 50.960 ;
        RECT 46.505 50.560 46.795 50.605 ;
        RECT 47.695 50.560 47.985 50.605 ;
        RECT 50.215 50.560 50.505 50.605 ;
        RECT 25.000 50.420 26.060 50.560 ;
        RECT 26.380 50.420 46.300 50.560 ;
        RECT 9.360 50.080 13.870 50.220 ;
        RECT 6.970 49.680 7.290 49.940 ;
        RECT 7.905 49.695 8.195 49.925 ;
        RECT 10.620 49.880 10.910 49.925 ;
        RECT 12.030 49.880 12.350 49.940 ;
        RECT 10.620 49.740 12.350 49.880 ;
        RECT 13.730 49.880 13.870 50.080 ;
        RECT 17.550 50.080 23.760 50.220 ;
        RECT 17.550 50.020 17.870 50.080 ;
        RECT 18.945 49.880 19.235 49.925 ;
        RECT 20.770 49.880 21.090 49.940 ;
        RECT 13.730 49.740 21.090 49.880 ;
        RECT 23.620 49.880 23.760 50.080 ;
        RECT 24.005 50.035 24.295 50.265 ;
        RECT 24.450 50.020 24.770 50.280 ;
        RECT 25.000 49.880 25.140 50.420 ;
        RECT 25.920 50.265 26.060 50.420 ;
        RECT 25.385 50.035 25.675 50.265 ;
        RECT 25.845 50.220 26.135 50.265 ;
        RECT 40.550 50.220 40.870 50.280 ;
        RECT 41.930 50.220 42.250 50.280 ;
        RECT 25.845 50.080 42.250 50.220 ;
        RECT 25.845 50.035 26.135 50.080 ;
        RECT 23.620 49.740 25.140 49.880 ;
        RECT 10.620 49.695 10.910 49.740 ;
        RECT 7.980 49.540 8.120 49.695 ;
        RECT 12.030 49.680 12.350 49.740 ;
        RECT 18.945 49.695 19.235 49.740 ;
        RECT 20.770 49.680 21.090 49.740 ;
        RECT 8.350 49.540 8.670 49.600 ;
        RECT 16.185 49.540 16.475 49.585 ;
        RECT 25.460 49.540 25.600 50.035 ;
        RECT 40.550 50.020 40.870 50.080 ;
        RECT 41.930 50.020 42.250 50.080 ;
        RECT 42.405 50.035 42.695 50.265 ;
        RECT 43.325 50.035 43.615 50.265 ;
        RECT 26.750 49.880 27.070 49.940 ;
        RECT 42.480 49.880 42.620 50.035 ;
        RECT 26.750 49.740 42.620 49.880 ;
        RECT 26.750 49.680 27.070 49.740 ;
        RECT 7.980 49.400 25.600 49.540 ;
        RECT 43.400 49.540 43.540 50.035 ;
        RECT 43.770 50.020 44.090 50.280 ;
        RECT 45.625 50.035 45.915 50.265 ;
        RECT 46.160 50.220 46.300 50.420 ;
        RECT 46.505 50.420 50.505 50.560 ;
        RECT 46.505 50.375 46.795 50.420 ;
        RECT 47.695 50.375 47.985 50.420 ;
        RECT 50.215 50.375 50.505 50.420 ;
        RECT 55.295 50.560 55.585 50.605 ;
        RECT 57.815 50.560 58.105 50.605 ;
        RECT 59.005 50.560 59.295 50.605 ;
        RECT 55.295 50.420 59.295 50.560 ;
        RECT 55.295 50.375 55.585 50.420 ;
        RECT 57.815 50.375 58.105 50.420 ;
        RECT 59.005 50.375 59.295 50.420 ;
        RECT 62.655 50.560 62.945 50.605 ;
        RECT 65.175 50.560 65.465 50.605 ;
        RECT 66.365 50.560 66.655 50.605 ;
        RECT 62.655 50.420 66.655 50.560 ;
        RECT 62.655 50.375 62.945 50.420 ;
        RECT 65.175 50.375 65.465 50.420 ;
        RECT 66.365 50.375 66.655 50.420 ;
        RECT 67.245 50.560 67.535 50.605 ;
        RECT 73.300 50.560 73.440 50.700 ;
        RECT 73.760 50.605 73.900 51.100 ;
        RECT 74.130 51.100 74.895 51.240 ;
        RECT 74.130 51.040 74.450 51.100 ;
        RECT 74.605 51.055 74.895 51.100 ;
        RECT 67.245 50.420 73.440 50.560 ;
        RECT 67.245 50.375 67.535 50.420 ;
        RECT 73.685 50.375 73.975 50.605 ;
        RECT 53.430 50.220 53.750 50.280 ;
        RECT 46.160 50.080 53.750 50.220 ;
        RECT 45.700 49.880 45.840 50.035 ;
        RECT 53.430 50.020 53.750 50.080 ;
        RECT 58.490 50.265 58.810 50.280 ;
        RECT 58.490 50.220 58.840 50.265 ;
        RECT 59.885 50.220 60.175 50.265 ;
        RECT 67.320 50.220 67.460 50.375 ;
        RECT 76.890 50.360 77.210 50.620 ;
        RECT 77.350 50.360 77.670 50.620 ;
        RECT 79.650 50.560 79.970 50.620 ;
        RECT 81.505 50.560 81.795 50.605 ;
        RECT 82.410 50.560 82.730 50.620 ;
        RECT 79.650 50.420 82.730 50.560 ;
        RECT 79.650 50.360 79.970 50.420 ;
        RECT 81.505 50.375 81.795 50.420 ;
        RECT 82.410 50.360 82.730 50.420 ;
        RECT 58.490 50.080 59.005 50.220 ;
        RECT 59.885 50.080 67.460 50.220 ;
        RECT 58.490 50.035 58.840 50.080 ;
        RECT 59.885 50.035 60.175 50.080 ;
        RECT 58.490 50.020 58.810 50.035 ;
        RECT 67.690 50.020 68.010 50.280 ;
        RECT 68.625 50.220 68.915 50.265 ;
        RECT 69.070 50.220 69.390 50.280 ;
        RECT 68.625 50.080 69.390 50.220 ;
        RECT 68.625 50.035 68.915 50.080 ;
        RECT 69.070 50.020 69.390 50.080 ;
        RECT 46.070 49.880 46.390 49.940 ;
        RECT 45.700 49.740 46.390 49.880 ;
        RECT 46.070 49.680 46.390 49.740 ;
        RECT 46.960 49.880 47.250 49.925 ;
        RECT 50.670 49.880 50.990 49.940 ;
        RECT 46.960 49.740 50.990 49.880 ;
        RECT 46.960 49.695 47.250 49.740 ;
        RECT 50.670 49.680 50.990 49.740 ;
        RECT 63.550 49.880 63.870 49.940 ;
        RECT 65.910 49.880 66.200 49.925 ;
        RECT 63.550 49.740 66.200 49.880 ;
        RECT 63.550 49.680 63.870 49.740 ;
        RECT 65.910 49.695 66.200 49.740 ;
        RECT 54.350 49.540 54.670 49.600 ;
        RECT 43.400 49.400 54.670 49.540 ;
        RECT 8.350 49.340 8.670 49.400 ;
        RECT 16.185 49.355 16.475 49.400 ;
        RECT 54.350 49.340 54.670 49.400 ;
        RECT 70.450 49.340 70.770 49.600 ;
        RECT 76.445 49.540 76.735 49.585 ;
        RECT 78.745 49.540 79.035 49.585 ;
        RECT 76.445 49.400 79.035 49.540 ;
        RECT 76.445 49.355 76.735 49.400 ;
        RECT 78.745 49.355 79.035 49.400 ;
        RECT 5.520 48.720 84.180 49.200 ;
        RECT 20.310 48.520 20.630 48.580 ;
        RECT 25.370 48.520 25.690 48.580 ;
        RECT 20.310 48.380 25.690 48.520 ;
        RECT 20.310 48.320 20.630 48.380 ;
        RECT 25.370 48.320 25.690 48.380 ;
        RECT 25.830 48.520 26.150 48.580 ;
        RECT 28.130 48.520 28.450 48.580 ;
        RECT 25.830 48.380 28.450 48.520 ;
        RECT 25.830 48.320 26.150 48.380 ;
        RECT 28.130 48.320 28.450 48.380 ;
        RECT 50.670 48.320 50.990 48.580 ;
        RECT 52.525 48.520 52.815 48.565 ;
        RECT 52.970 48.520 53.290 48.580 ;
        RECT 52.525 48.380 53.290 48.520 ;
        RECT 52.525 48.335 52.815 48.380 ;
        RECT 52.970 48.320 53.290 48.380 ;
        RECT 53.430 48.520 53.750 48.580 ;
        RECT 69.990 48.520 70.310 48.580 ;
        RECT 53.430 48.380 70.310 48.520 ;
        RECT 53.430 48.320 53.750 48.380 ;
        RECT 69.990 48.320 70.310 48.380 ;
        RECT 16.645 48.180 16.935 48.225 ;
        RECT 18.930 48.180 19.250 48.240 ;
        RECT 16.645 48.040 19.250 48.180 ;
        RECT 16.645 47.995 16.935 48.040 ;
        RECT 18.930 47.980 19.250 48.040 ;
        RECT 23.545 48.180 23.835 48.225 ;
        RECT 31.810 48.180 32.130 48.240 ;
        RECT 44.690 48.225 45.010 48.240 ;
        RECT 44.660 48.180 45.010 48.225 ;
        RECT 23.545 48.040 32.130 48.180 ;
        RECT 44.495 48.040 45.010 48.180 ;
        RECT 23.545 47.995 23.835 48.040 ;
        RECT 31.810 47.980 32.130 48.040 ;
        RECT 44.660 47.995 45.010 48.040 ;
        RECT 44.690 47.980 45.010 47.995 ;
        RECT 69.530 48.180 69.850 48.240 ;
        RECT 70.925 48.180 71.215 48.225 ;
        RECT 69.530 48.040 71.215 48.180 ;
        RECT 69.530 47.980 69.850 48.040 ;
        RECT 70.925 47.995 71.215 48.040 ;
        RECT 8.350 47.640 8.670 47.900 ;
        RECT 10.205 47.840 10.495 47.885 ;
        RECT 12.490 47.840 12.810 47.900 ;
        RECT 10.205 47.700 12.810 47.840 ;
        RECT 10.205 47.655 10.495 47.700 ;
        RECT 12.490 47.640 12.810 47.700 ;
        RECT 17.565 47.655 17.855 47.885 ;
        RECT 19.020 47.840 19.160 47.980 ;
        RECT 24.005 47.840 24.295 47.885 ;
        RECT 19.020 47.700 24.295 47.840 ;
        RECT 24.005 47.655 24.295 47.700 ;
        RECT 24.925 47.840 25.215 47.885 ;
        RECT 26.750 47.840 27.070 47.900 ;
        RECT 24.925 47.700 27.070 47.840 ;
        RECT 24.925 47.655 25.215 47.700 ;
        RECT 5.130 47.160 5.450 47.220 ;
        RECT 9.285 47.160 9.575 47.205 ;
        RECT 17.640 47.160 17.780 47.655 ;
        RECT 26.750 47.640 27.070 47.700 ;
        RECT 30.445 47.655 30.735 47.885 ;
        RECT 19.865 47.500 20.155 47.545 ;
        RECT 20.770 47.500 21.090 47.560 ;
        RECT 23.070 47.500 23.390 47.560 ;
        RECT 19.865 47.360 23.390 47.500 ;
        RECT 19.865 47.315 20.155 47.360 ;
        RECT 20.770 47.300 21.090 47.360 ;
        RECT 23.070 47.300 23.390 47.360 ;
        RECT 23.530 47.500 23.850 47.560 ;
        RECT 25.845 47.500 26.135 47.545 ;
        RECT 23.530 47.360 26.135 47.500 ;
        RECT 30.520 47.500 30.660 47.655 ;
        RECT 33.190 47.640 33.510 47.900 ;
        RECT 33.650 47.640 33.970 47.900 ;
        RECT 34.570 47.640 34.890 47.900 ;
        RECT 35.045 47.840 35.335 47.885 ;
        RECT 36.410 47.840 36.730 47.900 ;
        RECT 37.330 47.885 37.650 47.900 ;
        RECT 35.045 47.700 36.730 47.840 ;
        RECT 35.045 47.655 35.335 47.700 ;
        RECT 36.410 47.640 36.730 47.700 ;
        RECT 37.300 47.655 37.650 47.885 ;
        RECT 43.325 47.840 43.615 47.885 ;
        RECT 46.070 47.840 46.390 47.900 ;
        RECT 43.325 47.700 46.390 47.840 ;
        RECT 43.325 47.655 43.615 47.700 ;
        RECT 37.330 47.640 37.650 47.655 ;
        RECT 46.070 47.640 46.390 47.700 ;
        RECT 70.450 47.640 70.770 47.900 ;
        RECT 82.410 47.640 82.730 47.900 ;
        RECT 30.520 47.360 34.800 47.500 ;
        RECT 23.530 47.300 23.850 47.360 ;
        RECT 25.845 47.315 26.135 47.360 ;
        RECT 34.660 47.220 34.800 47.360 ;
        RECT 35.965 47.315 36.255 47.545 ;
        RECT 36.845 47.500 37.135 47.545 ;
        RECT 38.035 47.500 38.325 47.545 ;
        RECT 40.555 47.500 40.845 47.545 ;
        RECT 36.845 47.360 40.845 47.500 ;
        RECT 36.845 47.315 37.135 47.360 ;
        RECT 38.035 47.315 38.325 47.360 ;
        RECT 40.555 47.315 40.845 47.360 ;
        RECT 44.205 47.500 44.495 47.545 ;
        RECT 45.395 47.500 45.685 47.545 ;
        RECT 47.915 47.500 48.205 47.545 ;
        RECT 44.205 47.360 48.205 47.500 ;
        RECT 44.205 47.315 44.495 47.360 ;
        RECT 45.395 47.315 45.685 47.360 ;
        RECT 47.915 47.315 48.205 47.360 ;
        RECT 33.650 47.160 33.970 47.220 ;
        RECT 5.130 47.020 9.575 47.160 ;
        RECT 5.130 46.960 5.450 47.020 ;
        RECT 9.285 46.975 9.575 47.020 ;
        RECT 13.730 47.020 33.970 47.160 ;
        RECT 6.510 46.820 6.830 46.880 ;
        RECT 7.445 46.820 7.735 46.865 ;
        RECT 6.510 46.680 7.735 46.820 ;
        RECT 6.510 46.620 6.830 46.680 ;
        RECT 7.445 46.635 7.735 46.680 ;
        RECT 8.350 46.820 8.670 46.880 ;
        RECT 13.730 46.820 13.870 47.020 ;
        RECT 33.650 46.960 33.970 47.020 ;
        RECT 34.570 47.160 34.890 47.220 ;
        RECT 36.040 47.160 36.180 47.315 ;
        RECT 52.970 47.300 53.290 47.560 ;
        RECT 53.445 47.315 53.735 47.545 ;
        RECT 34.570 47.020 36.180 47.160 ;
        RECT 36.450 47.160 36.740 47.205 ;
        RECT 38.550 47.160 38.840 47.205 ;
        RECT 40.120 47.160 40.410 47.205 ;
        RECT 36.450 47.020 40.410 47.160 ;
        RECT 34.570 46.960 34.890 47.020 ;
        RECT 36.450 46.975 36.740 47.020 ;
        RECT 38.550 46.975 38.840 47.020 ;
        RECT 40.120 46.975 40.410 47.020 ;
        RECT 42.850 46.960 43.170 47.220 ;
        RECT 43.810 47.160 44.100 47.205 ;
        RECT 45.910 47.160 46.200 47.205 ;
        RECT 47.480 47.160 47.770 47.205 ;
        RECT 43.810 47.020 47.770 47.160 ;
        RECT 43.810 46.975 44.100 47.020 ;
        RECT 45.910 46.975 46.200 47.020 ;
        RECT 47.480 46.975 47.770 47.020 ;
        RECT 50.225 47.160 50.515 47.205 ;
        RECT 51.130 47.160 51.450 47.220 ;
        RECT 50.225 47.020 51.450 47.160 ;
        RECT 50.225 46.975 50.515 47.020 ;
        RECT 51.130 46.960 51.450 47.020 ;
        RECT 8.350 46.680 13.870 46.820 ;
        RECT 18.485 46.820 18.775 46.865 ;
        RECT 20.310 46.820 20.630 46.880 ;
        RECT 18.485 46.680 20.630 46.820 ;
        RECT 8.350 46.620 8.670 46.680 ;
        RECT 18.485 46.635 18.775 46.680 ;
        RECT 20.310 46.620 20.630 46.680 ;
        RECT 32.285 46.820 32.575 46.865 ;
        RECT 39.630 46.820 39.950 46.880 ;
        RECT 32.285 46.680 39.950 46.820 ;
        RECT 32.285 46.635 32.575 46.680 ;
        RECT 39.630 46.620 39.950 46.680 ;
        RECT 41.470 46.820 41.790 46.880 ;
        RECT 47.910 46.820 48.230 46.880 ;
        RECT 53.520 46.820 53.660 47.315 ;
        RECT 81.030 47.160 81.350 47.220 ;
        RECT 81.505 47.160 81.795 47.205 ;
        RECT 81.030 47.020 81.795 47.160 ;
        RECT 81.030 46.960 81.350 47.020 ;
        RECT 81.505 46.975 81.795 47.020 ;
        RECT 41.470 46.680 53.660 46.820 ;
        RECT 41.470 46.620 41.790 46.680 ;
        RECT 47.910 46.620 48.230 46.680 ;
        RECT 5.520 46.000 84.180 46.480 ;
        RECT 22.150 45.800 22.470 45.860 ;
        RECT 29.510 45.800 29.830 45.860 ;
        RECT 22.150 45.660 29.830 45.800 ;
        RECT 22.150 45.600 22.470 45.660 ;
        RECT 29.510 45.600 29.830 45.660 ;
        RECT 29.985 45.800 30.275 45.845 ;
        RECT 33.650 45.800 33.970 45.860 ;
        RECT 29.985 45.660 33.970 45.800 ;
        RECT 29.985 45.615 30.275 45.660 ;
        RECT 33.650 45.600 33.970 45.660 ;
        RECT 37.330 45.800 37.650 45.860 ;
        RECT 37.805 45.800 38.095 45.845 ;
        RECT 37.330 45.660 38.095 45.800 ;
        RECT 37.330 45.600 37.650 45.660 ;
        RECT 37.805 45.615 38.095 45.660 ;
        RECT 45.150 45.800 45.470 45.860 ;
        RECT 49.305 45.800 49.595 45.845 ;
        RECT 45.150 45.660 49.595 45.800 ;
        RECT 45.150 45.600 45.470 45.660 ;
        RECT 49.305 45.615 49.595 45.660 ;
        RECT 54.350 45.600 54.670 45.860 ;
        RECT 55.270 45.800 55.590 45.860 ;
        RECT 64.010 45.800 64.330 45.860 ;
        RECT 55.270 45.660 64.330 45.800 ;
        RECT 55.270 45.600 55.590 45.660 ;
        RECT 64.010 45.600 64.330 45.660 ;
        RECT 4.210 45.460 4.530 45.520 ;
        RECT 7.445 45.460 7.735 45.505 ;
        RECT 13.870 45.460 14.190 45.520 ;
        RECT 17.550 45.460 17.870 45.520 ;
        RECT 4.210 45.320 7.735 45.460 ;
        RECT 4.210 45.260 4.530 45.320 ;
        RECT 7.445 45.275 7.735 45.320 ;
        RECT 9.820 45.320 17.870 45.460 ;
        RECT 8.350 44.580 8.670 44.840 ;
        RECT 9.820 44.825 9.960 45.320 ;
        RECT 13.870 45.260 14.190 45.320 ;
        RECT 17.550 45.260 17.870 45.320 ;
        RECT 23.570 45.460 23.860 45.505 ;
        RECT 25.670 45.460 25.960 45.505 ;
        RECT 27.240 45.460 27.530 45.505 ;
        RECT 23.570 45.320 27.530 45.460 ;
        RECT 23.570 45.275 23.860 45.320 ;
        RECT 25.670 45.275 25.960 45.320 ;
        RECT 27.240 45.275 27.530 45.320 ;
        RECT 30.930 45.460 31.220 45.505 ;
        RECT 33.030 45.460 33.320 45.505 ;
        RECT 34.600 45.460 34.890 45.505 ;
        RECT 30.930 45.320 34.890 45.460 ;
        RECT 30.930 45.275 31.220 45.320 ;
        RECT 33.030 45.275 33.320 45.320 ;
        RECT 34.600 45.275 34.890 45.320 ;
        RECT 36.410 45.460 36.730 45.520 ;
        RECT 64.945 45.460 65.235 45.505 ;
        RECT 36.410 45.320 65.235 45.460 ;
        RECT 36.410 45.260 36.730 45.320 ;
        RECT 64.945 45.275 65.235 45.320 ;
        RECT 12.950 45.120 13.270 45.180 ;
        RECT 21.690 45.120 22.010 45.180 ;
        RECT 11.200 44.980 22.010 45.120 ;
        RECT 9.745 44.595 10.035 44.825 ;
        RECT 10.190 44.780 10.510 44.840 ;
        RECT 11.200 44.825 11.340 44.980 ;
        RECT 12.950 44.920 13.270 44.980 ;
        RECT 10.665 44.780 10.955 44.825 ;
        RECT 10.190 44.640 10.955 44.780 ;
        RECT 10.190 44.580 10.510 44.640 ;
        RECT 10.665 44.595 10.955 44.640 ;
        RECT 11.125 44.595 11.415 44.825 ;
        RECT 11.570 44.580 11.890 44.840 ;
        RECT 14.790 44.580 15.110 44.840 ;
        RECT 18.470 44.780 18.790 44.840 ;
        RECT 19.405 44.780 19.695 44.825 ;
        RECT 18.470 44.640 19.695 44.780 ;
        RECT 18.470 44.580 18.790 44.640 ;
        RECT 19.405 44.595 19.695 44.640 ;
        RECT 12.950 43.900 13.270 44.160 ;
        RECT 13.870 43.900 14.190 44.160 ;
        RECT 19.480 44.100 19.620 44.595 ;
        RECT 20.310 44.580 20.630 44.840 ;
        RECT 20.860 44.825 21.000 44.980 ;
        RECT 21.690 44.920 22.010 44.980 ;
        RECT 23.070 44.920 23.390 45.180 ;
        RECT 23.965 45.120 24.255 45.165 ;
        RECT 25.155 45.120 25.445 45.165 ;
        RECT 27.675 45.120 27.965 45.165 ;
        RECT 23.965 44.980 27.965 45.120 ;
        RECT 23.965 44.935 24.255 44.980 ;
        RECT 25.155 44.935 25.445 44.980 ;
        RECT 27.675 44.935 27.965 44.980 ;
        RECT 31.325 45.120 31.615 45.165 ;
        RECT 32.515 45.120 32.805 45.165 ;
        RECT 35.035 45.120 35.325 45.165 ;
        RECT 31.325 44.980 35.325 45.120 ;
        RECT 31.325 44.935 31.615 44.980 ;
        RECT 32.515 44.935 32.805 44.980 ;
        RECT 35.035 44.935 35.325 44.980 ;
        RECT 39.630 45.120 39.950 45.180 ;
        RECT 40.105 45.120 40.395 45.165 ;
        RECT 39.630 44.980 40.395 45.120 ;
        RECT 39.630 44.920 39.950 44.980 ;
        RECT 40.105 44.935 40.395 44.980 ;
        RECT 41.025 45.120 41.315 45.165 ;
        RECT 41.470 45.120 41.790 45.180 ;
        RECT 41.025 44.980 41.790 45.120 ;
        RECT 41.025 44.935 41.315 44.980 ;
        RECT 41.470 44.920 41.790 44.980 ;
        RECT 42.850 45.120 43.170 45.180 ;
        RECT 47.465 45.120 47.755 45.165 ;
        RECT 42.850 44.980 47.755 45.120 ;
        RECT 42.850 44.920 43.170 44.980 ;
        RECT 47.465 44.935 47.755 44.980 ;
        RECT 47.910 45.120 48.230 45.180 ;
        RECT 66.310 45.120 66.630 45.180 ;
        RECT 47.910 44.980 50.440 45.120 ;
        RECT 47.910 44.920 48.230 44.980 ;
        RECT 20.785 44.595 21.075 44.825 ;
        RECT 21.245 44.780 21.535 44.825 ;
        RECT 23.530 44.780 23.850 44.840 ;
        RECT 27.210 44.780 27.530 44.840 ;
        RECT 21.245 44.640 27.530 44.780 ;
        RECT 21.245 44.595 21.535 44.640 ;
        RECT 23.530 44.580 23.850 44.640 ;
        RECT 27.210 44.580 27.530 44.640 ;
        RECT 30.445 44.780 30.735 44.825 ;
        RECT 34.570 44.780 34.890 44.840 ;
        RECT 30.445 44.640 34.890 44.780 ;
        RECT 30.445 44.595 30.735 44.640 ;
        RECT 34.570 44.580 34.890 44.640 ;
        RECT 35.120 44.640 49.980 44.780 ;
        RECT 22.625 44.440 22.915 44.485 ;
        RECT 24.310 44.440 24.600 44.485 ;
        RECT 22.625 44.300 24.600 44.440 ;
        RECT 22.625 44.255 22.915 44.300 ;
        RECT 24.310 44.255 24.600 44.300 ;
        RECT 25.370 44.440 25.690 44.500 ;
        RECT 26.750 44.440 27.070 44.500 ;
        RECT 25.370 44.300 27.070 44.440 ;
        RECT 25.370 44.240 25.690 44.300 ;
        RECT 26.750 44.240 27.070 44.300 ;
        RECT 31.780 44.440 32.070 44.485 ;
        RECT 32.270 44.440 32.590 44.500 ;
        RECT 35.120 44.440 35.260 44.640 ;
        RECT 31.780 44.300 32.590 44.440 ;
        RECT 31.780 44.255 32.070 44.300 ;
        RECT 32.270 44.240 32.590 44.300 ;
        RECT 32.820 44.300 35.260 44.440 ;
        RECT 39.645 44.440 39.935 44.485 ;
        RECT 44.705 44.440 44.995 44.485 ;
        RECT 39.645 44.300 44.995 44.440 ;
        RECT 32.820 44.100 32.960 44.300 ;
        RECT 39.645 44.255 39.935 44.300 ;
        RECT 44.705 44.255 44.995 44.300 ;
        RECT 48.370 44.240 48.690 44.500 ;
        RECT 19.480 43.960 32.960 44.100 ;
        RECT 33.190 44.100 33.510 44.160 ;
        RECT 37.330 44.100 37.650 44.160 ;
        RECT 33.190 43.960 37.650 44.100 ;
        RECT 33.190 43.900 33.510 43.960 ;
        RECT 37.330 43.900 37.650 43.960 ;
        RECT 49.290 43.900 49.610 44.160 ;
        RECT 49.840 44.100 49.980 44.640 ;
        RECT 50.300 44.440 50.440 44.980 ;
        RECT 55.820 44.980 66.630 45.120 ;
        RECT 50.685 44.780 50.975 44.825 ;
        RECT 55.270 44.780 55.590 44.840 ;
        RECT 55.820 44.825 55.960 44.980 ;
        RECT 66.310 44.920 66.630 44.980 ;
        RECT 50.685 44.640 55.590 44.780 ;
        RECT 50.685 44.595 50.975 44.640 ;
        RECT 55.270 44.580 55.590 44.640 ;
        RECT 55.745 44.595 56.035 44.825 ;
        RECT 57.110 44.580 57.430 44.840 ;
        RECT 57.585 44.780 57.875 44.825 ;
        RECT 58.965 44.780 59.255 44.825 ;
        RECT 60.790 44.780 61.110 44.840 ;
        RECT 57.585 44.640 58.260 44.780 ;
        RECT 57.585 44.595 57.875 44.640 ;
        RECT 51.605 44.440 51.895 44.485 ;
        RECT 50.300 44.300 51.895 44.440 ;
        RECT 51.605 44.255 51.895 44.300 ;
        RECT 52.525 44.440 52.815 44.485 ;
        RECT 54.810 44.440 55.130 44.500 ;
        RECT 56.205 44.440 56.495 44.485 ;
        RECT 52.525 44.300 56.495 44.440 ;
        RECT 52.525 44.255 52.815 44.300 ;
        RECT 54.810 44.240 55.130 44.300 ;
        RECT 56.205 44.255 56.495 44.300 ;
        RECT 58.120 44.100 58.260 44.640 ;
        RECT 58.965 44.640 61.110 44.780 ;
        RECT 58.965 44.595 59.255 44.640 ;
        RECT 60.790 44.580 61.110 44.640 ;
        RECT 62.185 44.780 62.475 44.825 ;
        RECT 62.630 44.780 62.950 44.840 ;
        RECT 62.185 44.640 62.950 44.780 ;
        RECT 62.185 44.595 62.475 44.640 ;
        RECT 62.630 44.580 62.950 44.640 ;
        RECT 64.010 44.580 64.330 44.840 ;
        RECT 70.465 44.780 70.755 44.825 ;
        RECT 65.480 44.640 70.755 44.780 ;
        RECT 58.490 44.440 58.810 44.500 ;
        RECT 63.105 44.440 63.395 44.485 ;
        RECT 58.490 44.300 63.395 44.440 ;
        RECT 58.490 44.240 58.810 44.300 ;
        RECT 63.105 44.255 63.395 44.300 ;
        RECT 63.565 44.440 63.855 44.485 ;
        RECT 64.470 44.440 64.790 44.500 ;
        RECT 65.480 44.440 65.620 44.640 ;
        RECT 70.465 44.595 70.755 44.640 ;
        RECT 63.565 44.300 64.790 44.440 ;
        RECT 63.565 44.255 63.855 44.300 ;
        RECT 64.470 44.240 64.790 44.300 ;
        RECT 65.020 44.300 65.620 44.440 ;
        RECT 49.840 43.960 58.260 44.100 ;
        RECT 60.790 44.100 61.110 44.160 ;
        RECT 65.020 44.100 65.160 44.300 ;
        RECT 66.310 44.240 66.630 44.500 ;
        RECT 67.230 44.240 67.550 44.500 ;
        RECT 70.540 44.440 70.680 44.595 ;
        RECT 71.370 44.580 71.690 44.840 ;
        RECT 71.830 44.580 72.150 44.840 ;
        RECT 72.290 44.580 72.610 44.840 ;
        RECT 76.890 44.440 77.210 44.500 ;
        RECT 70.540 44.300 77.210 44.440 ;
        RECT 76.890 44.240 77.210 44.300 ;
        RECT 60.790 43.960 65.160 44.100 ;
        RECT 60.790 43.900 61.110 43.960 ;
        RECT 65.390 43.900 65.710 44.160 ;
        RECT 73.670 43.900 73.990 44.160 ;
        RECT 5.520 43.280 84.180 43.760 ;
        RECT 10.190 42.880 10.510 43.140 ;
        RECT 15.710 43.080 16.030 43.140 ;
        RECT 17.565 43.080 17.855 43.125 ;
        RECT 30.890 43.080 31.210 43.140 ;
        RECT 11.660 42.940 17.855 43.080 ;
        RECT 6.970 42.740 7.290 42.800 ;
        RECT 8.365 42.740 8.655 42.785 ;
        RECT 6.970 42.600 8.655 42.740 ;
        RECT 6.970 42.540 7.290 42.600 ;
        RECT 8.365 42.555 8.655 42.600 ;
        RECT 9.285 42.740 9.575 42.785 ;
        RECT 11.660 42.740 11.800 42.940 ;
        RECT 15.710 42.880 16.030 42.940 ;
        RECT 17.565 42.895 17.855 42.940 ;
        RECT 19.480 42.940 31.210 43.080 ;
        RECT 9.285 42.600 11.800 42.740 ;
        RECT 12.000 42.740 12.290 42.785 ;
        RECT 12.950 42.740 13.270 42.800 ;
        RECT 12.000 42.600 13.270 42.740 ;
        RECT 9.285 42.555 9.575 42.600 ;
        RECT 12.000 42.555 12.290 42.600 ;
        RECT 8.440 42.400 8.580 42.555 ;
        RECT 12.950 42.540 13.270 42.600 ;
        RECT 14.790 42.740 15.110 42.800 ;
        RECT 18.985 42.740 19.275 42.785 ;
        RECT 19.480 42.740 19.620 42.940 ;
        RECT 30.890 42.880 31.210 42.940 ;
        RECT 66.310 43.080 66.630 43.140 ;
        RECT 73.225 43.080 73.515 43.125 ;
        RECT 75.970 43.080 76.290 43.140 ;
        RECT 66.310 42.940 76.290 43.080 ;
        RECT 66.310 42.880 66.630 42.940 ;
        RECT 73.225 42.895 73.515 42.940 ;
        RECT 75.970 42.880 76.290 42.940 ;
        RECT 14.790 42.600 19.620 42.740 ;
        RECT 19.865 42.740 20.155 42.785 ;
        RECT 19.865 42.600 21.460 42.740 ;
        RECT 14.790 42.540 15.110 42.600 ;
        RECT 18.985 42.555 19.275 42.600 ;
        RECT 19.865 42.555 20.155 42.600 ;
        RECT 18.025 42.400 18.315 42.445 ;
        RECT 19.390 42.400 19.710 42.460 ;
        RECT 21.320 42.445 21.460 42.600 ;
        RECT 24.080 42.600 26.060 42.740 ;
        RECT 8.440 42.260 19.710 42.400 ;
        RECT 18.025 42.215 18.315 42.260 ;
        RECT 19.390 42.200 19.710 42.260 ;
        RECT 20.325 42.215 20.615 42.445 ;
        RECT 21.245 42.215 21.535 42.445 ;
        RECT 8.810 42.060 9.130 42.120 ;
        RECT 10.665 42.060 10.955 42.105 ;
        RECT 8.810 41.920 10.955 42.060 ;
        RECT 8.810 41.860 9.130 41.920 ;
        RECT 10.665 41.875 10.955 41.920 ;
        RECT 11.545 42.060 11.835 42.105 ;
        RECT 12.735 42.060 13.025 42.105 ;
        RECT 15.255 42.060 15.545 42.105 ;
        RECT 11.545 41.920 15.545 42.060 ;
        RECT 11.545 41.875 11.835 41.920 ;
        RECT 12.735 41.875 13.025 41.920 ;
        RECT 15.255 41.875 15.545 41.920 ;
        RECT 17.550 42.060 17.870 42.120 ;
        RECT 18.930 42.060 19.250 42.120 ;
        RECT 20.400 42.060 20.540 42.215 ;
        RECT 21.690 42.200 22.010 42.460 ;
        RECT 22.150 42.200 22.470 42.460 ;
        RECT 24.080 42.445 24.220 42.600 ;
        RECT 24.005 42.215 24.295 42.445 ;
        RECT 25.285 42.400 25.575 42.445 ;
        RECT 24.540 42.260 25.575 42.400 ;
        RECT 25.920 42.400 26.060 42.600 ;
        RECT 31.810 42.540 32.130 42.800 ;
        RECT 33.650 42.740 33.970 42.800 ;
        RECT 36.885 42.740 37.175 42.785 ;
        RECT 46.545 42.740 46.835 42.785 ;
        RECT 47.910 42.740 48.230 42.800 ;
        RECT 33.650 42.600 37.175 42.740 ;
        RECT 33.650 42.540 33.970 42.600 ;
        RECT 36.885 42.555 37.175 42.600 ;
        RECT 41.560 42.600 48.230 42.740 ;
        RECT 34.570 42.400 34.890 42.460 ;
        RECT 37.330 42.400 37.650 42.460 ;
        RECT 39.645 42.400 39.935 42.445 ;
        RECT 41.025 42.400 41.315 42.445 ;
        RECT 25.920 42.260 35.720 42.400 ;
        RECT 17.550 41.920 20.540 42.060 ;
        RECT 21.780 42.060 21.920 42.200 ;
        RECT 23.070 42.060 23.390 42.120 ;
        RECT 21.780 41.920 23.390 42.060 ;
        RECT 17.550 41.860 17.870 41.920 ;
        RECT 18.930 41.860 19.250 41.920 ;
        RECT 23.070 41.860 23.390 41.920 ;
        RECT 23.545 42.060 23.835 42.105 ;
        RECT 24.540 42.060 24.680 42.260 ;
        RECT 25.285 42.215 25.575 42.260 ;
        RECT 34.570 42.200 34.890 42.260 ;
        RECT 35.580 42.105 35.720 42.260 ;
        RECT 37.330 42.260 41.315 42.400 ;
        RECT 37.330 42.200 37.650 42.260 ;
        RECT 39.645 42.215 39.935 42.260 ;
        RECT 41.025 42.215 41.315 42.260 ;
        RECT 23.545 41.920 24.680 42.060 ;
        RECT 24.885 42.060 25.175 42.105 ;
        RECT 26.075 42.060 26.365 42.105 ;
        RECT 28.595 42.060 28.885 42.105 ;
        RECT 24.885 41.920 28.885 42.060 ;
        RECT 23.545 41.875 23.835 41.920 ;
        RECT 24.885 41.875 25.175 41.920 ;
        RECT 26.075 41.875 26.365 41.920 ;
        RECT 28.595 41.875 28.885 41.920 ;
        RECT 35.505 42.060 35.795 42.105 ;
        RECT 36.870 42.060 37.190 42.120 ;
        RECT 35.505 41.920 37.190 42.060 ;
        RECT 35.505 41.875 35.795 41.920 ;
        RECT 36.870 41.860 37.190 41.920 ;
        RECT 11.150 41.720 11.440 41.765 ;
        RECT 13.250 41.720 13.540 41.765 ;
        RECT 14.820 41.720 15.110 41.765 ;
        RECT 11.150 41.580 15.110 41.720 ;
        RECT 11.150 41.535 11.440 41.580 ;
        RECT 13.250 41.535 13.540 41.580 ;
        RECT 14.820 41.535 15.110 41.580 ;
        RECT 24.490 41.720 24.780 41.765 ;
        RECT 26.590 41.720 26.880 41.765 ;
        RECT 28.160 41.720 28.450 41.765 ;
        RECT 24.490 41.580 28.450 41.720 ;
        RECT 24.490 41.535 24.780 41.580 ;
        RECT 26.590 41.535 26.880 41.580 ;
        RECT 28.160 41.535 28.450 41.580 ;
        RECT 30.890 41.520 31.210 41.780 ;
        RECT 15.250 41.380 15.570 41.440 ;
        RECT 41.560 41.380 41.700 42.600 ;
        RECT 46.545 42.555 46.835 42.600 ;
        RECT 47.910 42.540 48.230 42.600 ;
        RECT 59.410 42.740 59.730 42.800 ;
        RECT 65.405 42.740 65.695 42.785 ;
        RECT 70.450 42.740 70.770 42.800 ;
        RECT 59.410 42.600 61.480 42.740 ;
        RECT 59.410 42.540 59.730 42.600 ;
        RECT 61.340 42.460 61.480 42.600 ;
        RECT 65.405 42.600 70.770 42.740 ;
        RECT 65.405 42.555 65.695 42.600 ;
        RECT 41.930 42.400 42.250 42.460 ;
        RECT 42.865 42.400 43.155 42.445 ;
        RECT 43.785 42.400 44.075 42.445 ;
        RECT 44.230 42.400 44.550 42.460 ;
        RECT 41.930 42.260 44.550 42.400 ;
        RECT 41.930 42.200 42.250 42.260 ;
        RECT 42.865 42.215 43.155 42.260 ;
        RECT 43.785 42.215 44.075 42.260 ;
        RECT 44.230 42.200 44.550 42.260 ;
        RECT 45.150 42.200 45.470 42.460 ;
        RECT 46.070 42.400 46.390 42.460 ;
        RECT 48.830 42.400 49.150 42.460 ;
        RECT 46.070 42.260 49.150 42.400 ;
        RECT 46.070 42.200 46.390 42.260 ;
        RECT 48.830 42.200 49.150 42.260 ;
        RECT 53.430 42.200 53.750 42.460 ;
        RECT 54.365 42.400 54.655 42.445 ;
        RECT 54.810 42.400 55.130 42.460 ;
        RECT 58.490 42.400 58.810 42.460 ;
        RECT 54.365 42.260 58.810 42.400 ;
        RECT 54.365 42.215 54.655 42.260 ;
        RECT 54.810 42.200 55.130 42.260 ;
        RECT 58.490 42.200 58.810 42.260 ;
        RECT 60.805 42.215 61.095 42.445 ;
        RECT 45.625 41.875 45.915 42.105 ;
        RECT 45.700 41.720 45.840 41.875 ;
        RECT 52.510 41.860 52.830 42.120 ;
        RECT 59.410 42.060 59.730 42.120 ;
        RECT 60.880 42.060 61.020 42.215 ;
        RECT 61.250 42.200 61.570 42.460 ;
        RECT 65.480 42.060 65.620 42.555 ;
        RECT 70.450 42.540 70.770 42.600 ;
        RECT 65.850 42.400 66.170 42.460 ;
        RECT 67.605 42.400 67.895 42.445 ;
        RECT 65.850 42.260 67.895 42.400 ;
        RECT 65.850 42.200 66.170 42.260 ;
        RECT 67.605 42.215 67.895 42.260 ;
        RECT 81.030 42.200 81.350 42.460 ;
        RECT 66.325 42.060 66.615 42.105 ;
        RECT 59.410 41.920 66.615 42.060 ;
        RECT 59.410 41.860 59.730 41.920 ;
        RECT 66.325 41.875 66.615 41.920 ;
        RECT 67.205 42.060 67.495 42.105 ;
        RECT 68.395 42.060 68.685 42.105 ;
        RECT 70.915 42.060 71.205 42.105 ;
        RECT 67.205 41.920 71.205 42.060 ;
        RECT 67.205 41.875 67.495 41.920 ;
        RECT 68.395 41.875 68.685 41.920 ;
        RECT 70.915 41.875 71.205 41.920 ;
        RECT 49.290 41.720 49.610 41.780 ;
        RECT 45.700 41.580 49.610 41.720 ;
        RECT 49.290 41.520 49.610 41.580 ;
        RECT 66.810 41.720 67.100 41.765 ;
        RECT 68.910 41.720 69.200 41.765 ;
        RECT 70.480 41.720 70.770 41.765 ;
        RECT 66.810 41.580 70.770 41.720 ;
        RECT 66.810 41.535 67.100 41.580 ;
        RECT 68.910 41.535 69.200 41.580 ;
        RECT 70.480 41.535 70.770 41.580 ;
        RECT 81.965 41.720 82.255 41.765 ;
        RECT 82.870 41.720 83.190 41.780 ;
        RECT 81.965 41.580 83.190 41.720 ;
        RECT 81.965 41.535 82.255 41.580 ;
        RECT 82.870 41.520 83.190 41.580 ;
        RECT 15.250 41.240 41.700 41.380 ;
        RECT 15.250 41.180 15.570 41.240 ;
        RECT 5.520 40.560 84.180 41.040 ;
        RECT 8.810 40.360 9.130 40.420 ;
        RECT 7.060 40.220 9.130 40.360 ;
        RECT 7.060 39.725 7.200 40.220 ;
        RECT 8.810 40.160 9.130 40.220 ;
        RECT 12.490 40.360 12.810 40.420 ;
        RECT 13.885 40.360 14.175 40.405 ;
        RECT 12.490 40.220 14.175 40.360 ;
        RECT 12.490 40.160 12.810 40.220 ;
        RECT 13.885 40.175 14.175 40.220 ;
        RECT 22.625 40.360 22.915 40.405 ;
        RECT 23.070 40.360 23.390 40.420 ;
        RECT 22.625 40.220 23.390 40.360 ;
        RECT 22.625 40.175 22.915 40.220 ;
        RECT 23.070 40.160 23.390 40.220 ;
        RECT 31.825 40.360 32.115 40.405 ;
        RECT 32.270 40.360 32.590 40.420 ;
        RECT 43.785 40.360 44.075 40.405 ;
        RECT 45.150 40.360 45.470 40.420 ;
        RECT 53.430 40.360 53.750 40.420 ;
        RECT 64.470 40.360 64.790 40.420 ;
        RECT 31.825 40.220 32.590 40.360 ;
        RECT 31.825 40.175 32.115 40.220 ;
        RECT 32.270 40.160 32.590 40.220 ;
        RECT 32.820 40.220 41.700 40.360 ;
        RECT 7.470 40.020 7.760 40.065 ;
        RECT 9.570 40.020 9.860 40.065 ;
        RECT 11.140 40.020 11.430 40.065 ;
        RECT 7.470 39.880 11.430 40.020 ;
        RECT 7.470 39.835 7.760 39.880 ;
        RECT 9.570 39.835 9.860 39.880 ;
        RECT 11.140 39.835 11.430 39.880 ;
        RECT 18.010 40.020 18.330 40.080 ;
        RECT 21.705 40.020 21.995 40.065 ;
        RECT 30.430 40.020 30.750 40.080 ;
        RECT 18.010 39.880 21.000 40.020 ;
        RECT 18.010 39.820 18.330 39.880 ;
        RECT 6.985 39.495 7.275 39.725 ;
        RECT 7.865 39.680 8.155 39.725 ;
        RECT 9.055 39.680 9.345 39.725 ;
        RECT 11.575 39.680 11.865 39.725 ;
        RECT 20.860 39.680 21.000 39.880 ;
        RECT 21.705 39.880 30.750 40.020 ;
        RECT 21.705 39.835 21.995 39.880 ;
        RECT 30.430 39.820 30.750 39.880 ;
        RECT 22.610 39.680 22.930 39.740 ;
        RECT 7.865 39.540 11.865 39.680 ;
        RECT 7.865 39.495 8.155 39.540 ;
        RECT 9.055 39.495 9.345 39.540 ;
        RECT 11.575 39.495 11.865 39.540 ;
        RECT 15.800 39.540 20.540 39.680 ;
        RECT 15.800 39.400 15.940 39.540 ;
        RECT 15.710 39.140 16.030 39.400 ;
        RECT 17.090 39.340 17.410 39.400 ;
        RECT 18.945 39.340 19.235 39.385 ;
        RECT 17.090 39.200 19.235 39.340 ;
        RECT 17.090 39.140 17.410 39.200 ;
        RECT 18.945 39.155 19.235 39.200 ;
        RECT 19.405 39.340 19.695 39.385 ;
        RECT 19.850 39.340 20.170 39.400 ;
        RECT 20.400 39.385 20.540 39.540 ;
        RECT 20.860 39.540 22.930 39.680 ;
        RECT 20.860 39.385 21.000 39.540 ;
        RECT 22.610 39.480 22.930 39.540 ;
        RECT 24.925 39.680 25.215 39.725 ;
        RECT 26.750 39.680 27.070 39.740 ;
        RECT 32.820 39.680 32.960 40.220 ;
        RECT 37.370 40.020 37.660 40.065 ;
        RECT 39.470 40.020 39.760 40.065 ;
        RECT 41.040 40.020 41.330 40.065 ;
        RECT 37.370 39.880 41.330 40.020 ;
        RECT 41.560 40.020 41.700 40.220 ;
        RECT 43.785 40.220 45.470 40.360 ;
        RECT 43.785 40.175 44.075 40.220 ;
        RECT 45.150 40.160 45.470 40.220 ;
        RECT 45.700 40.220 64.790 40.360 ;
        RECT 45.700 40.020 45.840 40.220 ;
        RECT 53.430 40.160 53.750 40.220 ;
        RECT 64.470 40.160 64.790 40.220 ;
        RECT 65.850 40.160 66.170 40.420 ;
        RECT 68.165 40.360 68.455 40.405 ;
        RECT 71.370 40.360 71.690 40.420 ;
        RECT 68.165 40.220 71.690 40.360 ;
        RECT 68.165 40.175 68.455 40.220 ;
        RECT 71.370 40.160 71.690 40.220 ;
        RECT 41.560 39.880 45.840 40.020 ;
        RECT 46.570 40.020 46.860 40.065 ;
        RECT 48.670 40.020 48.960 40.065 ;
        RECT 50.240 40.020 50.530 40.065 ;
        RECT 46.570 39.880 50.530 40.020 ;
        RECT 37.370 39.835 37.660 39.880 ;
        RECT 39.470 39.835 39.760 39.880 ;
        RECT 41.040 39.835 41.330 39.880 ;
        RECT 46.570 39.835 46.860 39.880 ;
        RECT 48.670 39.835 48.960 39.880 ;
        RECT 50.240 39.835 50.530 39.880 ;
        RECT 54.850 40.020 55.140 40.065 ;
        RECT 56.950 40.020 57.240 40.065 ;
        RECT 58.520 40.020 58.810 40.065 ;
        RECT 54.850 39.880 58.810 40.020 ;
        RECT 54.850 39.835 55.140 39.880 ;
        RECT 56.950 39.835 57.240 39.880 ;
        RECT 58.520 39.835 58.810 39.880 ;
        RECT 70.950 40.020 71.240 40.065 ;
        RECT 73.050 40.020 73.340 40.065 ;
        RECT 74.620 40.020 74.910 40.065 ;
        RECT 70.950 39.880 74.910 40.020 ;
        RECT 70.950 39.835 71.240 39.880 ;
        RECT 73.050 39.835 73.340 39.880 ;
        RECT 74.620 39.835 74.910 39.880 ;
        RECT 34.125 39.680 34.415 39.725 ;
        RECT 24.925 39.540 32.960 39.680 ;
        RECT 33.280 39.540 34.415 39.680 ;
        RECT 24.925 39.495 25.215 39.540 ;
        RECT 26.750 39.480 27.070 39.540 ;
        RECT 19.405 39.200 20.170 39.340 ;
        RECT 19.405 39.155 19.695 39.200 ;
        RECT 19.850 39.140 20.170 39.200 ;
        RECT 20.325 39.155 20.615 39.385 ;
        RECT 20.785 39.155 21.075 39.385 ;
        RECT 21.230 39.340 21.550 39.400 ;
        RECT 24.005 39.340 24.295 39.385 ;
        RECT 24.465 39.340 24.755 39.385 ;
        RECT 26.290 39.340 26.610 39.400 ;
        RECT 21.230 39.200 26.610 39.340 ;
        RECT 21.230 39.140 21.550 39.200 ;
        RECT 24.005 39.155 24.295 39.200 ;
        RECT 24.465 39.155 24.755 39.200 ;
        RECT 26.290 39.140 26.610 39.200 ;
        RECT 29.970 39.340 30.290 39.400 ;
        RECT 33.280 39.340 33.420 39.540 ;
        RECT 34.125 39.495 34.415 39.540 ;
        RECT 35.045 39.680 35.335 39.725 ;
        RECT 37.765 39.680 38.055 39.725 ;
        RECT 38.955 39.680 39.245 39.725 ;
        RECT 41.475 39.680 41.765 39.725 ;
        RECT 35.045 39.540 37.560 39.680 ;
        RECT 35.045 39.495 35.335 39.540 ;
        RECT 29.970 39.200 33.420 39.340 ;
        RECT 29.970 39.140 30.290 39.200 ;
        RECT 33.650 39.140 33.970 39.400 ;
        RECT 36.870 39.140 37.190 39.400 ;
        RECT 37.420 39.340 37.560 39.540 ;
        RECT 37.765 39.540 41.765 39.680 ;
        RECT 37.765 39.495 38.055 39.540 ;
        RECT 38.955 39.495 39.245 39.540 ;
        RECT 41.475 39.495 41.765 39.540 ;
        RECT 46.965 39.680 47.255 39.725 ;
        RECT 48.155 39.680 48.445 39.725 ;
        RECT 50.675 39.680 50.965 39.725 ;
        RECT 46.965 39.540 50.965 39.680 ;
        RECT 46.965 39.495 47.255 39.540 ;
        RECT 48.155 39.495 48.445 39.540 ;
        RECT 50.675 39.495 50.965 39.540 ;
        RECT 55.245 39.680 55.535 39.725 ;
        RECT 56.435 39.680 56.725 39.725 ;
        RECT 58.955 39.680 59.245 39.725 ;
        RECT 65.390 39.680 65.710 39.740 ;
        RECT 55.245 39.540 59.245 39.680 ;
        RECT 55.245 39.495 55.535 39.540 ;
        RECT 56.435 39.495 56.725 39.540 ;
        RECT 58.955 39.495 59.245 39.540 ;
        RECT 63.640 39.540 65.710 39.680 ;
        RECT 44.230 39.340 44.550 39.400 ;
        RECT 44.705 39.340 44.995 39.385 ;
        RECT 37.420 39.200 41.700 39.340 ;
        RECT 41.560 39.060 41.700 39.200 ;
        RECT 44.230 39.200 44.995 39.340 ;
        RECT 44.230 39.140 44.550 39.200 ;
        RECT 44.705 39.155 44.995 39.200 ;
        RECT 46.085 39.340 46.375 39.385 ;
        RECT 48.830 39.340 49.150 39.400 ;
        RECT 54.365 39.340 54.655 39.385 ;
        RECT 59.410 39.340 59.730 39.400 ;
        RECT 46.085 39.200 50.900 39.340 ;
        RECT 46.085 39.155 46.375 39.200 ;
        RECT 48.830 39.140 49.150 39.200 ;
        RECT 50.760 39.060 50.900 39.200 ;
        RECT 54.365 39.200 59.730 39.340 ;
        RECT 54.365 39.155 54.655 39.200 ;
        RECT 59.410 39.140 59.730 39.200 ;
        RECT 60.790 39.340 61.110 39.400 ;
        RECT 63.640 39.385 63.780 39.540 ;
        RECT 65.390 39.480 65.710 39.540 ;
        RECT 71.345 39.680 71.635 39.725 ;
        RECT 72.535 39.680 72.825 39.725 ;
        RECT 75.055 39.680 75.345 39.725 ;
        RECT 71.345 39.540 75.345 39.680 ;
        RECT 71.345 39.495 71.635 39.540 ;
        RECT 72.535 39.495 72.825 39.540 ;
        RECT 75.055 39.495 75.345 39.540 ;
        RECT 62.645 39.340 62.935 39.385 ;
        RECT 60.790 39.200 62.935 39.340 ;
        RECT 60.790 39.140 61.110 39.200 ;
        RECT 62.645 39.155 62.935 39.200 ;
        RECT 63.565 39.155 63.855 39.385 ;
        RECT 64.010 39.140 64.330 39.400 ;
        RECT 64.485 39.155 64.775 39.385 ;
        RECT 64.930 39.340 65.250 39.400 ;
        RECT 67.245 39.340 67.535 39.385 ;
        RECT 64.930 39.200 67.535 39.340 ;
        RECT 8.350 39.045 8.670 39.060 ;
        RECT 8.320 38.815 8.670 39.045 ;
        RECT 8.350 38.800 8.670 38.815 ;
        RECT 23.070 39.000 23.390 39.060 ;
        RECT 38.220 39.000 38.510 39.045 ;
        RECT 40.090 39.000 40.410 39.060 ;
        RECT 23.070 38.860 37.100 39.000 ;
        RECT 23.070 38.800 23.390 38.860 ;
        RECT 14.790 38.460 15.110 38.720 ;
        RECT 36.960 38.660 37.100 38.860 ;
        RECT 38.220 38.860 40.410 39.000 ;
        RECT 38.220 38.815 38.510 38.860 ;
        RECT 40.090 38.800 40.410 38.860 ;
        RECT 41.470 39.000 41.790 39.060 ;
        RECT 43.310 39.000 43.630 39.060 ;
        RECT 47.450 39.045 47.770 39.060 ;
        RECT 41.470 38.860 43.630 39.000 ;
        RECT 41.470 38.800 41.790 38.860 ;
        RECT 43.310 38.800 43.630 38.860 ;
        RECT 47.420 38.815 47.770 39.045 ;
        RECT 47.450 38.800 47.770 38.815 ;
        RECT 50.670 38.800 50.990 39.060 ;
        RECT 55.700 39.000 55.990 39.045 ;
        RECT 57.570 39.000 57.890 39.060 ;
        RECT 55.700 38.860 57.890 39.000 ;
        RECT 55.700 38.815 55.990 38.860 ;
        RECT 57.570 38.800 57.890 38.860 ;
        RECT 62.170 39.000 62.490 39.060 ;
        RECT 64.560 39.000 64.700 39.155 ;
        RECT 64.930 39.140 65.250 39.200 ;
        RECT 67.245 39.155 67.535 39.200 ;
        RECT 70.450 39.340 70.770 39.400 ;
        RECT 75.510 39.340 75.830 39.400 ;
        RECT 70.450 39.200 75.830 39.340 ;
        RECT 62.170 38.860 64.700 39.000 ;
        RECT 66.325 39.000 66.615 39.045 ;
        RECT 66.325 38.860 67.000 39.000 ;
        RECT 62.170 38.800 62.490 38.860 ;
        RECT 66.325 38.815 66.615 38.860 ;
        RECT 66.860 38.720 67.000 38.860 ;
        RECT 45.165 38.660 45.455 38.705 ;
        RECT 46.530 38.660 46.850 38.720 ;
        RECT 48.370 38.660 48.690 38.720 ;
        RECT 36.960 38.520 48.690 38.660 ;
        RECT 45.165 38.475 45.455 38.520 ;
        RECT 46.530 38.460 46.850 38.520 ;
        RECT 48.370 38.460 48.690 38.520 ;
        RECT 52.985 38.660 53.275 38.705 ;
        RECT 54.350 38.660 54.670 38.720 ;
        RECT 52.985 38.520 54.670 38.660 ;
        RECT 52.985 38.475 53.275 38.520 ;
        RECT 54.350 38.460 54.670 38.520 ;
        RECT 61.265 38.660 61.555 38.705 ;
        RECT 63.090 38.660 63.410 38.720 ;
        RECT 61.265 38.520 63.410 38.660 ;
        RECT 61.265 38.475 61.555 38.520 ;
        RECT 63.090 38.460 63.410 38.520 ;
        RECT 64.010 38.660 64.330 38.720 ;
        RECT 65.390 38.660 65.710 38.720 ;
        RECT 64.010 38.520 65.710 38.660 ;
        RECT 64.010 38.460 64.330 38.520 ;
        RECT 65.390 38.460 65.710 38.520 ;
        RECT 66.770 38.460 67.090 38.720 ;
        RECT 67.320 38.660 67.460 39.155 ;
        RECT 70.450 39.140 70.770 39.200 ;
        RECT 75.510 39.140 75.830 39.200 ;
        RECT 71.800 39.000 72.090 39.045 ;
        RECT 73.670 39.000 73.990 39.060 ;
        RECT 71.800 38.860 73.990 39.000 ;
        RECT 71.800 38.815 72.090 38.860 ;
        RECT 73.670 38.800 73.990 38.860 ;
        RECT 77.365 38.660 77.655 38.705 ;
        RECT 81.030 38.660 81.350 38.720 ;
        RECT 67.320 38.520 81.350 38.660 ;
        RECT 77.365 38.475 77.655 38.520 ;
        RECT 81.030 38.460 81.350 38.520 ;
        RECT 5.520 37.840 84.180 38.320 ;
        RECT 7.905 37.640 8.195 37.685 ;
        RECT 8.350 37.640 8.670 37.700 ;
        RECT 7.905 37.500 8.670 37.640 ;
        RECT 7.905 37.455 8.195 37.500 ;
        RECT 8.350 37.440 8.670 37.500 ;
        RECT 16.645 37.640 16.935 37.685 ;
        RECT 23.990 37.640 24.310 37.700 ;
        RECT 16.645 37.500 24.310 37.640 ;
        RECT 16.645 37.455 16.935 37.500 ;
        RECT 23.990 37.440 24.310 37.500 ;
        RECT 40.090 37.440 40.410 37.700 ;
        RECT 41.945 37.640 42.235 37.685 ;
        RECT 45.150 37.640 45.470 37.700 ;
        RECT 41.945 37.500 45.470 37.640 ;
        RECT 41.945 37.455 42.235 37.500 ;
        RECT 45.150 37.440 45.470 37.500 ;
        RECT 45.625 37.640 45.915 37.685 ;
        RECT 46.990 37.640 47.310 37.700 ;
        RECT 47.925 37.640 48.215 37.685 ;
        RECT 56.650 37.640 56.970 37.700 ;
        RECT 45.625 37.500 48.215 37.640 ;
        RECT 45.625 37.455 45.915 37.500 ;
        RECT 46.990 37.440 47.310 37.500 ;
        RECT 47.925 37.455 48.215 37.500 ;
        RECT 53.060 37.500 56.970 37.640 ;
        RECT 11.585 37.300 11.875 37.345 ;
        RECT 10.280 37.160 11.875 37.300 ;
        RECT 9.285 36.775 9.575 37.005 ;
        RECT 9.360 35.940 9.500 36.775 ;
        RECT 9.730 36.760 10.050 37.020 ;
        RECT 10.280 37.005 10.420 37.160 ;
        RECT 11.585 37.115 11.875 37.160 ;
        RECT 12.490 37.300 12.810 37.360 ;
        RECT 14.330 37.300 14.650 37.360 ;
        RECT 15.265 37.300 15.555 37.345 ;
        RECT 20.770 37.300 21.090 37.360 ;
        RECT 21.705 37.300 21.995 37.345 ;
        RECT 12.490 37.160 14.100 37.300 ;
        RECT 12.490 37.100 12.810 37.160 ;
        RECT 10.205 36.775 10.495 37.005 ;
        RECT 11.125 36.775 11.415 37.005 ;
        RECT 12.950 36.960 13.270 37.020 ;
        RECT 13.960 37.005 14.100 37.160 ;
        RECT 14.330 37.160 15.555 37.300 ;
        RECT 14.330 37.100 14.650 37.160 ;
        RECT 15.265 37.115 15.555 37.160 ;
        RECT 15.800 37.160 19.160 37.300 ;
        RECT 13.425 36.960 13.715 37.005 ;
        RECT 12.950 36.820 13.715 36.960 ;
        RECT 9.820 36.280 9.960 36.760 ;
        RECT 11.200 36.620 11.340 36.775 ;
        RECT 12.950 36.760 13.270 36.820 ;
        RECT 13.425 36.775 13.715 36.820 ;
        RECT 13.885 36.775 14.175 37.005 ;
        RECT 14.790 36.760 15.110 37.020 ;
        RECT 15.800 37.005 15.940 37.160 ;
        RECT 15.800 36.820 16.135 37.005 ;
        RECT 19.020 36.960 19.160 37.160 ;
        RECT 20.770 37.160 21.995 37.300 ;
        RECT 20.770 37.100 21.090 37.160 ;
        RECT 21.705 37.115 21.995 37.160 ;
        RECT 22.610 37.300 22.930 37.360 ;
        RECT 30.890 37.300 31.210 37.360 ;
        RECT 22.610 37.160 27.440 37.300 ;
        RECT 22.610 37.100 22.930 37.160 ;
        RECT 19.020 36.820 21.000 36.960 ;
        RECT 15.845 36.775 16.135 36.820 ;
        RECT 18.470 36.620 18.790 36.680 ;
        RECT 11.200 36.480 18.790 36.620 ;
        RECT 20.860 36.620 21.000 36.820 ;
        RECT 21.230 36.760 21.550 37.020 ;
        RECT 22.165 36.960 22.455 37.005 ;
        RECT 23.070 36.960 23.390 37.020 ;
        RECT 22.165 36.820 23.390 36.960 ;
        RECT 22.165 36.775 22.455 36.820 ;
        RECT 23.070 36.760 23.390 36.820 ;
        RECT 24.925 36.775 25.215 37.005 ;
        RECT 25.845 36.960 26.135 37.005 ;
        RECT 26.750 36.960 27.070 37.020 ;
        RECT 25.845 36.820 27.070 36.960 ;
        RECT 27.300 36.960 27.440 37.160 ;
        RECT 30.890 37.160 35.260 37.300 ;
        RECT 30.890 37.100 31.210 37.160 ;
        RECT 35.120 37.005 35.260 37.160 ;
        RECT 46.530 37.100 46.850 37.360 ;
        RECT 53.060 37.300 53.200 37.500 ;
        RECT 56.650 37.440 56.970 37.500 ;
        RECT 57.570 37.440 57.890 37.700 ;
        RECT 75.985 37.455 76.275 37.685 ;
        RECT 48.000 37.160 53.200 37.300 ;
        RECT 53.445 37.300 53.735 37.345 ;
        RECT 61.250 37.300 61.570 37.360 ;
        RECT 53.445 37.160 61.570 37.300 ;
        RECT 34.585 36.960 34.875 37.005 ;
        RECT 27.300 36.820 34.875 36.960 ;
        RECT 25.845 36.775 26.135 36.820 ;
        RECT 25.000 36.620 25.140 36.775 ;
        RECT 26.750 36.760 27.070 36.820 ;
        RECT 34.585 36.775 34.875 36.820 ;
        RECT 35.045 36.775 35.335 37.005 ;
        RECT 35.950 36.760 36.270 37.020 ;
        RECT 36.425 36.960 36.715 37.005 ;
        RECT 48.000 36.960 48.140 37.160 ;
        RECT 53.445 37.115 53.735 37.160 ;
        RECT 61.250 37.100 61.570 37.160 ;
        RECT 63.550 37.300 63.870 37.360 ;
        RECT 76.060 37.300 76.200 37.455 ;
        RECT 63.550 37.160 67.460 37.300 ;
        RECT 63.550 37.100 63.870 37.160 ;
        RECT 36.425 36.820 48.140 36.960 ;
        RECT 48.385 36.960 48.675 37.005 ;
        RECT 49.290 36.960 49.610 37.020 ;
        RECT 54.350 36.960 54.670 37.020 ;
        RECT 48.385 36.820 54.670 36.960 ;
        RECT 36.425 36.775 36.715 36.820 ;
        RECT 48.385 36.775 48.675 36.820 ;
        RECT 49.290 36.760 49.610 36.820 ;
        RECT 54.350 36.760 54.670 36.820 ;
        RECT 54.810 36.760 55.130 37.020 ;
        RECT 58.950 36.760 59.270 37.020 ;
        RECT 59.425 36.775 59.715 37.005 ;
        RECT 59.885 36.775 60.175 37.005 ;
        RECT 27.210 36.620 27.530 36.680 ;
        RECT 20.860 36.480 27.530 36.620 ;
        RECT 18.470 36.420 18.790 36.480 ;
        RECT 27.210 36.420 27.530 36.480 ;
        RECT 41.930 36.620 42.250 36.680 ;
        RECT 42.405 36.620 42.695 36.665 ;
        RECT 41.930 36.480 42.695 36.620 ;
        RECT 41.930 36.420 42.250 36.480 ;
        RECT 42.405 36.435 42.695 36.480 ;
        RECT 43.310 36.420 43.630 36.680 ;
        RECT 49.765 36.620 50.055 36.665 ;
        RECT 50.670 36.620 50.990 36.680 ;
        RECT 49.765 36.480 50.990 36.620 ;
        RECT 49.765 36.435 50.055 36.480 ;
        RECT 50.670 36.420 50.990 36.480 ;
        RECT 53.430 36.620 53.750 36.680 ;
        RECT 53.905 36.620 54.195 36.665 ;
        RECT 59.500 36.620 59.640 36.775 ;
        RECT 53.430 36.480 54.195 36.620 ;
        RECT 53.430 36.420 53.750 36.480 ;
        RECT 53.905 36.435 54.195 36.480 ;
        RECT 54.440 36.480 59.640 36.620 ;
        RECT 59.960 36.620 60.100 36.775 ;
        RECT 60.790 36.760 61.110 37.020 ;
        RECT 61.710 36.760 62.030 37.020 ;
        RECT 62.645 36.960 62.935 37.005 ;
        RECT 63.090 36.960 63.410 37.020 ;
        RECT 64.100 37.005 64.240 37.160 ;
        RECT 62.645 36.820 63.410 36.960 ;
        RECT 62.645 36.775 62.935 36.820 ;
        RECT 63.090 36.760 63.410 36.820 ;
        RECT 64.025 36.775 64.315 37.005 ;
        RECT 64.470 36.960 64.790 37.020 ;
        RECT 67.320 37.005 67.460 37.160 ;
        RECT 72.380 37.160 76.200 37.300 ;
        RECT 64.945 36.960 65.235 37.005 ;
        RECT 66.325 36.960 66.615 37.005 ;
        RECT 64.470 36.820 66.615 36.960 ;
        RECT 64.470 36.760 64.790 36.820 ;
        RECT 64.945 36.775 65.235 36.820 ;
        RECT 66.325 36.775 66.615 36.820 ;
        RECT 67.245 36.960 67.535 37.005 ;
        RECT 67.690 36.960 68.010 37.020 ;
        RECT 67.245 36.820 68.010 36.960 ;
        RECT 67.245 36.775 67.535 36.820 ;
        RECT 67.690 36.760 68.010 36.820 ;
        RECT 71.370 36.960 71.690 37.020 ;
        RECT 72.380 37.005 72.520 37.160 ;
        RECT 72.305 36.960 72.595 37.005 ;
        RECT 71.370 36.820 72.595 36.960 ;
        RECT 71.370 36.760 71.690 36.820 ;
        RECT 72.305 36.775 72.595 36.820 ;
        RECT 73.210 36.760 73.530 37.020 ;
        RECT 73.685 36.775 73.975 37.005 ;
        RECT 74.145 36.960 74.435 37.005 ;
        RECT 74.590 36.960 74.910 37.020 ;
        RECT 74.145 36.820 74.910 36.960 ;
        RECT 74.145 36.775 74.435 36.820 ;
        RECT 63.565 36.620 63.855 36.665 ;
        RECT 59.960 36.480 63.855 36.620 ;
        RECT 33.665 36.280 33.955 36.325 ;
        RECT 52.970 36.280 53.290 36.340 ;
        RECT 9.820 36.140 33.420 36.280 ;
        RECT 13.410 35.940 13.730 36.000 ;
        RECT 14.790 35.940 15.110 36.000 ;
        RECT 9.360 35.800 15.110 35.940 ;
        RECT 13.410 35.740 13.730 35.800 ;
        RECT 14.790 35.740 15.110 35.800 ;
        RECT 23.070 35.940 23.390 36.000 ;
        RECT 24.005 35.940 24.295 35.985 ;
        RECT 23.070 35.800 24.295 35.940 ;
        RECT 33.280 35.940 33.420 36.140 ;
        RECT 33.665 36.140 53.290 36.280 ;
        RECT 33.665 36.095 33.955 36.140 ;
        RECT 52.970 36.080 53.290 36.140 ;
        RECT 42.850 35.940 43.170 36.000 ;
        RECT 33.280 35.800 43.170 35.940 ;
        RECT 23.070 35.740 23.390 35.800 ;
        RECT 24.005 35.755 24.295 35.800 ;
        RECT 42.850 35.740 43.170 35.800 ;
        RECT 44.690 35.740 45.010 36.000 ;
        RECT 45.150 35.940 45.470 36.000 ;
        RECT 45.625 35.940 45.915 35.985 ;
        RECT 45.150 35.800 45.915 35.940 ;
        RECT 45.150 35.740 45.470 35.800 ;
        RECT 45.625 35.755 45.915 35.800 ;
        RECT 52.510 35.940 52.830 36.000 ;
        RECT 54.440 35.940 54.580 36.480 ;
        RECT 63.565 36.435 63.855 36.480 ;
        RECT 65.390 36.620 65.710 36.680 ;
        RECT 71.830 36.620 72.150 36.680 ;
        RECT 73.760 36.620 73.900 36.775 ;
        RECT 74.590 36.760 74.910 36.820 ;
        RECT 76.890 36.760 77.210 37.020 ;
        RECT 65.390 36.480 73.900 36.620 ;
        RECT 65.390 36.420 65.710 36.480 ;
        RECT 71.830 36.420 72.150 36.480 ;
        RECT 61.710 36.280 62.030 36.340 ;
        RECT 72.290 36.280 72.610 36.340 ;
        RECT 55.820 36.140 62.030 36.280 ;
        RECT 52.510 35.800 54.580 35.940 ;
        RECT 55.270 35.940 55.590 36.000 ;
        RECT 55.820 35.985 55.960 36.140 ;
        RECT 61.710 36.080 62.030 36.140 ;
        RECT 64.100 36.140 72.610 36.280 ;
        RECT 55.745 35.940 56.035 35.985 ;
        RECT 55.270 35.800 56.035 35.940 ;
        RECT 52.510 35.740 52.830 35.800 ;
        RECT 55.270 35.740 55.590 35.800 ;
        RECT 55.745 35.755 56.035 35.800 ;
        RECT 58.950 35.940 59.270 36.000 ;
        RECT 64.100 35.940 64.240 36.140 ;
        RECT 72.290 36.080 72.610 36.140 ;
        RECT 75.525 36.280 75.815 36.325 ;
        RECT 76.890 36.280 77.210 36.340 ;
        RECT 75.525 36.140 77.210 36.280 ;
        RECT 75.525 36.095 75.815 36.140 ;
        RECT 76.890 36.080 77.210 36.140 ;
        RECT 58.950 35.800 64.240 35.940 ;
        RECT 58.950 35.740 59.270 35.800 ;
        RECT 64.470 35.740 64.790 36.000 ;
        RECT 67.230 35.940 67.550 36.000 ;
        RECT 68.165 35.940 68.455 35.985 ;
        RECT 67.230 35.800 68.455 35.940 ;
        RECT 67.230 35.740 67.550 35.800 ;
        RECT 68.165 35.755 68.455 35.800 ;
        RECT 5.520 35.120 84.180 35.600 ;
        RECT 13.870 34.920 14.190 34.980 ;
        RECT 15.250 34.920 15.570 34.980 ;
        RECT 27.225 34.920 27.515 34.965 ;
        RECT 13.870 34.780 15.570 34.920 ;
        RECT 13.870 34.720 14.190 34.780 ;
        RECT 15.250 34.720 15.570 34.780 ;
        RECT 23.160 34.780 27.515 34.920 ;
        RECT 10.690 34.580 10.980 34.625 ;
        RECT 12.790 34.580 13.080 34.625 ;
        RECT 14.360 34.580 14.650 34.625 ;
        RECT 10.690 34.440 14.650 34.580 ;
        RECT 10.690 34.395 10.980 34.440 ;
        RECT 12.790 34.395 13.080 34.440 ;
        RECT 14.360 34.395 14.650 34.440 ;
        RECT 8.810 34.240 9.130 34.300 ;
        RECT 10.190 34.240 10.510 34.300 ;
        RECT 8.810 34.100 10.510 34.240 ;
        RECT 8.810 34.040 9.130 34.100 ;
        RECT 10.190 34.040 10.510 34.100 ;
        RECT 11.085 34.240 11.375 34.285 ;
        RECT 12.275 34.240 12.565 34.285 ;
        RECT 14.795 34.240 15.085 34.285 ;
        RECT 11.085 34.100 15.085 34.240 ;
        RECT 23.160 34.240 23.300 34.780 ;
        RECT 23.160 34.100 23.760 34.240 ;
        RECT 11.085 34.055 11.375 34.100 ;
        RECT 12.275 34.055 12.565 34.100 ;
        RECT 14.795 34.055 15.085 34.100 ;
        RECT 18.930 33.900 19.250 33.960 ;
        RECT 22.150 33.900 22.470 33.960 ;
        RECT 18.930 33.760 22.470 33.900 ;
        RECT 18.930 33.700 19.250 33.760 ;
        RECT 22.150 33.700 22.470 33.760 ;
        RECT 22.610 33.900 22.930 33.960 ;
        RECT 23.620 33.945 23.760 34.100 ;
        RECT 26.840 33.960 26.980 34.780 ;
        RECT 27.225 34.735 27.515 34.780 ;
        RECT 47.450 34.720 47.770 34.980 ;
        RECT 69.545 34.920 69.835 34.965 ;
        RECT 73.210 34.920 73.530 34.980 ;
        RECT 69.545 34.780 73.530 34.920 ;
        RECT 69.545 34.735 69.835 34.780 ;
        RECT 73.210 34.720 73.530 34.780 ;
        RECT 32.730 34.580 33.020 34.625 ;
        RECT 34.300 34.580 34.590 34.625 ;
        RECT 36.400 34.580 36.690 34.625 ;
        RECT 32.730 34.440 36.690 34.580 ;
        RECT 32.730 34.395 33.020 34.440 ;
        RECT 34.300 34.395 34.590 34.440 ;
        RECT 36.400 34.395 36.690 34.440 ;
        RECT 41.930 34.580 42.250 34.640 ;
        RECT 66.770 34.580 67.090 34.640 ;
        RECT 41.930 34.440 67.090 34.580 ;
        RECT 41.930 34.380 42.250 34.440 ;
        RECT 66.770 34.380 67.090 34.440 ;
        RECT 75.550 34.580 75.840 34.625 ;
        RECT 77.650 34.580 77.940 34.625 ;
        RECT 79.220 34.580 79.510 34.625 ;
        RECT 75.550 34.440 79.510 34.580 ;
        RECT 75.550 34.395 75.840 34.440 ;
        RECT 77.650 34.395 77.940 34.440 ;
        RECT 79.220 34.395 79.510 34.440 ;
        RECT 32.295 34.240 32.585 34.285 ;
        RECT 34.815 34.240 35.105 34.285 ;
        RECT 36.005 34.240 36.295 34.285 ;
        RECT 32.295 34.100 36.295 34.240 ;
        RECT 32.295 34.055 32.585 34.100 ;
        RECT 34.815 34.055 35.105 34.100 ;
        RECT 36.005 34.055 36.295 34.100 ;
        RECT 43.310 34.240 43.630 34.300 ;
        RECT 50.225 34.240 50.515 34.285 ;
        RECT 43.310 34.100 50.515 34.240 ;
        RECT 43.310 34.040 43.630 34.100 ;
        RECT 50.225 34.055 50.515 34.100 ;
        RECT 54.350 34.040 54.670 34.300 ;
        RECT 74.590 34.240 74.910 34.300 ;
        RECT 73.300 34.100 74.910 34.240 ;
        RECT 23.085 33.900 23.375 33.945 ;
        RECT 22.610 33.760 23.375 33.900 ;
        RECT 22.610 33.700 22.930 33.760 ;
        RECT 23.085 33.715 23.375 33.760 ;
        RECT 23.545 33.715 23.835 33.945 ;
        RECT 23.990 33.700 24.310 33.960 ;
        RECT 26.290 33.700 26.610 33.960 ;
        RECT 26.750 33.700 27.070 33.960 ;
        RECT 27.210 33.900 27.530 33.960 ;
        RECT 27.685 33.900 27.975 33.945 ;
        RECT 32.730 33.900 33.050 33.960 ;
        RECT 36.870 33.900 37.190 33.960 ;
        RECT 27.210 33.760 33.050 33.900 ;
        RECT 27.210 33.700 27.530 33.760 ;
        RECT 27.685 33.715 27.975 33.760 ;
        RECT 32.730 33.700 33.050 33.760 ;
        RECT 34.660 33.760 37.190 33.900 ;
        RECT 11.540 33.560 11.830 33.605 ;
        RECT 13.410 33.560 13.730 33.620 ;
        RECT 19.865 33.560 20.155 33.605 ;
        RECT 11.540 33.420 13.730 33.560 ;
        RECT 11.540 33.375 11.830 33.420 ;
        RECT 13.410 33.360 13.730 33.420 ;
        RECT 17.180 33.420 20.155 33.560 ;
        RECT 14.330 33.220 14.650 33.280 ;
        RECT 17.180 33.265 17.320 33.420 ;
        RECT 19.865 33.375 20.155 33.420 ;
        RECT 20.770 33.360 21.090 33.620 ;
        RECT 24.080 33.560 24.220 33.700 ;
        RECT 34.660 33.620 34.800 33.760 ;
        RECT 36.870 33.700 37.190 33.760 ;
        RECT 38.725 33.715 39.015 33.945 ;
        RECT 24.080 33.420 30.660 33.560 ;
        RECT 17.105 33.220 17.395 33.265 ;
        RECT 14.330 33.080 17.395 33.220 ;
        RECT 14.330 33.020 14.650 33.080 ;
        RECT 17.105 33.035 17.395 33.080 ;
        RECT 18.930 33.020 19.250 33.280 ;
        RECT 20.860 33.220 21.000 33.360 ;
        RECT 23.070 33.220 23.390 33.280 ;
        RECT 20.860 33.080 23.390 33.220 ;
        RECT 23.070 33.020 23.390 33.080 ;
        RECT 23.530 33.220 23.850 33.280 ;
        RECT 25.385 33.220 25.675 33.265 ;
        RECT 23.530 33.080 25.675 33.220 ;
        RECT 23.530 33.020 23.850 33.080 ;
        RECT 25.385 33.035 25.675 33.080 ;
        RECT 29.970 33.020 30.290 33.280 ;
        RECT 30.520 33.220 30.660 33.420 ;
        RECT 34.570 33.360 34.890 33.620 ;
        RECT 35.660 33.560 35.950 33.605 ;
        RECT 37.345 33.560 37.635 33.605 ;
        RECT 35.660 33.420 37.635 33.560 ;
        RECT 35.660 33.375 35.950 33.420 ;
        RECT 37.345 33.375 37.635 33.420 ;
        RECT 38.800 33.560 38.940 33.715 ;
        RECT 39.170 33.700 39.490 33.960 ;
        RECT 39.630 33.700 39.950 33.960 ;
        RECT 40.090 33.900 40.410 33.960 ;
        RECT 40.565 33.900 40.855 33.945 ;
        RECT 58.950 33.900 59.270 33.960 ;
        RECT 40.090 33.760 40.855 33.900 ;
        RECT 40.090 33.700 40.410 33.760 ;
        RECT 40.565 33.715 40.855 33.760 ;
        RECT 48.920 33.760 59.270 33.900 ;
        RECT 48.920 33.560 49.060 33.760 ;
        RECT 58.950 33.700 59.270 33.760 ;
        RECT 71.370 33.700 71.690 33.960 ;
        RECT 72.290 33.700 72.610 33.960 ;
        RECT 73.300 33.945 73.440 34.100 ;
        RECT 74.590 34.040 74.910 34.100 ;
        RECT 75.945 34.240 76.235 34.285 ;
        RECT 77.135 34.240 77.425 34.285 ;
        RECT 79.655 34.240 79.945 34.285 ;
        RECT 75.945 34.100 79.945 34.240 ;
        RECT 75.945 34.055 76.235 34.100 ;
        RECT 77.135 34.055 77.425 34.100 ;
        RECT 79.655 34.055 79.945 34.100 ;
        RECT 72.765 33.715 73.055 33.945 ;
        RECT 73.225 33.715 73.515 33.945 ;
        RECT 75.065 33.900 75.355 33.945 ;
        RECT 75.510 33.900 75.830 33.960 ;
        RECT 75.065 33.760 75.830 33.900 ;
        RECT 75.065 33.715 75.355 33.760 ;
        RECT 38.800 33.420 49.060 33.560 ;
        RECT 49.305 33.560 49.595 33.605 ;
        RECT 51.605 33.560 51.895 33.605 ;
        RECT 49.305 33.420 51.895 33.560 ;
        RECT 38.800 33.220 38.940 33.420 ;
        RECT 49.305 33.375 49.595 33.420 ;
        RECT 51.605 33.375 51.895 33.420 ;
        RECT 55.730 33.360 56.050 33.620 ;
        RECT 67.230 33.560 67.550 33.620 ;
        RECT 67.705 33.560 67.995 33.605 ;
        RECT 67.230 33.420 67.995 33.560 ;
        RECT 67.230 33.360 67.550 33.420 ;
        RECT 67.705 33.375 67.995 33.420 ;
        RECT 68.625 33.560 68.915 33.605 ;
        RECT 71.830 33.560 72.150 33.620 ;
        RECT 68.625 33.420 72.150 33.560 ;
        RECT 68.625 33.375 68.915 33.420 ;
        RECT 71.830 33.360 72.150 33.420 ;
        RECT 30.520 33.080 38.940 33.220 ;
        RECT 49.765 33.220 50.055 33.265 ;
        RECT 50.210 33.220 50.530 33.280 ;
        RECT 49.765 33.080 50.530 33.220 ;
        RECT 49.765 33.035 50.055 33.080 ;
        RECT 50.210 33.020 50.530 33.080 ;
        RECT 56.190 33.020 56.510 33.280 ;
        RECT 66.310 33.220 66.630 33.280 ;
        RECT 72.840 33.220 72.980 33.715 ;
        RECT 75.510 33.700 75.830 33.760 ;
        RECT 74.605 33.560 74.895 33.605 ;
        RECT 76.290 33.560 76.580 33.605 ;
        RECT 74.605 33.420 76.580 33.560 ;
        RECT 74.605 33.375 74.895 33.420 ;
        RECT 76.290 33.375 76.580 33.420 ;
        RECT 66.310 33.080 72.980 33.220 ;
        RECT 79.190 33.220 79.510 33.280 ;
        RECT 81.965 33.220 82.255 33.265 ;
        RECT 79.190 33.080 82.255 33.220 ;
        RECT 66.310 33.020 66.630 33.080 ;
        RECT 79.190 33.020 79.510 33.080 ;
        RECT 81.965 33.035 82.255 33.080 ;
        RECT 5.520 32.400 84.180 32.880 ;
        RECT 13.410 32.000 13.730 32.260 ;
        RECT 22.610 32.000 22.930 32.260 ;
        RECT 23.070 32.200 23.390 32.260 ;
        RECT 26.290 32.200 26.610 32.260 ;
        RECT 23.070 32.060 26.610 32.200 ;
        RECT 23.070 32.000 23.390 32.060 ;
        RECT 26.290 32.000 26.610 32.060 ;
        RECT 34.585 32.200 34.875 32.245 ;
        RECT 35.030 32.200 35.350 32.260 ;
        RECT 34.585 32.060 35.350 32.200 ;
        RECT 34.585 32.015 34.875 32.060 ;
        RECT 35.030 32.000 35.350 32.060 ;
        RECT 36.885 32.200 37.175 32.245 ;
        RECT 39.630 32.200 39.950 32.260 ;
        RECT 36.885 32.060 39.950 32.200 ;
        RECT 36.885 32.015 37.175 32.060 ;
        RECT 39.630 32.000 39.950 32.060 ;
        RECT 43.310 32.200 43.630 32.260 ;
        RECT 45.165 32.200 45.455 32.245 ;
        RECT 55.730 32.200 56.050 32.260 ;
        RECT 43.310 32.060 56.050 32.200 ;
        RECT 43.310 32.000 43.630 32.060 ;
        RECT 45.165 32.015 45.455 32.060 ;
        RECT 55.730 32.000 56.050 32.060 ;
        RECT 59.410 32.200 59.730 32.260 ;
        RECT 70.925 32.200 71.215 32.245 ;
        RECT 72.290 32.200 72.610 32.260 ;
        RECT 81.030 32.200 81.350 32.260 ;
        RECT 82.425 32.200 82.715 32.245 ;
        RECT 59.410 32.060 67.920 32.200 ;
        RECT 59.410 32.000 59.730 32.060 ;
        RECT 67.780 31.920 67.920 32.060 ;
        RECT 70.925 32.060 72.610 32.200 ;
        RECT 70.925 32.015 71.215 32.060 ;
        RECT 72.290 32.000 72.610 32.060 ;
        RECT 72.840 32.060 82.715 32.200 ;
        RECT 18.930 31.860 19.250 31.920 ;
        RECT 22.150 31.860 22.470 31.920 ;
        RECT 27.210 31.860 27.530 31.920 ;
        RECT 15.800 31.720 19.250 31.860 ;
        RECT 14.790 31.320 15.110 31.580 ;
        RECT 15.250 31.320 15.570 31.580 ;
        RECT 15.800 31.565 15.940 31.720 ;
        RECT 18.930 31.660 19.250 31.720 ;
        RECT 19.480 31.720 22.470 31.860 ;
        RECT 15.725 31.335 16.015 31.565 ;
        RECT 16.645 31.335 16.935 31.565 ;
        RECT 17.105 31.520 17.395 31.565 ;
        RECT 19.480 31.520 19.620 31.720 ;
        RECT 22.150 31.660 22.470 31.720 ;
        RECT 23.160 31.720 27.530 31.860 ;
        RECT 17.105 31.380 19.620 31.520 ;
        RECT 17.105 31.335 17.395 31.380 ;
        RECT 16.720 31.180 16.860 31.335 ;
        RECT 20.770 31.320 21.090 31.580 ;
        RECT 23.160 31.565 23.300 31.720 ;
        RECT 27.210 31.660 27.530 31.720 ;
        RECT 29.970 31.860 30.290 31.920 ;
        RECT 33.205 31.860 33.495 31.905 ;
        RECT 35.965 31.860 36.255 31.905 ;
        RECT 29.970 31.720 36.255 31.860 ;
        RECT 29.970 31.660 30.290 31.720 ;
        RECT 33.205 31.675 33.495 31.720 ;
        RECT 35.965 31.675 36.255 31.720 ;
        RECT 47.910 31.860 48.230 31.920 ;
        RECT 61.710 31.860 62.030 31.920 ;
        RECT 47.910 31.720 62.030 31.860 ;
        RECT 47.910 31.660 48.230 31.720 ;
        RECT 61.710 31.660 62.030 31.720 ;
        RECT 67.690 31.860 68.010 31.920 ;
        RECT 71.830 31.860 72.150 31.920 ;
        RECT 72.840 31.905 72.980 32.060 ;
        RECT 81.030 32.000 81.350 32.060 ;
        RECT 82.425 32.015 82.715 32.060 ;
        RECT 76.890 31.905 77.210 31.920 ;
        RECT 72.765 31.860 73.055 31.905 ;
        RECT 76.860 31.860 77.210 31.905 ;
        RECT 67.690 31.720 70.680 31.860 ;
        RECT 67.690 31.660 68.010 31.720 ;
        RECT 21.705 31.520 21.995 31.565 ;
        RECT 21.705 31.380 22.840 31.520 ;
        RECT 21.705 31.335 21.995 31.380 ;
        RECT 16.720 31.040 18.240 31.180 ;
        RECT 18.100 30.545 18.240 31.040 ;
        RECT 18.025 30.500 18.315 30.545 ;
        RECT 19.390 30.500 19.710 30.560 ;
        RECT 18.025 30.360 19.710 30.500 ;
        RECT 22.700 30.500 22.840 31.380 ;
        RECT 23.085 31.335 23.375 31.565 ;
        RECT 23.530 31.520 23.850 31.580 ;
        RECT 24.365 31.520 24.655 31.565 ;
        RECT 31.825 31.520 32.115 31.565 ;
        RECT 23.530 31.380 24.655 31.520 ;
        RECT 23.530 31.320 23.850 31.380 ;
        RECT 24.365 31.335 24.655 31.380 ;
        RECT 30.060 31.380 32.115 31.520 ;
        RECT 23.965 31.180 24.255 31.225 ;
        RECT 25.155 31.180 25.445 31.225 ;
        RECT 27.675 31.180 27.965 31.225 ;
        RECT 23.965 31.040 27.965 31.180 ;
        RECT 23.965 30.995 24.255 31.040 ;
        RECT 25.155 30.995 25.445 31.040 ;
        RECT 27.675 30.995 27.965 31.040 ;
        RECT 23.570 30.840 23.860 30.885 ;
        RECT 25.670 30.840 25.960 30.885 ;
        RECT 27.240 30.840 27.530 30.885 ;
        RECT 23.570 30.700 27.530 30.840 ;
        RECT 23.570 30.655 23.860 30.700 ;
        RECT 25.670 30.655 25.960 30.700 ;
        RECT 27.240 30.655 27.530 30.700 ;
        RECT 23.990 30.500 24.310 30.560 ;
        RECT 30.060 30.545 30.200 31.380 ;
        RECT 31.825 31.335 32.115 31.380 ;
        RECT 32.730 31.320 33.050 31.580 ;
        RECT 33.665 31.335 33.955 31.565 ;
        RECT 32.820 30.840 32.960 31.320 ;
        RECT 33.740 31.180 33.880 31.335 ;
        RECT 35.030 31.320 35.350 31.580 ;
        RECT 44.230 31.520 44.550 31.580 ;
        RECT 44.705 31.520 44.995 31.565 ;
        RECT 44.230 31.380 44.995 31.520 ;
        RECT 44.230 31.320 44.550 31.380 ;
        RECT 44.705 31.335 44.995 31.380 ;
        RECT 45.150 31.520 45.470 31.580 ;
        RECT 46.085 31.520 46.375 31.565 ;
        RECT 45.150 31.380 46.375 31.520 ;
        RECT 45.150 31.320 45.470 31.380 ;
        RECT 46.085 31.335 46.375 31.380 ;
        RECT 46.990 31.320 47.310 31.580 ;
        RECT 49.290 31.520 49.610 31.580 ;
        RECT 51.045 31.520 51.335 31.565 ;
        RECT 49.290 31.380 51.335 31.520 ;
        RECT 49.290 31.320 49.610 31.380 ;
        RECT 51.045 31.335 51.335 31.380 ;
        RECT 56.190 31.520 56.510 31.580 ;
        RECT 63.105 31.520 63.395 31.565 ;
        RECT 64.485 31.520 64.775 31.565 ;
        RECT 56.190 31.380 64.775 31.520 ;
        RECT 56.190 31.320 56.510 31.380 ;
        RECT 35.490 31.180 35.810 31.240 ;
        RECT 33.740 31.040 35.810 31.180 ;
        RECT 35.490 30.980 35.810 31.040 ;
        RECT 49.765 30.995 50.055 31.225 ;
        RECT 50.645 31.180 50.935 31.225 ;
        RECT 51.835 31.180 52.125 31.225 ;
        RECT 54.355 31.180 54.645 31.225 ;
        RECT 50.645 31.040 54.645 31.180 ;
        RECT 50.645 30.995 50.935 31.040 ;
        RECT 51.835 30.995 52.125 31.040 ;
        RECT 54.355 30.995 54.645 31.040 ;
        RECT 44.690 30.840 45.010 30.900 ;
        RECT 32.820 30.700 45.010 30.840 ;
        RECT 44.690 30.640 45.010 30.700 ;
        RECT 29.985 30.500 30.275 30.545 ;
        RECT 22.700 30.360 30.275 30.500 ;
        RECT 49.840 30.500 49.980 30.995 ;
        RECT 50.250 30.840 50.540 30.885 ;
        RECT 52.350 30.840 52.640 30.885 ;
        RECT 53.920 30.840 54.210 30.885 ;
        RECT 50.250 30.700 54.210 30.840 ;
        RECT 50.250 30.655 50.540 30.700 ;
        RECT 52.350 30.655 52.640 30.700 ;
        RECT 53.920 30.655 54.210 30.700 ;
        RECT 50.670 30.500 50.990 30.560 ;
        RECT 49.840 30.360 50.990 30.500 ;
        RECT 18.025 30.315 18.315 30.360 ;
        RECT 19.390 30.300 19.710 30.360 ;
        RECT 23.990 30.300 24.310 30.360 ;
        RECT 29.985 30.315 30.275 30.360 ;
        RECT 50.670 30.300 50.990 30.360 ;
        RECT 51.130 30.500 51.450 30.560 ;
        RECT 56.665 30.500 56.955 30.545 ;
        RECT 57.110 30.500 57.430 30.560 ;
        RECT 51.130 30.360 57.430 30.500 ;
        RECT 61.800 30.500 61.940 31.380 ;
        RECT 63.105 31.335 63.395 31.380 ;
        RECT 64.485 31.335 64.775 31.380 ;
        RECT 65.405 31.335 65.695 31.565 ;
        RECT 69.085 31.335 69.375 31.565 ;
        RECT 69.530 31.520 69.850 31.580 ;
        RECT 70.005 31.520 70.295 31.565 ;
        RECT 69.530 31.380 70.295 31.520 ;
        RECT 70.540 31.520 70.680 31.720 ;
        RECT 71.830 31.720 73.055 31.860 ;
        RECT 76.695 31.720 77.210 31.860 ;
        RECT 71.830 31.660 72.150 31.720 ;
        RECT 72.765 31.675 73.055 31.720 ;
        RECT 76.860 31.675 77.210 31.720 ;
        RECT 76.890 31.660 77.210 31.675 ;
        RECT 72.290 31.520 72.610 31.580 ;
        RECT 70.540 31.380 72.610 31.520 ;
        RECT 64.010 31.180 64.330 31.240 ;
        RECT 65.480 31.180 65.620 31.335 ;
        RECT 64.010 31.040 65.620 31.180 ;
        RECT 64.010 30.980 64.330 31.040 ;
        RECT 66.310 30.980 66.630 31.240 ;
        RECT 69.160 30.900 69.300 31.335 ;
        RECT 69.530 31.320 69.850 31.380 ;
        RECT 70.005 31.335 70.295 31.380 ;
        RECT 72.290 31.320 72.610 31.380 ;
        RECT 73.210 31.320 73.530 31.580 ;
        RECT 74.130 31.520 74.450 31.580 ;
        RECT 79.190 31.520 79.510 31.580 ;
        RECT 74.130 31.380 79.510 31.520 ;
        RECT 74.130 31.320 74.450 31.380 ;
        RECT 79.190 31.320 79.510 31.380 ;
        RECT 75.510 30.980 75.830 31.240 ;
        RECT 76.405 31.180 76.695 31.225 ;
        RECT 77.595 31.180 77.885 31.225 ;
        RECT 80.115 31.180 80.405 31.225 ;
        RECT 76.405 31.040 80.405 31.180 ;
        RECT 76.405 30.995 76.695 31.040 ;
        RECT 77.595 30.995 77.885 31.040 ;
        RECT 80.115 30.995 80.405 31.040 ;
        RECT 62.185 30.840 62.475 30.885 ;
        RECT 69.070 30.840 69.390 30.900 ;
        RECT 62.185 30.700 69.390 30.840 ;
        RECT 62.185 30.655 62.475 30.700 ;
        RECT 69.070 30.640 69.390 30.700 ;
        RECT 69.990 30.840 70.310 30.900 ;
        RECT 71.385 30.840 71.675 30.885 ;
        RECT 69.990 30.700 71.675 30.840 ;
        RECT 69.990 30.640 70.310 30.700 ;
        RECT 71.385 30.655 71.675 30.700 ;
        RECT 72.290 30.840 72.610 30.900 ;
        RECT 74.590 30.840 74.910 30.900 ;
        RECT 72.290 30.700 74.910 30.840 ;
        RECT 72.290 30.640 72.610 30.700 ;
        RECT 74.590 30.640 74.910 30.700 ;
        RECT 76.010 30.840 76.300 30.885 ;
        RECT 78.110 30.840 78.400 30.885 ;
        RECT 79.680 30.840 79.970 30.885 ;
        RECT 76.010 30.700 79.970 30.840 ;
        RECT 76.010 30.655 76.300 30.700 ;
        RECT 78.110 30.655 78.400 30.700 ;
        RECT 79.680 30.655 79.970 30.700 ;
        RECT 73.210 30.500 73.530 30.560 ;
        RECT 61.800 30.360 73.530 30.500 ;
        RECT 51.130 30.300 51.450 30.360 ;
        RECT 56.665 30.315 56.955 30.360 ;
        RECT 57.110 30.300 57.430 30.360 ;
        RECT 73.210 30.300 73.530 30.360 ;
        RECT 5.520 29.680 84.180 30.160 ;
        RECT 13.730 29.340 43.540 29.480 ;
        RECT 11.110 29.140 11.430 29.200 ;
        RECT 12.950 29.140 13.270 29.200 ;
        RECT 13.730 29.140 13.870 29.340 ;
        RECT 11.110 29.000 13.870 29.140 ;
        RECT 15.250 29.140 15.570 29.200 ;
        RECT 15.250 29.000 15.940 29.140 ;
        RECT 11.110 28.940 11.430 29.000 ;
        RECT 12.950 28.940 13.270 29.000 ;
        RECT 15.250 28.940 15.570 29.000 ;
        RECT 14.330 28.800 14.650 28.860 ;
        RECT 8.440 28.660 14.650 28.800 ;
        RECT 8.440 28.505 8.580 28.660 ;
        RECT 14.330 28.600 14.650 28.660 ;
        RECT 15.800 28.800 15.940 29.000 ;
        RECT 35.030 28.940 35.350 29.200 ;
        RECT 43.400 29.140 43.540 29.340 ;
        RECT 43.770 29.280 44.090 29.540 ;
        RECT 49.290 29.280 49.610 29.540 ;
        RECT 60.880 29.340 68.840 29.480 ;
        RECT 52.550 29.140 52.840 29.185 ;
        RECT 54.650 29.140 54.940 29.185 ;
        RECT 56.220 29.140 56.510 29.185 ;
        RECT 43.400 29.000 50.440 29.140 ;
        RECT 26.750 28.800 27.070 28.860 ;
        RECT 35.120 28.800 35.260 28.940 ;
        RECT 41.930 28.800 42.250 28.860 ;
        RECT 44.230 28.800 44.550 28.860 ;
        RECT 49.765 28.800 50.055 28.845 ;
        RECT 15.800 28.660 27.070 28.800 ;
        RECT 8.365 28.275 8.655 28.505 ;
        RECT 8.810 28.460 9.130 28.520 ;
        RECT 11.110 28.460 11.430 28.520 ;
        RECT 8.810 28.320 11.430 28.460 ;
        RECT 8.810 28.260 9.130 28.320 ;
        RECT 11.110 28.260 11.430 28.320 ;
        RECT 11.570 28.460 11.890 28.520 ;
        RECT 15.800 28.505 15.940 28.660 ;
        RECT 26.750 28.600 27.070 28.660 ;
        RECT 34.660 28.660 42.250 28.800 ;
        RECT 15.265 28.460 15.555 28.505 ;
        RECT 11.570 28.320 15.555 28.460 ;
        RECT 11.570 28.260 11.890 28.320 ;
        RECT 15.265 28.275 15.555 28.320 ;
        RECT 15.725 28.275 16.015 28.505 ;
        RECT 16.170 28.260 16.490 28.520 ;
        RECT 17.105 28.460 17.395 28.505 ;
        RECT 17.550 28.460 17.870 28.520 ;
        RECT 19.390 28.460 19.710 28.520 ;
        RECT 17.105 28.320 19.710 28.460 ;
        RECT 17.105 28.275 17.395 28.320 ;
        RECT 17.550 28.260 17.870 28.320 ;
        RECT 19.390 28.260 19.710 28.320 ;
        RECT 10.205 28.120 10.495 28.165 ;
        RECT 10.650 28.120 10.970 28.180 ;
        RECT 10.205 27.980 10.970 28.120 ;
        RECT 34.660 28.120 34.800 28.660 ;
        RECT 41.930 28.600 42.250 28.660 ;
        RECT 42.480 28.660 44.550 28.800 ;
        RECT 35.030 28.460 35.350 28.520 ;
        RECT 41.025 28.460 41.315 28.505 ;
        RECT 35.030 28.320 41.315 28.460 ;
        RECT 35.030 28.260 35.350 28.320 ;
        RECT 41.025 28.275 41.315 28.320 ;
        RECT 36.425 28.120 36.715 28.165 ;
        RECT 34.660 27.980 36.715 28.120 ;
        RECT 10.205 27.935 10.495 27.980 ;
        RECT 10.650 27.920 10.970 27.980 ;
        RECT 36.425 27.935 36.715 27.980 ;
        RECT 37.345 28.120 37.635 28.165 ;
        RECT 37.790 28.120 38.110 28.180 ;
        RECT 42.480 28.165 42.620 28.660 ;
        RECT 44.230 28.600 44.550 28.660 ;
        RECT 47.080 28.660 50.055 28.800 ;
        RECT 42.865 28.460 43.155 28.505 ;
        RECT 43.770 28.460 44.090 28.520 ;
        RECT 42.865 28.320 44.090 28.460 ;
        RECT 42.865 28.275 43.155 28.320 ;
        RECT 43.770 28.260 44.090 28.320 ;
        RECT 46.070 28.260 46.390 28.520 ;
        RECT 47.080 28.505 47.220 28.660 ;
        RECT 49.765 28.615 50.055 28.660 ;
        RECT 47.005 28.275 47.295 28.505 ;
        RECT 47.465 28.275 47.755 28.505 ;
        RECT 37.345 27.980 38.110 28.120 ;
        RECT 37.345 27.935 37.635 27.980 ;
        RECT 37.790 27.920 38.110 27.980 ;
        RECT 41.945 27.935 42.235 28.165 ;
        RECT 42.405 27.935 42.695 28.165 ;
        RECT 43.310 28.120 43.630 28.180 ;
        RECT 47.540 28.120 47.680 28.275 ;
        RECT 47.910 28.260 48.230 28.520 ;
        RECT 50.300 28.460 50.440 29.000 ;
        RECT 52.550 29.000 56.510 29.140 ;
        RECT 52.550 28.955 52.840 29.000 ;
        RECT 54.650 28.955 54.940 29.000 ;
        RECT 56.220 28.955 56.510 29.000 ;
        RECT 50.670 28.800 50.990 28.860 ;
        RECT 52.065 28.800 52.355 28.845 ;
        RECT 50.670 28.660 52.355 28.800 ;
        RECT 50.670 28.600 50.990 28.660 ;
        RECT 52.065 28.615 52.355 28.660 ;
        RECT 52.945 28.800 53.235 28.845 ;
        RECT 54.135 28.800 54.425 28.845 ;
        RECT 56.655 28.800 56.945 28.845 ;
        RECT 52.945 28.660 56.945 28.800 ;
        RECT 52.945 28.615 53.235 28.660 ;
        RECT 54.135 28.615 54.425 28.660 ;
        RECT 56.655 28.615 56.945 28.660 ;
        RECT 51.605 28.460 51.895 28.505 ;
        RECT 55.270 28.460 55.590 28.520 ;
        RECT 56.190 28.460 56.510 28.520 ;
        RECT 50.300 28.320 56.510 28.460 ;
        RECT 51.605 28.275 51.895 28.320 ;
        RECT 55.270 28.260 55.590 28.320 ;
        RECT 56.190 28.260 56.510 28.320 ;
        RECT 59.870 28.460 60.190 28.520 ;
        RECT 60.345 28.460 60.635 28.505 ;
        RECT 60.880 28.460 61.020 29.340 ;
        RECT 68.700 29.185 68.840 29.340 ;
        RECT 62.210 29.140 62.500 29.185 ;
        RECT 64.310 29.140 64.600 29.185 ;
        RECT 65.880 29.140 66.170 29.185 ;
        RECT 62.210 29.000 66.170 29.140 ;
        RECT 62.210 28.955 62.500 29.000 ;
        RECT 64.310 28.955 64.600 29.000 ;
        RECT 65.880 28.955 66.170 29.000 ;
        RECT 68.625 29.140 68.915 29.185 ;
        RECT 75.970 29.140 76.290 29.200 ;
        RECT 68.625 29.000 76.290 29.140 ;
        RECT 68.625 28.955 68.915 29.000 ;
        RECT 75.970 28.940 76.290 29.000 ;
        RECT 62.605 28.800 62.895 28.845 ;
        RECT 63.795 28.800 64.085 28.845 ;
        RECT 66.315 28.800 66.605 28.845 ;
        RECT 62.605 28.660 66.605 28.800 ;
        RECT 62.605 28.615 62.895 28.660 ;
        RECT 63.795 28.615 64.085 28.660 ;
        RECT 66.315 28.615 66.605 28.660 ;
        RECT 59.870 28.320 61.020 28.460 ;
        RECT 61.725 28.460 62.015 28.505 ;
        RECT 65.390 28.460 65.710 28.520 ;
        RECT 61.725 28.320 65.710 28.460 ;
        RECT 59.870 28.260 60.190 28.320 ;
        RECT 60.345 28.275 60.635 28.320 ;
        RECT 61.725 28.275 62.015 28.320 ;
        RECT 65.390 28.260 65.710 28.320 ;
        RECT 81.030 28.260 81.350 28.520 ;
        RECT 43.310 27.980 47.680 28.120 ;
        RECT 7.445 27.780 7.735 27.825 ;
        RECT 7.890 27.780 8.210 27.840 ;
        RECT 7.445 27.640 8.210 27.780 ;
        RECT 7.445 27.595 7.735 27.640 ;
        RECT 7.890 27.580 8.210 27.640 ;
        RECT 9.285 27.780 9.575 27.825 ;
        RECT 9.730 27.780 10.050 27.840 ;
        RECT 9.285 27.640 10.050 27.780 ;
        RECT 9.285 27.595 9.575 27.640 ;
        RECT 9.730 27.580 10.050 27.640 ;
        RECT 13.870 27.580 14.190 27.840 ;
        RECT 38.250 27.580 38.570 27.840 ;
        RECT 42.020 27.780 42.160 27.935 ;
        RECT 43.310 27.920 43.630 27.980 ;
        RECT 44.690 27.780 45.010 27.840 ;
        RECT 42.020 27.640 45.010 27.780 ;
        RECT 47.540 27.780 47.680 27.980 ;
        RECT 49.750 28.120 50.070 28.180 ;
        RECT 50.685 28.120 50.975 28.165 ;
        RECT 51.130 28.120 51.450 28.180 ;
        RECT 49.750 27.980 51.450 28.120 ;
        RECT 49.750 27.920 50.070 27.980 ;
        RECT 50.685 27.935 50.975 27.980 ;
        RECT 51.130 27.920 51.450 27.980 ;
        RECT 52.050 28.120 52.370 28.180 ;
        RECT 53.290 28.120 53.580 28.165 ;
        RECT 52.050 27.980 53.580 28.120 ;
        RECT 52.050 27.920 52.370 27.980 ;
        RECT 53.290 27.935 53.580 27.980 ;
        RECT 61.265 28.120 61.555 28.165 ;
        RECT 63.060 28.120 63.350 28.165 ;
        RECT 64.930 28.120 65.250 28.180 ;
        RECT 61.265 27.980 62.860 28.120 ;
        RECT 61.265 27.935 61.555 27.980 ;
        RECT 52.510 27.780 52.830 27.840 ;
        RECT 47.540 27.640 52.830 27.780 ;
        RECT 44.690 27.580 45.010 27.640 ;
        RECT 52.510 27.580 52.830 27.640 ;
        RECT 55.270 27.780 55.590 27.840 ;
        RECT 58.965 27.780 59.255 27.825 ;
        RECT 55.270 27.640 59.255 27.780 ;
        RECT 55.270 27.580 55.590 27.640 ;
        RECT 58.965 27.595 59.255 27.640 ;
        RECT 59.425 27.780 59.715 27.825 ;
        RECT 62.170 27.780 62.490 27.840 ;
        RECT 59.425 27.640 62.490 27.780 ;
        RECT 62.720 27.780 62.860 27.980 ;
        RECT 63.060 27.980 65.250 28.120 ;
        RECT 63.060 27.935 63.350 27.980 ;
        RECT 64.930 27.920 65.250 27.980 ;
        RECT 67.230 28.120 67.550 28.180 ;
        RECT 70.925 28.120 71.215 28.165 ;
        RECT 67.230 27.980 71.215 28.120 ;
        RECT 67.230 27.920 67.550 27.980 ;
        RECT 70.925 27.935 71.215 27.980 ;
        RECT 71.830 27.920 72.150 28.180 ;
        RECT 67.320 27.780 67.460 27.920 ;
        RECT 62.720 27.640 67.460 27.780 ;
        RECT 59.425 27.595 59.715 27.640 ;
        RECT 62.170 27.580 62.490 27.640 ;
        RECT 72.750 27.580 73.070 27.840 ;
        RECT 81.965 27.780 82.255 27.825 ;
        RECT 82.870 27.780 83.190 27.840 ;
        RECT 81.965 27.640 83.190 27.780 ;
        RECT 81.965 27.595 82.255 27.640 ;
        RECT 82.870 27.580 83.190 27.640 ;
        RECT 5.520 26.960 84.180 27.440 ;
        RECT 11.570 26.760 11.890 26.820 ;
        RECT 9.360 26.620 11.890 26.760 ;
        RECT 9.360 26.420 9.500 26.620 ;
        RECT 11.570 26.560 11.890 26.620 ;
        RECT 16.170 26.760 16.490 26.820 ;
        RECT 18.485 26.760 18.775 26.805 ;
        RECT 16.170 26.620 18.775 26.760 ;
        RECT 16.170 26.560 16.490 26.620 ;
        RECT 18.485 26.575 18.775 26.620 ;
        RECT 19.390 26.760 19.710 26.820 ;
        RECT 40.090 26.760 40.410 26.820 ;
        RECT 56.650 26.760 56.970 26.820 ;
        RECT 58.505 26.760 58.795 26.805 ;
        RECT 61.710 26.760 62.030 26.820 ;
        RECT 19.390 26.620 40.410 26.760 ;
        RECT 19.390 26.560 19.710 26.620 ;
        RECT 8.900 26.280 9.500 26.420 ;
        RECT 12.460 26.420 12.750 26.465 ;
        RECT 13.870 26.420 14.190 26.480 ;
        RECT 12.460 26.280 14.190 26.420 ;
        RECT 8.900 26.125 9.040 26.280 ;
        RECT 12.460 26.235 12.750 26.280 ;
        RECT 13.870 26.220 14.190 26.280 ;
        RECT 8.825 25.895 9.115 26.125 ;
        RECT 9.270 25.880 9.590 26.140 ;
        RECT 9.730 25.880 10.050 26.140 ;
        RECT 10.665 26.080 10.955 26.125 ;
        RECT 12.120 26.080 12.720 26.095 ;
        RECT 17.550 26.080 17.870 26.140 ;
        RECT 19.405 26.080 19.695 26.125 ;
        RECT 10.665 25.955 17.870 26.080 ;
        RECT 10.665 25.940 12.260 25.955 ;
        RECT 12.580 25.940 17.870 25.955 ;
        RECT 10.665 25.895 10.955 25.940 ;
        RECT 17.550 25.880 17.870 25.940 ;
        RECT 18.100 25.940 19.695 26.080 ;
        RECT 10.190 25.740 10.510 25.800 ;
        RECT 11.125 25.740 11.415 25.785 ;
        RECT 10.190 25.600 11.415 25.740 ;
        RECT 10.190 25.540 10.510 25.600 ;
        RECT 11.125 25.555 11.415 25.600 ;
        RECT 12.005 25.740 12.295 25.785 ;
        RECT 13.195 25.740 13.485 25.785 ;
        RECT 15.715 25.740 16.005 25.785 ;
        RECT 12.005 25.600 16.005 25.740 ;
        RECT 12.005 25.555 12.295 25.600 ;
        RECT 13.195 25.555 13.485 25.600 ;
        RECT 15.715 25.555 16.005 25.600 ;
        RECT 11.610 25.400 11.900 25.445 ;
        RECT 13.710 25.400 14.000 25.445 ;
        RECT 15.280 25.400 15.570 25.445 ;
        RECT 11.610 25.260 15.570 25.400 ;
        RECT 11.610 25.215 11.900 25.260 ;
        RECT 13.710 25.215 14.000 25.260 ;
        RECT 15.280 25.215 15.570 25.260 ;
        RECT 7.430 24.860 7.750 25.120 ;
        RECT 14.790 25.060 15.110 25.120 ;
        RECT 18.100 25.105 18.240 25.940 ;
        RECT 19.405 25.895 19.695 25.940 ;
        RECT 20.310 25.880 20.630 26.140 ;
        RECT 22.625 25.895 22.915 26.125 ;
        RECT 23.085 25.895 23.375 26.125 ;
        RECT 22.700 25.400 22.840 25.895 ;
        RECT 23.160 25.740 23.300 25.895 ;
        RECT 23.530 25.880 23.850 26.140 ;
        RECT 24.540 26.125 24.680 26.620 ;
        RECT 40.090 26.560 40.410 26.620 ;
        RECT 42.940 26.620 56.420 26.760 ;
        RECT 30.905 26.420 31.195 26.465 ;
        RECT 26.380 26.280 31.195 26.420 ;
        RECT 24.465 25.895 24.755 26.125 ;
        RECT 25.385 26.080 25.675 26.125 ;
        RECT 25.830 26.080 26.150 26.140 ;
        RECT 26.380 26.125 26.520 26.280 ;
        RECT 30.905 26.235 31.195 26.280 ;
        RECT 34.110 26.420 34.430 26.480 ;
        RECT 42.940 26.420 43.080 26.620 ;
        RECT 50.670 26.420 50.990 26.480 ;
        RECT 34.110 26.280 43.080 26.420 ;
        RECT 43.400 26.280 50.990 26.420 ;
        RECT 34.110 26.220 34.430 26.280 ;
        RECT 25.385 25.940 26.150 26.080 ;
        RECT 25.385 25.895 25.675 25.940 ;
        RECT 25.830 25.880 26.150 25.940 ;
        RECT 26.305 25.895 26.595 26.125 ;
        RECT 26.750 25.880 27.070 26.140 ;
        RECT 27.225 26.080 27.515 26.125 ;
        RECT 27.670 26.080 27.990 26.140 ;
        RECT 27.225 25.940 27.990 26.080 ;
        RECT 27.225 25.895 27.515 25.940 ;
        RECT 27.670 25.880 27.990 25.940 ;
        RECT 29.050 25.880 29.370 26.140 ;
        RECT 29.985 26.080 30.275 26.125 ;
        RECT 35.030 26.080 35.350 26.140 ;
        RECT 35.950 26.125 36.270 26.140 ;
        RECT 43.400 26.125 43.540 26.280 ;
        RECT 50.670 26.220 50.990 26.280 ;
        RECT 44.690 26.125 45.010 26.140 ;
        RECT 29.985 25.940 35.350 26.080 ;
        RECT 29.985 25.895 30.275 25.940 ;
        RECT 35.030 25.880 35.350 25.940 ;
        RECT 35.920 25.895 36.270 26.125 ;
        RECT 43.325 25.895 43.615 26.125 ;
        RECT 44.660 25.895 45.010 26.125 ;
        RECT 35.950 25.880 36.270 25.895 ;
        RECT 44.690 25.880 45.010 25.895 ;
        RECT 46.070 26.080 46.390 26.140 ;
        RECT 52.600 26.125 52.740 26.620 ;
        RECT 54.825 26.420 55.115 26.465 ;
        RECT 53.520 26.280 55.115 26.420 ;
        RECT 56.280 26.420 56.420 26.620 ;
        RECT 56.650 26.620 58.795 26.760 ;
        RECT 56.650 26.560 56.970 26.620 ;
        RECT 58.505 26.575 58.795 26.620 ;
        RECT 59.500 26.620 62.030 26.760 ;
        RECT 59.500 26.420 59.640 26.620 ;
        RECT 61.710 26.560 62.030 26.620 ;
        RECT 64.930 26.560 65.250 26.820 ;
        RECT 71.830 26.760 72.150 26.820 ;
        RECT 74.605 26.760 74.895 26.805 ;
        RECT 71.830 26.620 76.660 26.760 ;
        RECT 71.830 26.560 72.150 26.620 ;
        RECT 74.605 26.575 74.895 26.620 ;
        RECT 56.280 26.280 59.640 26.420 ;
        RECT 46.070 25.940 48.600 26.080 ;
        RECT 46.070 25.880 46.390 25.940 ;
        RECT 26.840 25.740 26.980 25.880 ;
        RECT 48.460 25.800 48.600 25.940 ;
        RECT 52.525 25.895 52.815 26.125 ;
        RECT 52.970 25.880 53.290 26.140 ;
        RECT 53.520 26.125 53.660 26.280 ;
        RECT 54.825 26.235 55.115 26.280 ;
        RECT 59.870 26.220 60.190 26.480 ;
        RECT 64.010 26.420 64.330 26.480 ;
        RECT 63.180 26.280 64.330 26.420 ;
        RECT 53.445 25.895 53.735 26.125 ;
        RECT 54.365 25.895 54.655 26.125 ;
        RECT 55.270 26.080 55.590 26.140 ;
        RECT 55.745 26.080 56.035 26.125 ;
        RECT 55.270 25.940 56.035 26.080 ;
        RECT 34.570 25.740 34.890 25.800 ;
        RECT 23.160 25.600 26.980 25.740 ;
        RECT 27.760 25.600 34.890 25.740 ;
        RECT 27.760 25.460 27.900 25.600 ;
        RECT 34.570 25.540 34.890 25.600 ;
        RECT 35.465 25.740 35.755 25.785 ;
        RECT 36.655 25.740 36.945 25.785 ;
        RECT 39.175 25.740 39.465 25.785 ;
        RECT 35.465 25.600 39.465 25.740 ;
        RECT 35.465 25.555 35.755 25.600 ;
        RECT 36.655 25.555 36.945 25.600 ;
        RECT 39.175 25.555 39.465 25.600 ;
        RECT 44.205 25.740 44.495 25.785 ;
        RECT 45.395 25.740 45.685 25.785 ;
        RECT 47.915 25.740 48.205 25.785 ;
        RECT 44.205 25.600 48.205 25.740 ;
        RECT 44.205 25.555 44.495 25.600 ;
        RECT 45.395 25.555 45.685 25.600 ;
        RECT 47.915 25.555 48.205 25.600 ;
        RECT 48.370 25.740 48.690 25.800 ;
        RECT 54.440 25.740 54.580 25.895 ;
        RECT 55.270 25.880 55.590 25.940 ;
        RECT 55.745 25.895 56.035 25.940 ;
        RECT 56.190 26.080 56.510 26.140 ;
        RECT 56.665 26.080 56.955 26.125 ;
        RECT 56.190 25.940 56.955 26.080 ;
        RECT 48.370 25.600 54.580 25.740 ;
        RECT 55.820 25.740 55.960 25.895 ;
        RECT 56.190 25.880 56.510 25.940 ;
        RECT 56.665 25.895 56.955 25.940 ;
        RECT 59.410 25.880 59.730 26.140 ;
        RECT 60.330 25.880 60.650 26.140 ;
        RECT 61.265 26.080 61.555 26.125 ;
        RECT 60.880 25.940 61.555 26.080 ;
        RECT 60.880 25.740 61.020 25.940 ;
        RECT 61.265 25.895 61.555 25.940 ;
        RECT 61.725 25.895 62.015 26.125 ;
        RECT 62.170 26.080 62.490 26.140 ;
        RECT 63.180 26.125 63.320 26.280 ;
        RECT 64.010 26.220 64.330 26.280 ;
        RECT 65.390 26.420 65.710 26.480 ;
        RECT 75.510 26.420 75.830 26.480 ;
        RECT 76.520 26.465 76.660 26.620 ;
        RECT 65.390 26.280 75.830 26.420 ;
        RECT 65.390 26.220 65.710 26.280 ;
        RECT 67.780 26.125 67.920 26.280 ;
        RECT 75.510 26.220 75.830 26.280 ;
        RECT 76.445 26.420 76.735 26.465 ;
        RECT 78.270 26.420 78.590 26.480 ;
        RECT 76.445 26.280 78.590 26.420 ;
        RECT 76.445 26.235 76.735 26.280 ;
        RECT 78.270 26.220 78.590 26.280 ;
        RECT 62.645 26.080 62.935 26.125 ;
        RECT 62.170 25.940 62.935 26.080 ;
        RECT 61.800 25.740 61.940 25.895 ;
        RECT 62.170 25.880 62.490 25.940 ;
        RECT 62.645 25.895 62.935 25.940 ;
        RECT 63.105 25.895 63.395 26.125 ;
        RECT 63.565 25.895 63.855 26.125 ;
        RECT 67.705 25.895 67.995 26.125 ;
        RECT 69.040 26.080 69.330 26.125 ;
        RECT 70.450 26.080 70.770 26.140 ;
        RECT 69.040 25.940 70.770 26.080 ;
        RECT 69.040 25.895 69.330 25.940 ;
        RECT 55.820 25.600 61.020 25.740 ;
        RECT 61.340 25.600 61.940 25.740 ;
        RECT 48.370 25.540 48.690 25.600 ;
        RECT 22.700 25.260 23.760 25.400 ;
        RECT 18.025 25.060 18.315 25.105 ;
        RECT 14.790 24.920 18.315 25.060 ;
        RECT 14.790 24.860 15.110 24.920 ;
        RECT 18.025 24.875 18.315 24.920 ;
        RECT 21.245 25.060 21.535 25.105 ;
        RECT 23.070 25.060 23.390 25.120 ;
        RECT 21.245 24.920 23.390 25.060 ;
        RECT 23.620 25.060 23.760 25.260 ;
        RECT 27.670 25.200 27.990 25.460 ;
        RECT 29.510 25.400 29.830 25.460 ;
        RECT 28.220 25.260 29.830 25.400 ;
        RECT 28.220 25.060 28.360 25.260 ;
        RECT 29.510 25.200 29.830 25.260 ;
        RECT 35.070 25.400 35.360 25.445 ;
        RECT 37.170 25.400 37.460 25.445 ;
        RECT 38.740 25.400 39.030 25.445 ;
        RECT 35.070 25.260 39.030 25.400 ;
        RECT 35.070 25.215 35.360 25.260 ;
        RECT 37.170 25.215 37.460 25.260 ;
        RECT 38.740 25.215 39.030 25.260 ;
        RECT 43.810 25.400 44.100 25.445 ;
        RECT 45.910 25.400 46.200 25.445 ;
        RECT 47.480 25.400 47.770 25.445 ;
        RECT 43.810 25.260 47.770 25.400 ;
        RECT 43.810 25.215 44.100 25.260 ;
        RECT 45.910 25.215 46.200 25.260 ;
        RECT 47.480 25.215 47.770 25.260 ;
        RECT 51.145 25.400 51.435 25.445 ;
        RECT 52.050 25.400 52.370 25.460 ;
        RECT 51.145 25.260 52.370 25.400 ;
        RECT 51.145 25.215 51.435 25.260 ;
        RECT 52.050 25.200 52.370 25.260 ;
        RECT 23.620 24.920 28.360 25.060 ;
        RECT 21.245 24.875 21.535 24.920 ;
        RECT 23.070 24.860 23.390 24.920 ;
        RECT 28.590 24.860 28.910 25.120 ;
        RECT 37.790 25.060 38.110 25.120 ;
        RECT 41.485 25.060 41.775 25.105 ;
        RECT 37.790 24.920 41.775 25.060 ;
        RECT 37.790 24.860 38.110 24.920 ;
        RECT 41.485 24.875 41.775 24.920 ;
        RECT 47.910 25.060 48.230 25.120 ;
        RECT 50.225 25.060 50.515 25.105 ;
        RECT 47.910 24.920 50.515 25.060 ;
        RECT 54.440 25.060 54.580 25.600 ;
        RECT 54.810 25.400 55.130 25.460 ;
        RECT 59.410 25.400 59.730 25.460 ;
        RECT 54.810 25.260 59.730 25.400 ;
        RECT 54.810 25.200 55.130 25.260 ;
        RECT 59.410 25.200 59.730 25.260 ;
        RECT 61.340 25.060 61.480 25.600 ;
        RECT 61.710 25.400 62.030 25.460 ;
        RECT 63.640 25.400 63.780 25.895 ;
        RECT 70.450 25.880 70.770 25.940 ;
        RECT 70.910 26.080 71.230 26.140 ;
        RECT 74.590 26.080 74.910 26.140 ;
        RECT 75.985 26.080 76.275 26.125 ;
        RECT 70.910 25.940 73.440 26.080 ;
        RECT 70.910 25.880 71.230 25.940 ;
        RECT 73.300 25.800 73.440 25.940 ;
        RECT 74.590 25.940 76.275 26.080 ;
        RECT 74.590 25.880 74.910 25.940 ;
        RECT 75.985 25.895 76.275 25.940 ;
        RECT 76.905 25.895 77.195 26.125 ;
        RECT 68.585 25.740 68.875 25.785 ;
        RECT 69.775 25.740 70.065 25.785 ;
        RECT 72.295 25.740 72.585 25.785 ;
        RECT 68.585 25.600 72.585 25.740 ;
        RECT 68.585 25.555 68.875 25.600 ;
        RECT 69.775 25.555 70.065 25.600 ;
        RECT 72.295 25.555 72.585 25.600 ;
        RECT 73.210 25.740 73.530 25.800 ;
        RECT 76.980 25.740 77.120 25.895 ;
        RECT 77.810 25.880 78.130 26.140 ;
        RECT 73.210 25.600 77.120 25.740 ;
        RECT 73.210 25.540 73.530 25.600 ;
        RECT 61.710 25.260 63.780 25.400 ;
        RECT 68.190 25.400 68.480 25.445 ;
        RECT 70.290 25.400 70.580 25.445 ;
        RECT 71.860 25.400 72.150 25.445 ;
        RECT 68.190 25.260 72.150 25.400 ;
        RECT 61.710 25.200 62.030 25.260 ;
        RECT 68.190 25.215 68.480 25.260 ;
        RECT 70.290 25.215 70.580 25.260 ;
        RECT 71.860 25.215 72.150 25.260 ;
        RECT 73.670 25.060 73.990 25.120 ;
        RECT 54.440 24.920 73.990 25.060 ;
        RECT 47.910 24.860 48.230 24.920 ;
        RECT 50.225 24.875 50.515 24.920 ;
        RECT 73.670 24.860 73.990 24.920 ;
        RECT 75.050 24.860 75.370 25.120 ;
        RECT 5.520 24.240 84.180 24.720 ;
        RECT 10.650 24.040 10.970 24.100 ;
        RECT 13.885 24.040 14.175 24.085 ;
        RECT 10.650 23.900 14.175 24.040 ;
        RECT 10.650 23.840 10.970 23.900 ;
        RECT 13.885 23.855 14.175 23.900 ;
        RECT 7.470 23.700 7.760 23.745 ;
        RECT 9.570 23.700 9.860 23.745 ;
        RECT 11.140 23.700 11.430 23.745 ;
        RECT 7.470 23.560 11.430 23.700 ;
        RECT 7.470 23.515 7.760 23.560 ;
        RECT 9.570 23.515 9.860 23.560 ;
        RECT 11.140 23.515 11.430 23.560 ;
        RECT 7.865 23.360 8.155 23.405 ;
        RECT 9.055 23.360 9.345 23.405 ;
        RECT 11.575 23.360 11.865 23.405 ;
        RECT 7.865 23.220 11.865 23.360 ;
        RECT 7.865 23.175 8.155 23.220 ;
        RECT 9.055 23.175 9.345 23.220 ;
        RECT 11.575 23.175 11.865 23.220 ;
        RECT 6.985 23.020 7.275 23.065 ;
        RECT 10.190 23.020 10.510 23.080 ;
        RECT 6.985 22.880 10.510 23.020 ;
        RECT 13.960 23.020 14.100 23.855 ;
        RECT 17.090 23.840 17.410 24.100 ;
        RECT 19.850 24.040 20.170 24.100 ;
        RECT 34.585 24.040 34.875 24.085 ;
        RECT 35.030 24.040 35.350 24.100 ;
        RECT 19.850 23.900 34.340 24.040 ;
        RECT 19.850 23.840 20.170 23.900 ;
        RECT 20.810 23.700 21.100 23.745 ;
        RECT 22.910 23.700 23.200 23.745 ;
        RECT 24.480 23.700 24.770 23.745 ;
        RECT 20.810 23.560 24.770 23.700 ;
        RECT 20.810 23.515 21.100 23.560 ;
        RECT 22.910 23.515 23.200 23.560 ;
        RECT 24.480 23.515 24.770 23.560 ;
        RECT 28.170 23.700 28.460 23.745 ;
        RECT 30.270 23.700 30.560 23.745 ;
        RECT 31.840 23.700 32.130 23.745 ;
        RECT 28.170 23.560 32.130 23.700 ;
        RECT 34.200 23.700 34.340 23.900 ;
        RECT 34.585 23.900 35.350 24.040 ;
        RECT 34.585 23.855 34.875 23.900 ;
        RECT 35.030 23.840 35.350 23.900 ;
        RECT 35.950 23.840 36.270 24.100 ;
        RECT 38.800 23.900 62.170 24.040 ;
        RECT 38.800 23.700 38.940 23.900 ;
        RECT 34.200 23.560 38.940 23.700 ;
        RECT 28.170 23.515 28.460 23.560 ;
        RECT 30.270 23.515 30.560 23.560 ;
        RECT 31.840 23.515 32.130 23.560 ;
        RECT 39.170 23.500 39.490 23.760 ;
        RECT 44.690 23.500 45.010 23.760 ;
        RECT 62.030 23.700 62.170 23.900 ;
        RECT 70.450 23.840 70.770 24.100 ;
        RECT 75.050 23.700 75.370 23.760 ;
        RECT 62.030 23.560 75.370 23.700 ;
        RECT 75.050 23.500 75.370 23.560 ;
        RECT 76.010 23.700 76.300 23.745 ;
        RECT 78.110 23.700 78.400 23.745 ;
        RECT 79.680 23.700 79.970 23.745 ;
        RECT 76.010 23.560 79.970 23.700 ;
        RECT 76.010 23.515 76.300 23.560 ;
        RECT 78.110 23.515 78.400 23.560 ;
        RECT 79.680 23.515 79.970 23.560 ;
        RECT 21.205 23.360 21.495 23.405 ;
        RECT 22.395 23.360 22.685 23.405 ;
        RECT 24.915 23.360 25.205 23.405 ;
        RECT 21.205 23.220 25.205 23.360 ;
        RECT 21.205 23.175 21.495 23.220 ;
        RECT 22.395 23.175 22.685 23.220 ;
        RECT 24.915 23.175 25.205 23.220 ;
        RECT 28.565 23.360 28.855 23.405 ;
        RECT 29.755 23.360 30.045 23.405 ;
        RECT 32.275 23.360 32.565 23.405 ;
        RECT 39.260 23.360 39.400 23.500 ;
        RECT 41.010 23.360 41.330 23.420 ;
        RECT 66.310 23.360 66.630 23.420 ;
        RECT 70.450 23.360 70.770 23.420 ;
        RECT 73.210 23.360 73.530 23.420 ;
        RECT 75.510 23.360 75.830 23.420 ;
        RECT 28.565 23.220 32.565 23.360 ;
        RECT 28.565 23.175 28.855 23.220 ;
        RECT 29.755 23.175 30.045 23.220 ;
        RECT 32.275 23.175 32.565 23.220 ;
        RECT 37.880 23.220 70.220 23.360 ;
        RECT 14.345 23.020 14.635 23.065 ;
        RECT 13.960 22.880 14.635 23.020 ;
        RECT 6.985 22.835 7.275 22.880 ;
        RECT 10.190 22.820 10.510 22.880 ;
        RECT 14.345 22.835 14.635 22.880 ;
        RECT 14.790 23.020 15.110 23.080 ;
        RECT 15.725 23.020 16.015 23.065 ;
        RECT 14.790 22.880 16.015 23.020 ;
        RECT 14.790 22.820 15.110 22.880 ;
        RECT 15.725 22.835 16.015 22.880 ;
        RECT 16.185 23.020 16.475 23.065 ;
        RECT 17.550 23.020 17.870 23.080 ;
        RECT 16.185 22.880 17.870 23.020 ;
        RECT 16.185 22.835 16.475 22.880 ;
        RECT 17.550 22.820 17.870 22.880 ;
        RECT 20.310 22.820 20.630 23.080 ;
        RECT 21.660 23.020 21.950 23.065 ;
        RECT 23.070 23.020 23.390 23.080 ;
        RECT 21.660 22.880 23.390 23.020 ;
        RECT 21.660 22.835 21.950 22.880 ;
        RECT 23.070 22.820 23.390 22.880 ;
        RECT 27.670 22.820 27.990 23.080 ;
        RECT 37.880 23.065 38.020 23.220 ;
        RECT 41.010 23.160 41.330 23.220 ;
        RECT 29.020 22.835 29.310 23.065 ;
        RECT 37.345 22.835 37.635 23.065 ;
        RECT 37.805 22.835 38.095 23.065 ;
        RECT 7.430 22.680 7.750 22.740 ;
        RECT 8.210 22.680 8.500 22.725 ;
        RECT 15.265 22.680 15.555 22.725 ;
        RECT 7.430 22.540 8.500 22.680 ;
        RECT 7.430 22.480 7.750 22.540 ;
        RECT 8.210 22.495 8.500 22.540 ;
        RECT 14.420 22.540 15.555 22.680 ;
        RECT 14.420 22.400 14.560 22.540 ;
        RECT 15.265 22.495 15.555 22.540 ;
        RECT 28.590 22.680 28.910 22.740 ;
        RECT 29.140 22.680 29.280 22.835 ;
        RECT 28.590 22.540 29.280 22.680 ;
        RECT 29.510 22.680 29.830 22.740 ;
        RECT 34.110 22.680 34.430 22.740 ;
        RECT 37.420 22.680 37.560 22.835 ;
        RECT 38.250 22.820 38.570 23.080 ;
        RECT 39.185 23.020 39.475 23.065 ;
        RECT 40.090 23.020 40.410 23.080 ;
        RECT 46.070 23.020 46.390 23.080 ;
        RECT 46.620 23.065 46.760 23.220 ;
        RECT 66.310 23.160 66.630 23.220 ;
        RECT 39.185 22.880 40.410 23.020 ;
        RECT 39.185 22.835 39.475 22.880 ;
        RECT 40.090 22.820 40.410 22.880 ;
        RECT 42.480 22.880 46.390 23.020 ;
        RECT 29.510 22.540 37.560 22.680 ;
        RECT 28.590 22.480 28.910 22.540 ;
        RECT 29.510 22.480 29.830 22.540 ;
        RECT 34.110 22.480 34.430 22.540 ;
        RECT 41.930 22.480 42.250 22.740 ;
        RECT 14.330 22.140 14.650 22.400 ;
        RECT 23.070 22.340 23.390 22.400 ;
        RECT 27.225 22.340 27.515 22.385 ;
        RECT 23.070 22.200 27.515 22.340 ;
        RECT 23.070 22.140 23.390 22.200 ;
        RECT 27.225 22.155 27.515 22.200 ;
        RECT 28.130 22.340 28.450 22.400 ;
        RECT 42.480 22.340 42.620 22.880 ;
        RECT 46.070 22.820 46.390 22.880 ;
        RECT 46.545 22.835 46.835 23.065 ;
        RECT 47.005 22.835 47.295 23.065 ;
        RECT 47.925 22.835 48.215 23.065 ;
        RECT 51.605 23.020 51.895 23.065 ;
        RECT 60.790 23.020 61.110 23.080 ;
        RECT 67.705 23.020 67.995 23.065 ;
        RECT 69.530 23.020 69.850 23.080 ;
        RECT 51.605 22.880 61.110 23.020 ;
        RECT 51.605 22.835 51.895 22.880 ;
        RECT 42.865 22.495 43.155 22.725 ;
        RECT 43.785 22.680 44.075 22.725 ;
        RECT 47.080 22.680 47.220 22.835 ;
        RECT 43.785 22.540 47.220 22.680 ;
        RECT 43.785 22.495 44.075 22.540 ;
        RECT 28.130 22.200 42.620 22.340 ;
        RECT 42.940 22.340 43.080 22.495 ;
        RECT 48.000 22.400 48.140 22.835 ;
        RECT 60.790 22.820 61.110 22.880 ;
        RECT 62.030 22.880 69.850 23.020 ;
        RECT 70.080 23.020 70.220 23.220 ;
        RECT 70.450 23.220 72.520 23.360 ;
        RECT 70.450 23.160 70.770 23.220 ;
        RECT 71.370 23.020 71.690 23.080 ;
        RECT 70.080 22.880 71.690 23.020 ;
        RECT 48.370 22.680 48.690 22.740 ;
        RECT 62.030 22.680 62.170 22.880 ;
        RECT 67.705 22.835 67.995 22.880 ;
        RECT 69.530 22.820 69.850 22.880 ;
        RECT 71.370 22.820 71.690 22.880 ;
        RECT 71.830 22.820 72.150 23.080 ;
        RECT 72.380 23.065 72.520 23.220 ;
        RECT 73.210 23.220 75.830 23.360 ;
        RECT 73.210 23.160 73.530 23.220 ;
        RECT 75.510 23.160 75.830 23.220 ;
        RECT 76.405 23.360 76.695 23.405 ;
        RECT 77.595 23.360 77.885 23.405 ;
        RECT 80.115 23.360 80.405 23.405 ;
        RECT 76.405 23.220 80.405 23.360 ;
        RECT 76.405 23.175 76.695 23.220 ;
        RECT 77.595 23.175 77.885 23.220 ;
        RECT 80.115 23.175 80.405 23.220 ;
        RECT 72.305 22.835 72.595 23.065 ;
        RECT 72.750 22.820 73.070 23.080 ;
        RECT 73.670 22.820 73.990 23.080 ;
        RECT 48.370 22.540 62.170 22.680 ;
        RECT 68.625 22.680 68.915 22.725 ;
        RECT 75.510 22.680 75.830 22.740 ;
        RECT 76.750 22.680 77.040 22.725 ;
        RECT 68.625 22.540 75.280 22.680 ;
        RECT 48.370 22.480 48.690 22.540 ;
        RECT 68.625 22.495 68.915 22.540 ;
        RECT 44.230 22.340 44.550 22.400 ;
        RECT 47.450 22.340 47.770 22.400 ;
        RECT 42.940 22.200 47.770 22.340 ;
        RECT 28.130 22.140 28.450 22.200 ;
        RECT 44.230 22.140 44.550 22.200 ;
        RECT 47.450 22.140 47.770 22.200 ;
        RECT 47.910 22.340 48.230 22.400 ;
        RECT 50.685 22.340 50.975 22.385 ;
        RECT 47.910 22.200 50.975 22.340 ;
        RECT 47.910 22.140 48.230 22.200 ;
        RECT 50.685 22.155 50.975 22.200 ;
        RECT 69.545 22.340 69.835 22.385 ;
        RECT 72.750 22.340 73.070 22.400 ;
        RECT 69.545 22.200 73.070 22.340 ;
        RECT 75.140 22.340 75.280 22.540 ;
        RECT 75.510 22.540 77.040 22.680 ;
        RECT 75.510 22.480 75.830 22.540 ;
        RECT 76.750 22.495 77.040 22.540 ;
        RECT 77.810 22.340 78.130 22.400 ;
        RECT 82.410 22.340 82.730 22.400 ;
        RECT 75.140 22.200 82.730 22.340 ;
        RECT 69.545 22.155 69.835 22.200 ;
        RECT 72.750 22.140 73.070 22.200 ;
        RECT 77.810 22.140 78.130 22.200 ;
        RECT 82.410 22.140 82.730 22.200 ;
        RECT 5.520 21.520 84.180 22.000 ;
        RECT 22.625 21.320 22.915 21.365 ;
        RECT 23.530 21.320 23.850 21.380 ;
        RECT 22.625 21.180 23.850 21.320 ;
        RECT 22.625 21.135 22.915 21.180 ;
        RECT 23.530 21.120 23.850 21.180 ;
        RECT 35.950 21.320 36.270 21.380 ;
        RECT 41.930 21.320 42.250 21.380 ;
        RECT 48.370 21.320 48.690 21.380 ;
        RECT 35.950 21.180 39.860 21.320 ;
        RECT 35.950 21.120 36.270 21.180 ;
        RECT 14.330 20.980 14.650 21.040 ;
        RECT 15.725 20.980 16.015 21.025 ;
        RECT 14.330 20.840 16.015 20.980 ;
        RECT 14.330 20.780 14.650 20.840 ;
        RECT 15.725 20.795 16.015 20.840 ;
        RECT 19.850 20.980 20.170 21.040 ;
        RECT 20.785 20.980 21.075 21.025 ;
        RECT 19.850 20.840 21.075 20.980 ;
        RECT 19.850 20.780 20.170 20.840 ;
        RECT 20.785 20.795 21.075 20.840 ;
        RECT 21.705 20.980 21.995 21.025 ;
        RECT 23.070 20.980 23.390 21.040 ;
        RECT 21.705 20.840 23.390 20.980 ;
        RECT 21.705 20.795 21.995 20.840 ;
        RECT 23.070 20.780 23.390 20.840 ;
        RECT 32.730 20.980 33.050 21.040 ;
        RECT 34.585 20.980 34.875 21.025 ;
        RECT 37.790 20.980 38.110 21.040 ;
        RECT 32.730 20.840 34.875 20.980 ;
        RECT 32.730 20.780 33.050 20.840 ;
        RECT 34.585 20.795 34.875 20.840 ;
        RECT 35.120 20.840 38.110 20.980 ;
        RECT 8.365 20.455 8.655 20.685 ;
        RECT 10.650 20.640 10.970 20.700 ;
        RECT 11.585 20.640 11.875 20.685 ;
        RECT 10.650 20.500 11.875 20.640 ;
        RECT 8.440 19.960 8.580 20.455 ;
        RECT 10.650 20.440 10.970 20.500 ;
        RECT 11.585 20.455 11.875 20.500 ;
        RECT 13.425 20.640 13.715 20.685 ;
        RECT 13.870 20.640 14.190 20.700 ;
        RECT 14.805 20.640 15.095 20.685 ;
        RECT 13.425 20.500 15.095 20.640 ;
        RECT 13.425 20.455 13.715 20.500 ;
        RECT 13.870 20.440 14.190 20.500 ;
        RECT 14.805 20.455 15.095 20.500 ;
        RECT 16.185 20.455 16.475 20.685 ;
        RECT 16.645 20.640 16.935 20.685 ;
        RECT 17.550 20.640 17.870 20.700 ;
        RECT 16.645 20.500 17.870 20.640 ;
        RECT 16.645 20.455 16.935 20.500 ;
        RECT 16.260 20.300 16.400 20.455 ;
        RECT 17.550 20.440 17.870 20.500 ;
        RECT 18.025 20.640 18.315 20.685 ;
        RECT 18.470 20.640 18.790 20.700 ;
        RECT 18.025 20.500 18.790 20.640 ;
        RECT 23.160 20.640 23.300 20.780 ;
        RECT 35.120 20.685 35.260 20.840 ;
        RECT 37.790 20.780 38.110 20.840 ;
        RECT 39.170 20.780 39.490 21.040 ;
        RECT 39.720 20.980 39.860 21.180 ;
        RECT 41.930 21.180 48.690 21.320 ;
        RECT 41.930 21.120 42.250 21.180 ;
        RECT 48.370 21.120 48.690 21.180 ;
        RECT 58.030 21.320 58.350 21.380 ;
        RECT 64.010 21.320 64.330 21.380 ;
        RECT 70.450 21.320 70.770 21.380 ;
        RECT 58.030 21.180 60.560 21.320 ;
        RECT 58.030 21.120 58.350 21.180 ;
        RECT 43.770 20.980 44.090 21.040 ;
        RECT 39.720 20.840 44.090 20.980 ;
        RECT 33.665 20.640 33.955 20.685 ;
        RECT 23.160 20.500 33.955 20.640 ;
        RECT 18.025 20.455 18.315 20.500 ;
        RECT 18.100 20.300 18.240 20.455 ;
        RECT 18.470 20.440 18.790 20.500 ;
        RECT 33.665 20.455 33.955 20.500 ;
        RECT 35.045 20.455 35.335 20.685 ;
        RECT 35.505 20.640 35.795 20.685 ;
        RECT 35.950 20.640 36.270 20.700 ;
        RECT 40.180 20.685 40.320 20.840 ;
        RECT 43.770 20.780 44.090 20.840 ;
        RECT 47.910 20.980 48.230 21.040 ;
        RECT 55.745 20.980 56.035 21.025 ;
        RECT 60.420 20.980 60.560 21.180 ;
        RECT 62.720 21.180 70.770 21.320 ;
        RECT 47.910 20.840 54.580 20.980 ;
        RECT 47.910 20.780 48.230 20.840 ;
        RECT 35.505 20.500 36.270 20.640 ;
        RECT 35.505 20.455 35.795 20.500 ;
        RECT 35.950 20.440 36.270 20.500 ;
        RECT 38.265 20.455 38.555 20.685 ;
        RECT 39.645 20.455 39.935 20.685 ;
        RECT 40.105 20.455 40.395 20.685 ;
        RECT 50.210 20.640 50.530 20.700 ;
        RECT 52.525 20.640 52.815 20.685 ;
        RECT 50.210 20.500 52.815 20.640 ;
        RECT 16.260 20.160 18.240 20.300 ;
        RECT 34.110 20.300 34.430 20.360 ;
        RECT 38.340 20.300 38.480 20.455 ;
        RECT 34.110 20.160 38.480 20.300 ;
        RECT 39.720 20.300 39.860 20.455 ;
        RECT 50.210 20.440 50.530 20.500 ;
        RECT 52.525 20.455 52.815 20.500 ;
        RECT 52.970 20.440 53.290 20.700 ;
        RECT 54.440 20.685 54.580 20.840 ;
        RECT 55.745 20.840 60.100 20.980 ;
        RECT 60.420 20.840 61.020 20.980 ;
        RECT 55.745 20.795 56.035 20.840 ;
        RECT 59.960 20.700 60.100 20.840 ;
        RECT 53.445 20.455 53.735 20.685 ;
        RECT 54.365 20.455 54.655 20.685 ;
        RECT 56.190 20.640 56.510 20.700 ;
        RECT 56.665 20.640 56.955 20.685 ;
        RECT 56.190 20.500 56.955 20.640 ;
        RECT 41.470 20.300 41.790 20.360 ;
        RECT 39.720 20.160 41.790 20.300 ;
        RECT 34.110 20.100 34.430 20.160 ;
        RECT 41.470 20.100 41.790 20.160 ;
        RECT 48.830 20.300 49.150 20.360 ;
        RECT 53.060 20.300 53.200 20.440 ;
        RECT 48.830 20.160 53.200 20.300 ;
        RECT 53.520 20.300 53.660 20.455 ;
        RECT 56.190 20.440 56.510 20.500 ;
        RECT 56.665 20.455 56.955 20.500 ;
        RECT 58.490 20.440 58.810 20.700 ;
        RECT 58.965 20.455 59.255 20.685 ;
        RECT 54.825 20.300 55.115 20.345 ;
        RECT 58.030 20.300 58.350 20.360 ;
        RECT 53.520 20.160 55.115 20.300 ;
        RECT 48.830 20.100 49.150 20.160 ;
        RECT 54.825 20.115 55.115 20.160 ;
        RECT 55.360 20.160 58.350 20.300 ;
        RECT 59.040 20.300 59.180 20.455 ;
        RECT 59.410 20.440 59.730 20.700 ;
        RECT 59.870 20.640 60.190 20.700 ;
        RECT 60.345 20.640 60.635 20.685 ;
        RECT 59.870 20.500 60.635 20.640 ;
        RECT 60.880 20.640 61.020 20.840 ;
        RECT 62.720 20.685 62.860 21.180 ;
        RECT 64.010 21.120 64.330 21.180 ;
        RECT 70.450 21.120 70.770 21.180 ;
        RECT 71.370 21.120 71.690 21.380 ;
        RECT 71.830 21.320 72.150 21.380 ;
        RECT 71.830 21.180 74.360 21.320 ;
        RECT 71.830 21.120 72.150 21.180 ;
        RECT 66.325 20.980 66.615 21.025 ;
        RECT 67.230 20.980 67.550 21.040 ;
        RECT 66.325 20.840 67.550 20.980 ;
        RECT 66.325 20.795 66.615 20.840 ;
        RECT 67.230 20.780 67.550 20.840 ;
        RECT 67.690 20.980 68.010 21.040 ;
        RECT 71.460 20.980 71.600 21.120 ;
        RECT 74.220 20.980 74.360 21.180 ;
        RECT 74.590 20.980 74.910 21.040 ;
        RECT 67.690 20.840 70.220 20.980 ;
        RECT 71.460 20.840 73.900 20.980 ;
        RECT 67.690 20.780 68.010 20.840 ;
        RECT 62.185 20.640 62.475 20.685 ;
        RECT 60.880 20.500 62.475 20.640 ;
        RECT 59.870 20.440 60.190 20.500 ;
        RECT 60.345 20.455 60.635 20.500 ;
        RECT 62.185 20.455 62.475 20.500 ;
        RECT 62.645 20.455 62.935 20.685 ;
        RECT 63.105 20.455 63.395 20.685 ;
        RECT 64.025 20.640 64.315 20.685 ;
        RECT 64.025 20.500 65.160 20.640 ;
        RECT 64.025 20.455 64.315 20.500 ;
        RECT 61.250 20.300 61.570 20.360 ;
        RECT 59.040 20.160 61.570 20.300 ;
        RECT 63.180 20.300 63.320 20.455 ;
        RECT 64.485 20.300 64.775 20.345 ;
        RECT 63.180 20.160 64.775 20.300 ;
        RECT 65.020 20.300 65.160 20.500 ;
        RECT 65.390 20.440 65.710 20.700 ;
        RECT 69.070 20.640 69.390 20.700 ;
        RECT 70.080 20.685 70.220 20.840 ;
        RECT 65.940 20.500 69.390 20.640 ;
        RECT 65.940 20.300 66.080 20.500 ;
        RECT 69.070 20.440 69.390 20.500 ;
        RECT 70.005 20.455 70.295 20.685 ;
        RECT 70.465 20.455 70.755 20.685 ;
        RECT 65.020 20.160 66.080 20.300 ;
        RECT 70.540 20.300 70.680 20.455 ;
        RECT 70.910 20.440 71.230 20.700 ;
        RECT 71.370 20.640 71.690 20.700 ;
        RECT 71.845 20.640 72.135 20.685 ;
        RECT 71.370 20.500 72.135 20.640 ;
        RECT 71.370 20.440 71.690 20.500 ;
        RECT 71.845 20.455 72.135 20.500 ;
        RECT 72.290 20.440 72.610 20.700 ;
        RECT 72.750 20.640 73.070 20.700 ;
        RECT 73.760 20.685 73.900 20.840 ;
        RECT 74.220 20.840 74.910 20.980 ;
        RECT 74.220 20.685 74.360 20.840 ;
        RECT 74.590 20.780 74.910 20.840 ;
        RECT 73.225 20.640 73.515 20.685 ;
        RECT 72.750 20.500 73.515 20.640 ;
        RECT 72.750 20.440 73.070 20.500 ;
        RECT 73.225 20.455 73.515 20.500 ;
        RECT 73.685 20.455 73.975 20.685 ;
        RECT 74.145 20.455 74.435 20.685 ;
        RECT 77.365 20.640 77.655 20.685 ;
        RECT 77.810 20.640 78.130 20.700 ;
        RECT 74.635 20.500 78.130 20.640 ;
        RECT 74.635 20.300 74.775 20.500 ;
        RECT 77.365 20.455 77.655 20.500 ;
        RECT 77.810 20.440 78.130 20.500 ;
        RECT 79.190 20.440 79.510 20.700 ;
        RECT 82.410 20.440 82.730 20.700 ;
        RECT 70.540 20.160 74.775 20.300 ;
        RECT 15.710 19.960 16.030 20.020 ;
        RECT 8.440 19.820 16.030 19.960 ;
        RECT 15.710 19.760 16.030 19.820 ;
        RECT 16.630 19.960 16.950 20.020 ;
        RECT 18.945 19.960 19.235 20.005 ;
        RECT 16.630 19.820 19.235 19.960 ;
        RECT 16.630 19.760 16.950 19.820 ;
        RECT 18.945 19.775 19.235 19.820 ;
        RECT 36.410 19.760 36.730 20.020 ;
        RECT 41.025 19.960 41.315 20.005 ;
        RECT 42.390 19.960 42.710 20.020 ;
        RECT 41.025 19.820 42.710 19.960 ;
        RECT 41.025 19.775 41.315 19.820 ;
        RECT 42.390 19.760 42.710 19.820 ;
        RECT 48.370 19.960 48.690 20.020 ;
        RECT 55.360 19.960 55.500 20.160 ;
        RECT 58.030 20.100 58.350 20.160 ;
        RECT 61.250 20.100 61.570 20.160 ;
        RECT 64.485 20.115 64.775 20.160 ;
        RECT 75.510 20.100 75.830 20.360 ;
        RECT 87.010 20.300 87.330 20.360 ;
        RECT 78.360 20.160 87.330 20.300 ;
        RECT 48.370 19.820 55.500 19.960 ;
        RECT 48.370 19.760 48.690 19.820 ;
        RECT 57.570 19.760 57.890 20.020 ;
        RECT 62.630 19.960 62.950 20.020 ;
        RECT 78.360 20.005 78.500 20.160 ;
        RECT 87.010 20.100 87.330 20.160 ;
        RECT 69.085 19.960 69.375 20.005 ;
        RECT 62.630 19.820 69.375 19.960 ;
        RECT 62.630 19.760 62.950 19.820 ;
        RECT 69.085 19.775 69.375 19.820 ;
        RECT 78.285 19.775 78.575 20.005 ;
        RECT 80.125 19.960 80.415 20.005 ;
        RECT 83.790 19.960 84.110 20.020 ;
        RECT 80.125 19.820 84.110 19.960 ;
        RECT 80.125 19.775 80.415 19.820 ;
        RECT 83.790 19.760 84.110 19.820 ;
        RECT 6.970 19.620 7.290 19.680 ;
        RECT 7.445 19.620 7.735 19.665 ;
        RECT 6.970 19.480 7.735 19.620 ;
        RECT 6.970 19.420 7.290 19.480 ;
        RECT 7.445 19.435 7.735 19.480 ;
        RECT 10.650 19.420 10.970 19.680 ;
        RECT 11.570 19.620 11.890 19.680 ;
        RECT 12.505 19.620 12.795 19.665 ;
        RECT 11.570 19.480 12.795 19.620 ;
        RECT 11.570 19.420 11.890 19.480 ;
        RECT 12.505 19.435 12.795 19.480 ;
        RECT 17.090 19.620 17.410 19.680 ;
        RECT 17.565 19.620 17.855 19.665 ;
        RECT 17.090 19.480 17.855 19.620 ;
        RECT 17.090 19.420 17.410 19.480 ;
        RECT 17.565 19.435 17.855 19.480 ;
        RECT 51.130 19.420 51.450 19.680 ;
        RECT 59.410 19.620 59.730 19.680 ;
        RECT 60.805 19.620 61.095 19.665 ;
        RECT 59.410 19.480 61.095 19.620 ;
        RECT 59.410 19.420 59.730 19.480 ;
        RECT 60.805 19.435 61.095 19.480 ;
        RECT 70.450 19.620 70.770 19.680 ;
        RECT 72.290 19.620 72.610 19.680 ;
        RECT 70.450 19.480 72.610 19.620 ;
        RECT 70.450 19.420 70.770 19.480 ;
        RECT 72.290 19.420 72.610 19.480 ;
        RECT 80.570 19.620 80.890 19.680 ;
        RECT 81.505 19.620 81.795 19.665 ;
        RECT 80.570 19.480 81.795 19.620 ;
        RECT 80.570 19.420 80.890 19.480 ;
        RECT 81.505 19.435 81.795 19.480 ;
        RECT 5.520 18.800 84.180 19.280 ;
        RECT 18.010 18.600 18.330 18.660 ;
        RECT 33.665 18.600 33.955 18.645 ;
        RECT 34.110 18.600 34.430 18.660 ;
        RECT 18.010 18.460 33.420 18.600 ;
        RECT 18.010 18.400 18.330 18.460 ;
        RECT 15.250 18.260 15.570 18.320 ;
        RECT 27.250 18.260 27.540 18.305 ;
        RECT 29.350 18.260 29.640 18.305 ;
        RECT 30.920 18.260 31.210 18.305 ;
        RECT 15.250 18.120 15.940 18.260 ;
        RECT 15.250 18.060 15.570 18.120 ;
        RECT 12.030 17.920 12.350 17.980 ;
        RECT 15.800 17.920 15.940 18.120 ;
        RECT 27.250 18.120 31.210 18.260 ;
        RECT 27.250 18.075 27.540 18.120 ;
        RECT 29.350 18.075 29.640 18.120 ;
        RECT 30.920 18.075 31.210 18.120 ;
        RECT 27.645 17.920 27.935 17.965 ;
        RECT 28.835 17.920 29.125 17.965 ;
        RECT 31.355 17.920 31.645 17.965 ;
        RECT 8.900 17.780 15.480 17.920 ;
        RECT 8.900 17.625 9.040 17.780 ;
        RECT 12.030 17.720 12.350 17.780 ;
        RECT 8.825 17.395 9.115 17.625 ;
        RECT 9.270 17.380 9.590 17.640 ;
        RECT 9.730 17.380 10.050 17.640 ;
        RECT 10.665 17.395 10.955 17.625 ;
        RECT 13.425 17.580 13.715 17.625 ;
        RECT 14.790 17.580 15.110 17.640 ;
        RECT 15.340 17.625 15.480 17.780 ;
        RECT 15.800 17.780 24.680 17.920 ;
        RECT 15.800 17.625 15.940 17.780 ;
        RECT 13.425 17.440 15.110 17.580 ;
        RECT 13.425 17.395 13.715 17.440 ;
        RECT 10.740 17.240 10.880 17.395 ;
        RECT 14.790 17.380 15.110 17.440 ;
        RECT 15.265 17.395 15.555 17.625 ;
        RECT 15.725 17.395 16.015 17.625 ;
        RECT 16.170 17.380 16.490 17.640 ;
        RECT 17.105 17.580 17.395 17.625 ;
        RECT 19.390 17.580 19.710 17.640 ;
        RECT 20.860 17.625 21.000 17.780 ;
        RECT 17.105 17.440 19.710 17.580 ;
        RECT 17.105 17.395 17.395 17.440 ;
        RECT 17.180 17.240 17.320 17.395 ;
        RECT 19.390 17.380 19.710 17.440 ;
        RECT 20.325 17.395 20.615 17.625 ;
        RECT 20.785 17.395 21.075 17.625 ;
        RECT 10.740 17.100 17.320 17.240 ;
        RECT 7.430 16.700 7.750 16.960 ;
        RECT 12.490 16.700 12.810 16.960 ;
        RECT 12.950 16.900 13.270 16.960 ;
        RECT 13.885 16.900 14.175 16.945 ;
        RECT 12.950 16.760 14.175 16.900 ;
        RECT 20.400 16.900 20.540 17.395 ;
        RECT 21.230 17.380 21.550 17.640 ;
        RECT 23.085 17.395 23.375 17.625 ;
        RECT 23.160 17.240 23.300 17.395 ;
        RECT 23.990 17.380 24.310 17.640 ;
        RECT 24.540 17.625 24.680 17.780 ;
        RECT 27.645 17.780 31.645 17.920 ;
        RECT 33.280 17.920 33.420 18.460 ;
        RECT 33.665 18.460 34.430 18.600 ;
        RECT 33.665 18.415 33.955 18.460 ;
        RECT 34.110 18.400 34.430 18.460 ;
        RECT 36.410 18.600 36.730 18.660 ;
        RECT 50.210 18.600 50.530 18.660 ;
        RECT 61.710 18.600 62.030 18.660 ;
        RECT 36.410 18.460 50.530 18.600 ;
        RECT 36.410 18.400 36.730 18.460 ;
        RECT 50.210 18.400 50.530 18.460 ;
        RECT 50.760 18.460 62.030 18.600 ;
        RECT 50.760 18.260 50.900 18.460 ;
        RECT 61.710 18.400 62.030 18.460 ;
        RECT 64.945 18.600 65.235 18.645 ;
        RECT 65.390 18.600 65.710 18.660 ;
        RECT 64.945 18.460 65.710 18.600 ;
        RECT 64.945 18.415 65.235 18.460 ;
        RECT 65.390 18.400 65.710 18.460 ;
        RECT 66.770 18.600 67.090 18.660 ;
        RECT 66.770 18.460 76.200 18.600 ;
        RECT 66.770 18.400 67.090 18.460 ;
        RECT 36.500 18.120 50.900 18.260 ;
        RECT 51.170 18.260 51.460 18.305 ;
        RECT 53.270 18.260 53.560 18.305 ;
        RECT 54.840 18.260 55.130 18.305 ;
        RECT 51.170 18.120 55.130 18.260 ;
        RECT 36.500 17.920 36.640 18.120 ;
        RECT 51.170 18.075 51.460 18.120 ;
        RECT 53.270 18.075 53.560 18.120 ;
        RECT 54.840 18.075 55.130 18.120 ;
        RECT 58.530 18.260 58.820 18.305 ;
        RECT 60.630 18.260 60.920 18.305 ;
        RECT 62.200 18.260 62.490 18.305 ;
        RECT 58.530 18.120 62.490 18.260 ;
        RECT 58.530 18.075 58.820 18.120 ;
        RECT 60.630 18.075 60.920 18.120 ;
        RECT 62.200 18.075 62.490 18.120 ;
        RECT 71.830 18.060 72.150 18.320 ;
        RECT 76.060 18.260 76.200 18.460 ;
        RECT 77.350 18.260 77.670 18.320 ;
        RECT 81.045 18.260 81.335 18.305 ;
        RECT 76.060 18.120 76.660 18.260 ;
        RECT 41.010 17.920 41.330 17.980 ;
        RECT 51.565 17.920 51.855 17.965 ;
        RECT 52.755 17.920 53.045 17.965 ;
        RECT 55.275 17.920 55.565 17.965 ;
        RECT 33.280 17.780 36.640 17.920 ;
        RECT 36.960 17.780 42.620 17.920 ;
        RECT 27.645 17.735 27.935 17.780 ;
        RECT 28.835 17.735 29.125 17.780 ;
        RECT 31.355 17.735 31.645 17.780 ;
        RECT 24.465 17.395 24.755 17.625 ;
        RECT 24.910 17.380 25.230 17.640 ;
        RECT 26.765 17.580 27.055 17.625 ;
        RECT 27.210 17.580 27.530 17.640 ;
        RECT 26.765 17.440 27.530 17.580 ;
        RECT 26.765 17.395 27.055 17.440 ;
        RECT 27.210 17.380 27.530 17.440 ;
        RECT 36.410 17.380 36.730 17.640 ;
        RECT 36.960 17.625 37.100 17.780 ;
        RECT 41.010 17.720 41.330 17.780 ;
        RECT 36.885 17.395 37.175 17.625 ;
        RECT 37.330 17.380 37.650 17.640 ;
        RECT 38.265 17.580 38.555 17.625 ;
        RECT 40.090 17.580 40.410 17.640 ;
        RECT 42.480 17.625 42.620 17.780 ;
        RECT 43.400 17.780 48.600 17.920 ;
        RECT 38.265 17.440 40.410 17.580 ;
        RECT 38.265 17.395 38.555 17.440 ;
        RECT 40.090 17.380 40.410 17.440 ;
        RECT 41.945 17.395 42.235 17.625 ;
        RECT 42.405 17.395 42.695 17.625 ;
        RECT 25.830 17.240 26.150 17.300 ;
        RECT 23.160 17.100 26.150 17.240 ;
        RECT 25.830 17.040 26.150 17.100 ;
        RECT 26.305 17.240 26.595 17.285 ;
        RECT 27.990 17.240 28.280 17.285 ;
        RECT 42.020 17.240 42.160 17.395 ;
        RECT 42.850 17.380 43.170 17.640 ;
        RECT 43.400 17.240 43.540 17.780 ;
        RECT 48.460 17.640 48.600 17.780 ;
        RECT 51.565 17.780 55.565 17.920 ;
        RECT 51.565 17.735 51.855 17.780 ;
        RECT 52.755 17.735 53.045 17.780 ;
        RECT 55.275 17.735 55.565 17.780 ;
        RECT 58.925 17.920 59.215 17.965 ;
        RECT 60.115 17.920 60.405 17.965 ;
        RECT 62.635 17.920 62.925 17.965 ;
        RECT 58.925 17.780 62.925 17.920 ;
        RECT 58.925 17.735 59.215 17.780 ;
        RECT 60.115 17.735 60.405 17.780 ;
        RECT 62.635 17.735 62.925 17.780 ;
        RECT 66.310 17.920 66.630 17.980 ;
        RECT 69.070 17.920 69.390 17.980 ;
        RECT 71.920 17.920 72.060 18.060 ;
        RECT 66.310 17.780 67.460 17.920 ;
        RECT 66.310 17.720 66.630 17.780 ;
        RECT 43.785 17.395 44.075 17.625 ;
        RECT 26.305 17.100 28.280 17.240 ;
        RECT 26.305 17.055 26.595 17.100 ;
        RECT 27.990 17.055 28.280 17.100 ;
        RECT 28.680 17.100 43.540 17.240 ;
        RECT 43.860 17.240 44.000 17.395 ;
        RECT 47.910 17.380 48.230 17.640 ;
        RECT 48.370 17.380 48.690 17.640 ;
        RECT 48.830 17.380 49.150 17.640 ;
        RECT 49.290 17.380 49.610 17.640 ;
        RECT 50.225 17.395 50.515 17.625 ;
        RECT 48.000 17.240 48.140 17.380 ;
        RECT 50.300 17.240 50.440 17.395 ;
        RECT 50.670 17.380 50.990 17.640 ;
        RECT 51.130 17.580 51.450 17.640 ;
        RECT 51.965 17.580 52.255 17.625 ;
        RECT 51.130 17.440 52.255 17.580 ;
        RECT 51.130 17.380 51.450 17.440 ;
        RECT 51.965 17.395 52.255 17.440 ;
        RECT 58.045 17.580 58.335 17.625 ;
        RECT 62.170 17.580 62.490 17.640 ;
        RECT 58.045 17.440 62.490 17.580 ;
        RECT 58.045 17.395 58.335 17.440 ;
        RECT 62.170 17.380 62.490 17.440 ;
        RECT 66.770 17.380 67.090 17.640 ;
        RECT 67.320 17.625 67.460 17.780 ;
        RECT 68.700 17.780 72.060 17.920 ;
        RECT 72.395 17.780 76.200 17.920 ;
        RECT 67.245 17.395 67.535 17.625 ;
        RECT 67.690 17.380 68.010 17.640 ;
        RECT 68.700 17.625 68.840 17.780 ;
        RECT 69.070 17.720 69.390 17.780 ;
        RECT 72.395 17.640 72.535 17.780 ;
        RECT 68.625 17.395 68.915 17.625 ;
        RECT 70.910 17.380 71.230 17.640 ;
        RECT 71.830 17.380 72.150 17.640 ;
        RECT 72.290 17.380 72.610 17.640 ;
        RECT 72.750 17.380 73.070 17.640 ;
        RECT 73.670 17.580 73.990 17.640 ;
        RECT 76.060 17.625 76.200 17.780 ;
        RECT 76.520 17.625 76.660 18.120 ;
        RECT 77.350 18.120 81.335 18.260 ;
        RECT 77.350 18.060 77.670 18.120 ;
        RECT 81.045 18.075 81.335 18.120 ;
        RECT 74.605 17.580 74.895 17.625 ;
        RECT 73.670 17.440 74.895 17.580 ;
        RECT 73.670 17.380 73.990 17.440 ;
        RECT 74.605 17.395 74.895 17.440 ;
        RECT 75.525 17.380 75.815 17.610 ;
        RECT 75.985 17.395 76.275 17.625 ;
        RECT 76.445 17.395 76.735 17.625 ;
        RECT 78.270 17.380 78.590 17.640 ;
        RECT 80.110 17.380 80.430 17.640 ;
        RECT 59.410 17.285 59.730 17.300 ;
        RECT 59.380 17.240 59.730 17.285 ;
        RECT 43.860 17.100 50.440 17.240 ;
        RECT 59.215 17.100 59.730 17.240 ;
        RECT 20.770 16.900 21.090 16.960 ;
        RECT 20.400 16.760 21.090 16.900 ;
        RECT 12.950 16.700 13.270 16.760 ;
        RECT 13.885 16.715 14.175 16.760 ;
        RECT 20.770 16.700 21.090 16.760 ;
        RECT 22.610 16.700 22.930 16.960 ;
        RECT 24.910 16.900 25.230 16.960 ;
        RECT 28.680 16.900 28.820 17.100 ;
        RECT 59.380 17.055 59.730 17.100 ;
        RECT 59.410 17.040 59.730 17.055 ;
        RECT 75.600 16.960 75.740 17.380 ;
        RECT 24.910 16.760 28.820 16.900 ;
        RECT 24.910 16.700 25.230 16.760 ;
        RECT 35.030 16.700 35.350 16.960 ;
        RECT 40.550 16.700 40.870 16.960 ;
        RECT 47.005 16.900 47.295 16.945 ;
        RECT 47.910 16.900 48.230 16.960 ;
        RECT 47.005 16.760 48.230 16.900 ;
        RECT 47.005 16.715 47.295 16.760 ;
        RECT 47.910 16.700 48.230 16.760 ;
        RECT 50.210 16.900 50.530 16.960 ;
        RECT 54.810 16.900 55.130 16.960 ;
        RECT 50.210 16.760 55.130 16.900 ;
        RECT 50.210 16.700 50.530 16.760 ;
        RECT 54.810 16.700 55.130 16.760 ;
        RECT 57.585 16.900 57.875 16.945 ;
        RECT 59.870 16.900 60.190 16.960 ;
        RECT 57.585 16.760 60.190 16.900 ;
        RECT 57.585 16.715 57.875 16.760 ;
        RECT 59.870 16.700 60.190 16.760 ;
        RECT 65.390 16.700 65.710 16.960 ;
        RECT 70.910 16.900 71.230 16.960 ;
        RECT 73.670 16.900 73.990 16.960 ;
        RECT 70.910 16.760 73.990 16.900 ;
        RECT 70.910 16.700 71.230 16.760 ;
        RECT 73.670 16.700 73.990 16.760 ;
        RECT 74.145 16.900 74.435 16.945 ;
        RECT 74.590 16.900 74.910 16.960 ;
        RECT 74.145 16.760 74.910 16.900 ;
        RECT 74.145 16.715 74.435 16.760 ;
        RECT 74.590 16.700 74.910 16.760 ;
        RECT 75.510 16.700 75.830 16.960 ;
        RECT 76.890 16.900 77.210 16.960 ;
        RECT 77.825 16.900 78.115 16.945 ;
        RECT 76.890 16.760 78.115 16.900 ;
        RECT 76.890 16.700 77.210 16.760 ;
        RECT 77.825 16.715 78.115 16.760 ;
        RECT 79.190 16.700 79.510 16.960 ;
        RECT 5.520 16.080 84.180 16.560 ;
        RECT 9.730 15.680 10.050 15.940 ;
        RECT 13.870 15.880 14.190 15.940 ;
        RECT 10.280 15.740 14.190 15.880 ;
        RECT 7.905 15.540 8.195 15.585 ;
        RECT 8.350 15.540 8.670 15.600 ;
        RECT 7.905 15.400 8.670 15.540 ;
        RECT 7.905 15.355 8.195 15.400 ;
        RECT 8.350 15.340 8.670 15.400 ;
        RECT 8.825 15.540 9.115 15.585 ;
        RECT 10.280 15.540 10.420 15.740 ;
        RECT 13.870 15.680 14.190 15.740 ;
        RECT 20.770 15.680 21.090 15.940 ;
        RECT 23.990 15.880 24.310 15.940 ;
        RECT 28.605 15.880 28.895 15.925 ;
        RECT 23.990 15.740 28.895 15.880 ;
        RECT 23.990 15.680 24.310 15.740 ;
        RECT 28.605 15.695 28.895 15.740 ;
        RECT 41.470 15.880 41.790 15.940 ;
        RECT 47.005 15.880 47.295 15.925 ;
        RECT 41.470 15.740 47.295 15.880 ;
        RECT 41.470 15.680 41.790 15.740 ;
        RECT 47.005 15.695 47.295 15.740 ;
        RECT 49.290 15.880 49.610 15.940 ;
        RECT 54.825 15.880 55.115 15.925 ;
        RECT 64.930 15.880 65.250 15.940 ;
        RECT 49.290 15.740 55.115 15.880 ;
        RECT 49.290 15.680 49.610 15.740 ;
        RECT 54.825 15.695 55.115 15.740 ;
        RECT 59.040 15.740 65.250 15.880 ;
        RECT 22.610 15.585 22.930 15.600 ;
        RECT 22.580 15.540 22.930 15.585 ;
        RECT 8.825 15.400 10.420 15.540 ;
        RECT 10.740 15.400 20.540 15.540 ;
        RECT 22.415 15.400 22.930 15.540 ;
        RECT 8.825 15.355 9.115 15.400 ;
        RECT 10.190 15.200 10.510 15.260 ;
        RECT 10.740 15.200 10.880 15.400 ;
        RECT 20.400 15.260 20.540 15.400 ;
        RECT 22.580 15.355 22.930 15.400 ;
        RECT 22.610 15.340 22.930 15.355 ;
        RECT 27.210 15.540 27.530 15.600 ;
        RECT 29.525 15.540 29.815 15.585 ;
        RECT 34.110 15.540 34.430 15.600 ;
        RECT 27.210 15.400 34.430 15.540 ;
        RECT 27.210 15.340 27.530 15.400 ;
        RECT 29.525 15.355 29.815 15.400 ;
        RECT 34.110 15.340 34.430 15.400 ;
        RECT 35.030 15.540 35.350 15.600 ;
        RECT 37.850 15.540 38.140 15.585 ;
        RECT 50.670 15.540 50.990 15.600 ;
        RECT 35.030 15.400 38.140 15.540 ;
        RECT 35.030 15.340 35.350 15.400 ;
        RECT 37.850 15.355 38.140 15.400 ;
        RECT 40.180 15.400 50.990 15.540 ;
        RECT 11.110 15.200 11.430 15.260 ;
        RECT 12.950 15.245 13.270 15.260 ;
        RECT 11.585 15.200 11.875 15.245 ;
        RECT 12.920 15.200 13.270 15.245 ;
        RECT 10.190 15.060 11.875 15.200 ;
        RECT 12.755 15.060 13.270 15.200 ;
        RECT 10.190 15.000 10.510 15.060 ;
        RECT 11.110 15.000 11.430 15.060 ;
        RECT 11.585 15.015 11.875 15.060 ;
        RECT 12.920 15.015 13.270 15.060 ;
        RECT 12.950 15.000 13.270 15.015 ;
        RECT 15.710 15.200 16.030 15.260 ;
        RECT 18.945 15.200 19.235 15.245 ;
        RECT 19.390 15.200 19.710 15.260 ;
        RECT 15.710 15.060 18.700 15.200 ;
        RECT 15.710 15.000 16.030 15.060 ;
        RECT 12.465 14.860 12.755 14.905 ;
        RECT 13.655 14.860 13.945 14.905 ;
        RECT 16.175 14.860 16.465 14.905 ;
        RECT 12.465 14.720 16.465 14.860 ;
        RECT 18.560 14.860 18.700 15.060 ;
        RECT 18.945 15.060 19.710 15.200 ;
        RECT 18.945 15.015 19.235 15.060 ;
        RECT 19.390 15.000 19.710 15.060 ;
        RECT 19.865 15.015 20.155 15.245 ;
        RECT 20.310 15.200 20.630 15.260 ;
        RECT 40.180 15.245 40.320 15.400 ;
        RECT 21.245 15.200 21.535 15.245 ;
        RECT 20.310 15.060 21.535 15.200 ;
        RECT 19.940 14.860 20.080 15.015 ;
        RECT 20.310 15.000 20.630 15.060 ;
        RECT 21.245 15.015 21.535 15.060 ;
        RECT 21.780 15.060 27.900 15.200 ;
        RECT 21.780 14.860 21.920 15.060 ;
        RECT 18.560 14.720 20.080 14.860 ;
        RECT 12.465 14.675 12.755 14.720 ;
        RECT 13.655 14.675 13.945 14.720 ;
        RECT 16.175 14.675 16.465 14.720 ;
        RECT 12.070 14.520 12.360 14.565 ;
        RECT 14.170 14.520 14.460 14.565 ;
        RECT 15.740 14.520 16.030 14.565 ;
        RECT 12.070 14.380 16.030 14.520 ;
        RECT 12.070 14.335 12.360 14.380 ;
        RECT 14.170 14.335 14.460 14.380 ;
        RECT 15.740 14.335 16.030 14.380 ;
        RECT 18.470 13.980 18.790 14.240 ;
        RECT 19.940 14.180 20.080 14.720 ;
        RECT 20.400 14.720 21.920 14.860 ;
        RECT 22.125 14.860 22.415 14.905 ;
        RECT 23.315 14.860 23.605 14.905 ;
        RECT 25.835 14.860 26.125 14.905 ;
        RECT 22.125 14.720 26.125 14.860 ;
        RECT 27.760 14.860 27.900 15.060 ;
        RECT 30.445 15.015 30.735 15.245 ;
        RECT 39.185 15.200 39.475 15.245 ;
        RECT 40.105 15.200 40.395 15.245 ;
        RECT 39.185 15.060 40.395 15.200 ;
        RECT 39.185 15.015 39.475 15.060 ;
        RECT 40.105 15.015 40.395 15.060 ;
        RECT 40.550 15.200 40.870 15.260 ;
        RECT 47.540 15.245 47.680 15.400 ;
        RECT 50.670 15.340 50.990 15.400 ;
        RECT 56.190 15.540 56.510 15.600 ;
        RECT 59.040 15.585 59.180 15.740 ;
        RECT 64.930 15.680 65.250 15.740 ;
        RECT 67.690 15.880 68.010 15.940 ;
        RECT 71.385 15.880 71.675 15.925 ;
        RECT 67.690 15.740 71.675 15.880 ;
        RECT 67.690 15.680 68.010 15.740 ;
        RECT 71.385 15.695 71.675 15.740 ;
        RECT 72.290 15.880 72.610 15.940 ;
        RECT 80.110 15.880 80.430 15.940 ;
        RECT 72.290 15.740 80.430 15.880 ;
        RECT 72.290 15.680 72.610 15.740 ;
        RECT 80.110 15.680 80.430 15.740 ;
        RECT 56.665 15.540 56.955 15.585 ;
        RECT 56.190 15.400 56.955 15.540 ;
        RECT 56.190 15.340 56.510 15.400 ;
        RECT 56.665 15.355 56.955 15.400 ;
        RECT 58.965 15.355 59.255 15.585 ;
        RECT 59.410 15.340 59.730 15.600 ;
        RECT 73.210 15.540 73.530 15.600 ;
        RECT 63.180 15.400 73.530 15.540 ;
        RECT 41.385 15.200 41.675 15.245 ;
        RECT 40.550 15.060 41.675 15.200 ;
        RECT 29.050 14.860 29.370 14.920 ;
        RECT 30.520 14.860 30.660 15.015 ;
        RECT 40.550 15.000 40.870 15.060 ;
        RECT 41.385 15.015 41.675 15.060 ;
        RECT 47.465 15.015 47.755 15.245 ;
        RECT 47.910 15.200 48.230 15.260 ;
        RECT 48.745 15.200 49.035 15.245 ;
        RECT 47.910 15.060 49.035 15.200 ;
        RECT 47.910 15.000 48.230 15.060 ;
        RECT 48.745 15.015 49.035 15.060 ;
        RECT 55.745 15.015 56.035 15.245 ;
        RECT 27.760 14.720 30.660 14.860 ;
        RECT 34.595 14.860 34.885 14.905 ;
        RECT 37.115 14.860 37.405 14.905 ;
        RECT 38.305 14.860 38.595 14.905 ;
        RECT 34.595 14.720 38.595 14.860 ;
        RECT 20.400 14.580 20.540 14.720 ;
        RECT 22.125 14.675 22.415 14.720 ;
        RECT 23.315 14.675 23.605 14.720 ;
        RECT 25.835 14.675 26.125 14.720 ;
        RECT 29.050 14.660 29.370 14.720 ;
        RECT 34.595 14.675 34.885 14.720 ;
        RECT 37.115 14.675 37.405 14.720 ;
        RECT 38.305 14.675 38.595 14.720 ;
        RECT 40.985 14.860 41.275 14.905 ;
        RECT 42.175 14.860 42.465 14.905 ;
        RECT 44.695 14.860 44.985 14.905 ;
        RECT 40.985 14.720 44.985 14.860 ;
        RECT 40.985 14.675 41.275 14.720 ;
        RECT 42.175 14.675 42.465 14.720 ;
        RECT 44.695 14.675 44.985 14.720 ;
        RECT 48.345 14.860 48.635 14.905 ;
        RECT 49.535 14.860 49.825 14.905 ;
        RECT 52.055 14.860 52.345 14.905 ;
        RECT 55.820 14.860 55.960 15.015 ;
        RECT 58.490 15.000 58.810 15.260 ;
        RECT 60.345 15.015 60.635 15.245 ;
        RECT 63.180 15.200 63.320 15.400 ;
        RECT 73.210 15.340 73.530 15.400 ;
        RECT 62.720 15.060 63.320 15.200 ;
        RECT 63.520 15.200 63.810 15.245 ;
        RECT 65.390 15.200 65.710 15.260 ;
        RECT 63.520 15.060 65.710 15.200 ;
        RECT 57.110 14.860 57.430 14.920 ;
        RECT 60.420 14.860 60.560 15.015 ;
        RECT 48.345 14.720 52.345 14.860 ;
        RECT 48.345 14.675 48.635 14.720 ;
        RECT 49.535 14.675 49.825 14.720 ;
        RECT 52.055 14.675 52.345 14.720 ;
        RECT 54.440 14.720 60.560 14.860 ;
        RECT 62.170 14.860 62.490 14.920 ;
        RECT 62.720 14.860 62.860 15.060 ;
        RECT 63.520 15.015 63.810 15.060 ;
        RECT 65.390 15.000 65.710 15.060 ;
        RECT 69.530 15.000 69.850 15.260 ;
        RECT 70.465 15.200 70.755 15.245 ;
        RECT 71.370 15.200 71.690 15.260 ;
        RECT 74.590 15.245 74.910 15.260 ;
        RECT 74.560 15.200 74.910 15.245 ;
        RECT 70.465 15.060 71.690 15.200 ;
        RECT 74.395 15.060 74.910 15.200 ;
        RECT 70.465 15.015 70.755 15.060 ;
        RECT 62.170 14.720 62.860 14.860 ;
        RECT 63.065 14.860 63.355 14.905 ;
        RECT 64.255 14.860 64.545 14.905 ;
        RECT 66.775 14.860 67.065 14.905 ;
        RECT 63.065 14.720 67.065 14.860 ;
        RECT 20.310 14.320 20.630 14.580 ;
        RECT 21.730 14.520 22.020 14.565 ;
        RECT 23.830 14.520 24.120 14.565 ;
        RECT 25.400 14.520 25.690 14.565 ;
        RECT 32.730 14.520 33.050 14.580 ;
        RECT 54.440 14.565 54.580 14.720 ;
        RECT 57.110 14.660 57.430 14.720 ;
        RECT 62.170 14.660 62.490 14.720 ;
        RECT 63.065 14.675 63.355 14.720 ;
        RECT 64.255 14.675 64.545 14.720 ;
        RECT 66.775 14.675 67.065 14.720 ;
        RECT 21.730 14.380 25.690 14.520 ;
        RECT 21.730 14.335 22.020 14.380 ;
        RECT 23.830 14.335 24.120 14.380 ;
        RECT 25.400 14.335 25.690 14.380 ;
        RECT 28.220 14.380 33.050 14.520 ;
        RECT 28.220 14.225 28.360 14.380 ;
        RECT 32.730 14.320 33.050 14.380 ;
        RECT 35.030 14.520 35.320 14.565 ;
        RECT 36.600 14.520 36.890 14.565 ;
        RECT 38.700 14.520 38.990 14.565 ;
        RECT 35.030 14.380 38.990 14.520 ;
        RECT 35.030 14.335 35.320 14.380 ;
        RECT 36.600 14.335 36.890 14.380 ;
        RECT 38.700 14.335 38.990 14.380 ;
        RECT 40.590 14.520 40.880 14.565 ;
        RECT 42.690 14.520 42.980 14.565 ;
        RECT 44.260 14.520 44.550 14.565 ;
        RECT 40.590 14.380 44.550 14.520 ;
        RECT 40.590 14.335 40.880 14.380 ;
        RECT 42.690 14.335 42.980 14.380 ;
        RECT 44.260 14.335 44.550 14.380 ;
        RECT 47.950 14.520 48.240 14.565 ;
        RECT 50.050 14.520 50.340 14.565 ;
        RECT 51.620 14.520 51.910 14.565 ;
        RECT 47.950 14.380 51.910 14.520 ;
        RECT 47.950 14.335 48.240 14.380 ;
        RECT 50.050 14.335 50.340 14.380 ;
        RECT 51.620 14.335 51.910 14.380 ;
        RECT 54.365 14.335 54.655 14.565 ;
        RECT 54.810 14.520 55.130 14.580 ;
        RECT 62.670 14.520 62.960 14.565 ;
        RECT 64.770 14.520 65.060 14.565 ;
        RECT 66.340 14.520 66.630 14.565 ;
        RECT 54.810 14.380 62.170 14.520 ;
        RECT 54.810 14.320 55.130 14.380 ;
        RECT 28.145 14.180 28.435 14.225 ;
        RECT 19.940 14.040 28.435 14.180 ;
        RECT 28.145 13.995 28.435 14.040 ;
        RECT 30.890 14.180 31.210 14.240 ;
        RECT 32.285 14.180 32.575 14.225 ;
        RECT 30.890 14.040 32.575 14.180 ;
        RECT 30.890 13.980 31.210 14.040 ;
        RECT 32.285 13.995 32.575 14.040 ;
        RECT 45.610 14.180 45.930 14.240 ;
        RECT 57.585 14.180 57.875 14.225 ;
        RECT 45.610 14.040 57.875 14.180 ;
        RECT 62.030 14.180 62.170 14.380 ;
        RECT 62.670 14.380 66.630 14.520 ;
        RECT 62.670 14.335 62.960 14.380 ;
        RECT 64.770 14.335 65.060 14.380 ;
        RECT 66.340 14.335 66.630 14.380 ;
        RECT 69.085 14.520 69.375 14.565 ;
        RECT 69.530 14.520 69.850 14.580 ;
        RECT 70.540 14.520 70.680 15.015 ;
        RECT 71.370 15.000 71.690 15.060 ;
        RECT 74.560 15.015 74.910 15.060 ;
        RECT 74.590 15.000 74.910 15.015 ;
        RECT 75.970 15.200 76.290 15.260 ;
        RECT 80.585 15.200 80.875 15.245 ;
        RECT 75.970 15.060 80.875 15.200 ;
        RECT 75.970 15.000 76.290 15.060 ;
        RECT 80.585 15.015 80.875 15.060 ;
        RECT 73.210 14.660 73.530 14.920 ;
        RECT 74.105 14.860 74.395 14.905 ;
        RECT 75.295 14.860 75.585 14.905 ;
        RECT 77.815 14.860 78.105 14.905 ;
        RECT 74.105 14.720 78.105 14.860 ;
        RECT 74.105 14.675 74.395 14.720 ;
        RECT 75.295 14.675 75.585 14.720 ;
        RECT 77.815 14.675 78.105 14.720 ;
        RECT 69.085 14.380 70.680 14.520 ;
        RECT 73.710 14.520 74.000 14.565 ;
        RECT 75.810 14.520 76.100 14.565 ;
        RECT 77.380 14.520 77.670 14.565 ;
        RECT 73.710 14.380 77.670 14.520 ;
        RECT 69.085 14.335 69.375 14.380 ;
        RECT 69.530 14.320 69.850 14.380 ;
        RECT 73.710 14.335 74.000 14.380 ;
        RECT 75.810 14.335 76.100 14.380 ;
        RECT 77.380 14.335 77.670 14.380 ;
        RECT 72.750 14.180 73.070 14.240 ;
        RECT 62.030 14.040 73.070 14.180 ;
        RECT 45.610 13.980 45.930 14.040 ;
        RECT 57.585 13.995 57.875 14.040 ;
        RECT 72.750 13.980 73.070 14.040 ;
        RECT 81.490 13.980 81.810 14.240 ;
        RECT 5.520 13.360 84.180 13.840 ;
        RECT 13.870 12.960 14.190 13.220 ;
        RECT 15.265 13.160 15.555 13.205 ;
        RECT 16.170 13.160 16.490 13.220 ;
        RECT 34.570 13.160 34.890 13.220 ;
        RECT 15.265 13.020 16.490 13.160 ;
        RECT 15.265 12.975 15.555 13.020 ;
        RECT 16.170 12.960 16.490 13.020 ;
        RECT 25.460 13.020 34.890 13.160 ;
        RECT 7.470 12.820 7.760 12.865 ;
        RECT 9.570 12.820 9.860 12.865 ;
        RECT 11.140 12.820 11.430 12.865 ;
        RECT 7.470 12.680 11.430 12.820 ;
        RECT 7.470 12.635 7.760 12.680 ;
        RECT 9.570 12.635 9.860 12.680 ;
        RECT 11.140 12.635 11.430 12.680 ;
        RECT 7.865 12.480 8.155 12.525 ;
        RECT 9.055 12.480 9.345 12.525 ;
        RECT 11.575 12.480 11.865 12.525 ;
        RECT 7.865 12.340 11.865 12.480 ;
        RECT 7.865 12.295 8.155 12.340 ;
        RECT 9.055 12.295 9.345 12.340 ;
        RECT 11.575 12.295 11.865 12.340 ;
        RECT 6.985 12.140 7.275 12.185 ;
        RECT 11.110 12.140 11.430 12.200 ;
        RECT 6.985 12.000 11.430 12.140 ;
        RECT 6.985 11.955 7.275 12.000 ;
        RECT 11.110 11.940 11.430 12.000 ;
        RECT 16.185 12.140 16.475 12.185 ;
        RECT 18.470 12.140 18.790 12.200 ;
        RECT 16.185 12.000 18.790 12.140 ;
        RECT 16.185 11.955 16.475 12.000 ;
        RECT 18.470 11.940 18.790 12.000 ;
        RECT 21.245 12.140 21.535 12.185 ;
        RECT 23.070 12.140 23.390 12.200 ;
        RECT 21.245 12.000 23.390 12.140 ;
        RECT 21.245 11.955 21.535 12.000 ;
        RECT 23.070 11.940 23.390 12.000 ;
        RECT 23.530 11.940 23.850 12.200 ;
        RECT 25.460 12.185 25.600 13.020 ;
        RECT 34.570 12.960 34.890 13.020 ;
        RECT 37.330 13.160 37.650 13.220 ;
        RECT 37.805 13.160 38.095 13.205 ;
        RECT 37.330 13.020 38.095 13.160 ;
        RECT 37.330 12.960 37.650 13.020 ;
        RECT 37.805 12.975 38.095 13.020 ;
        RECT 42.850 13.160 43.170 13.220 ;
        RECT 43.785 13.160 44.075 13.205 ;
        RECT 42.850 13.020 44.075 13.160 ;
        RECT 42.850 12.960 43.170 13.020 ;
        RECT 43.785 12.975 44.075 13.020 ;
        RECT 71.830 13.160 72.150 13.220 ;
        RECT 72.305 13.160 72.595 13.205 ;
        RECT 71.830 13.020 72.595 13.160 ;
        RECT 71.830 12.960 72.150 13.020 ;
        RECT 72.305 12.975 72.595 13.020 ;
        RECT 74.605 13.160 74.895 13.205 ;
        RECT 75.510 13.160 75.830 13.220 ;
        RECT 74.605 13.020 75.830 13.160 ;
        RECT 74.605 12.975 74.895 13.020 ;
        RECT 75.510 12.960 75.830 13.020 ;
        RECT 26.305 12.820 26.595 12.865 ;
        RECT 29.050 12.820 29.370 12.880 ;
        RECT 26.305 12.680 29.370 12.820 ;
        RECT 26.305 12.635 26.595 12.680 ;
        RECT 29.050 12.620 29.370 12.680 ;
        RECT 35.505 12.820 35.795 12.865 ;
        RECT 40.090 12.820 40.410 12.880 ;
        RECT 35.505 12.680 40.410 12.820 ;
        RECT 35.505 12.635 35.795 12.680 ;
        RECT 40.090 12.620 40.410 12.680 ;
        RECT 76.010 12.820 76.300 12.865 ;
        RECT 78.110 12.820 78.400 12.865 ;
        RECT 79.680 12.820 79.970 12.865 ;
        RECT 76.010 12.680 79.970 12.820 ;
        RECT 76.010 12.635 76.300 12.680 ;
        RECT 78.110 12.635 78.400 12.680 ;
        RECT 79.680 12.635 79.970 12.680 ;
        RECT 47.450 12.480 47.770 12.540 ;
        RECT 61.250 12.480 61.570 12.540 ;
        RECT 72.290 12.480 72.610 12.540 ;
        RECT 30.980 12.340 37.100 12.480 ;
        RECT 30.980 12.200 31.120 12.340 ;
        RECT 25.385 11.955 25.675 12.185 ;
        RECT 27.210 11.940 27.530 12.200 ;
        RECT 29.065 12.140 29.355 12.185 ;
        RECT 29.970 12.140 30.290 12.200 ;
        RECT 29.065 12.000 30.290 12.140 ;
        RECT 29.065 11.955 29.355 12.000 ;
        RECT 29.970 11.940 30.290 12.000 ;
        RECT 30.890 11.940 31.210 12.200 ;
        RECT 32.730 11.940 33.050 12.200 ;
        RECT 33.190 12.140 33.510 12.200 ;
        RECT 34.200 12.185 34.340 12.340 ;
        RECT 33.665 12.140 33.955 12.185 ;
        RECT 33.190 12.000 33.955 12.140 ;
        RECT 33.190 11.940 33.510 12.000 ;
        RECT 33.665 11.955 33.955 12.000 ;
        RECT 34.125 11.955 34.415 12.185 ;
        RECT 34.585 12.140 34.875 12.185 ;
        RECT 36.410 12.140 36.730 12.200 ;
        RECT 36.960 12.185 37.100 12.340 ;
        RECT 47.450 12.340 52.280 12.480 ;
        RECT 47.450 12.280 47.770 12.340 ;
        RECT 34.585 12.000 36.730 12.140 ;
        RECT 34.585 11.955 34.875 12.000 ;
        RECT 36.410 11.940 36.730 12.000 ;
        RECT 36.885 11.955 37.175 12.185 ;
        RECT 37.790 12.140 38.110 12.200 ;
        RECT 39.645 12.140 39.935 12.185 ;
        RECT 37.790 12.000 39.935 12.140 ;
        RECT 37.790 11.940 38.110 12.000 ;
        RECT 39.645 11.955 39.935 12.000 ;
        RECT 40.105 12.140 40.395 12.185 ;
        RECT 41.470 12.140 41.790 12.200 ;
        RECT 42.865 12.140 43.155 12.185 ;
        RECT 40.105 12.000 43.155 12.140 ;
        RECT 40.105 11.955 40.395 12.000 ;
        RECT 41.470 11.940 41.790 12.000 ;
        RECT 42.865 11.955 43.155 12.000 ;
        RECT 47.005 12.140 47.295 12.185 ;
        RECT 49.750 12.140 50.070 12.200 ;
        RECT 52.140 12.185 52.280 12.340 ;
        RECT 61.250 12.340 72.610 12.480 ;
        RECT 61.250 12.280 61.570 12.340 ;
        RECT 47.005 12.000 50.070 12.140 ;
        RECT 47.005 11.955 47.295 12.000 ;
        RECT 49.750 11.940 50.070 12.000 ;
        RECT 50.225 11.955 50.515 12.185 ;
        RECT 52.065 11.955 52.355 12.185 ;
        RECT 56.665 12.140 56.955 12.185 ;
        RECT 57.110 12.140 57.430 12.200 ;
        RECT 56.665 12.000 57.430 12.140 ;
        RECT 56.665 11.955 56.955 12.000 ;
        RECT 7.430 11.800 7.750 11.860 ;
        RECT 8.210 11.800 8.500 11.845 ;
        RECT 7.430 11.660 8.500 11.800 ;
        RECT 7.430 11.600 7.750 11.660 ;
        RECT 8.210 11.615 8.500 11.660 ;
        RECT 17.105 11.800 17.395 11.845 ;
        RECT 18.930 11.800 19.250 11.860 ;
        RECT 32.270 11.800 32.590 11.860 ;
        RECT 17.105 11.660 19.250 11.800 ;
        RECT 17.105 11.615 17.395 11.660 ;
        RECT 18.930 11.600 19.250 11.660 ;
        RECT 28.220 11.660 32.590 11.800 ;
        RECT 19.390 11.460 19.710 11.520 ;
        RECT 20.325 11.460 20.615 11.505 ;
        RECT 19.390 11.320 20.615 11.460 ;
        RECT 19.390 11.260 19.710 11.320 ;
        RECT 20.325 11.275 20.615 11.320 ;
        RECT 22.610 11.260 22.930 11.520 ;
        RECT 24.465 11.460 24.755 11.505 ;
        RECT 25.830 11.460 26.150 11.520 ;
        RECT 28.220 11.505 28.360 11.660 ;
        RECT 32.270 11.600 32.590 11.660 ;
        RECT 35.965 11.800 36.255 11.845 ;
        RECT 41.930 11.800 42.250 11.860 ;
        RECT 35.965 11.660 42.250 11.800 ;
        RECT 50.300 11.800 50.440 11.955 ;
        RECT 57.110 11.940 57.430 12.000 ;
        RECT 59.870 11.940 60.190 12.200 ;
        RECT 63.090 11.940 63.410 12.200 ;
        RECT 64.930 11.940 65.250 12.200 ;
        RECT 69.530 11.940 69.850 12.200 ;
        RECT 71.460 12.185 71.600 12.340 ;
        RECT 72.290 12.280 72.610 12.340 ;
        RECT 73.210 12.480 73.530 12.540 ;
        RECT 75.525 12.480 75.815 12.525 ;
        RECT 73.210 12.340 75.815 12.480 ;
        RECT 73.210 12.280 73.530 12.340 ;
        RECT 75.525 12.295 75.815 12.340 ;
        RECT 76.405 12.480 76.695 12.525 ;
        RECT 77.595 12.480 77.885 12.525 ;
        RECT 80.115 12.480 80.405 12.525 ;
        RECT 76.405 12.340 80.405 12.480 ;
        RECT 76.405 12.295 76.695 12.340 ;
        RECT 77.595 12.295 77.885 12.340 ;
        RECT 80.115 12.295 80.405 12.340 ;
        RECT 76.890 12.185 77.210 12.200 ;
        RECT 71.385 11.955 71.675 12.185 ;
        RECT 76.860 12.140 77.210 12.185 ;
        RECT 76.695 12.000 77.210 12.140 ;
        RECT 76.860 11.955 77.210 12.000 ;
        RECT 76.890 11.940 77.210 11.955 ;
        RECT 55.270 11.800 55.590 11.860 ;
        RECT 50.300 11.660 55.590 11.800 ;
        RECT 35.965 11.615 36.255 11.660 ;
        RECT 41.930 11.600 42.250 11.660 ;
        RECT 55.270 11.600 55.590 11.660 ;
        RECT 66.310 11.800 66.630 11.860 ;
        RECT 70.465 11.800 70.755 11.845 ;
        RECT 72.765 11.800 73.055 11.845 ;
        RECT 66.310 11.660 73.055 11.800 ;
        RECT 66.310 11.600 66.630 11.660 ;
        RECT 70.465 11.615 70.755 11.660 ;
        RECT 72.765 11.615 73.055 11.660 ;
        RECT 73.685 11.800 73.975 11.845 ;
        RECT 77.810 11.800 78.130 11.860 ;
        RECT 73.685 11.660 82.640 11.800 ;
        RECT 73.685 11.615 73.975 11.660 ;
        RECT 77.810 11.600 78.130 11.660 ;
        RECT 24.465 11.320 26.150 11.460 ;
        RECT 24.465 11.275 24.755 11.320 ;
        RECT 25.830 11.260 26.150 11.320 ;
        RECT 28.145 11.275 28.435 11.505 ;
        RECT 29.985 11.460 30.275 11.505 ;
        RECT 35.030 11.460 35.350 11.520 ;
        RECT 29.985 11.320 35.350 11.460 ;
        RECT 29.985 11.275 30.275 11.320 ;
        RECT 35.030 11.260 35.350 11.320 ;
        RECT 38.710 11.260 39.030 11.520 ;
        RECT 41.025 11.460 41.315 11.505 ;
        RECT 41.470 11.460 41.790 11.520 ;
        RECT 41.025 11.320 41.790 11.460 ;
        RECT 41.025 11.275 41.315 11.320 ;
        RECT 41.470 11.260 41.790 11.320 ;
        RECT 45.150 11.460 45.470 11.520 ;
        RECT 46.085 11.460 46.375 11.505 ;
        RECT 45.150 11.320 46.375 11.460 ;
        RECT 45.150 11.260 45.470 11.320 ;
        RECT 46.085 11.275 46.375 11.320 ;
        RECT 48.370 11.460 48.690 11.520 ;
        RECT 49.305 11.460 49.595 11.505 ;
        RECT 48.370 11.320 49.595 11.460 ;
        RECT 48.370 11.260 48.690 11.320 ;
        RECT 49.305 11.275 49.595 11.320 ;
        RECT 51.590 11.460 51.910 11.520 ;
        RECT 52.985 11.460 53.275 11.505 ;
        RECT 51.590 11.320 53.275 11.460 ;
        RECT 51.590 11.260 51.910 11.320 ;
        RECT 52.985 11.275 53.275 11.320 ;
        RECT 54.810 11.460 55.130 11.520 ;
        RECT 55.745 11.460 56.035 11.505 ;
        RECT 54.810 11.320 56.035 11.460 ;
        RECT 54.810 11.260 55.130 11.320 ;
        RECT 55.745 11.275 56.035 11.320 ;
        RECT 58.030 11.460 58.350 11.520 ;
        RECT 58.965 11.460 59.255 11.505 ;
        RECT 58.030 11.320 59.255 11.460 ;
        RECT 58.030 11.260 58.350 11.320 ;
        RECT 58.965 11.275 59.255 11.320 ;
        RECT 61.250 11.460 61.570 11.520 ;
        RECT 62.185 11.460 62.475 11.505 ;
        RECT 61.250 11.320 62.475 11.460 ;
        RECT 61.250 11.260 61.570 11.320 ;
        RECT 62.185 11.275 62.475 11.320 ;
        RECT 64.470 11.460 64.790 11.520 ;
        RECT 65.865 11.460 66.155 11.505 ;
        RECT 64.470 11.320 66.155 11.460 ;
        RECT 64.470 11.260 64.790 11.320 ;
        RECT 65.865 11.275 66.155 11.320 ;
        RECT 67.690 11.460 68.010 11.520 ;
        RECT 82.500 11.505 82.640 11.660 ;
        RECT 68.625 11.460 68.915 11.505 ;
        RECT 67.690 11.320 68.915 11.460 ;
        RECT 67.690 11.260 68.010 11.320 ;
        RECT 68.625 11.275 68.915 11.320 ;
        RECT 82.425 11.275 82.715 11.505 ;
        RECT 5.520 10.640 84.180 11.120 ;
        RECT 0.070 6.700 0.390 6.760 ;
        RECT 7.890 6.700 8.210 6.760 ;
        RECT 0.070 6.560 8.210 6.700 ;
        RECT 0.070 6.500 0.390 6.560 ;
        RECT 7.890 6.500 8.210 6.560 ;
        RECT 70.910 6.700 71.230 6.760 ;
        RECT 81.490 6.700 81.810 6.760 ;
        RECT 70.910 6.560 81.810 6.700 ;
        RECT 70.910 6.500 71.230 6.560 ;
        RECT 81.490 6.500 81.810 6.560 ;
        RECT 3.290 6.360 3.610 6.420 ;
        RECT 11.570 6.360 11.890 6.420 ;
        RECT 3.290 6.220 11.890 6.360 ;
        RECT 3.290 6.160 3.610 6.220 ;
        RECT 11.570 6.160 11.890 6.220 ;
        RECT 74.130 5.680 74.450 5.740 ;
        RECT 79.190 5.680 79.510 5.740 ;
        RECT 74.130 5.540 79.510 5.680 ;
        RECT 74.130 5.480 74.450 5.540 ;
        RECT 79.190 5.480 79.510 5.540 ;
      LAYER met2 ;
        RECT 21.070 198.375 22.610 198.745 ;
        RECT 43.340 197.890 43.600 198.210 ;
        RECT 41.040 196.530 41.300 196.850 ;
        RECT 0.550 195.315 0.830 195.685 ;
        RECT 24.370 195.655 25.910 196.025 ;
        RECT 0.620 109.810 0.760 195.315 ;
        RECT 35.060 194.830 35.320 195.150 ;
        RECT 36.900 194.830 37.160 195.150 ;
        RECT 34.600 194.490 34.860 194.810 ;
        RECT 30.460 194.150 30.720 194.470 ;
        RECT 21.070 192.935 22.610 193.305 ;
        RECT 30.520 192.090 30.660 194.150 ;
        RECT 30.460 191.770 30.720 192.090 ;
        RECT 24.370 190.215 25.910 190.585 ;
        RECT 21.070 187.495 22.610 187.865 ;
        RECT 24.370 184.775 25.910 185.145 ;
        RECT 14.820 183.950 15.080 184.270 ;
        RECT 10.220 183.270 10.480 183.590 ;
        RECT 10.280 181.890 10.420 183.270 ;
        RECT 13.900 182.590 14.160 182.910 ;
        RECT 10.220 181.570 10.480 181.890 ;
        RECT 13.960 180.870 14.100 182.590 ;
        RECT 10.680 180.550 10.940 180.870 ;
        RECT 13.900 180.550 14.160 180.870 ;
        RECT 10.740 178.490 10.880 180.550 ;
        RECT 14.880 179.170 15.020 183.950 ;
        RECT 30.520 183.930 30.660 191.770 ;
        RECT 33.220 191.090 33.480 191.410 ;
        RECT 33.280 190.050 33.420 191.090 ;
        RECT 33.220 189.730 33.480 190.050 ;
        RECT 34.660 188.350 34.800 194.490 ;
        RECT 35.120 189.710 35.260 194.830 ;
        RECT 35.520 194.720 35.780 194.810 ;
        RECT 35.520 194.580 36.180 194.720 ;
        RECT 35.520 194.490 35.780 194.580 ;
        RECT 35.520 193.470 35.780 193.790 ;
        RECT 35.580 190.050 35.720 193.470 ;
        RECT 36.040 190.050 36.180 194.580 ;
        RECT 36.960 192.430 37.100 194.830 ;
        RECT 41.100 194.810 41.240 196.530 ;
        RECT 41.040 194.490 41.300 194.810 ;
        RECT 39.660 193.470 39.920 193.790 ;
        RECT 39.720 192.770 39.860 193.470 ;
        RECT 38.740 192.450 39.000 192.770 ;
        RECT 39.660 192.450 39.920 192.770 ;
        RECT 36.900 192.110 37.160 192.430 ;
        RECT 37.820 190.750 38.080 191.070 ;
        RECT 38.280 190.750 38.540 191.070 ;
        RECT 35.520 189.730 35.780 190.050 ;
        RECT 35.980 189.730 36.240 190.050 ;
        RECT 35.060 189.390 35.320 189.710 ;
        RECT 34.140 188.030 34.400 188.350 ;
        RECT 34.600 188.030 34.860 188.350 ;
        RECT 34.200 187.330 34.340 188.030 ;
        RECT 34.140 187.010 34.400 187.330 ;
        RECT 33.680 185.310 33.940 185.630 ;
        RECT 33.740 184.270 33.880 185.310 ;
        RECT 33.680 183.950 33.940 184.270 ;
        RECT 20.340 183.610 20.600 183.930 ;
        RECT 30.460 183.610 30.720 183.930 ;
        RECT 18.040 183.270 18.300 183.590 ;
        RECT 18.100 180.870 18.240 183.270 ;
        RECT 19.880 182.590 20.140 182.910 ;
        RECT 19.940 181.290 20.080 182.590 ;
        RECT 20.400 181.890 20.540 183.610 ;
        RECT 26.780 182.590 27.040 182.910 ;
        RECT 21.070 182.055 22.610 182.425 ;
        RECT 20.340 181.570 20.600 181.890 ;
        RECT 20.800 181.570 21.060 181.890 ;
        RECT 20.860 181.290 21.000 181.570 ;
        RECT 19.940 181.150 21.000 181.290 ;
        RECT 18.040 180.550 18.300 180.870 ;
        RECT 16.200 179.870 16.460 180.190 ;
        RECT 14.820 178.850 15.080 179.170 ;
        RECT 16.260 178.830 16.400 179.870 ;
        RECT 16.200 178.510 16.460 178.830 ;
        RECT 10.680 178.170 10.940 178.490 ;
        RECT 10.740 176.450 10.880 178.170 ;
        RECT 10.680 176.130 10.940 176.450 ;
        RECT 10.740 173.390 10.880 176.130 ;
        RECT 18.100 175.430 18.240 180.550 ;
        RECT 20.860 177.890 21.000 181.150 ;
        RECT 23.560 180.890 23.820 181.210 ;
        RECT 24.080 181.150 25.140 181.290 ;
        RECT 22.640 180.550 22.900 180.870 ;
        RECT 22.700 178.830 22.840 180.550 ;
        RECT 23.100 179.870 23.360 180.190 ;
        RECT 22.640 178.510 22.900 178.830 ;
        RECT 19.940 177.750 21.000 177.890 ;
        RECT 18.040 175.110 18.300 175.430 ;
        RECT 19.940 175.170 20.080 177.750 ;
        RECT 20.800 177.380 21.060 177.470 ;
        RECT 20.400 177.240 21.060 177.380 ;
        RECT 20.400 176.110 20.540 177.240 ;
        RECT 20.800 177.150 21.060 177.240 ;
        RECT 21.070 176.615 22.610 176.985 ;
        RECT 23.160 176.450 23.300 179.870 ;
        RECT 23.620 178.400 23.760 180.890 ;
        RECT 24.080 180.870 24.220 181.150 ;
        RECT 24.020 180.550 24.280 180.870 ;
        RECT 24.480 180.550 24.740 180.870 ;
        RECT 24.540 180.100 24.680 180.550 ;
        RECT 25.000 180.190 25.140 181.150 ;
        RECT 26.840 180.870 26.980 182.590 ;
        RECT 26.780 180.550 27.040 180.870 ;
        RECT 28.160 180.550 28.420 180.870 ;
        RECT 29.540 180.550 29.800 180.870 ;
        RECT 25.860 180.440 26.120 180.530 ;
        RECT 25.860 180.300 26.520 180.440 ;
        RECT 25.860 180.210 26.120 180.300 ;
        RECT 24.080 179.960 24.680 180.100 ;
        RECT 24.080 179.170 24.220 179.960 ;
        RECT 24.940 179.870 25.200 180.190 ;
        RECT 24.370 179.335 25.910 179.705 ;
        RECT 26.380 179.170 26.520 180.300 ;
        RECT 26.780 179.870 27.040 180.190 ;
        RECT 24.020 178.850 24.280 179.170 ;
        RECT 26.320 178.850 26.580 179.170 ;
        RECT 24.020 178.400 24.280 178.490 ;
        RECT 23.620 178.260 24.280 178.400 ;
        RECT 24.020 178.170 24.280 178.260 ;
        RECT 26.840 178.150 26.980 179.870 ;
        RECT 27.700 178.850 27.960 179.170 ;
        RECT 27.760 178.490 27.900 178.850 ;
        RECT 28.220 178.490 28.360 180.550 ;
        RECT 27.700 178.170 27.960 178.490 ;
        RECT 28.160 178.170 28.420 178.490 ;
        RECT 28.620 178.170 28.880 178.490 ;
        RECT 26.780 177.830 27.040 178.150 ;
        RECT 23.560 177.150 23.820 177.470 ;
        RECT 26.780 177.150 27.040 177.470 ;
        RECT 23.100 176.130 23.360 176.450 ;
        RECT 20.340 175.790 20.600 176.110 ;
        RECT 15.280 174.770 15.540 175.090 ;
        RECT 15.340 173.730 15.480 174.770 ;
        RECT 15.280 173.410 15.540 173.730 ;
        RECT 10.680 173.070 10.940 173.390 ;
        RECT 14.360 172.050 14.620 172.370 ;
        RECT 14.420 159.020 14.560 172.050 ;
        RECT 18.100 167.950 18.240 175.110 ;
        RECT 19.940 175.030 21.000 175.170 ;
        RECT 20.860 174.750 21.000 175.030 ;
        RECT 20.800 174.430 21.060 174.750 ;
        RECT 20.860 172.370 21.000 174.430 ;
        RECT 20.800 172.050 21.060 172.370 ;
        RECT 21.070 171.175 22.610 171.545 ;
        RECT 22.640 170.690 22.900 171.010 ;
        RECT 20.800 170.350 21.060 170.670 ;
        RECT 19.880 169.330 20.140 169.650 ;
        RECT 18.040 167.630 18.300 167.950 ;
        RECT 14.820 167.290 15.080 167.610 ;
        RECT 14.880 165.570 15.020 167.290 ;
        RECT 19.420 166.270 19.680 166.590 ;
        RECT 14.820 165.250 15.080 165.570 ;
        RECT 19.480 164.550 19.620 166.270 ;
        RECT 19.420 164.230 19.680 164.550 ;
        RECT 19.940 163.870 20.080 169.330 ;
        RECT 20.860 166.500 21.000 170.350 ;
        RECT 22.180 170.010 22.440 170.330 ;
        RECT 21.720 169.670 21.980 169.990 ;
        RECT 21.780 167.610 21.920 169.670 ;
        RECT 22.240 167.610 22.380 170.010 ;
        RECT 22.700 168.290 22.840 170.690 ;
        RECT 23.620 169.990 23.760 177.150 ;
        RECT 24.370 173.895 25.910 174.265 ;
        RECT 23.560 169.670 23.820 169.990 ;
        RECT 23.100 168.990 23.360 169.310 ;
        RECT 24.020 168.990 24.280 169.310 ;
        RECT 23.160 168.370 23.300 168.990 ;
        RECT 22.640 167.970 22.900 168.290 ;
        RECT 23.160 168.230 23.760 168.370 ;
        RECT 23.100 167.630 23.360 167.950 ;
        RECT 21.720 167.290 21.980 167.610 ;
        RECT 22.180 167.290 22.440 167.610 ;
        RECT 21.780 166.590 21.920 167.290 ;
        RECT 20.400 166.360 21.000 166.500 ;
        RECT 20.400 165.230 20.540 166.360 ;
        RECT 21.720 166.270 21.980 166.590 ;
        RECT 21.070 165.735 22.610 166.105 ;
        RECT 20.340 164.970 20.600 165.230 ;
        RECT 20.340 164.910 21.000 164.970 ;
        RECT 20.400 164.830 21.000 164.910 ;
        RECT 17.580 163.550 17.840 163.870 ;
        RECT 19.880 163.550 20.140 163.870 ;
        RECT 20.340 163.550 20.600 163.870 ;
        RECT 14.820 159.020 15.080 159.110 ;
        RECT 14.420 158.880 15.080 159.020 ;
        RECT 14.820 158.790 15.080 158.880 ;
        RECT 14.880 151.630 15.020 158.790 ;
        RECT 15.740 152.670 16.000 152.990 ;
        RECT 14.820 151.310 15.080 151.630 ;
        RECT 11.140 147.910 11.400 148.230 ;
        RECT 11.200 137.690 11.340 147.910 ;
        RECT 12.520 147.570 12.780 147.890 ;
        RECT 12.580 146.530 12.720 147.570 ;
        RECT 14.880 146.530 15.020 151.310 ;
        RECT 15.800 150.270 15.940 152.670 ;
        RECT 15.740 149.950 16.000 150.270 ;
        RECT 12.520 146.210 12.780 146.530 ;
        RECT 14.820 146.210 15.080 146.530 ;
        RECT 11.140 137.370 11.400 137.690 ;
        RECT 13.440 136.690 13.700 137.010 ;
        RECT 13.500 135.650 13.640 136.690 ;
        RECT 14.880 136.670 15.020 146.210 ;
        RECT 16.200 144.850 16.460 145.170 ;
        RECT 16.260 140.410 16.400 144.850 ;
        RECT 16.200 140.090 16.460 140.410 ;
        RECT 15.280 137.030 15.540 137.350 ;
        RECT 14.820 136.350 15.080 136.670 ;
        RECT 14.880 135.650 15.020 136.350 ;
        RECT 13.440 135.330 13.700 135.650 ;
        RECT 14.820 135.330 15.080 135.650 ;
        RECT 4.240 133.805 4.500 133.950 ;
        RECT 4.230 133.435 4.510 133.805 ;
        RECT 15.340 118.650 15.480 137.030 ;
        RECT 17.640 137.010 17.780 163.550 ;
        RECT 20.400 162.250 20.540 163.550 ;
        RECT 20.860 162.510 21.000 164.830 ;
        RECT 23.160 164.550 23.300 167.630 ;
        RECT 21.260 164.230 21.520 164.550 ;
        RECT 23.100 164.230 23.360 164.550 ;
        RECT 21.320 162.850 21.460 164.230 ;
        RECT 21.720 163.890 21.980 164.210 ;
        RECT 21.260 162.530 21.520 162.850 ;
        RECT 19.940 162.170 20.540 162.250 ;
        RECT 20.800 162.190 21.060 162.510 ;
        RECT 21.780 162.170 21.920 163.890 ;
        RECT 19.880 162.110 20.540 162.170 ;
        RECT 19.880 161.850 20.140 162.110 ;
        RECT 21.720 161.850 21.980 162.170 ;
        RECT 23.160 161.830 23.300 164.230 ;
        RECT 23.100 161.510 23.360 161.830 ;
        RECT 18.040 160.830 18.300 161.150 ;
        RECT 18.500 160.830 18.760 161.150 ;
        RECT 18.100 160.130 18.240 160.830 ;
        RECT 18.040 159.810 18.300 160.130 ;
        RECT 18.560 159.790 18.700 160.830 ;
        RECT 21.070 160.295 22.610 160.665 ;
        RECT 18.500 159.470 18.760 159.790 ;
        RECT 18.560 154.010 18.700 159.470 ;
        RECT 21.720 158.110 21.980 158.430 ;
        RECT 21.780 157.070 21.920 158.110 ;
        RECT 21.720 156.750 21.980 157.070 ;
        RECT 23.160 156.810 23.300 161.510 ;
        RECT 23.620 160.130 23.760 168.230 ;
        RECT 24.080 167.520 24.220 168.990 ;
        RECT 24.370 168.455 25.910 168.825 ;
        RECT 24.480 167.520 24.740 167.610 ;
        RECT 24.080 167.380 24.740 167.520 ;
        RECT 24.480 167.290 24.740 167.380 ;
        RECT 24.020 166.270 24.280 166.590 ;
        RECT 24.080 164.890 24.220 166.270 ;
        RECT 24.020 164.570 24.280 164.890 ;
        RECT 24.080 162.250 24.220 164.570 ;
        RECT 24.370 163.015 25.910 163.385 ;
        RECT 25.860 162.530 26.120 162.850 ;
        RECT 24.080 162.110 24.680 162.250 ;
        RECT 24.020 161.170 24.280 161.490 ;
        RECT 23.560 159.810 23.820 160.130 ;
        RECT 24.080 159.530 24.220 161.170 ;
        RECT 23.620 159.390 24.220 159.530 ;
        RECT 23.620 157.410 23.760 159.390 ;
        RECT 24.540 159.110 24.680 162.110 ;
        RECT 24.940 160.830 25.200 161.150 ;
        RECT 25.000 159.110 25.140 160.830 ;
        RECT 25.920 159.790 26.060 162.530 ;
        RECT 26.320 161.850 26.580 162.170 ;
        RECT 25.860 159.470 26.120 159.790 ;
        RECT 24.480 158.790 24.740 159.110 ;
        RECT 24.940 158.790 25.200 159.110 ;
        RECT 24.020 158.450 24.280 158.770 ;
        RECT 24.080 157.410 24.220 158.450 ;
        RECT 24.370 157.575 25.910 157.945 ;
        RECT 23.560 157.090 23.820 157.410 ;
        RECT 24.020 157.090 24.280 157.410 ;
        RECT 23.160 156.670 23.760 156.810 ;
        RECT 23.620 156.390 23.760 156.670 ;
        RECT 25.860 156.410 26.120 156.730 ;
        RECT 23.560 156.070 23.820 156.390 ;
        RECT 21.070 154.855 22.610 155.225 ;
        RECT 18.500 153.690 18.760 154.010 ;
        RECT 18.560 151.630 18.700 153.690 ;
        RECT 19.420 153.350 19.680 153.670 ;
        RECT 19.480 151.970 19.620 153.350 ;
        RECT 19.420 151.650 19.680 151.970 ;
        RECT 18.500 151.310 18.760 151.630 ;
        RECT 18.560 148.570 18.700 151.310 ;
        RECT 18.500 148.250 18.760 148.570 ;
        RECT 18.040 147.230 18.300 147.550 ;
        RECT 18.100 146.190 18.240 147.230 ;
        RECT 18.560 146.530 18.700 148.250 ;
        RECT 19.480 147.550 19.620 151.650 ;
        RECT 23.620 151.630 23.760 156.070 ;
        RECT 25.920 154.010 26.060 156.410 ;
        RECT 25.860 153.690 26.120 154.010 ;
        RECT 24.020 152.670 24.280 152.990 ;
        RECT 23.560 151.310 23.820 151.630 ;
        RECT 21.070 149.415 22.610 149.785 ;
        RECT 23.560 148.250 23.820 148.570 ;
        RECT 18.960 147.230 19.220 147.550 ;
        RECT 19.420 147.230 19.680 147.550 ;
        RECT 18.500 146.210 18.760 146.530 ;
        RECT 18.040 145.870 18.300 146.190 ;
        RECT 19.020 145.170 19.160 147.230 ;
        RECT 18.960 144.850 19.220 145.170 ;
        RECT 19.480 144.830 19.620 147.230 ;
        RECT 23.620 146.530 23.760 148.250 ;
        RECT 23.560 146.210 23.820 146.530 ;
        RECT 24.080 146.440 24.220 152.670 ;
        RECT 24.370 152.135 25.910 152.505 ;
        RECT 24.370 146.695 25.910 147.065 ;
        RECT 24.080 146.300 24.680 146.440 ;
        RECT 19.420 144.510 19.680 144.830 ;
        RECT 21.070 143.975 22.610 144.345 ;
        RECT 21.260 143.150 21.520 143.470 ;
        RECT 19.880 142.810 20.140 143.130 ;
        RECT 18.500 141.790 18.760 142.110 ;
        RECT 18.040 140.770 18.300 141.090 ;
        RECT 17.580 136.690 17.840 137.010 ;
        RECT 17.640 130.210 17.780 136.690 ;
        RECT 18.100 135.310 18.240 140.770 ;
        RECT 18.560 139.730 18.700 141.790 ;
        RECT 19.940 140.490 20.080 142.810 ;
        RECT 21.320 142.790 21.460 143.150 ;
        RECT 23.620 142.790 23.760 146.210 ;
        RECT 24.540 145.850 24.680 146.300 ;
        RECT 24.020 145.530 24.280 145.850 ;
        RECT 24.480 145.530 24.740 145.850 ;
        RECT 24.080 143.810 24.220 145.530 ;
        RECT 24.020 143.490 24.280 143.810 ;
        RECT 20.340 142.470 20.600 142.790 ;
        RECT 21.260 142.470 21.520 142.790 ;
        RECT 21.720 142.470 21.980 142.790 ;
        RECT 23.560 142.470 23.820 142.790 ;
        RECT 20.400 141.090 20.540 142.470 ;
        RECT 20.340 140.770 20.600 141.090 ;
        RECT 21.320 140.750 21.460 142.470 ;
        RECT 19.480 140.410 20.080 140.490 ;
        RECT 21.260 140.430 21.520 140.750 ;
        RECT 21.780 140.410 21.920 142.470 ;
        RECT 24.020 141.790 24.280 142.110 ;
        RECT 19.420 140.350 20.080 140.410 ;
        RECT 19.420 140.090 19.680 140.350 ;
        RECT 18.960 139.750 19.220 140.070 ;
        RECT 18.500 139.410 18.760 139.730 ;
        RECT 18.040 134.990 18.300 135.310 ;
        RECT 18.560 134.290 18.700 139.410 ;
        RECT 19.020 134.970 19.160 139.750 ;
        RECT 19.940 139.390 20.080 140.350 ;
        RECT 21.720 140.090 21.980 140.410 ;
        RECT 23.100 139.750 23.360 140.070 ;
        RECT 19.420 139.070 19.680 139.390 ;
        RECT 19.880 139.070 20.140 139.390 ;
        RECT 18.960 134.650 19.220 134.970 ;
        RECT 18.500 133.970 18.760 134.290 ;
        RECT 19.480 133.950 19.620 139.070 ;
        RECT 19.940 138.370 20.080 139.070 ;
        RECT 21.070 138.535 22.610 138.905 ;
        RECT 19.880 138.050 20.140 138.370 ;
        RECT 20.340 137.710 20.600 138.030 ;
        RECT 20.400 136.670 20.540 137.710 ;
        RECT 23.160 137.350 23.300 139.750 ;
        RECT 23.560 139.070 23.820 139.390 ;
        RECT 23.100 137.030 23.360 137.350 ;
        RECT 20.340 136.350 20.600 136.670 ;
        RECT 20.400 135.310 20.540 136.350 ;
        RECT 20.340 134.990 20.600 135.310 ;
        RECT 23.160 134.970 23.300 137.030 ;
        RECT 23.100 134.650 23.360 134.970 ;
        RECT 20.340 134.310 20.600 134.630 ;
        RECT 19.420 133.630 19.680 133.950 ;
        RECT 20.400 132.330 20.540 134.310 ;
        RECT 21.070 133.095 22.610 133.465 ;
        RECT 20.400 132.190 21.000 132.330 ;
        RECT 17.580 129.890 17.840 130.210 ;
        RECT 20.860 128.930 21.000 132.190 ;
        RECT 23.160 131.910 23.300 134.650 ;
        RECT 23.100 131.590 23.360 131.910 ;
        RECT 23.620 131.650 23.760 139.070 ;
        RECT 24.080 136.670 24.220 141.790 ;
        RECT 24.370 141.255 25.910 141.625 ;
        RECT 26.380 140.750 26.520 161.850 ;
        RECT 26.840 159.450 26.980 177.150 ;
        RECT 28.680 176.450 28.820 178.170 ;
        RECT 28.620 176.130 28.880 176.450 ;
        RECT 29.600 176.110 29.740 180.550 ;
        RECT 30.000 177.830 30.260 178.150 ;
        RECT 30.060 176.450 30.200 177.830 ;
        RECT 30.000 176.130 30.260 176.450 ;
        RECT 29.540 175.790 29.800 176.110 ;
        RECT 30.520 175.430 30.660 183.610 ;
        RECT 34.660 181.210 34.800 188.030 ;
        RECT 35.120 186.310 35.260 189.390 ;
        RECT 37.880 189.370 38.020 190.750 ;
        RECT 38.340 190.050 38.480 190.750 ;
        RECT 38.280 189.730 38.540 190.050 ;
        RECT 38.270 189.450 38.550 189.565 ;
        RECT 38.800 189.450 38.940 192.450 ;
        RECT 40.580 191.430 40.840 191.750 ;
        RECT 39.200 190.750 39.460 191.070 ;
        RECT 39.260 189.710 39.400 190.750 ;
        RECT 40.640 190.050 40.780 191.430 ;
        RECT 41.100 191.410 41.240 194.490 ;
        RECT 41.500 193.470 41.760 193.790 ;
        RECT 41.040 191.090 41.300 191.410 ;
        RECT 40.580 189.730 40.840 190.050 ;
        RECT 37.820 189.050 38.080 189.370 ;
        RECT 38.270 189.310 38.940 189.450 ;
        RECT 39.200 189.390 39.460 189.710 ;
        RECT 38.270 189.195 38.550 189.310 ;
        RECT 38.280 189.050 38.540 189.195 ;
        RECT 35.060 185.990 35.320 186.310 ;
        RECT 35.060 185.310 35.320 185.630 ;
        RECT 35.120 181.890 35.260 185.310 ;
        RECT 36.440 182.650 36.700 182.910 ;
        RECT 36.040 182.590 36.700 182.650 ;
        RECT 36.040 182.510 36.640 182.590 ;
        RECT 35.060 181.570 35.320 181.890 ;
        RECT 34.600 180.890 34.860 181.210 ;
        RECT 33.680 178.170 33.940 178.490 ;
        RECT 30.460 175.110 30.720 175.430 ;
        RECT 27.700 174.770 27.960 175.090 ;
        RECT 27.240 169.330 27.500 169.650 ;
        RECT 27.300 161.830 27.440 169.330 ;
        RECT 27.760 164.550 27.900 174.770 ;
        RECT 29.540 170.690 29.800 171.010 ;
        RECT 29.600 166.590 29.740 170.690 ;
        RECT 30.520 170.330 30.660 175.110 ;
        RECT 33.740 175.090 33.880 178.170 ;
        RECT 34.140 175.790 34.400 176.110 ;
        RECT 33.680 174.770 33.940 175.090 ;
        RECT 30.460 170.010 30.720 170.330 ;
        RECT 30.520 167.950 30.660 170.010 ;
        RECT 30.460 167.630 30.720 167.950 ;
        RECT 29.540 166.270 29.800 166.590 ;
        RECT 27.700 164.230 27.960 164.550 ;
        RECT 27.240 161.510 27.500 161.830 ;
        RECT 27.240 159.470 27.500 159.790 ;
        RECT 26.780 159.130 27.040 159.450 ;
        RECT 26.780 158.450 27.040 158.770 ;
        RECT 26.840 153.670 26.980 158.450 ;
        RECT 26.780 153.350 27.040 153.670 ;
        RECT 26.780 151.650 27.040 151.970 ;
        RECT 26.840 147.550 26.980 151.650 ;
        RECT 26.780 147.230 27.040 147.550 ;
        RECT 26.780 145.530 27.040 145.850 ;
        RECT 26.840 143.470 26.980 145.530 ;
        RECT 27.300 145.510 27.440 159.470 ;
        RECT 27.760 158.770 27.900 164.230 ;
        RECT 29.080 163.610 29.340 163.870 ;
        RECT 29.600 163.610 29.740 166.270 ;
        RECT 30.520 164.550 30.660 167.630 ;
        RECT 34.200 167.610 34.340 175.790 ;
        RECT 34.660 169.900 34.800 180.890 ;
        RECT 36.040 180.870 36.180 182.510 ;
        RECT 35.980 180.550 36.240 180.870 ;
        RECT 35.520 180.210 35.780 180.530 ;
        RECT 35.060 169.900 35.320 169.990 ;
        RECT 34.660 169.760 35.320 169.900 ;
        RECT 35.060 169.670 35.320 169.760 ;
        RECT 34.600 168.990 34.860 169.310 ;
        RECT 35.580 169.050 35.720 180.210 ;
        RECT 36.040 178.490 36.180 180.550 ;
        RECT 37.360 179.870 37.620 180.190 ;
        RECT 37.420 178.490 37.560 179.870 ;
        RECT 35.980 178.170 36.240 178.490 ;
        RECT 37.360 178.170 37.620 178.490 ;
        RECT 37.880 175.430 38.020 189.050 ;
        RECT 41.100 183.250 41.240 191.090 ;
        RECT 41.560 191.070 41.700 193.470 ;
        RECT 43.400 192.770 43.540 197.890 ;
        RECT 54.900 197.190 55.040 206.000 ;
        RECT 64.560 197.190 64.700 206.000 ;
        RECT 54.840 196.870 55.100 197.190 ;
        RECT 64.500 196.870 64.760 197.190 ;
        RECT 50.240 196.190 50.500 196.510 ;
        RECT 53.920 196.190 54.180 196.510 ;
        RECT 56.680 196.190 56.940 196.510 ;
        RECT 63.120 196.190 63.380 196.510 ;
        RECT 50.300 195.490 50.440 196.190 ;
        RECT 50.240 195.170 50.500 195.490 ;
        RECT 48.860 194.150 49.120 194.470 ;
        RECT 43.340 192.450 43.600 192.770 ;
        RECT 42.420 191.430 42.680 191.750 ;
        RECT 41.500 190.750 41.760 191.070 ;
        RECT 41.560 188.690 41.700 190.750 ;
        RECT 41.500 188.370 41.760 188.690 ;
        RECT 39.660 182.930 39.920 183.250 ;
        RECT 41.040 182.930 41.300 183.250 ;
        RECT 39.200 177.490 39.460 177.810 ;
        RECT 39.260 175.430 39.400 177.490 ;
        RECT 37.820 175.110 38.080 175.430 ;
        RECT 39.200 175.110 39.460 175.430 ;
        RECT 37.360 172.730 37.620 173.050 ;
        RECT 36.440 172.050 36.700 172.370 ;
        RECT 35.980 171.710 36.240 172.030 ;
        RECT 36.040 169.650 36.180 171.710 ;
        RECT 36.500 171.010 36.640 172.050 ;
        RECT 36.440 170.690 36.700 171.010 ;
        RECT 36.900 170.350 37.160 170.670 ;
        RECT 36.960 169.650 37.100 170.350 ;
        RECT 35.980 169.330 36.240 169.650 ;
        RECT 36.900 169.330 37.160 169.650 ;
        RECT 34.140 167.290 34.400 167.610 ;
        RECT 34.200 165.570 34.340 167.290 ;
        RECT 34.140 165.250 34.400 165.570 ;
        RECT 34.660 164.550 34.800 168.990 ;
        RECT 35.120 168.910 35.720 169.050 ;
        RECT 30.460 164.230 30.720 164.550 ;
        RECT 32.300 164.230 32.560 164.550 ;
        RECT 34.600 164.230 34.860 164.550 ;
        RECT 29.080 163.550 29.740 163.610 ;
        RECT 31.380 163.550 31.640 163.870 ;
        RECT 29.140 163.470 29.740 163.550 ;
        RECT 29.600 162.170 29.740 163.470 ;
        RECT 31.440 162.510 31.580 163.550 ;
        RECT 31.380 162.190 31.640 162.510 ;
        RECT 29.540 161.850 29.800 162.170 ;
        RECT 29.600 160.130 29.740 161.850 ;
        RECT 30.000 161.510 30.260 161.830 ;
        RECT 29.540 159.810 29.800 160.130 ;
        RECT 29.600 159.450 29.740 159.810 ;
        RECT 29.540 159.130 29.800 159.450 ;
        RECT 30.060 159.110 30.200 161.510 ;
        RECT 30.920 159.470 31.180 159.790 ;
        RECT 30.000 158.790 30.260 159.110 ;
        RECT 27.760 158.630 28.360 158.770 ;
        RECT 28.220 156.390 28.360 158.630 ;
        RECT 30.980 156.730 31.120 159.470 ;
        RECT 31.440 159.110 31.580 162.190 ;
        RECT 31.380 158.790 31.640 159.110 ;
        RECT 30.920 156.410 31.180 156.730 ;
        RECT 28.160 156.070 28.420 156.390 ;
        RECT 27.700 155.390 27.960 155.710 ;
        RECT 27.760 151.970 27.900 155.390 ;
        RECT 27.700 151.650 27.960 151.970 ;
        RECT 28.220 150.610 28.360 156.070 ;
        RECT 31.440 153.410 31.580 158.790 ;
        RECT 32.360 156.730 32.500 164.230 ;
        RECT 35.120 164.210 35.260 168.910 ;
        RECT 36.960 164.550 37.100 169.330 ;
        RECT 37.420 169.310 37.560 172.730 ;
        RECT 39.260 171.010 39.400 175.110 ;
        RECT 39.200 170.690 39.460 171.010 ;
        RECT 39.260 169.900 39.400 170.690 ;
        RECT 39.720 170.670 39.860 182.930 ;
        RECT 41.040 179.870 41.300 180.190 ;
        RECT 40.120 177.830 40.380 178.150 ;
        RECT 40.180 176.450 40.320 177.830 ;
        RECT 41.100 177.470 41.240 179.870 ;
        RECT 40.580 177.150 40.840 177.470 ;
        RECT 41.040 177.150 41.300 177.470 ;
        RECT 40.120 176.130 40.380 176.450 ;
        RECT 40.640 175.770 40.780 177.150 ;
        RECT 40.580 175.450 40.840 175.770 ;
        RECT 39.660 170.350 39.920 170.670 ;
        RECT 40.120 169.900 40.380 169.990 ;
        RECT 39.260 169.760 40.380 169.900 ;
        RECT 40.120 169.670 40.380 169.760 ;
        RECT 37.360 168.990 37.620 169.310 ;
        RECT 36.900 164.230 37.160 164.550 ;
        RECT 37.420 164.210 37.560 168.990 ;
        RECT 38.280 166.610 38.540 166.930 ;
        RECT 35.060 163.890 35.320 164.210 ;
        RECT 37.360 163.890 37.620 164.210 ;
        RECT 35.120 160.130 35.260 163.890 ;
        RECT 38.340 162.850 38.480 166.610 ;
        RECT 40.180 165.570 40.320 169.670 ;
        RECT 40.640 169.310 40.780 175.450 ;
        RECT 41.560 175.090 41.700 188.370 ;
        RECT 41.960 176.130 42.220 176.450 ;
        RECT 41.500 174.770 41.760 175.090 ;
        RECT 42.020 173.730 42.160 176.130 ;
        RECT 41.960 173.410 42.220 173.730 ;
        RECT 41.040 172.730 41.300 173.050 ;
        RECT 41.100 171.010 41.240 172.730 ;
        RECT 41.040 170.690 41.300 171.010 ;
        RECT 40.580 168.990 40.840 169.310 ;
        RECT 42.480 167.610 42.620 191.430 ;
        RECT 42.880 190.750 43.140 191.070 ;
        RECT 42.940 189.030 43.080 190.750 ;
        RECT 42.880 188.710 43.140 189.030 ;
        RECT 43.400 187.330 43.540 192.450 ;
        RECT 48.920 191.750 49.060 194.150 ;
        RECT 53.980 192.770 54.120 196.190 ;
        RECT 55.300 193.470 55.560 193.790 ;
        RECT 53.920 192.450 54.180 192.770 ;
        RECT 55.360 191.750 55.500 193.470 ;
        RECT 48.860 191.430 49.120 191.750 ;
        RECT 53.000 191.430 53.260 191.750 ;
        RECT 55.300 191.430 55.560 191.750 ;
        RECT 51.620 190.750 51.880 191.070 ;
        RECT 51.680 190.050 51.820 190.750 ;
        RECT 53.060 190.050 53.200 191.430 ;
        RECT 43.800 189.730 44.060 190.050 ;
        RECT 49.780 189.730 50.040 190.050 ;
        RECT 51.620 189.730 51.880 190.050 ;
        RECT 53.000 189.730 53.260 190.050 ;
        RECT 43.860 189.565 44.000 189.730 ;
        RECT 43.790 189.195 44.070 189.565 ;
        RECT 43.800 189.050 44.060 189.195 ;
        RECT 43.340 187.010 43.600 187.330 ;
        RECT 42.880 180.210 43.140 180.530 ;
        RECT 42.940 179.170 43.080 180.210 ;
        RECT 42.880 178.850 43.140 179.170 ;
        RECT 43.400 172.370 43.540 187.010 ;
        RECT 49.840 186.310 49.980 189.730 ;
        RECT 55.360 189.370 55.500 191.430 ;
        RECT 55.300 189.050 55.560 189.370 ;
        RECT 54.380 188.030 54.640 188.350 ;
        RECT 54.440 186.990 54.580 188.030 ;
        RECT 53.000 186.670 53.260 186.990 ;
        RECT 54.380 186.670 54.640 186.990 ;
        RECT 49.320 185.990 49.580 186.310 ;
        RECT 49.780 185.990 50.040 186.310 ;
        RECT 45.180 183.950 45.440 184.270 ;
        RECT 45.240 180.190 45.380 183.950 ;
        RECT 49.380 183.590 49.520 185.990 ;
        RECT 49.840 184.610 49.980 185.990 ;
        RECT 50.240 185.310 50.500 185.630 ;
        RECT 49.780 184.290 50.040 184.610 ;
        RECT 50.300 183.930 50.440 185.310 ;
        RECT 50.240 183.610 50.500 183.930 ;
        RECT 52.080 183.610 52.340 183.930 ;
        RECT 49.320 183.270 49.580 183.590 ;
        RECT 50.300 181.890 50.440 183.610 ;
        RECT 51.160 183.270 51.420 183.590 ;
        RECT 50.240 181.570 50.500 181.890 ;
        RECT 45.640 180.550 45.900 180.870 ;
        RECT 49.780 180.550 50.040 180.870 ;
        RECT 45.180 179.870 45.440 180.190 ;
        RECT 44.720 177.830 44.980 178.150 ;
        RECT 44.780 176.450 44.920 177.830 ;
        RECT 44.720 176.130 44.980 176.450 ;
        RECT 43.340 172.050 43.600 172.370 ;
        RECT 45.240 172.030 45.380 179.870 ;
        RECT 45.700 179.170 45.840 180.550 ;
        RECT 49.840 179.170 49.980 180.550 ;
        RECT 51.220 179.170 51.360 183.270 ;
        RECT 45.640 178.850 45.900 179.170 ;
        RECT 49.780 178.850 50.040 179.170 ;
        RECT 51.160 178.850 51.420 179.170 ;
        RECT 51.620 178.510 51.880 178.830 ;
        RECT 47.480 178.170 47.740 178.490 ;
        RECT 49.780 178.170 50.040 178.490 ;
        RECT 51.160 178.170 51.420 178.490 ;
        RECT 46.560 175.790 46.820 176.110 ;
        RECT 46.100 172.050 46.360 172.370 ;
        RECT 45.180 171.710 45.440 172.030 ;
        RECT 45.240 169.990 45.380 171.710 ;
        RECT 45.180 169.670 45.440 169.990 ;
        RECT 46.160 169.650 46.300 172.050 ;
        RECT 46.100 169.330 46.360 169.650 ;
        RECT 41.500 167.290 41.760 167.610 ;
        RECT 42.420 167.290 42.680 167.610 ;
        RECT 43.340 167.290 43.600 167.610 ;
        RECT 40.120 165.250 40.380 165.570 ;
        RECT 41.560 165.230 41.700 167.290 ;
        RECT 43.400 165.570 43.540 167.290 ;
        RECT 43.800 166.270 44.060 166.590 ;
        RECT 43.340 165.250 43.600 165.570 ;
        RECT 41.500 164.910 41.760 165.230 ;
        RECT 43.860 164.550 44.000 166.270 ;
        RECT 41.500 164.290 41.760 164.550 ;
        RECT 41.500 164.230 43.080 164.290 ;
        RECT 43.800 164.230 44.060 164.550 ;
        RECT 45.180 164.290 45.440 164.550 ;
        RECT 46.160 164.290 46.300 169.330 ;
        RECT 46.620 165.570 46.760 175.790 ;
        RECT 47.540 175.430 47.680 178.170 ;
        RECT 48.400 177.830 48.660 178.150 ;
        RECT 48.860 177.830 49.120 178.150 ;
        RECT 48.460 175.430 48.600 177.830 ;
        RECT 48.920 176.450 49.060 177.830 ;
        RECT 49.320 177.150 49.580 177.470 ;
        RECT 48.860 176.130 49.120 176.450 ;
        RECT 49.380 175.850 49.520 177.150 ;
        RECT 49.840 176.450 49.980 178.170 ;
        RECT 51.220 176.450 51.360 178.170 ;
        RECT 49.780 176.130 50.040 176.450 ;
        RECT 51.160 176.130 51.420 176.450 ;
        RECT 49.380 175.770 49.980 175.850 ;
        RECT 49.380 175.710 50.040 175.770 ;
        RECT 47.480 175.110 47.740 175.430 ;
        RECT 48.400 175.110 48.660 175.430 ;
        RECT 47.540 166.590 47.680 175.110 ;
        RECT 49.380 169.990 49.520 175.710 ;
        RECT 49.780 175.450 50.040 175.710 ;
        RECT 51.680 175.090 51.820 178.510 ;
        RECT 52.140 176.110 52.280 183.610 ;
        RECT 52.540 182.590 52.800 182.910 ;
        RECT 52.600 178.490 52.740 182.590 ;
        RECT 53.060 180.870 53.200 186.670 ;
        RECT 53.920 186.220 54.180 186.310 ;
        RECT 54.440 186.220 54.580 186.670 ;
        RECT 55.360 186.310 55.500 189.050 ;
        RECT 56.220 188.710 56.480 189.030 ;
        RECT 55.760 188.030 56.020 188.350 ;
        RECT 53.920 186.080 54.580 186.220 ;
        RECT 53.920 185.990 54.180 186.080 ;
        RECT 53.920 182.590 54.180 182.910 ;
        RECT 53.980 181.550 54.120 182.590 ;
        RECT 53.920 181.230 54.180 181.550 ;
        RECT 53.000 180.725 53.260 180.870 ;
        RECT 52.990 180.355 53.270 180.725 ;
        RECT 53.000 179.870 53.260 180.190 ;
        RECT 53.060 178.490 53.200 179.870 ;
        RECT 52.540 178.170 52.800 178.490 ;
        RECT 53.000 178.170 53.260 178.490 ;
        RECT 53.980 176.110 54.120 181.230 ;
        RECT 54.440 177.810 54.580 186.080 ;
        RECT 55.300 185.990 55.560 186.310 ;
        RECT 55.820 184.270 55.960 188.030 ;
        RECT 56.280 186.310 56.420 188.710 ;
        RECT 56.220 185.990 56.480 186.310 ;
        RECT 56.280 185.630 56.420 185.990 ;
        RECT 56.220 185.310 56.480 185.630 ;
        RECT 55.760 183.950 56.020 184.270 ;
        RECT 56.280 183.930 56.420 185.310 ;
        RECT 56.220 183.610 56.480 183.930 ;
        RECT 56.740 181.290 56.880 196.190 ;
        RECT 60.360 193.470 60.620 193.790 ;
        RECT 57.600 191.430 57.860 191.750 ;
        RECT 57.660 187.330 57.800 191.430 ;
        RECT 59.440 191.090 59.700 191.410 ;
        RECT 58.520 188.370 58.780 188.690 ;
        RECT 58.580 187.330 58.720 188.370 ;
        RECT 59.500 188.350 59.640 191.090 ;
        RECT 60.420 189.370 60.560 193.470 ;
        RECT 60.820 192.680 61.080 192.770 ;
        RECT 60.820 192.540 61.480 192.680 ;
        RECT 60.820 192.450 61.080 192.540 ;
        RECT 60.820 191.430 61.080 191.750 ;
        RECT 60.360 189.050 60.620 189.370 ;
        RECT 59.440 188.030 59.700 188.350 ;
        RECT 57.600 187.010 57.860 187.330 ;
        RECT 58.520 187.010 58.780 187.330 ;
        RECT 58.580 186.650 58.720 187.010 ;
        RECT 58.520 186.330 58.780 186.650 ;
        RECT 58.580 183.590 58.720 186.330 ;
        RECT 60.420 185.970 60.560 189.050 ;
        RECT 60.880 188.690 61.020 191.430 ;
        RECT 61.340 190.050 61.480 192.540 ;
        RECT 61.740 190.750 62.000 191.070 ;
        RECT 61.280 189.730 61.540 190.050 ;
        RECT 60.820 188.370 61.080 188.690 ;
        RECT 60.360 185.650 60.620 185.970 ;
        RECT 58.520 183.270 58.780 183.590 ;
        RECT 60.820 182.930 61.080 183.250 ;
        RECT 60.880 181.890 61.020 182.930 ;
        RECT 57.140 181.570 57.400 181.890 ;
        RECT 60.820 181.570 61.080 181.890 ;
        RECT 56.280 181.150 56.880 181.290 ;
        RECT 57.200 181.210 57.340 181.570 ;
        RECT 60.360 181.230 60.620 181.550 ;
        RECT 55.760 180.725 56.020 180.870 ;
        RECT 55.750 180.355 56.030 180.725 ;
        RECT 55.300 179.870 55.560 180.190 ;
        RECT 55.360 178.830 55.500 179.870 ;
        RECT 55.300 178.510 55.560 178.830 ;
        RECT 54.840 178.060 55.100 178.150 ;
        RECT 56.280 178.060 56.420 181.150 ;
        RECT 57.140 180.890 57.400 181.210 ;
        RECT 57.600 180.550 57.860 180.870 ;
        RECT 56.680 180.210 56.940 180.530 ;
        RECT 54.840 177.920 56.420 178.060 ;
        RECT 54.840 177.830 55.100 177.920 ;
        RECT 54.380 177.490 54.640 177.810 ;
        RECT 52.080 175.790 52.340 176.110 ;
        RECT 53.920 175.790 54.180 176.110 ;
        RECT 52.540 175.110 52.800 175.430 ;
        RECT 54.440 175.170 54.580 177.490 ;
        RECT 51.160 174.770 51.420 175.090 ;
        RECT 51.620 174.770 51.880 175.090 ;
        RECT 52.080 174.770 52.340 175.090 ;
        RECT 50.240 170.010 50.500 170.330 ;
        RECT 49.320 169.670 49.580 169.990 ;
        RECT 49.780 169.670 50.040 169.990 ;
        RECT 49.840 168.290 49.980 169.670 ;
        RECT 49.780 167.970 50.040 168.290 ;
        RECT 49.780 167.290 50.040 167.610 ;
        RECT 47.480 166.270 47.740 166.590 ;
        RECT 46.560 165.250 46.820 165.570 ;
        RECT 49.320 165.250 49.580 165.570 ;
        RECT 47.020 164.910 47.280 165.230 ;
        RECT 45.180 164.230 46.300 164.290 ;
        RECT 41.560 164.210 43.080 164.230 ;
        RECT 41.560 164.150 43.140 164.210 ;
        RECT 45.240 164.150 46.300 164.230 ;
        RECT 42.880 163.890 43.140 164.150 ;
        RECT 46.160 163.870 46.300 164.150 ;
        RECT 45.640 163.550 45.900 163.870 ;
        RECT 46.100 163.550 46.360 163.870 ;
        RECT 38.280 162.530 38.540 162.850 ;
        RECT 35.060 159.810 35.320 160.130 ;
        RECT 35.060 159.130 35.320 159.450 ;
        RECT 34.600 158.790 34.860 159.110 ;
        RECT 34.140 158.450 34.400 158.770 ;
        RECT 32.760 158.110 33.020 158.430 ;
        RECT 31.840 156.410 32.100 156.730 ;
        RECT 32.300 156.410 32.560 156.730 ;
        RECT 30.980 153.270 31.580 153.410 ;
        RECT 28.160 150.290 28.420 150.610 ;
        RECT 29.080 148.250 29.340 148.570 ;
        RECT 27.700 147.230 27.960 147.550 ;
        RECT 27.760 146.190 27.900 147.230 ;
        RECT 27.700 145.870 27.960 146.190 ;
        RECT 27.240 145.190 27.500 145.510 ;
        RECT 29.140 143.810 29.280 148.250 ;
        RECT 30.980 148.230 31.120 153.270 ;
        RECT 31.900 151.630 32.040 156.410 ;
        RECT 32.820 154.010 32.960 158.110 ;
        RECT 34.200 157.070 34.340 158.450 ;
        RECT 34.660 157.070 34.800 158.790 ;
        RECT 35.120 157.410 35.260 159.130 ;
        RECT 42.420 158.790 42.680 159.110 ;
        RECT 39.660 158.110 39.920 158.430 ;
        RECT 40.580 158.110 40.840 158.430 ;
        RECT 35.060 157.090 35.320 157.410 ;
        RECT 34.140 156.750 34.400 157.070 ;
        RECT 34.600 156.750 34.860 157.070 ;
        RECT 33.680 156.410 33.940 156.730 ;
        RECT 33.740 154.690 33.880 156.410 ;
        RECT 33.680 154.370 33.940 154.690 ;
        RECT 32.760 153.690 33.020 154.010 ;
        RECT 31.840 151.310 32.100 151.630 ;
        RECT 31.380 150.290 31.640 150.610 ;
        RECT 31.440 148.230 31.580 150.290 ;
        RECT 31.900 148.230 32.040 151.310 ;
        RECT 34.200 148.230 34.340 156.750 ;
        RECT 39.720 152.990 39.860 158.110 ;
        RECT 40.120 153.580 40.380 153.670 ;
        RECT 40.640 153.580 40.780 158.110 ;
        RECT 42.480 157.410 42.620 158.790 ;
        RECT 45.700 158.770 45.840 163.550 ;
        RECT 46.560 158.790 46.820 159.110 ;
        RECT 45.700 158.630 46.300 158.770 ;
        RECT 45.640 158.110 45.900 158.430 ;
        RECT 42.420 157.090 42.680 157.410 ;
        RECT 41.040 156.410 41.300 156.730 ;
        RECT 41.100 154.690 41.240 156.410 ;
        RECT 41.040 154.370 41.300 154.690 ;
        RECT 40.120 153.440 40.780 153.580 ;
        RECT 40.120 153.350 40.380 153.440 ;
        RECT 41.960 153.010 42.220 153.330 ;
        RECT 35.060 152.670 35.320 152.990 ;
        RECT 39.660 152.670 39.920 152.990 ;
        RECT 35.120 149.330 35.260 152.670 ;
        RECT 41.500 150.970 41.760 151.290 ;
        RECT 34.660 149.190 35.260 149.330 ;
        RECT 30.920 147.910 31.180 148.230 ;
        RECT 31.380 147.910 31.640 148.230 ;
        RECT 31.840 147.910 32.100 148.230 ;
        RECT 34.140 147.910 34.400 148.230 ;
        RECT 31.900 146.530 32.040 147.910 ;
        RECT 31.840 146.210 32.100 146.530 ;
        RECT 33.680 144.850 33.940 145.170 ;
        RECT 29.080 143.490 29.340 143.810 ;
        RECT 26.780 143.150 27.040 143.470 ;
        RECT 31.380 141.790 31.640 142.110 ;
        RECT 31.440 140.750 31.580 141.790 ;
        RECT 26.320 140.490 26.580 140.750 ;
        RECT 26.320 140.430 27.900 140.490 ;
        RECT 31.380 140.430 31.640 140.750 ;
        RECT 26.380 140.350 27.900 140.430 ;
        RECT 33.740 140.410 33.880 144.850 ;
        RECT 34.660 143.130 34.800 149.190 ;
        RECT 35.060 148.250 35.320 148.570 ;
        RECT 35.120 143.130 35.260 148.250 ;
        RECT 36.900 147.910 37.160 148.230 ;
        RECT 35.980 145.530 36.240 145.850 ;
        RECT 36.040 143.810 36.180 145.530 ;
        RECT 35.980 143.490 36.240 143.810 ;
        RECT 34.600 142.810 34.860 143.130 ;
        RECT 35.060 142.810 35.320 143.130 ;
        RECT 36.960 140.410 37.100 147.910 ;
        RECT 41.560 145.850 41.700 150.970 ;
        RECT 41.500 145.530 41.760 145.850 ;
        RECT 38.740 145.190 39.000 145.510 ;
        RECT 38.800 140.750 38.940 145.190 ;
        RECT 39.200 143.150 39.460 143.470 ;
        RECT 38.740 140.430 39.000 140.750 ;
        RECT 24.020 136.350 24.280 136.670 ;
        RECT 24.370 135.815 25.910 136.185 ;
        RECT 27.760 135.310 27.900 140.350 ;
        RECT 31.840 140.090 32.100 140.410 ;
        RECT 33.680 140.090 33.940 140.410 ;
        RECT 36.900 140.090 37.160 140.410 ;
        RECT 28.620 139.750 28.880 140.070 ;
        RECT 28.680 138.370 28.820 139.750 ;
        RECT 31.380 139.070 31.640 139.390 ;
        RECT 28.620 138.050 28.880 138.370 ;
        RECT 31.440 137.350 31.580 139.070 ;
        RECT 31.900 137.690 32.040 140.090 ;
        RECT 34.600 139.070 34.860 139.390 ;
        RECT 37.820 139.070 38.080 139.390 ;
        RECT 31.840 137.370 32.100 137.690 ;
        RECT 29.080 137.030 29.340 137.350 ;
        RECT 31.380 137.030 31.640 137.350 ;
        RECT 27.700 134.990 27.960 135.310 ;
        RECT 29.140 134.630 29.280 137.030 ;
        RECT 29.080 134.310 29.340 134.630 ;
        RECT 26.320 132.270 26.580 132.590 ;
        RECT 24.020 131.650 24.280 131.910 ;
        RECT 23.620 131.590 24.280 131.650 ;
        RECT 23.620 131.510 24.220 131.590 ;
        RECT 21.260 130.910 21.520 131.230 ;
        RECT 20.400 128.790 21.000 128.930 ;
        RECT 20.400 127.060 20.540 128.790 ;
        RECT 21.320 128.510 21.460 130.910 ;
        RECT 23.620 130.210 23.760 131.510 ;
        RECT 24.370 130.375 25.910 130.745 ;
        RECT 23.560 129.890 23.820 130.210 ;
        RECT 23.100 128.870 23.360 129.190 ;
        RECT 21.260 128.190 21.520 128.510 ;
        RECT 21.070 127.655 22.610 128.025 ;
        RECT 20.400 126.920 21.000 127.060 ;
        RECT 20.860 126.130 21.000 126.920 ;
        RECT 20.800 125.810 21.060 126.130 ;
        RECT 18.960 125.470 19.220 125.790 ;
        RECT 19.020 121.370 19.160 125.470 ;
        RECT 20.860 124.770 21.000 125.810 ;
        RECT 20.800 124.450 21.060 124.770 ;
        RECT 21.070 122.215 22.610 122.585 ;
        RECT 18.960 121.050 19.220 121.370 ;
        RECT 23.160 119.330 23.300 128.870 ;
        RECT 23.560 128.190 23.820 128.510 ;
        RECT 23.100 119.010 23.360 119.330 ;
        RECT 15.280 118.330 15.540 118.650 ;
        RECT 15.740 118.330 16.000 118.650 ;
        RECT 15.340 115.930 15.480 118.330 ;
        RECT 15.800 116.610 15.940 118.330 ;
        RECT 21.070 116.775 22.610 117.145 ;
        RECT 23.620 116.610 23.760 128.190 ;
        RECT 26.380 126.810 26.520 132.270 ;
        RECT 29.140 131.910 29.280 134.310 ;
        RECT 34.660 131.910 34.800 139.070 ;
        RECT 37.360 136.690 37.620 137.010 ;
        RECT 37.420 135.650 37.560 136.690 ;
        RECT 37.360 135.330 37.620 135.650 ;
        RECT 37.880 134.970 38.020 139.070 ;
        RECT 39.260 135.650 39.400 143.150 ;
        RECT 41.040 142.470 41.300 142.790 ;
        RECT 39.660 142.130 39.920 142.450 ;
        RECT 39.720 139.390 39.860 142.130 ;
        RECT 39.660 139.070 39.920 139.390 ;
        RECT 39.720 135.650 39.860 139.070 ;
        RECT 41.100 136.670 41.240 142.470 ;
        RECT 42.020 142.450 42.160 153.010 ;
        RECT 42.480 151.970 42.620 157.090 ;
        RECT 45.700 156.730 45.840 158.110 ;
        RECT 45.640 156.410 45.900 156.730 ;
        RECT 44.720 155.730 44.980 156.050 ;
        RECT 44.780 154.350 44.920 155.730 ;
        RECT 44.720 154.030 44.980 154.350 ;
        RECT 42.420 151.880 42.680 151.970 ;
        RECT 42.420 151.740 43.080 151.880 ;
        RECT 42.420 151.650 42.680 151.740 ;
        RECT 42.420 149.950 42.680 150.270 ;
        RECT 42.480 149.250 42.620 149.950 ;
        RECT 42.420 148.930 42.680 149.250 ;
        RECT 42.940 148.230 43.080 151.740 ;
        RECT 45.700 151.290 45.840 156.410 ;
        RECT 45.640 150.970 45.900 151.290 ;
        RECT 43.800 149.950 44.060 150.270 ;
        RECT 43.860 148.570 44.000 149.950 ;
        RECT 43.800 148.250 44.060 148.570 ;
        RECT 42.880 147.910 43.140 148.230 ;
        RECT 43.340 147.570 43.600 147.890 ;
        RECT 42.420 145.530 42.680 145.850 ;
        RECT 41.960 142.130 42.220 142.450 ;
        RECT 42.480 140.750 42.620 145.530 ;
        RECT 43.400 141.090 43.540 147.570 ;
        RECT 43.340 140.770 43.600 141.090 ;
        RECT 42.420 140.430 42.680 140.750 ;
        RECT 41.500 140.090 41.760 140.410 ;
        RECT 41.560 138.030 41.700 140.090 ;
        RECT 41.960 139.410 42.220 139.730 ;
        RECT 41.500 137.710 41.760 138.030 ;
        RECT 41.040 136.350 41.300 136.670 ;
        RECT 39.200 135.330 39.460 135.650 ;
        RECT 39.660 135.330 39.920 135.650 ;
        RECT 37.820 134.650 38.080 134.970 ;
        RECT 39.260 132.930 39.400 135.330 ;
        RECT 41.100 134.630 41.240 136.350 ;
        RECT 42.020 135.650 42.160 139.410 ;
        RECT 42.480 138.370 42.620 140.430 ;
        RECT 42.420 138.050 42.680 138.370 ;
        RECT 42.480 135.650 42.620 138.050 ;
        RECT 43.400 137.690 43.540 140.770 ;
        RECT 45.640 139.070 45.900 139.390 ;
        RECT 44.720 137.710 44.980 138.030 ;
        RECT 43.340 137.370 43.600 137.690 ;
        RECT 42.880 136.690 43.140 137.010 ;
        RECT 41.960 135.330 42.220 135.650 ;
        RECT 42.420 135.330 42.680 135.650 ;
        RECT 42.940 135.050 43.080 136.690 ;
        RECT 42.480 134.970 43.080 135.050 ;
        RECT 43.400 134.970 43.540 137.370 ;
        RECT 44.780 134.970 44.920 137.710 ;
        RECT 45.700 137.350 45.840 139.070 ;
        RECT 45.640 137.030 45.900 137.350 ;
        RECT 45.180 136.690 45.440 137.010 ;
        RECT 45.240 135.650 45.380 136.690 ;
        RECT 45.180 135.330 45.440 135.650 ;
        RECT 45.700 135.050 45.840 137.030 ;
        RECT 42.420 134.910 43.080 134.970 ;
        RECT 42.420 134.650 42.680 134.910 ;
        RECT 43.340 134.650 43.600 134.970 ;
        RECT 44.720 134.650 44.980 134.970 ;
        RECT 45.240 134.910 45.840 135.050 ;
        RECT 41.040 134.310 41.300 134.630 ;
        RECT 35.060 132.610 35.320 132.930 ;
        RECT 39.200 132.610 39.460 132.930 ;
        RECT 29.080 131.590 29.340 131.910 ;
        RECT 34.600 131.590 34.860 131.910 ;
        RECT 26.780 131.250 27.040 131.570 ;
        RECT 26.840 128.510 26.980 131.250 ;
        RECT 28.160 128.870 28.420 129.190 ;
        RECT 26.780 128.190 27.040 128.510 ;
        RECT 26.320 126.490 26.580 126.810 ;
        RECT 24.370 124.935 25.910 125.305 ;
        RECT 28.220 124.770 28.360 128.870 ;
        RECT 29.140 126.470 29.280 131.590 ;
        RECT 31.840 131.250 32.100 131.570 ;
        RECT 31.900 128.850 32.040 131.250 ;
        RECT 35.120 129.530 35.260 132.610 ;
        RECT 41.100 132.250 41.240 134.310 ;
        RECT 41.960 133.630 42.220 133.950 ;
        RECT 41.040 131.930 41.300 132.250 ;
        RECT 39.660 130.910 39.920 131.230 ;
        RECT 39.720 129.530 39.860 130.910 ;
        RECT 41.100 129.870 41.240 131.930 ;
        RECT 41.040 129.550 41.300 129.870 ;
        RECT 35.060 129.210 35.320 129.530 ;
        RECT 39.200 129.210 39.460 129.530 ;
        RECT 39.660 129.210 39.920 129.530 ;
        RECT 31.840 128.530 32.100 128.850 ;
        RECT 30.000 128.190 30.260 128.510 ;
        RECT 35.060 128.190 35.320 128.510 ;
        RECT 37.820 128.190 38.080 128.510 ;
        RECT 30.060 126.470 30.200 128.190 ;
        RECT 34.600 126.830 34.860 127.150 ;
        RECT 29.080 126.150 29.340 126.470 ;
        RECT 30.000 126.150 30.260 126.470 ;
        RECT 32.760 126.210 33.020 126.470 ;
        RECT 32.760 126.150 33.420 126.210 ;
        RECT 28.160 124.450 28.420 124.770 ;
        RECT 27.240 123.770 27.500 124.090 ;
        RECT 27.300 122.050 27.440 123.770 ;
        RECT 29.140 123.410 29.280 126.150 ;
        RECT 32.820 126.070 33.420 126.150 ;
        RECT 32.760 125.470 33.020 125.790 ;
        RECT 29.540 123.430 29.800 123.750 ;
        RECT 32.300 123.430 32.560 123.750 ;
        RECT 29.080 123.090 29.340 123.410 ;
        RECT 29.600 122.130 29.740 123.430 ;
        RECT 31.840 122.750 32.100 123.070 ;
        RECT 27.240 121.730 27.500 122.050 ;
        RECT 29.140 121.990 29.740 122.130 ;
        RECT 29.140 121.370 29.280 121.990 ;
        RECT 29.540 121.390 29.800 121.710 ;
        RECT 31.900 121.450 32.040 122.750 ;
        RECT 32.360 122.050 32.500 123.430 ;
        RECT 32.300 121.730 32.560 122.050 ;
        RECT 29.080 121.050 29.340 121.370 ;
        RECT 24.020 120.030 24.280 120.350 ;
        RECT 15.740 116.290 16.000 116.610 ;
        RECT 16.660 116.290 16.920 116.610 ;
        RECT 23.560 116.290 23.820 116.610 ;
        RECT 15.280 115.610 15.540 115.930 ;
        RECT 10.220 114.590 10.480 114.910 ;
        RECT 4.230 113.035 4.510 113.405 ;
        RECT 4.240 112.890 4.500 113.035 ;
        RECT 8.840 112.210 9.100 112.530 ;
        RECT 4.240 110.005 4.500 110.150 ;
        RECT 0.560 109.490 0.820 109.810 ;
        RECT 4.230 109.635 4.510 110.005 ;
        RECT 8.900 107.770 9.040 112.210 ;
        RECT 9.300 109.830 9.560 110.150 ;
        RECT 8.840 107.450 9.100 107.770 ;
        RECT 6.530 105.555 6.810 105.925 ;
        RECT 6.600 101.650 6.740 105.555 ;
        RECT 8.900 104.370 9.040 107.450 ;
        RECT 7.460 104.050 7.720 104.370 ;
        RECT 8.840 104.050 9.100 104.370 ;
        RECT 7.520 103.010 7.660 104.050 ;
        RECT 7.460 102.690 7.720 103.010 ;
        RECT 8.900 102.670 9.040 104.050 ;
        RECT 9.360 102.670 9.500 109.830 ;
        RECT 10.280 107.770 10.420 114.590 ;
        RECT 15.340 110.150 15.480 115.610 ;
        RECT 16.720 115.590 16.860 116.290 ;
        RECT 16.660 115.270 16.920 115.590 ;
        RECT 17.120 115.270 17.380 115.590 ;
        RECT 16.200 114.930 16.460 115.250 ;
        RECT 16.260 113.550 16.400 114.930 ;
        RECT 16.660 114.590 16.920 114.910 ;
        RECT 16.200 113.230 16.460 113.550 ;
        RECT 13.900 109.830 14.160 110.150 ;
        RECT 15.280 109.830 15.540 110.150 ;
        RECT 11.600 109.150 11.860 109.470 ;
        RECT 10.220 107.450 10.480 107.770 ;
        RECT 9.760 107.110 10.020 107.430 ;
        RECT 8.840 102.350 9.100 102.670 ;
        RECT 9.300 102.350 9.560 102.670 ;
        RECT 9.820 101.990 9.960 107.110 ;
        RECT 9.760 101.670 10.020 101.990 ;
        RECT 6.540 101.330 6.800 101.650 ;
        RECT 4.230 99.435 4.510 99.805 ;
        RECT 4.300 99.270 4.440 99.435 ;
        RECT 10.280 99.270 10.420 107.450 ;
        RECT 10.680 106.430 10.940 106.750 ;
        RECT 10.740 102.330 10.880 106.430 ;
        RECT 11.660 102.670 11.800 109.150 ;
        RECT 13.960 108.360 14.100 109.830 ;
        RECT 15.340 108.450 15.480 109.830 ;
        RECT 13.500 108.220 14.100 108.360 ;
        RECT 13.500 105.730 13.640 108.220 ;
        RECT 14.360 108.130 14.620 108.450 ;
        RECT 15.280 108.130 15.540 108.450 ;
        RECT 13.900 107.450 14.160 107.770 ;
        RECT 13.440 105.410 13.700 105.730 ;
        RECT 11.600 102.350 11.860 102.670 ;
        RECT 13.500 102.330 13.640 105.410 ;
        RECT 13.960 104.710 14.100 107.450 ;
        RECT 13.900 104.390 14.160 104.710 ;
        RECT 14.420 102.670 14.560 108.130 ;
        RECT 15.280 107.450 15.540 107.770 ;
        RECT 15.340 105.730 15.480 107.450 ;
        RECT 15.280 105.410 15.540 105.730 ;
        RECT 15.740 104.730 16.000 105.050 ;
        RECT 14.820 104.390 15.080 104.710 ;
        RECT 14.360 102.350 14.620 102.670 ;
        RECT 10.680 102.010 10.940 102.330 ;
        RECT 13.440 102.010 13.700 102.330 ;
        RECT 14.880 100.290 15.020 104.390 ;
        RECT 15.800 103.010 15.940 104.730 ;
        RECT 16.720 104.710 16.860 114.590 ;
        RECT 17.180 113.210 17.320 115.270 ;
        RECT 18.500 114.930 18.760 115.250 ;
        RECT 17.120 112.890 17.380 113.210 ;
        RECT 18.560 112.530 18.700 114.930 ;
        RECT 23.100 114.590 23.360 114.910 ;
        RECT 19.420 113.230 19.680 113.550 ;
        RECT 19.480 112.870 19.620 113.230 ;
        RECT 19.420 112.550 19.680 112.870 ;
        RECT 18.500 112.210 18.760 112.530 ;
        RECT 18.960 109.490 19.220 109.810 ;
        RECT 18.500 105.070 18.760 105.390 ;
        RECT 16.660 104.390 16.920 104.710 ;
        RECT 18.040 104.390 18.300 104.710 ;
        RECT 18.100 103.090 18.240 104.390 ;
        RECT 15.740 102.690 16.000 103.010 ;
        RECT 16.260 102.950 18.240 103.090 ;
        RECT 15.270 102.155 15.550 102.525 ;
        RECT 15.280 102.010 15.540 102.155 ;
        RECT 15.740 101.670 16.000 101.990 ;
        RECT 13.900 99.970 14.160 100.290 ;
        RECT 14.820 99.970 15.080 100.290 ;
        RECT 4.240 98.950 4.500 99.270 ;
        RECT 10.220 98.950 10.480 99.270 ;
        RECT 11.600 98.950 11.860 99.270 ;
        RECT 10.680 98.270 10.940 98.590 ;
        RECT 7.000 96.570 7.260 96.890 ;
        RECT 7.060 88.730 7.200 96.570 ;
        RECT 10.740 94.850 10.880 98.270 ;
        RECT 11.660 94.850 11.800 98.950 ;
        RECT 13.960 96.290 14.100 99.970 ;
        RECT 15.800 99.610 15.940 101.670 ;
        RECT 16.260 99.950 16.400 102.950 ;
        RECT 17.580 102.350 17.840 102.670 ;
        RECT 16.660 101.330 16.920 101.650 ;
        RECT 16.200 99.630 16.460 99.950 ;
        RECT 15.740 99.290 16.000 99.610 ;
        RECT 15.740 98.610 16.000 98.930 ;
        RECT 14.360 98.270 14.620 98.590 ;
        RECT 14.420 96.890 14.560 98.270 ;
        RECT 15.800 97.570 15.940 98.610 ;
        RECT 16.260 97.570 16.400 99.630 ;
        RECT 15.740 97.250 16.000 97.570 ;
        RECT 16.200 97.250 16.460 97.570 ;
        RECT 14.360 96.570 14.620 96.890 ;
        RECT 16.720 96.670 16.860 101.330 ;
        RECT 13.500 96.150 14.100 96.290 ;
        RECT 16.260 96.530 16.860 96.670 ;
        RECT 17.640 96.550 17.780 102.350 ;
        RECT 18.100 101.990 18.240 102.950 ;
        RECT 18.560 102.330 18.700 105.070 ;
        RECT 19.020 104.370 19.160 109.490 ;
        RECT 19.480 107.770 19.620 112.550 ;
        RECT 23.160 112.530 23.300 114.590 ;
        RECT 24.080 113.210 24.220 120.030 ;
        RECT 24.370 119.495 25.910 119.865 ;
        RECT 26.320 114.590 26.580 114.910 ;
        RECT 24.370 114.055 25.910 114.425 ;
        RECT 26.380 113.550 26.520 114.590 ;
        RECT 26.320 113.230 26.580 113.550 ;
        RECT 24.020 112.890 24.280 113.210 ;
        RECT 23.100 112.210 23.360 112.530 ;
        RECT 21.070 111.335 22.610 111.705 ;
        RECT 23.160 107.770 23.300 112.210 ;
        RECT 24.080 112.190 24.220 112.890 ;
        RECT 29.080 112.550 29.340 112.870 ;
        RECT 29.600 112.610 29.740 121.390 ;
        RECT 30.520 121.310 32.040 121.450 ;
        RECT 30.000 120.940 30.260 121.030 ;
        RECT 30.520 120.940 30.660 121.310 ;
        RECT 31.900 121.030 32.040 121.310 ;
        RECT 30.000 120.800 30.660 120.940 ;
        RECT 30.000 120.710 30.260 120.800 ;
        RECT 30.000 114.590 30.260 114.910 ;
        RECT 30.060 113.210 30.200 114.590 ;
        RECT 30.000 112.890 30.260 113.210 ;
        RECT 24.020 111.870 24.280 112.190 ;
        RECT 28.160 111.870 28.420 112.190 ;
        RECT 23.560 109.830 23.820 110.150 ;
        RECT 23.620 107.770 23.760 109.830 ;
        RECT 24.370 108.615 25.910 108.985 ;
        RECT 28.220 108.110 28.360 111.870 ;
        RECT 29.140 109.890 29.280 112.550 ;
        RECT 29.600 112.470 30.200 112.610 ;
        RECT 29.540 111.870 29.800 112.190 ;
        RECT 28.680 109.750 29.280 109.890 ;
        RECT 28.160 107.790 28.420 108.110 ;
        RECT 28.680 107.770 28.820 109.750 ;
        RECT 29.080 109.150 29.340 109.470 ;
        RECT 19.420 107.450 19.680 107.770 ;
        RECT 23.100 107.450 23.360 107.770 ;
        RECT 23.560 107.450 23.820 107.770 ;
        RECT 28.620 107.450 28.880 107.770 ;
        RECT 19.480 105.730 19.620 107.450 ;
        RECT 19.880 106.430 20.140 106.750 ;
        RECT 20.340 106.430 20.600 106.750 ;
        RECT 19.940 105.730 20.080 106.430 ;
        RECT 19.420 105.410 19.680 105.730 ;
        RECT 19.880 105.410 20.140 105.730 ;
        RECT 20.400 105.390 20.540 106.430 ;
        RECT 21.070 105.895 22.610 106.265 ;
        RECT 20.340 105.070 20.600 105.390 ;
        RECT 23.160 104.710 23.300 107.450 ;
        RECT 28.680 105.730 28.820 107.450 ;
        RECT 28.620 105.410 28.880 105.730 ;
        RECT 29.140 105.050 29.280 109.150 ;
        RECT 29.080 104.730 29.340 105.050 ;
        RECT 29.600 104.710 29.740 111.870 ;
        RECT 23.100 104.390 23.360 104.710 ;
        RECT 29.540 104.390 29.800 104.710 ;
        RECT 18.960 104.050 19.220 104.370 ;
        RECT 23.560 104.050 23.820 104.370 ;
        RECT 18.500 102.010 18.760 102.330 ;
        RECT 18.960 102.010 19.220 102.330 ;
        RECT 18.040 101.670 18.300 101.990 ;
        RECT 18.040 100.990 18.300 101.310 ;
        RECT 18.500 100.990 18.760 101.310 ;
        RECT 10.680 94.530 10.940 94.850 ;
        RECT 11.600 94.530 11.860 94.850 ;
        RECT 10.740 91.790 10.880 94.530 ;
        RECT 10.680 91.470 10.940 91.790 ;
        RECT 13.500 91.110 13.640 96.150 ;
        RECT 13.900 95.550 14.160 95.870 ;
        RECT 14.360 95.550 14.620 95.870 ;
        RECT 13.960 93.830 14.100 95.550 ;
        RECT 13.900 93.510 14.160 93.830 ;
        RECT 11.140 90.790 11.400 91.110 ;
        RECT 13.440 90.790 13.700 91.110 ;
        RECT 8.380 90.110 8.640 90.430 ;
        RECT 7.000 88.410 7.260 88.730 ;
        RECT 8.440 88.050 8.580 90.110 ;
        RECT 11.200 88.810 11.340 90.790 ;
        RECT 13.960 90.430 14.100 93.510 ;
        RECT 13.900 90.110 14.160 90.430 ;
        RECT 10.740 88.670 11.340 88.810 ;
        RECT 8.380 87.730 8.640 88.050 ;
        RECT 10.740 86.690 10.880 88.670 ;
        RECT 13.900 88.070 14.160 88.390 ;
        RECT 11.140 87.730 11.400 88.050 ;
        RECT 10.680 86.370 10.940 86.690 ;
        RECT 11.200 86.010 11.340 87.730 ;
        RECT 13.960 86.350 14.100 88.070 ;
        RECT 14.420 87.710 14.560 95.550 ;
        RECT 14.820 93.170 15.080 93.490 ;
        RECT 14.880 91.450 15.020 93.170 ;
        RECT 15.280 91.810 15.540 92.130 ;
        RECT 14.820 91.130 15.080 91.450 ;
        RECT 14.820 90.450 15.080 90.770 ;
        RECT 14.880 89.410 15.020 90.450 ;
        RECT 14.820 89.090 15.080 89.410 ;
        RECT 15.340 88.810 15.480 91.810 ;
        RECT 15.340 88.730 15.940 88.810 ;
        RECT 15.280 88.670 15.940 88.730 ;
        RECT 15.280 88.410 15.540 88.670 ;
        RECT 15.280 87.730 15.540 88.050 ;
        RECT 14.360 87.620 14.620 87.710 ;
        RECT 14.360 87.480 15.020 87.620 ;
        RECT 14.360 87.390 14.620 87.480 ;
        RECT 13.900 86.030 14.160 86.350 ;
        RECT 11.140 85.690 11.400 86.010 ;
        RECT 12.520 81.950 12.780 82.270 ;
        RECT 12.580 77.510 12.720 81.950 ;
        RECT 12.520 77.420 12.780 77.510 ;
        RECT 12.520 77.280 13.180 77.420 ;
        RECT 12.520 77.190 12.780 77.280 ;
        RECT 13.040 76.830 13.180 77.280 ;
        RECT 13.440 76.850 13.700 77.170 ;
        RECT 10.680 76.510 10.940 76.830 ;
        RECT 12.980 76.510 13.240 76.830 ;
        RECT 9.300 74.810 9.560 75.130 ;
        RECT 9.360 73.090 9.500 74.810 ;
        RECT 9.300 72.770 9.560 73.090 ;
        RECT 10.220 72.090 10.480 72.410 ;
        RECT 10.280 69.350 10.420 72.090 ;
        RECT 10.740 72.070 10.880 76.510 ;
        RECT 10.680 71.750 10.940 72.070 ;
        RECT 13.040 71.730 13.180 76.510 ;
        RECT 13.500 72.410 13.640 76.850 ;
        RECT 13.960 75.470 14.100 86.030 ;
        RECT 14.360 85.690 14.620 86.010 ;
        RECT 14.420 83.970 14.560 85.690 ;
        RECT 14.360 83.650 14.620 83.970 ;
        RECT 14.360 82.290 14.620 82.610 ;
        RECT 14.420 81.330 14.560 82.290 ;
        RECT 14.880 82.270 15.020 87.480 ;
        RECT 15.340 84.990 15.480 87.730 ;
        RECT 15.280 84.670 15.540 84.990 ;
        RECT 14.820 81.950 15.080 82.270 ;
        RECT 15.340 81.330 15.480 84.670 ;
        RECT 15.800 83.630 15.940 88.670 ;
        RECT 15.740 83.310 16.000 83.630 ;
        RECT 15.740 82.630 16.000 82.950 ;
        RECT 14.420 81.190 15.480 81.330 ;
        RECT 14.420 78.190 14.560 81.190 ;
        RECT 14.820 78.210 15.080 78.530 ;
        RECT 14.360 77.870 14.620 78.190 ;
        RECT 14.880 77.510 15.020 78.210 ;
        RECT 15.800 77.850 15.940 82.630 ;
        RECT 15.740 77.530 16.000 77.850 ;
        RECT 14.820 77.190 15.080 77.510 ;
        RECT 14.880 75.810 15.020 77.190 ;
        RECT 15.740 76.850 16.000 77.170 ;
        RECT 14.820 75.490 15.080 75.810 ;
        RECT 13.900 75.150 14.160 75.470 ;
        RECT 13.440 72.090 13.700 72.410 ;
        RECT 12.980 71.410 13.240 71.730 ;
        RECT 13.960 70.030 14.100 75.150 ;
        RECT 14.880 73.090 15.020 75.490 ;
        RECT 15.800 75.130 15.940 76.850 ;
        RECT 15.740 74.810 16.000 75.130 ;
        RECT 15.800 73.090 15.940 74.810 ;
        RECT 14.820 72.770 15.080 73.090 ;
        RECT 15.740 72.770 16.000 73.090 ;
        RECT 14.880 72.070 15.020 72.770 ;
        RECT 14.820 71.750 15.080 72.070 ;
        RECT 14.360 71.070 14.620 71.390 ;
        RECT 13.900 69.710 14.160 70.030 ;
        RECT 13.440 69.370 13.700 69.690 ;
        RECT 10.220 69.030 10.480 69.350 ;
        RECT 12.980 68.690 13.240 69.010 ;
        RECT 7.460 68.350 7.720 68.670 ;
        RECT 11.140 68.350 11.400 68.670 ;
        RECT 7.520 66.290 7.660 68.350 ;
        RECT 7.460 65.970 7.720 66.290 ;
        RECT 6.530 64.755 6.810 65.125 ;
        RECT 6.540 64.610 6.800 64.755 ;
        RECT 11.200 64.250 11.340 68.350 ;
        RECT 13.040 67.650 13.180 68.690 ;
        RECT 11.600 67.330 11.860 67.650 ;
        RECT 12.980 67.330 13.240 67.650 ;
        RECT 11.140 63.930 11.400 64.250 ;
        RECT 11.660 63.230 11.800 67.330 ;
        RECT 13.500 67.310 13.640 69.370 ;
        RECT 13.440 66.990 13.700 67.310 ;
        RECT 13.500 63.650 13.640 66.990 ;
        RECT 13.960 66.630 14.100 69.710 ;
        RECT 14.420 69.350 14.560 71.070 ;
        RECT 14.820 70.050 15.080 70.370 ;
        RECT 14.880 69.690 15.020 70.050 ;
        RECT 14.820 69.370 15.080 69.690 ;
        RECT 14.360 69.030 14.620 69.350 ;
        RECT 13.900 66.310 14.160 66.630 ;
        RECT 13.960 64.590 14.100 66.310 ;
        RECT 13.900 64.270 14.160 64.590 ;
        RECT 13.040 63.510 13.640 63.650 ;
        RECT 11.600 62.910 11.860 63.230 ;
        RECT 4.230 60.675 4.510 61.045 ;
        RECT 8.380 60.870 8.640 61.190 ;
        RECT 4.300 60.510 4.440 60.675 ;
        RECT 4.240 60.190 4.500 60.510 ;
        RECT 5.610 57.955 5.890 58.325 ;
        RECT 8.440 58.130 8.580 60.870 ;
        RECT 9.300 60.190 9.560 60.510 ;
        RECT 5.680 56.770 5.820 57.955 ;
        RECT 8.380 57.810 8.640 58.130 ;
        RECT 5.620 56.450 5.880 56.770 ;
        RECT 8.840 55.430 9.100 55.750 ;
        RECT 6.530 51.155 6.810 51.525 ;
        RECT 5.150 47.755 5.430 48.125 ;
        RECT 5.220 47.250 5.360 47.755 ;
        RECT 5.160 46.930 5.420 47.250 ;
        RECT 6.600 46.910 6.740 51.155 ;
        RECT 8.900 50.650 9.040 55.430 ;
        RECT 9.360 54.925 9.500 60.190 ;
        RECT 10.680 57.470 10.940 57.790 ;
        RECT 10.220 55.090 10.480 55.410 ;
        RECT 9.290 54.555 9.570 54.925 ;
        RECT 10.280 54.050 10.420 55.090 ;
        RECT 10.220 53.730 10.480 54.050 ;
        RECT 10.740 53.370 10.880 57.470 ;
        RECT 11.140 55.090 11.400 55.410 ;
        RECT 11.200 53.370 11.340 55.090 ;
        RECT 11.600 54.750 11.860 55.070 ;
        RECT 10.680 53.050 10.940 53.370 ;
        RECT 11.140 53.050 11.400 53.370 ;
        RECT 8.840 50.330 9.100 50.650 ;
        RECT 7.000 49.650 7.260 49.970 ;
        RECT 6.540 46.590 6.800 46.910 ;
        RECT 4.240 45.405 4.500 45.550 ;
        RECT 4.230 45.035 4.510 45.405 ;
        RECT 7.060 42.830 7.200 49.650 ;
        RECT 8.380 49.310 8.640 49.630 ;
        RECT 8.440 47.930 8.580 49.310 ;
        RECT 8.380 47.610 8.640 47.930 ;
        RECT 8.380 46.590 8.640 46.910 ;
        RECT 8.440 44.870 8.580 46.590 ;
        RECT 8.380 44.550 8.640 44.870 ;
        RECT 7.000 42.510 7.260 42.830 ;
        RECT 8.900 42.150 9.040 50.330 ;
        RECT 11.660 44.870 11.800 54.750 ;
        RECT 13.040 54.130 13.180 63.510 ;
        RECT 13.440 62.910 13.700 63.230 ;
        RECT 13.500 55.070 13.640 62.910 ;
        RECT 13.960 58.810 14.100 64.270 ;
        RECT 14.820 60.870 15.080 61.190 ;
        RECT 14.360 58.830 14.620 59.150 ;
        RECT 13.900 58.490 14.160 58.810 ;
        RECT 14.420 56.430 14.560 58.830 ;
        RECT 14.880 58.470 15.020 60.870 ;
        RECT 15.280 60.190 15.540 60.510 ;
        RECT 14.820 58.150 15.080 58.470 ;
        RECT 14.880 56.770 15.020 58.150 ;
        RECT 14.820 56.450 15.080 56.770 ;
        RECT 14.360 56.110 14.620 56.430 ;
        RECT 14.420 55.750 14.560 56.110 ;
        RECT 14.360 55.430 14.620 55.750 ;
        RECT 15.340 55.410 15.480 60.190 ;
        RECT 16.260 58.470 16.400 96.530 ;
        RECT 17.580 96.230 17.840 96.550 ;
        RECT 17.640 93.490 17.780 96.230 ;
        RECT 17.580 93.170 17.840 93.490 ;
        RECT 17.580 90.790 17.840 91.110 ;
        RECT 17.120 90.450 17.380 90.770 ;
        RECT 16.660 89.090 16.920 89.410 ;
        RECT 16.720 86.690 16.860 89.090 ;
        RECT 16.660 86.370 16.920 86.690 ;
        RECT 16.720 85.330 16.860 86.370 ;
        RECT 16.660 85.010 16.920 85.330 ;
        RECT 16.720 78.530 16.860 85.010 ;
        RECT 16.660 78.210 16.920 78.530 ;
        RECT 17.180 75.040 17.320 90.450 ;
        RECT 17.640 88.390 17.780 90.790 ;
        RECT 18.100 89.410 18.240 100.990 ;
        RECT 18.560 99.270 18.700 100.990 ;
        RECT 19.020 99.610 19.160 102.010 ;
        RECT 21.070 100.455 22.610 100.825 ;
        RECT 18.960 99.290 19.220 99.610 ;
        RECT 18.500 98.950 18.760 99.270 ;
        RECT 18.500 96.230 18.760 96.550 ;
        RECT 18.560 92.130 18.700 96.230 ;
        RECT 19.020 94.170 19.160 99.290 ;
        RECT 21.070 95.015 22.610 95.385 ;
        RECT 18.960 93.850 19.220 94.170 ;
        RECT 18.500 91.810 18.760 92.130 ;
        RECT 19.020 91.450 19.160 93.850 ;
        RECT 18.960 91.130 19.220 91.450 ;
        RECT 19.880 91.130 20.140 91.450 ;
        RECT 18.040 89.090 18.300 89.410 ;
        RECT 17.580 88.070 17.840 88.390 ;
        RECT 18.500 86.370 18.760 86.690 ;
        RECT 18.560 84.990 18.700 86.370 ;
        RECT 19.020 85.670 19.160 91.130 ;
        RECT 19.940 89.410 20.080 91.130 ;
        RECT 21.070 89.575 22.610 89.945 ;
        RECT 19.880 89.090 20.140 89.410 ;
        RECT 19.880 88.070 20.140 88.390 ;
        RECT 19.420 86.030 19.680 86.350 ;
        RECT 18.960 85.350 19.220 85.670 ;
        RECT 18.500 84.670 18.760 84.990 ;
        RECT 19.020 83.290 19.160 85.350 ;
        RECT 19.480 83.970 19.620 86.030 ;
        RECT 19.420 83.650 19.680 83.970 ;
        RECT 17.580 82.970 17.840 83.290 ;
        RECT 18.960 82.970 19.220 83.290 ;
        RECT 16.720 74.900 17.320 75.040 ;
        RECT 16.200 58.150 16.460 58.470 ;
        RECT 15.280 55.090 15.540 55.410 ;
        RECT 13.440 54.750 13.700 55.070 ;
        RECT 12.120 53.990 13.640 54.130 ;
        RECT 12.120 53.370 12.260 53.990 ;
        RECT 12.980 53.565 13.240 53.710 ;
        RECT 12.060 53.050 12.320 53.370 ;
        RECT 12.970 53.195 13.250 53.565 ;
        RECT 12.060 52.030 12.320 52.350 ;
        RECT 12.520 52.030 12.780 52.350 ;
        RECT 12.120 49.970 12.260 52.030 ;
        RECT 12.060 49.650 12.320 49.970 ;
        RECT 12.580 49.370 12.720 52.030 ;
        RECT 12.120 49.230 12.720 49.370 ;
        RECT 10.220 44.550 10.480 44.870 ;
        RECT 11.600 44.550 11.860 44.870 ;
        RECT 10.280 43.170 10.420 44.550 ;
        RECT 10.220 42.850 10.480 43.170 ;
        RECT 8.840 41.830 9.100 42.150 ;
        RECT 8.900 40.450 9.040 41.830 ;
        RECT 8.840 40.130 9.100 40.450 ;
        RECT 8.380 38.770 8.640 39.090 ;
        RECT 8.440 37.730 8.580 38.770 ;
        RECT 8.380 37.410 8.640 37.730 ;
        RECT 8.900 34.330 9.040 40.130 ;
        RECT 9.760 36.960 10.020 37.050 ;
        RECT 9.360 36.820 10.020 36.960 ;
        RECT 8.840 34.010 9.100 34.330 ;
        RECT 8.840 28.290 9.100 28.550 ;
        RECT 8.440 28.230 9.100 28.290 ;
        RECT 8.440 28.150 9.040 28.230 ;
        RECT 7.920 27.550 8.180 27.870 ;
        RECT 7.460 24.830 7.720 25.150 ;
        RECT 7.520 22.770 7.660 24.830 ;
        RECT 7.460 22.450 7.720 22.770 ;
        RECT 7.000 19.390 7.260 19.710 ;
        RECT 0.100 6.470 0.360 6.790 ;
        RECT 7.060 6.530 7.200 19.390 ;
        RECT 7.460 16.670 7.720 16.990 ;
        RECT 7.520 11.890 7.660 16.670 ;
        RECT 7.460 11.570 7.720 11.890 ;
        RECT 7.980 6.790 8.120 27.550 ;
        RECT 8.440 15.630 8.580 28.150 ;
        RECT 9.360 26.170 9.500 36.820 ;
        RECT 9.760 36.730 10.020 36.820 ;
        RECT 10.220 34.010 10.480 34.330 ;
        RECT 9.760 27.550 10.020 27.870 ;
        RECT 9.820 26.170 9.960 27.550 ;
        RECT 9.300 25.850 9.560 26.170 ;
        RECT 9.760 25.850 10.020 26.170 ;
        RECT 9.360 17.670 9.500 25.850 ;
        RECT 10.280 25.830 10.420 34.010 ;
        RECT 11.140 28.910 11.400 29.230 ;
        RECT 11.200 28.550 11.340 28.910 ;
        RECT 11.660 28.550 11.800 44.550 ;
        RECT 12.120 36.565 12.260 49.230 ;
        RECT 12.520 47.610 12.780 47.930 ;
        RECT 12.580 40.450 12.720 47.610 ;
        RECT 13.040 45.210 13.180 53.195 ;
        RECT 12.980 44.890 13.240 45.210 ;
        RECT 12.980 43.870 13.240 44.190 ;
        RECT 13.040 42.830 13.180 43.870 ;
        RECT 12.980 42.510 13.240 42.830 ;
        RECT 12.520 40.130 12.780 40.450 ;
        RECT 12.580 37.390 12.720 40.130 ;
        RECT 12.520 37.070 12.780 37.390 ;
        RECT 12.980 36.730 13.240 37.050 ;
        RECT 12.050 36.195 12.330 36.565 ;
        RECT 11.140 28.230 11.400 28.550 ;
        RECT 11.600 28.230 11.860 28.550 ;
        RECT 10.680 27.890 10.940 28.210 ;
        RECT 10.220 25.510 10.480 25.830 ;
        RECT 10.280 23.110 10.420 25.510 ;
        RECT 10.740 24.130 10.880 27.890 ;
        RECT 11.660 26.850 11.800 28.230 ;
        RECT 11.600 26.530 11.860 26.850 ;
        RECT 10.680 23.810 10.940 24.130 ;
        RECT 10.220 22.790 10.480 23.110 ;
        RECT 9.300 17.350 9.560 17.670 ;
        RECT 9.760 17.350 10.020 17.670 ;
        RECT 9.820 15.970 9.960 17.350 ;
        RECT 9.760 15.650 10.020 15.970 ;
        RECT 8.380 15.310 8.640 15.630 ;
        RECT 10.280 15.290 10.420 22.790 ;
        RECT 10.740 20.730 10.880 23.810 ;
        RECT 10.680 20.410 10.940 20.730 ;
        RECT 10.680 19.390 10.940 19.710 ;
        RECT 11.600 19.390 11.860 19.710 ;
        RECT 10.220 14.970 10.480 15.290 ;
        RECT 10.740 13.870 10.880 19.390 ;
        RECT 11.140 14.970 11.400 15.290 ;
        RECT 10.280 13.730 10.880 13.870 ;
        RECT 10.280 9.930 10.420 13.730 ;
        RECT 11.200 12.230 11.340 14.970 ;
        RECT 11.140 11.910 11.400 12.230 ;
        RECT 9.820 9.790 10.420 9.930 ;
        RECT 0.160 4.000 0.300 6.470 ;
        RECT 3.320 6.130 3.580 6.450 ;
        RECT 6.600 6.390 7.200 6.530 ;
        RECT 7.920 6.470 8.180 6.790 ;
        RECT 3.380 4.000 3.520 6.130 ;
        RECT 6.600 4.000 6.740 6.390 ;
        RECT 9.820 4.000 9.960 9.790 ;
        RECT 11.660 6.450 11.800 19.390 ;
        RECT 12.120 18.010 12.260 36.195 ;
        RECT 13.040 29.230 13.180 36.730 ;
        RECT 13.500 36.030 13.640 53.990 ;
        RECT 13.900 53.730 14.160 54.050 ;
        RECT 13.960 53.565 14.100 53.730 ;
        RECT 13.890 53.370 14.170 53.565 ;
        RECT 15.340 53.370 15.480 55.090 ;
        RECT 16.720 54.130 16.860 74.900 ;
        RECT 17.120 74.130 17.380 74.450 ;
        RECT 17.180 69.350 17.320 74.130 ;
        RECT 17.640 74.110 17.780 82.970 ;
        RECT 19.940 80.910 20.080 88.070 ;
        RECT 23.100 84.670 23.360 84.990 ;
        RECT 21.070 84.135 22.610 84.505 ;
        RECT 20.340 82.290 20.600 82.610 ;
        RECT 20.400 81.250 20.540 82.290 ;
        RECT 20.340 80.930 20.600 81.250 ;
        RECT 19.880 80.590 20.140 80.910 ;
        RECT 19.940 77.510 20.080 80.590 ;
        RECT 23.160 80.230 23.300 84.670 ;
        RECT 23.620 83.370 23.760 104.050 ;
        RECT 28.620 103.710 28.880 104.030 ;
        RECT 24.370 103.175 25.910 103.545 ;
        RECT 28.680 102.670 28.820 103.710 ;
        RECT 28.620 102.350 28.880 102.670 ;
        RECT 24.370 97.735 25.910 98.105 ;
        RECT 26.320 95.550 26.580 95.870 ;
        RECT 24.370 92.295 25.910 92.665 ;
        RECT 26.380 92.130 26.520 95.550 ;
        RECT 30.060 94.850 30.200 112.470 ;
        RECT 30.000 94.530 30.260 94.850 ;
        RECT 27.700 93.170 27.960 93.490 ;
        RECT 27.760 92.130 27.900 93.170 ;
        RECT 26.320 91.810 26.580 92.130 ;
        RECT 27.700 91.810 27.960 92.130 ;
        RECT 26.380 88.050 26.520 91.810 ;
        RECT 30.060 91.790 30.200 94.530 ;
        RECT 30.000 91.470 30.260 91.790 ;
        RECT 30.520 91.110 30.660 120.800 ;
        RECT 31.380 120.710 31.640 121.030 ;
        RECT 31.840 120.710 32.100 121.030 ;
        RECT 31.440 113.890 31.580 120.710 ;
        RECT 32.820 120.690 32.960 125.470 ;
        RECT 32.760 120.370 33.020 120.690 ;
        RECT 33.280 117.970 33.420 126.070 ;
        RECT 34.140 123.430 34.400 123.750 ;
        RECT 34.200 123.070 34.340 123.430 ;
        RECT 34.140 122.750 34.400 123.070 ;
        RECT 33.680 121.450 33.940 121.710 ;
        RECT 34.660 121.450 34.800 126.830 ;
        RECT 35.120 122.050 35.260 128.190 ;
        RECT 37.880 126.470 38.020 128.190 ;
        RECT 35.520 126.150 35.780 126.470 ;
        RECT 37.820 126.150 38.080 126.470 ;
        RECT 35.060 121.730 35.320 122.050 ;
        RECT 33.680 121.390 34.800 121.450 ;
        RECT 33.740 121.310 34.800 121.390 ;
        RECT 33.220 117.650 33.480 117.970 ;
        RECT 33.280 116.010 33.420 117.650 ;
        RECT 32.820 115.870 33.420 116.010 ;
        RECT 31.380 113.570 31.640 113.890 ;
        RECT 32.820 113.210 32.960 115.870 ;
        RECT 33.220 115.270 33.480 115.590 ;
        RECT 32.760 112.890 33.020 113.210 ;
        RECT 32.760 109.150 33.020 109.470 ;
        RECT 32.820 106.750 32.960 109.150 ;
        RECT 33.280 107.770 33.420 115.270 ;
        RECT 34.140 112.890 34.400 113.210 ;
        RECT 33.680 112.550 33.940 112.870 ;
        RECT 33.740 109.470 33.880 112.550 ;
        RECT 33.680 109.150 33.940 109.470 ;
        RECT 33.740 108.110 33.880 109.150 ;
        RECT 33.680 107.790 33.940 108.110 ;
        RECT 33.220 107.450 33.480 107.770 ;
        RECT 32.300 106.430 32.560 106.750 ;
        RECT 32.760 106.430 33.020 106.750 ;
        RECT 31.840 105.070 32.100 105.390 ;
        RECT 32.360 105.300 32.500 106.430 ;
        RECT 32.760 105.300 33.020 105.390 ;
        RECT 32.360 105.160 33.020 105.300 ;
        RECT 32.760 105.070 33.020 105.160 ;
        RECT 34.200 105.130 34.340 112.890 ;
        RECT 35.060 112.210 35.320 112.530 ;
        RECT 35.120 110.150 35.260 112.210 ;
        RECT 35.060 109.830 35.320 110.150 ;
        RECT 35.120 108.450 35.260 109.830 ;
        RECT 35.060 108.130 35.320 108.450 ;
        RECT 34.600 107.450 34.860 107.770 ;
        RECT 34.660 105.730 34.800 107.450 ;
        RECT 34.600 105.410 34.860 105.730 ;
        RECT 30.920 104.050 31.180 104.370 ;
        RECT 30.980 103.010 31.120 104.050 ;
        RECT 31.900 103.010 32.040 105.070 ;
        RECT 33.740 104.990 34.340 105.130 ;
        RECT 30.920 102.690 31.180 103.010 ;
        RECT 31.840 102.690 32.100 103.010 ;
        RECT 31.840 102.010 32.100 102.330 ;
        RECT 31.900 100.290 32.040 102.010 ;
        RECT 31.840 99.970 32.100 100.290 ;
        RECT 33.220 98.950 33.480 99.270 ;
        RECT 33.280 97.570 33.420 98.950 ;
        RECT 33.740 98.590 33.880 104.990 ;
        RECT 34.140 104.390 34.400 104.710 ;
        RECT 34.200 103.010 34.340 104.390 ;
        RECT 34.140 102.690 34.400 103.010 ;
        RECT 34.200 99.270 34.340 102.690 ;
        RECT 35.060 102.010 35.320 102.330 ;
        RECT 35.120 99.690 35.260 102.010 ;
        RECT 35.580 100.290 35.720 126.150 ;
        RECT 37.360 125.810 37.620 126.130 ;
        RECT 37.420 124.090 37.560 125.810 ;
        RECT 37.880 124.430 38.020 126.150 ;
        RECT 38.280 125.470 38.540 125.790 ;
        RECT 37.820 124.110 38.080 124.430 ;
        RECT 38.340 124.090 38.480 125.470 ;
        RECT 37.360 123.770 37.620 124.090 ;
        RECT 38.280 123.770 38.540 124.090 ;
        RECT 36.440 123.490 36.700 123.750 ;
        RECT 36.440 123.430 37.560 123.490 ;
        RECT 37.820 123.430 38.080 123.750 ;
        RECT 38.740 123.430 39.000 123.750 ;
        RECT 36.500 123.350 37.560 123.430 ;
        RECT 35.980 122.750 36.240 123.070 ;
        RECT 36.900 122.750 37.160 123.070 ;
        RECT 36.040 120.690 36.180 122.750 ;
        RECT 36.960 121.030 37.100 122.750 ;
        RECT 37.420 122.050 37.560 123.350 ;
        RECT 37.880 123.070 38.020 123.430 ;
        RECT 37.820 122.750 38.080 123.070 ;
        RECT 37.360 121.730 37.620 122.050 ;
        RECT 36.900 120.710 37.160 121.030 ;
        RECT 35.980 120.370 36.240 120.690 ;
        RECT 36.440 112.890 36.700 113.210 ;
        RECT 35.980 111.870 36.240 112.190 ;
        RECT 36.040 110.150 36.180 111.870 ;
        RECT 36.500 110.150 36.640 112.890 ;
        RECT 36.960 110.490 37.100 120.710 ;
        RECT 38.800 120.350 38.940 123.430 ;
        RECT 39.260 122.050 39.400 129.210 ;
        RECT 39.720 126.810 39.860 129.210 ;
        RECT 41.100 128.850 41.240 129.550 ;
        RECT 42.020 129.530 42.160 133.630 ;
        RECT 41.960 129.210 42.220 129.530 ;
        RECT 42.480 129.190 42.620 134.650 ;
        RECT 45.240 129.870 45.380 134.910 ;
        RECT 45.640 133.970 45.900 134.290 ;
        RECT 45.700 131.910 45.840 133.970 ;
        RECT 45.640 131.590 45.900 131.910 ;
        RECT 45.180 129.550 45.440 129.870 ;
        RECT 42.420 128.870 42.680 129.190 ;
        RECT 41.040 128.530 41.300 128.850 ;
        RECT 39.660 126.490 39.920 126.810 ;
        RECT 41.100 123.070 41.240 128.530 ;
        RECT 41.500 126.150 41.760 126.470 ;
        RECT 41.040 122.750 41.300 123.070 ;
        RECT 39.200 121.730 39.460 122.050 ;
        RECT 40.580 121.730 40.840 122.050 ;
        RECT 38.740 120.030 39.000 120.350 ;
        RECT 38.800 119.330 38.940 120.030 ;
        RECT 38.740 119.010 39.000 119.330 ;
        RECT 40.640 118.650 40.780 121.730 ;
        RECT 41.560 121.370 41.700 126.150 ;
        RECT 41.960 125.470 42.220 125.790 ;
        RECT 41.500 121.050 41.760 121.370 ;
        RECT 41.040 120.710 41.300 121.030 ;
        RECT 41.100 119.330 41.240 120.710 ;
        RECT 41.040 119.010 41.300 119.330 ;
        RECT 42.020 118.650 42.160 125.470 ;
        RECT 45.700 123.410 45.840 131.590 ;
        RECT 45.640 123.090 45.900 123.410 ;
        RECT 43.340 120.030 43.600 120.350 ;
        RECT 40.580 118.330 40.840 118.650 ;
        RECT 41.960 118.330 42.220 118.650 ;
        RECT 37.360 117.310 37.620 117.630 ;
        RECT 37.420 113.210 37.560 117.310 ;
        RECT 42.420 115.270 42.680 115.590 ;
        RECT 42.480 113.210 42.620 115.270 ;
        RECT 37.360 112.890 37.620 113.210 ;
        RECT 42.420 112.890 42.680 113.210 ;
        RECT 41.960 112.550 42.220 112.870 ;
        RECT 37.360 112.210 37.620 112.530 ;
        RECT 36.900 110.170 37.160 110.490 ;
        RECT 35.980 109.830 36.240 110.150 ;
        RECT 36.440 109.830 36.700 110.150 ;
        RECT 36.500 107.770 36.640 109.830 ;
        RECT 36.900 109.490 37.160 109.810 ;
        RECT 36.440 107.450 36.700 107.770 ;
        RECT 36.960 107.170 37.100 109.490 ;
        RECT 37.420 107.770 37.560 112.210 ;
        RECT 37.820 111.870 38.080 112.190 ;
        RECT 37.360 107.450 37.620 107.770 ;
        RECT 37.880 107.430 38.020 111.870 ;
        RECT 42.020 110.830 42.160 112.550 ;
        RECT 41.960 110.510 42.220 110.830 ;
        RECT 38.280 109.490 38.540 109.810 ;
        RECT 38.340 108.450 38.480 109.490 ;
        RECT 38.280 108.130 38.540 108.450 ;
        RECT 36.500 107.030 37.100 107.170 ;
        RECT 37.820 107.110 38.080 107.430 ;
        RECT 36.500 104.710 36.640 107.030 ;
        RECT 36.900 106.430 37.160 106.750 ;
        RECT 36.440 104.390 36.700 104.710 ;
        RECT 35.980 101.670 36.240 101.990 ;
        RECT 35.520 99.970 35.780 100.290 ;
        RECT 35.120 99.550 35.720 99.690 ;
        RECT 34.140 98.950 34.400 99.270 ;
        RECT 35.060 98.950 35.320 99.270 ;
        RECT 33.680 98.270 33.940 98.590 ;
        RECT 33.220 97.250 33.480 97.570 ;
        RECT 34.140 91.130 34.400 91.450 ;
        RECT 30.460 90.790 30.720 91.110 ;
        RECT 26.320 87.730 26.580 88.050 ;
        RECT 24.370 86.855 25.910 87.225 ;
        RECT 23.620 83.230 24.220 83.370 ;
        RECT 23.560 80.250 23.820 80.570 ;
        RECT 23.100 79.910 23.360 80.230 ;
        RECT 21.070 78.695 22.610 79.065 ;
        RECT 19.880 77.190 20.140 77.510 ;
        RECT 17.580 73.790 17.840 74.110 ;
        RECT 17.640 72.070 17.780 73.790 ;
        RECT 17.580 71.750 17.840 72.070 ;
        RECT 18.040 71.070 18.300 71.390 ;
        RECT 17.120 69.030 17.380 69.350 ;
        RECT 17.120 66.990 17.380 67.310 ;
        RECT 17.180 64.590 17.320 66.990 ;
        RECT 17.120 64.270 17.380 64.590 ;
        RECT 18.100 63.910 18.240 71.070 ;
        RECT 19.940 70.370 20.080 77.190 ;
        RECT 21.260 76.510 21.520 76.830 ;
        RECT 21.320 75.130 21.460 76.510 ;
        RECT 21.260 74.810 21.520 75.130 ;
        RECT 21.070 73.255 22.610 73.625 ;
        RECT 20.340 71.410 20.600 71.730 ;
        RECT 20.400 70.370 20.540 71.410 ;
        RECT 19.880 70.050 20.140 70.370 ;
        RECT 20.340 70.050 20.600 70.370 ;
        RECT 18.960 69.710 19.220 70.030 ;
        RECT 19.020 66.970 19.160 69.710 ;
        RECT 18.960 66.650 19.220 66.970 ;
        RECT 19.940 64.930 20.080 70.050 ;
        RECT 21.070 67.815 22.610 68.185 ;
        RECT 21.260 65.970 21.520 66.290 ;
        RECT 21.320 64.930 21.460 65.970 ;
        RECT 19.880 64.610 20.140 64.930 ;
        RECT 21.260 64.610 21.520 64.930 ;
        RECT 23.620 64.330 23.760 80.250 ;
        RECT 23.160 64.190 23.760 64.330 ;
        RECT 18.040 63.590 18.300 63.910 ;
        RECT 20.340 63.590 20.600 63.910 ;
        RECT 20.400 62.210 20.540 63.590 ;
        RECT 21.070 62.375 22.610 62.745 ;
        RECT 20.340 62.170 20.600 62.210 ;
        RECT 19.480 62.030 20.600 62.170 ;
        RECT 19.480 61.530 19.620 62.030 ;
        RECT 20.340 61.890 20.600 62.030 ;
        RECT 19.420 61.210 19.680 61.530 ;
        RECT 22.180 60.870 22.440 61.190 ;
        RECT 19.420 60.530 19.680 60.850 ;
        RECT 18.040 60.190 18.300 60.510 ;
        RECT 18.100 58.810 18.240 60.190 ;
        RECT 18.960 59.170 19.220 59.490 ;
        RECT 18.040 58.490 18.300 58.810 ;
        RECT 18.500 56.450 18.760 56.770 ;
        RECT 17.120 56.110 17.380 56.430 ;
        RECT 16.260 53.990 16.860 54.130 ;
        RECT 13.885 53.195 14.170 53.370 ;
        RECT 13.885 53.050 14.145 53.195 ;
        RECT 15.280 53.050 15.540 53.370 ;
        RECT 14.820 52.370 15.080 52.690 ;
        RECT 14.880 51.330 15.020 52.370 ;
        RECT 14.820 51.010 15.080 51.330 ;
        RECT 15.340 48.370 15.480 53.050 ;
        RECT 16.260 52.350 16.400 53.990 ;
        RECT 17.180 53.370 17.320 56.110 ;
        RECT 18.560 53.370 18.700 56.450 ;
        RECT 19.020 55.750 19.160 59.170 ;
        RECT 18.960 55.430 19.220 55.750 ;
        RECT 16.660 53.050 16.920 53.370 ;
        RECT 17.120 53.050 17.380 53.370 ;
        RECT 17.580 53.050 17.840 53.370 ;
        RECT 18.500 53.050 18.760 53.370 ;
        RECT 16.200 52.030 16.460 52.350 ;
        RECT 13.960 48.230 15.480 48.370 ;
        RECT 13.960 45.550 14.100 48.230 ;
        RECT 13.900 45.230 14.160 45.550 ;
        RECT 14.820 44.550 15.080 44.870 ;
        RECT 13.900 43.870 14.160 44.190 ;
        RECT 13.960 41.325 14.100 43.870 ;
        RECT 14.880 42.830 15.020 44.550 ;
        RECT 15.740 42.850 16.000 43.170 ;
        RECT 14.820 42.510 15.080 42.830 ;
        RECT 13.890 40.955 14.170 41.325 ;
        RECT 15.280 41.150 15.540 41.470 ;
        RECT 14.820 38.430 15.080 38.750 ;
        RECT 14.880 37.925 15.020 38.430 ;
        RECT 14.810 37.555 15.090 37.925 ;
        RECT 14.360 37.070 14.620 37.390 ;
        RECT 13.440 35.710 13.700 36.030 ;
        RECT 13.900 34.690 14.160 35.010 ;
        RECT 13.440 33.330 13.700 33.650 ;
        RECT 13.500 32.290 13.640 33.330 ;
        RECT 13.440 31.970 13.700 32.290 ;
        RECT 12.980 28.910 13.240 29.230 ;
        RECT 13.960 28.290 14.100 34.690 ;
        RECT 14.420 33.310 14.560 37.070 ;
        RECT 14.820 36.960 15.080 37.050 ;
        RECT 15.340 36.960 15.480 41.150 ;
        RECT 15.800 39.430 15.940 42.850 ;
        RECT 15.740 39.110 16.000 39.430 ;
        RECT 14.820 36.820 15.480 36.960 ;
        RECT 14.820 36.730 15.080 36.820 ;
        RECT 14.820 35.710 15.080 36.030 ;
        RECT 14.360 32.990 14.620 33.310 ;
        RECT 14.420 28.890 14.560 32.990 ;
        RECT 14.880 31.610 15.020 35.710 ;
        RECT 15.340 35.010 15.480 36.820 ;
        RECT 15.280 34.690 15.540 35.010 ;
        RECT 14.820 31.290 15.080 31.610 ;
        RECT 15.280 31.290 15.540 31.610 ;
        RECT 15.340 29.230 15.480 31.290 ;
        RECT 15.280 28.910 15.540 29.230 ;
        RECT 14.360 28.570 14.620 28.890 ;
        RECT 13.960 28.150 14.560 28.290 ;
        RECT 13.900 27.550 14.160 27.870 ;
        RECT 13.960 26.510 14.100 27.550 ;
        RECT 13.900 26.190 14.160 26.510 ;
        RECT 14.420 22.430 14.560 28.150 ;
        RECT 14.820 24.830 15.080 25.150 ;
        RECT 14.880 23.110 15.020 24.830 ;
        RECT 14.820 22.790 15.080 23.110 ;
        RECT 14.360 22.110 14.620 22.430 ;
        RECT 14.420 21.070 14.560 22.110 ;
        RECT 14.360 20.750 14.620 21.070 ;
        RECT 13.900 20.410 14.160 20.730 ;
        RECT 12.060 17.690 12.320 18.010 ;
        RECT 12.520 16.670 12.780 16.990 ;
        RECT 12.980 16.670 13.240 16.990 ;
        RECT 12.580 8.570 12.720 16.670 ;
        RECT 13.040 15.290 13.180 16.670 ;
        RECT 13.960 15.970 14.100 20.410 ;
        RECT 14.880 17.670 15.020 22.790 ;
        RECT 15.340 18.350 15.480 28.910 ;
        RECT 16.200 28.230 16.460 28.550 ;
        RECT 16.260 26.850 16.400 28.230 ;
        RECT 16.200 26.530 16.460 26.850 ;
        RECT 16.720 20.810 16.860 53.050 ;
        RECT 17.120 52.370 17.380 52.690 ;
        RECT 17.180 39.850 17.320 52.370 ;
        RECT 17.640 50.310 17.780 53.050 ;
        RECT 17.580 49.990 17.840 50.310 ;
        RECT 17.640 48.370 17.780 49.990 ;
        RECT 17.640 48.230 18.240 48.370 ;
        RECT 17.580 45.230 17.840 45.550 ;
        RECT 17.640 42.150 17.780 45.230 ;
        RECT 17.580 41.830 17.840 42.150 ;
        RECT 18.100 40.110 18.240 48.230 ;
        RECT 18.560 44.870 18.700 53.050 ;
        RECT 19.020 48.270 19.160 55.430 ;
        RECT 19.480 53.710 19.620 60.530 ;
        RECT 20.340 60.190 20.600 60.510 ;
        RECT 21.720 60.190 21.980 60.510 ;
        RECT 19.880 57.470 20.140 57.790 ;
        RECT 19.940 55.750 20.080 57.470 ;
        RECT 20.400 56.770 20.540 60.190 ;
        RECT 21.780 59.490 21.920 60.190 ;
        RECT 21.720 59.170 21.980 59.490 ;
        RECT 22.240 57.700 22.380 60.870 ;
        RECT 23.160 58.040 23.300 64.190 ;
        RECT 23.560 63.590 23.820 63.910 ;
        RECT 23.620 61.190 23.760 63.590 ;
        RECT 24.080 62.170 24.220 83.230 ;
        RECT 24.370 81.415 25.910 81.785 ;
        RECT 26.380 78.610 26.520 87.730 ;
        RECT 29.080 85.350 29.340 85.670 ;
        RECT 26.780 81.950 27.040 82.270 ;
        RECT 26.840 80.570 26.980 81.950 ;
        RECT 26.780 80.250 27.040 80.570 ;
        RECT 26.840 79.550 26.980 80.250 ;
        RECT 26.780 79.230 27.040 79.550 ;
        RECT 26.380 78.470 26.980 78.610 ;
        RECT 24.370 75.975 25.910 76.345 ;
        RECT 24.370 70.535 25.910 70.905 ;
        RECT 26.320 65.630 26.580 65.950 ;
        RECT 24.370 65.095 25.910 65.465 ;
        RECT 26.380 62.210 26.520 65.630 ;
        RECT 24.080 62.030 26.060 62.170 ;
        RECT 23.560 60.870 23.820 61.190 ;
        RECT 23.620 59.490 23.760 60.870 ;
        RECT 25.920 60.760 26.060 62.030 ;
        RECT 26.320 61.890 26.580 62.210 ;
        RECT 26.840 62.170 26.980 78.470 ;
        RECT 27.700 77.870 27.960 78.190 ;
        RECT 27.760 76.830 27.900 77.870 ;
        RECT 27.700 76.510 27.960 76.830 ;
        RECT 27.760 75.810 27.900 76.510 ;
        RECT 27.700 75.490 27.960 75.810 ;
        RECT 26.840 62.030 27.440 62.170 ;
        RECT 26.780 61.550 27.040 61.870 ;
        RECT 25.920 60.620 26.520 60.760 ;
        RECT 24.020 60.190 24.280 60.510 ;
        RECT 23.560 59.170 23.820 59.490 ;
        RECT 23.160 57.900 23.760 58.040 ;
        RECT 22.240 57.560 23.300 57.700 ;
        RECT 21.070 56.935 22.610 57.305 ;
        RECT 20.340 56.450 20.600 56.770 ;
        RECT 23.160 56.430 23.300 57.560 ;
        RECT 23.100 56.110 23.360 56.430 ;
        RECT 19.880 55.430 20.140 55.750 ;
        RECT 21.260 55.090 21.520 55.410 ;
        RECT 20.800 54.750 21.060 55.070 ;
        RECT 19.420 53.390 19.680 53.710 ;
        RECT 20.860 53.370 21.000 54.750 ;
        RECT 21.320 53.710 21.460 55.090 ;
        RECT 23.620 55.070 23.760 57.900 ;
        RECT 24.080 56.090 24.220 60.190 ;
        RECT 24.370 59.655 25.910 60.025 ;
        RECT 24.480 58.830 24.740 59.150 ;
        RECT 24.020 55.770 24.280 56.090 ;
        RECT 24.540 55.750 24.680 58.830 ;
        RECT 25.400 58.490 25.660 58.810 ;
        RECT 25.460 56.770 25.600 58.490 ;
        RECT 25.400 56.450 25.660 56.770 ;
        RECT 24.480 55.430 24.740 55.750 ;
        RECT 23.560 54.750 23.820 55.070 ;
        RECT 24.370 54.215 25.910 54.585 ;
        RECT 21.260 53.390 21.520 53.710 ;
        RECT 20.800 53.280 21.060 53.370 ;
        RECT 20.400 53.140 21.060 53.280 ;
        RECT 20.400 48.610 20.540 53.140 ;
        RECT 20.800 53.050 21.060 53.140 ;
        RECT 23.100 53.050 23.360 53.370 ;
        RECT 21.070 51.495 22.610 51.865 ;
        RECT 20.800 49.650 21.060 49.970 ;
        RECT 20.340 48.290 20.600 48.610 ;
        RECT 18.960 47.950 19.220 48.270 ;
        RECT 19.020 45.290 19.160 47.950 ;
        RECT 20.860 47.590 21.000 49.650 ;
        RECT 23.160 47.590 23.300 53.050 ;
        RECT 23.560 52.030 23.820 52.350 ;
        RECT 23.620 47.590 23.760 52.030 ;
        RECT 24.480 50.050 24.740 50.310 ;
        RECT 24.080 49.990 24.740 50.050 ;
        RECT 24.080 49.910 24.680 49.990 ;
        RECT 20.800 47.270 21.060 47.590 ;
        RECT 23.100 47.270 23.360 47.590 ;
        RECT 23.560 47.270 23.820 47.590 ;
        RECT 20.340 46.590 20.600 46.910 ;
        RECT 19.020 45.150 19.620 45.290 ;
        RECT 18.500 44.550 18.760 44.870 ;
        RECT 17.180 39.710 17.780 39.850 ;
        RECT 18.040 39.790 18.300 40.110 ;
        RECT 17.120 39.110 17.380 39.430 ;
        RECT 17.180 24.130 17.320 39.110 ;
        RECT 17.640 28.970 17.780 39.710 ;
        RECT 18.560 36.710 18.700 44.550 ;
        RECT 19.480 42.490 19.620 45.150 ;
        RECT 20.400 44.870 20.540 46.590 ;
        RECT 21.070 46.055 22.610 46.425 ;
        RECT 22.180 45.570 22.440 45.890 ;
        RECT 21.720 44.890 21.980 45.210 ;
        RECT 20.340 44.550 20.600 44.870 ;
        RECT 21.780 42.490 21.920 44.890 ;
        RECT 22.240 42.490 22.380 45.570 ;
        RECT 23.160 45.210 23.300 47.270 ;
        RECT 23.100 44.890 23.360 45.210 ;
        RECT 23.560 44.550 23.820 44.870 ;
        RECT 19.420 42.170 19.680 42.490 ;
        RECT 21.720 42.170 21.980 42.490 ;
        RECT 22.180 42.170 22.440 42.490 ;
        RECT 18.960 41.830 19.220 42.150 ;
        RECT 18.500 36.390 18.760 36.710 ;
        RECT 19.020 33.990 19.160 41.830 ;
        RECT 19.480 40.360 19.620 42.170 ;
        RECT 23.100 41.830 23.360 42.150 ;
        RECT 21.070 40.615 22.610 40.985 ;
        RECT 23.160 40.450 23.300 41.830 ;
        RECT 19.480 40.220 21.000 40.360 ;
        RECT 19.880 39.110 20.140 39.430 ;
        RECT 18.960 33.670 19.220 33.990 ;
        RECT 18.960 32.990 19.220 33.310 ;
        RECT 19.020 31.950 19.160 32.990 ;
        RECT 18.960 31.630 19.220 31.950 ;
        RECT 19.420 30.270 19.680 30.590 ;
        RECT 17.640 28.830 18.240 28.970 ;
        RECT 17.580 28.230 17.840 28.550 ;
        RECT 17.640 26.170 17.780 28.230 ;
        RECT 17.580 25.850 17.840 26.170 ;
        RECT 17.120 23.810 17.380 24.130 ;
        RECT 17.580 22.790 17.840 23.110 ;
        RECT 17.640 20.925 17.780 22.790 ;
        RECT 16.720 20.670 17.320 20.810 ;
        RECT 15.740 19.730 16.000 20.050 ;
        RECT 16.660 19.730 16.920 20.050 ;
        RECT 15.280 18.030 15.540 18.350 ;
        RECT 14.820 17.350 15.080 17.670 ;
        RECT 13.900 15.650 14.160 15.970 ;
        RECT 12.980 14.970 13.240 15.290 ;
        RECT 13.960 13.250 14.100 15.650 ;
        RECT 15.800 15.290 15.940 19.730 ;
        RECT 16.200 17.350 16.460 17.670 ;
        RECT 15.740 14.970 16.000 15.290 ;
        RECT 16.260 13.250 16.400 17.350 ;
        RECT 13.900 12.930 14.160 13.250 ;
        RECT 16.200 12.930 16.460 13.250 ;
        RECT 16.720 9.930 16.860 19.730 ;
        RECT 17.180 19.710 17.320 20.670 ;
        RECT 17.570 20.555 17.850 20.925 ;
        RECT 17.580 20.410 17.840 20.555 ;
        RECT 17.120 19.390 17.380 19.710 ;
        RECT 18.100 18.690 18.240 28.830 ;
        RECT 19.480 28.550 19.620 30.270 ;
        RECT 19.420 28.230 19.680 28.550 ;
        RECT 19.480 26.850 19.620 28.230 ;
        RECT 19.420 26.530 19.680 26.850 ;
        RECT 18.500 20.410 18.760 20.730 ;
        RECT 18.040 18.370 18.300 18.690 ;
        RECT 18.560 14.270 18.700 20.410 ;
        RECT 19.480 17.670 19.620 26.530 ;
        RECT 19.940 24.130 20.080 39.110 ;
        RECT 20.860 37.390 21.000 40.220 ;
        RECT 23.100 40.130 23.360 40.450 ;
        RECT 22.640 39.450 22.900 39.770 ;
        RECT 21.260 39.110 21.520 39.430 ;
        RECT 20.800 37.070 21.060 37.390 ;
        RECT 21.320 37.050 21.460 39.110 ;
        RECT 22.700 37.390 22.840 39.450 ;
        RECT 23.100 38.770 23.360 39.090 ;
        RECT 22.640 37.070 22.900 37.390 ;
        RECT 23.160 37.050 23.300 38.770 ;
        RECT 21.260 36.730 21.520 37.050 ;
        RECT 23.100 36.730 23.360 37.050 ;
        RECT 23.100 35.710 23.360 36.030 ;
        RECT 21.070 35.175 22.610 35.545 ;
        RECT 22.180 33.670 22.440 33.990 ;
        RECT 22.640 33.670 22.900 33.990 ;
        RECT 20.800 33.330 21.060 33.650 ;
        RECT 20.860 31.610 21.000 33.330 ;
        RECT 22.240 31.950 22.380 33.670 ;
        RECT 22.700 32.290 22.840 33.670 ;
        RECT 23.160 33.310 23.300 35.710 ;
        RECT 23.620 33.900 23.760 44.550 ;
        RECT 24.080 37.730 24.220 49.910 ;
        RECT 24.370 48.775 25.910 49.145 ;
        RECT 25.400 48.290 25.660 48.610 ;
        RECT 25.860 48.290 26.120 48.610 ;
        RECT 25.460 44.530 25.600 48.290 ;
        RECT 25.920 44.725 26.060 48.290 ;
        RECT 25.400 44.210 25.660 44.530 ;
        RECT 25.850 44.355 26.130 44.725 ;
        RECT 24.370 43.335 25.910 43.705 ;
        RECT 26.380 39.430 26.520 60.620 ;
        RECT 26.840 52.260 26.980 61.550 ;
        RECT 27.300 52.770 27.440 62.030 ;
        RECT 27.760 59.150 27.900 75.490 ;
        RECT 28.620 65.630 28.880 65.950 ;
        RECT 28.680 60.850 28.820 65.630 ;
        RECT 28.620 60.530 28.880 60.850 ;
        RECT 27.700 59.060 27.960 59.150 ;
        RECT 27.700 58.920 28.360 59.060 ;
        RECT 27.700 58.830 27.960 58.920 ;
        RECT 27.700 57.470 27.960 57.790 ;
        RECT 27.760 53.710 27.900 57.470 ;
        RECT 27.700 53.390 27.960 53.710 ;
        RECT 27.300 52.630 27.900 52.770 ;
        RECT 27.240 52.260 27.500 52.350 ;
        RECT 26.840 52.120 27.500 52.260 ;
        RECT 26.840 49.970 26.980 52.120 ;
        RECT 27.240 52.030 27.500 52.120 ;
        RECT 27.760 51.410 27.900 52.630 ;
        RECT 27.300 51.270 27.900 51.410 ;
        RECT 26.780 49.650 27.040 49.970 ;
        RECT 26.840 47.930 26.980 49.650 ;
        RECT 26.780 47.610 27.040 47.930 ;
        RECT 27.300 44.870 27.440 51.270 ;
        RECT 28.220 48.610 28.360 58.920 ;
        RECT 29.140 54.050 29.280 85.350 ;
        RECT 30.520 77.850 30.660 90.790 ;
        RECT 34.200 88.730 34.340 91.130 ;
        RECT 30.920 88.410 31.180 88.730 ;
        RECT 34.140 88.410 34.400 88.730 ;
        RECT 30.980 86.690 31.120 88.410 ;
        RECT 33.680 87.390 33.940 87.710 ;
        RECT 33.740 86.690 33.880 87.390 ;
        RECT 35.120 86.690 35.260 98.950 ;
        RECT 35.580 96.670 35.720 99.550 ;
        RECT 36.040 97.230 36.180 101.670 ;
        RECT 35.980 96.910 36.240 97.230 ;
        RECT 36.500 96.670 36.640 104.390 ;
        RECT 36.960 99.610 37.100 106.430 ;
        RECT 37.360 104.390 37.620 104.710 ;
        RECT 37.820 104.390 38.080 104.710 ;
        RECT 37.420 103.010 37.560 104.390 ;
        RECT 37.360 102.690 37.620 103.010 ;
        RECT 36.900 99.290 37.160 99.610 ;
        RECT 37.420 99.270 37.560 102.690 ;
        RECT 37.880 99.270 38.020 104.390 ;
        RECT 39.200 104.050 39.460 104.370 ;
        RECT 41.960 104.050 42.220 104.370 ;
        RECT 38.740 102.010 39.000 102.330 ;
        RECT 38.800 100.290 38.940 102.010 ;
        RECT 38.740 99.970 39.000 100.290 ;
        RECT 37.360 98.950 37.620 99.270 ;
        RECT 37.820 98.950 38.080 99.270 ;
        RECT 37.420 96.670 37.560 98.950 ;
        RECT 35.580 96.530 36.640 96.670 ;
        RECT 36.500 91.790 36.640 96.530 ;
        RECT 36.960 96.530 37.560 96.670 ;
        RECT 38.280 96.570 38.540 96.890 ;
        RECT 36.440 91.470 36.700 91.790 ;
        RECT 30.920 86.370 31.180 86.690 ;
        RECT 33.680 86.370 33.940 86.690 ;
        RECT 35.060 86.370 35.320 86.690 ;
        RECT 36.500 86.010 36.640 91.470 ;
        RECT 36.960 90.340 37.100 96.530 ;
        RECT 37.360 93.850 37.620 94.170 ;
        RECT 37.420 92.130 37.560 93.850 ;
        RECT 37.360 91.810 37.620 92.130 ;
        RECT 37.360 90.340 37.620 90.430 ;
        RECT 36.960 90.200 37.620 90.340 ;
        RECT 37.360 90.110 37.620 90.200 ;
        RECT 36.440 85.690 36.700 86.010 ;
        RECT 36.500 83.630 36.640 85.690 ;
        RECT 37.420 83.970 37.560 90.110 ;
        RECT 37.360 83.650 37.620 83.970 ;
        RECT 36.440 83.310 36.700 83.630 ;
        RECT 37.820 82.290 38.080 82.610 ;
        RECT 32.300 81.950 32.560 82.270 ;
        RECT 32.360 77.850 32.500 81.950 ;
        RECT 37.880 81.250 38.020 82.290 ;
        RECT 37.820 80.930 38.080 81.250 ;
        RECT 34.600 80.590 34.860 80.910 ;
        RECT 33.220 80.250 33.480 80.570 ;
        RECT 33.280 78.530 33.420 80.250 ;
        RECT 33.220 78.210 33.480 78.530 ;
        RECT 30.460 77.530 30.720 77.850 ;
        RECT 32.300 77.530 32.560 77.850 ;
        RECT 34.140 77.190 34.400 77.510 ;
        RECT 33.220 74.810 33.480 75.130 ;
        RECT 33.280 73.090 33.420 74.810 ;
        RECT 33.220 72.770 33.480 73.090 ;
        RECT 34.200 72.750 34.340 77.190 ;
        RECT 34.660 75.470 34.800 80.590 ;
        RECT 38.340 77.850 38.480 96.570 ;
        RECT 39.260 96.210 39.400 104.050 ;
        RECT 42.020 101.310 42.160 104.050 ;
        RECT 42.880 103.710 43.140 104.030 ;
        RECT 41.960 100.990 42.220 101.310 ;
        RECT 42.940 100.290 43.080 103.710 ;
        RECT 42.880 99.970 43.140 100.290 ;
        RECT 41.040 96.910 41.300 97.230 ;
        RECT 40.580 96.570 40.840 96.890 ;
        RECT 39.200 95.890 39.460 96.210 ;
        RECT 39.260 88.050 39.400 95.890 ;
        RECT 40.640 94.850 40.780 96.570 ;
        RECT 40.580 94.530 40.840 94.850 ;
        RECT 40.580 90.110 40.840 90.430 ;
        RECT 40.640 88.390 40.780 90.110 ;
        RECT 40.580 88.070 40.840 88.390 ;
        RECT 39.200 87.730 39.460 88.050 ;
        RECT 38.740 81.950 39.000 82.270 ;
        RECT 38.800 80.230 38.940 81.950 ;
        RECT 39.260 80.570 39.400 87.730 ;
        RECT 40.120 85.690 40.380 86.010 ;
        RECT 40.180 81.250 40.320 85.690 ;
        RECT 40.580 83.310 40.840 83.630 ;
        RECT 40.120 80.930 40.380 81.250 ;
        RECT 39.200 80.250 39.460 80.570 ;
        RECT 38.740 79.910 39.000 80.230 ;
        RECT 40.640 77.850 40.780 83.310 ;
        RECT 41.100 80.910 41.240 96.910 ;
        RECT 42.880 94.190 43.140 94.510 ;
        RECT 41.500 89.090 41.760 89.410 ;
        RECT 41.560 86.690 41.700 89.090 ;
        RECT 41.960 87.390 42.220 87.710 ;
        RECT 41.500 86.370 41.760 86.690 ;
        RECT 42.020 86.010 42.160 87.390 ;
        RECT 41.960 85.690 42.220 86.010 ;
        RECT 41.500 85.010 41.760 85.330 ;
        RECT 41.560 83.630 41.700 85.010 ;
        RECT 42.420 84.670 42.680 84.990 ;
        RECT 42.480 83.970 42.620 84.670 ;
        RECT 42.420 83.650 42.680 83.970 ;
        RECT 41.500 83.310 41.760 83.630 ;
        RECT 42.480 82.610 42.620 83.650 ;
        RECT 42.420 82.290 42.680 82.610 ;
        RECT 41.500 81.950 41.760 82.270 ;
        RECT 41.560 80.910 41.700 81.950 ;
        RECT 41.040 80.590 41.300 80.910 ;
        RECT 41.500 80.590 41.760 80.910 ;
        RECT 41.100 80.230 41.240 80.590 ;
        RECT 41.040 79.910 41.300 80.230 ;
        RECT 41.500 79.230 41.760 79.550 ;
        RECT 41.560 78.530 41.700 79.230 ;
        RECT 41.500 78.210 41.760 78.530 ;
        RECT 38.280 77.530 38.540 77.850 ;
        RECT 40.580 77.530 40.840 77.850 ;
        RECT 35.060 76.510 35.320 76.830 ;
        RECT 36.900 76.510 37.160 76.830 ;
        RECT 34.600 75.150 34.860 75.470 ;
        RECT 34.140 72.430 34.400 72.750 ;
        RECT 34.660 72.070 34.800 75.150 ;
        RECT 34.600 71.750 34.860 72.070 ;
        RECT 30.000 71.410 30.260 71.730 ;
        RECT 30.060 69.350 30.200 71.410 ;
        RECT 34.660 70.030 34.800 71.750 ;
        RECT 31.840 69.710 32.100 70.030 ;
        RECT 33.220 69.710 33.480 70.030 ;
        RECT 34.600 69.710 34.860 70.030 ;
        RECT 30.000 69.030 30.260 69.350 ;
        RECT 29.080 53.730 29.340 54.050 ;
        RECT 28.160 48.290 28.420 48.610 ;
        RECT 29.540 45.800 29.800 45.890 ;
        RECT 30.060 45.800 30.200 69.030 ;
        RECT 30.460 65.630 30.720 65.950 ;
        RECT 30.920 65.630 31.180 65.950 ;
        RECT 30.520 64.930 30.660 65.630 ;
        RECT 30.460 64.610 30.720 64.930 ;
        RECT 30.980 62.170 31.120 65.630 ;
        RECT 29.540 45.660 30.200 45.800 ;
        RECT 29.540 45.570 29.800 45.660 ;
        RECT 27.240 44.550 27.500 44.870 ;
        RECT 26.780 44.210 27.040 44.530 ;
        RECT 26.840 40.360 26.980 44.210 ;
        RECT 26.840 40.220 27.440 40.360 ;
        RECT 26.780 39.450 27.040 39.770 ;
        RECT 26.320 39.110 26.580 39.430 ;
        RECT 24.370 37.895 25.910 38.265 ;
        RECT 24.020 37.410 24.280 37.730 ;
        RECT 26.840 37.050 26.980 39.450 ;
        RECT 27.300 37.130 27.440 40.220 ;
        RECT 30.060 39.430 30.200 45.660 ;
        RECT 30.520 62.030 31.120 62.170 ;
        RECT 30.520 40.110 30.660 62.030 ;
        RECT 31.380 55.090 31.640 55.410 ;
        RECT 31.440 54.050 31.580 55.090 ;
        RECT 31.380 53.730 31.640 54.050 ;
        RECT 31.900 48.270 32.040 69.710 ;
        RECT 33.280 66.630 33.420 69.710 ;
        RECT 33.220 66.310 33.480 66.630 ;
        RECT 32.760 61.890 33.020 62.210 ;
        RECT 32.820 56.430 32.960 61.890 ;
        RECT 33.280 61.190 33.420 66.310 ;
        RECT 33.220 60.870 33.480 61.190 ;
        RECT 33.280 58.810 33.420 60.870 ;
        RECT 33.220 58.490 33.480 58.810 ;
        RECT 32.760 56.110 33.020 56.430 ;
        RECT 33.280 55.750 33.420 58.490 ;
        RECT 35.120 56.770 35.260 76.510 ;
        RECT 36.960 72.410 37.100 76.510 ;
        RECT 38.340 75.810 38.480 77.530 ;
        RECT 40.640 75.810 40.780 77.530 ;
        RECT 38.280 75.490 38.540 75.810 ;
        RECT 40.580 75.490 40.840 75.810 ;
        RECT 36.900 72.090 37.160 72.410 ;
        RECT 39.660 71.750 39.920 72.070 ;
        RECT 35.520 64.610 35.780 64.930 ;
        RECT 35.580 64.250 35.720 64.610 ;
        RECT 35.520 63.930 35.780 64.250 ;
        RECT 35.980 63.930 36.240 64.250 ;
        RECT 36.900 63.930 37.160 64.250 ;
        RECT 35.580 62.210 35.720 63.930 ;
        RECT 36.040 63.085 36.180 63.930 ;
        RECT 35.970 62.715 36.250 63.085 ;
        RECT 35.520 61.890 35.780 62.210 ;
        RECT 36.960 62.170 37.100 63.930 ;
        RECT 39.720 63.230 39.860 71.750 ;
        RECT 40.580 71.070 40.840 71.390 ;
        RECT 40.640 64.930 40.780 71.070 ;
        RECT 41.040 66.310 41.300 66.630 ;
        RECT 40.580 64.610 40.840 64.930 ;
        RECT 40.580 63.590 40.840 63.910 ;
        RECT 39.660 62.910 39.920 63.230 ;
        RECT 36.960 62.030 38.940 62.170 ;
        RECT 36.900 60.190 37.160 60.510 ;
        RECT 36.960 59.150 37.100 60.190 ;
        RECT 36.900 58.830 37.160 59.150 ;
        RECT 35.060 56.450 35.320 56.770 ;
        RECT 33.220 55.430 33.480 55.750 ;
        RECT 36.440 54.750 36.700 55.070 ;
        RECT 36.500 53.370 36.640 54.750 ;
        RECT 36.440 53.050 36.700 53.370 ;
        RECT 34.140 52.710 34.400 53.030 ;
        RECT 34.200 51.330 34.340 52.710 ;
        RECT 34.140 51.010 34.400 51.330 ;
        RECT 31.840 47.950 32.100 48.270 ;
        RECT 30.920 42.850 31.180 43.170 ;
        RECT 30.980 41.810 31.120 42.850 ;
        RECT 31.900 42.830 32.040 47.950 ;
        RECT 33.220 47.610 33.480 47.930 ;
        RECT 33.680 47.610 33.940 47.930 ;
        RECT 34.600 47.840 34.860 47.930 ;
        RECT 34.600 47.700 35.260 47.840 ;
        RECT 34.600 47.610 34.860 47.700 ;
        RECT 32.300 44.210 32.560 44.530 ;
        RECT 31.840 42.510 32.100 42.830 ;
        RECT 30.920 41.490 31.180 41.810 ;
        RECT 30.460 39.790 30.720 40.110 ;
        RECT 30.000 39.340 30.260 39.430 ;
        RECT 29.600 39.200 30.260 39.340 ;
        RECT 26.780 36.730 27.040 37.050 ;
        RECT 27.300 36.990 27.900 37.130 ;
        RECT 26.840 34.410 26.980 36.730 ;
        RECT 27.240 36.390 27.500 36.710 ;
        RECT 26.380 34.270 26.980 34.410 ;
        RECT 26.380 33.990 26.520 34.270 ;
        RECT 27.300 33.990 27.440 36.390 ;
        RECT 24.020 33.900 24.280 33.990 ;
        RECT 23.620 33.760 24.280 33.900 ;
        RECT 24.020 33.670 24.280 33.760 ;
        RECT 26.320 33.670 26.580 33.990 ;
        RECT 26.780 33.670 27.040 33.990 ;
        RECT 27.240 33.670 27.500 33.990 ;
        RECT 23.100 32.990 23.360 33.310 ;
        RECT 23.560 32.990 23.820 33.310 ;
        RECT 22.640 31.970 22.900 32.290 ;
        RECT 23.100 31.970 23.360 32.290 ;
        RECT 22.180 31.690 22.440 31.950 ;
        RECT 23.160 31.690 23.300 31.970 ;
        RECT 22.180 31.630 23.300 31.690 ;
        RECT 20.800 31.290 21.060 31.610 ;
        RECT 22.240 31.550 23.300 31.630 ;
        RECT 23.620 31.610 23.760 32.990 ;
        RECT 24.370 32.455 25.910 32.825 ;
        RECT 26.320 31.970 26.580 32.290 ;
        RECT 23.560 31.290 23.820 31.610 ;
        RECT 20.860 31.010 21.000 31.290 ;
        RECT 20.400 30.870 21.000 31.010 ;
        RECT 20.400 26.170 20.540 30.870 ;
        RECT 24.020 30.270 24.280 30.590 ;
        RECT 21.070 29.735 22.610 30.105 ;
        RECT 20.340 25.850 20.600 26.170 ;
        RECT 23.560 25.850 23.820 26.170 ;
        RECT 19.880 23.810 20.140 24.130 ;
        RECT 20.400 23.530 20.540 25.850 ;
        RECT 23.100 24.830 23.360 25.150 ;
        RECT 21.070 24.295 22.610 24.665 ;
        RECT 19.940 23.390 20.540 23.530 ;
        RECT 19.940 21.070 20.080 23.390 ;
        RECT 23.160 23.110 23.300 24.830 ;
        RECT 20.340 22.790 20.600 23.110 ;
        RECT 23.100 22.790 23.360 23.110 ;
        RECT 19.880 20.750 20.140 21.070 ;
        RECT 19.420 17.350 19.680 17.670 ;
        RECT 19.420 14.970 19.680 15.290 ;
        RECT 19.480 14.690 19.620 14.970 ;
        RECT 19.940 14.690 20.080 20.750 ;
        RECT 20.400 15.290 20.540 22.790 ;
        RECT 23.100 22.110 23.360 22.430 ;
        RECT 23.160 21.070 23.300 22.110 ;
        RECT 23.620 21.410 23.760 25.850 ;
        RECT 23.560 21.090 23.820 21.410 ;
        RECT 23.100 20.750 23.360 21.070 ;
        RECT 24.080 20.810 24.220 30.270 ;
        RECT 24.370 27.015 25.910 27.385 ;
        RECT 25.860 26.080 26.120 26.170 ;
        RECT 26.380 26.080 26.520 31.970 ;
        RECT 26.840 28.890 26.980 33.670 ;
        RECT 27.240 31.630 27.500 31.950 ;
        RECT 26.780 28.570 27.040 28.890 ;
        RECT 26.840 26.170 26.980 28.570 ;
        RECT 25.860 25.940 26.520 26.080 ;
        RECT 25.860 25.850 26.120 25.940 ;
        RECT 24.370 21.575 25.910 21.945 ;
        RECT 21.070 18.855 22.610 19.225 ;
        RECT 21.250 17.835 21.530 18.205 ;
        RECT 21.320 17.670 21.460 17.835 ;
        RECT 21.260 17.350 21.520 17.670 ;
        RECT 20.800 16.670 21.060 16.990 ;
        RECT 22.640 16.670 22.900 16.990 ;
        RECT 20.860 15.970 21.000 16.670 ;
        RECT 20.800 15.650 21.060 15.970 ;
        RECT 22.700 15.630 22.840 16.670 ;
        RECT 22.640 15.310 22.900 15.630 ;
        RECT 20.340 14.970 20.600 15.290 ;
        RECT 19.480 14.610 20.540 14.690 ;
        RECT 19.480 14.550 20.600 14.610 ;
        RECT 18.500 13.950 18.760 14.270 ;
        RECT 18.560 12.230 18.700 13.950 ;
        RECT 19.480 13.870 19.620 14.550 ;
        RECT 20.340 14.290 20.600 14.550 ;
        RECT 19.020 13.730 19.620 13.870 ;
        RECT 18.500 11.910 18.760 12.230 ;
        RECT 19.020 11.890 19.160 13.730 ;
        RECT 21.070 13.415 22.610 13.785 ;
        RECT 23.160 12.230 23.300 20.750 ;
        RECT 23.620 20.670 24.220 20.810 ;
        RECT 23.620 12.230 23.760 20.670 ;
        RECT 24.020 17.350 24.280 17.670 ;
        RECT 24.940 17.350 25.200 17.670 ;
        RECT 24.080 15.970 24.220 17.350 ;
        RECT 25.000 16.990 25.140 17.350 ;
        RECT 25.860 17.240 26.120 17.330 ;
        RECT 26.380 17.240 26.520 25.940 ;
        RECT 26.780 25.850 27.040 26.170 ;
        RECT 27.300 24.890 27.440 31.630 ;
        RECT 27.760 26.170 27.900 36.990 ;
        RECT 27.700 26.080 27.960 26.170 ;
        RECT 27.700 25.940 28.360 26.080 ;
        RECT 27.700 25.850 27.960 25.940 ;
        RECT 27.700 25.170 27.960 25.490 ;
        RECT 27.760 24.890 27.900 25.170 ;
        RECT 27.300 24.750 27.900 24.890 ;
        RECT 27.300 22.850 27.440 24.750 ;
        RECT 27.700 22.850 27.960 23.110 ;
        RECT 27.300 22.790 27.960 22.850 ;
        RECT 27.300 22.710 27.900 22.790 ;
        RECT 27.300 17.670 27.440 22.710 ;
        RECT 28.220 22.430 28.360 25.940 ;
        RECT 29.080 25.850 29.340 26.170 ;
        RECT 28.620 24.830 28.880 25.150 ;
        RECT 28.680 22.770 28.820 24.830 ;
        RECT 28.620 22.450 28.880 22.770 ;
        RECT 28.160 22.110 28.420 22.430 ;
        RECT 27.240 17.350 27.500 17.670 ;
        RECT 25.860 17.100 26.520 17.240 ;
        RECT 25.860 17.010 26.120 17.100 ;
        RECT 24.940 16.670 25.200 16.990 ;
        RECT 24.370 16.135 25.910 16.505 ;
        RECT 24.020 15.650 24.280 15.970 ;
        RECT 27.240 15.310 27.500 15.630 ;
        RECT 27.300 12.230 27.440 15.310 ;
        RECT 29.140 14.950 29.280 25.850 ;
        RECT 29.600 25.490 29.740 39.200 ;
        RECT 30.000 39.110 30.260 39.200 ;
        RECT 30.980 37.390 31.120 41.490 ;
        RECT 32.360 40.450 32.500 44.210 ;
        RECT 33.280 44.190 33.420 47.610 ;
        RECT 33.740 47.250 33.880 47.610 ;
        RECT 33.680 46.930 33.940 47.250 ;
        RECT 34.600 46.930 34.860 47.250 ;
        RECT 33.740 45.890 33.880 46.930 ;
        RECT 33.680 45.570 33.940 45.890 ;
        RECT 34.660 44.870 34.800 46.930 ;
        RECT 34.600 44.550 34.860 44.870 ;
        RECT 33.220 43.870 33.480 44.190 ;
        RECT 33.680 42.510 33.940 42.830 ;
        RECT 32.300 40.130 32.560 40.450 ;
        RECT 33.740 39.430 33.880 42.510 ;
        RECT 34.660 42.490 34.800 44.550 ;
        RECT 34.600 42.170 34.860 42.490 ;
        RECT 33.680 39.110 33.940 39.430 ;
        RECT 30.920 37.070 31.180 37.390 ;
        RECT 32.760 33.670 33.020 33.990 ;
        RECT 30.000 32.990 30.260 33.310 ;
        RECT 30.060 31.950 30.200 32.990 ;
        RECT 30.000 31.630 30.260 31.950 ;
        RECT 29.540 25.170 29.800 25.490 ;
        RECT 29.600 22.770 29.740 25.170 ;
        RECT 29.540 22.450 29.800 22.770 ;
        RECT 29.080 14.630 29.340 14.950 ;
        RECT 29.080 12.590 29.340 12.910 ;
        RECT 23.100 11.910 23.360 12.230 ;
        RECT 23.560 11.910 23.820 12.230 ;
        RECT 27.240 11.910 27.500 12.230 ;
        RECT 18.960 11.570 19.220 11.890 ;
        RECT 19.420 11.230 19.680 11.550 ;
        RECT 22.640 11.230 22.900 11.550 ;
        RECT 25.860 11.460 26.120 11.550 ;
        RECT 25.860 11.320 26.520 11.460 ;
        RECT 25.860 11.230 26.120 11.320 ;
        RECT 16.260 9.790 16.860 9.930 ;
        RECT 12.580 8.430 13.180 8.570 ;
        RECT 11.600 6.130 11.860 6.450 ;
        RECT 13.040 4.000 13.180 8.430 ;
        RECT 16.260 4.000 16.400 9.790 ;
        RECT 19.480 4.000 19.620 11.230 ;
        RECT 22.700 4.000 22.840 11.230 ;
        RECT 24.370 10.695 25.910 11.065 ;
        RECT 26.380 5.850 26.520 11.320 ;
        RECT 25.920 5.710 26.520 5.850 ;
        RECT 25.920 4.000 26.060 5.710 ;
        RECT 29.140 4.000 29.280 12.590 ;
        RECT 30.060 12.230 30.200 31.630 ;
        RECT 32.820 31.610 32.960 33.670 ;
        RECT 34.600 33.330 34.860 33.650 ;
        RECT 32.760 31.290 33.020 31.610 ;
        RECT 32.820 21.070 32.960 31.290 ;
        RECT 34.140 26.190 34.400 26.510 ;
        RECT 34.200 22.770 34.340 26.190 ;
        RECT 34.660 25.830 34.800 33.330 ;
        RECT 35.120 32.290 35.260 47.700 ;
        RECT 36.440 47.610 36.700 47.930 ;
        RECT 37.360 47.610 37.620 47.930 ;
        RECT 36.500 45.550 36.640 47.610 ;
        RECT 37.420 45.890 37.560 47.610 ;
        RECT 37.360 45.570 37.620 45.890 ;
        RECT 36.440 45.230 36.700 45.550 ;
        RECT 37.360 43.870 37.620 44.190 ;
        RECT 37.420 42.490 37.560 43.870 ;
        RECT 37.360 42.170 37.620 42.490 ;
        RECT 36.900 41.830 37.160 42.150 ;
        RECT 36.960 39.430 37.100 41.830 ;
        RECT 36.900 39.110 37.160 39.430 ;
        RECT 35.980 36.960 36.240 37.050 ;
        RECT 35.980 36.820 36.640 36.960 ;
        RECT 35.980 36.730 36.240 36.820 ;
        RECT 35.060 31.970 35.320 32.290 ;
        RECT 35.060 31.290 35.320 31.610 ;
        RECT 35.120 29.230 35.260 31.290 ;
        RECT 35.520 30.950 35.780 31.270 ;
        RECT 35.060 28.910 35.320 29.230 ;
        RECT 35.060 28.230 35.320 28.550 ;
        RECT 35.120 26.170 35.260 28.230 ;
        RECT 35.060 25.850 35.320 26.170 ;
        RECT 34.600 25.510 34.860 25.830 ;
        RECT 35.120 24.130 35.260 25.850 ;
        RECT 35.060 23.810 35.320 24.130 ;
        RECT 34.140 22.450 34.400 22.770 ;
        RECT 32.760 20.925 33.020 21.070 ;
        RECT 32.750 20.810 33.030 20.925 ;
        RECT 32.750 20.670 33.420 20.810 ;
        RECT 32.750 20.555 33.030 20.670 ;
        RECT 32.760 14.290 33.020 14.610 ;
        RECT 30.920 13.950 31.180 14.270 ;
        RECT 30.980 12.230 31.120 13.950 ;
        RECT 32.820 12.230 32.960 14.290 ;
        RECT 33.280 12.230 33.420 20.670 ;
        RECT 34.140 20.070 34.400 20.390 ;
        RECT 34.200 18.690 34.340 20.070 ;
        RECT 34.140 18.370 34.400 18.690 ;
        RECT 34.200 15.630 34.340 18.370 ;
        RECT 35.120 17.920 35.260 23.810 ;
        RECT 35.580 21.320 35.720 30.950 ;
        RECT 35.980 25.850 36.240 26.170 ;
        RECT 36.040 24.130 36.180 25.850 ;
        RECT 35.980 23.810 36.240 24.130 ;
        RECT 35.980 21.320 36.240 21.410 ;
        RECT 35.580 21.180 36.240 21.320 ;
        RECT 35.980 21.090 36.240 21.180 ;
        RECT 36.040 20.730 36.180 21.090 ;
        RECT 35.980 20.410 36.240 20.730 ;
        RECT 34.660 17.780 35.260 17.920 ;
        RECT 34.140 15.310 34.400 15.630 ;
        RECT 34.660 13.250 34.800 17.780 ;
        RECT 35.060 16.670 35.320 16.990 ;
        RECT 35.120 15.630 35.260 16.670 ;
        RECT 35.060 15.310 35.320 15.630 ;
        RECT 34.600 12.930 34.860 13.250 ;
        RECT 30.000 11.910 30.260 12.230 ;
        RECT 30.920 11.910 31.180 12.230 ;
        RECT 32.760 11.910 33.020 12.230 ;
        RECT 33.220 11.910 33.480 12.230 ;
        RECT 36.040 12.140 36.180 20.410 ;
        RECT 36.500 20.050 36.640 36.820 ;
        RECT 36.960 33.990 37.100 39.110 ;
        RECT 36.900 33.670 37.160 33.990 ;
        RECT 37.820 27.890 38.080 28.210 ;
        RECT 37.880 25.150 38.020 27.890 ;
        RECT 38.280 27.550 38.540 27.870 ;
        RECT 37.820 24.830 38.080 25.150 ;
        RECT 37.880 21.070 38.020 24.830 ;
        RECT 38.340 23.110 38.480 27.550 ;
        RECT 38.280 22.790 38.540 23.110 ;
        RECT 37.820 20.750 38.080 21.070 ;
        RECT 36.440 19.730 36.700 20.050 ;
        RECT 36.440 18.370 36.700 18.690 ;
        RECT 36.500 18.205 36.640 18.370 ;
        RECT 36.430 17.835 36.710 18.205 ;
        RECT 36.500 17.670 36.640 17.835 ;
        RECT 36.440 17.350 36.700 17.670 ;
        RECT 37.360 17.350 37.620 17.670 ;
        RECT 37.420 13.250 37.560 17.350 ;
        RECT 37.360 12.930 37.620 13.250 ;
        RECT 37.880 12.230 38.020 20.750 ;
        RECT 38.800 13.870 38.940 62.030 ;
        RECT 39.200 60.190 39.460 60.510 ;
        RECT 39.260 54.050 39.400 60.190 ;
        RECT 39.720 56.090 39.860 62.910 ;
        RECT 40.640 61.190 40.780 63.590 ;
        RECT 41.100 61.610 41.240 66.310 ;
        RECT 41.960 65.630 42.220 65.950 ;
        RECT 41.500 63.930 41.760 64.250 ;
        RECT 41.560 62.210 41.700 63.930 ;
        RECT 41.500 61.890 41.760 62.210 ;
        RECT 41.100 61.530 41.700 61.610 ;
        RECT 41.040 61.470 41.700 61.530 ;
        RECT 41.040 61.210 41.300 61.470 ;
        RECT 40.580 60.870 40.840 61.190 ;
        RECT 41.560 60.510 41.700 61.470 ;
        RECT 41.500 60.190 41.760 60.510 ;
        RECT 42.020 56.770 42.160 65.630 ;
        RECT 42.420 61.890 42.680 62.210 ;
        RECT 41.960 56.450 42.220 56.770 ;
        RECT 42.480 56.170 42.620 61.890 ;
        RECT 39.660 55.770 39.920 56.090 ;
        RECT 42.020 56.030 42.620 56.170 ;
        RECT 39.200 53.730 39.460 54.050 ;
        RECT 40.580 53.050 40.840 53.370 ;
        RECT 40.640 50.310 40.780 53.050 ;
        RECT 41.500 52.710 41.760 53.030 ;
        RECT 40.580 49.990 40.840 50.310 ;
        RECT 41.560 46.910 41.700 52.710 ;
        RECT 42.020 50.310 42.160 56.030 ;
        RECT 42.420 53.050 42.680 53.370 ;
        RECT 41.960 49.990 42.220 50.310 ;
        RECT 39.660 46.590 39.920 46.910 ;
        RECT 41.500 46.590 41.760 46.910 ;
        RECT 39.720 45.210 39.860 46.590 ;
        RECT 41.560 45.210 41.700 46.590 ;
        RECT 39.660 44.890 39.920 45.210 ;
        RECT 41.500 44.890 41.760 45.210 ;
        RECT 41.560 39.090 41.700 44.890 ;
        RECT 42.020 42.490 42.160 49.990 ;
        RECT 41.960 42.170 42.220 42.490 ;
        RECT 40.120 38.770 40.380 39.090 ;
        RECT 41.500 38.770 41.760 39.090 ;
        RECT 40.180 37.730 40.320 38.770 ;
        RECT 40.120 37.410 40.380 37.730 ;
        RECT 41.960 36.565 42.220 36.710 ;
        RECT 41.950 36.195 42.230 36.565 ;
        RECT 42.020 34.670 42.160 36.195 ;
        RECT 41.960 34.350 42.220 34.670 ;
        RECT 39.200 33.670 39.460 33.990 ;
        RECT 39.660 33.670 39.920 33.990 ;
        RECT 40.120 33.670 40.380 33.990 ;
        RECT 39.260 23.790 39.400 33.670 ;
        RECT 39.720 32.290 39.860 33.670 ;
        RECT 39.660 31.970 39.920 32.290 ;
        RECT 40.180 26.850 40.320 33.670 ;
        RECT 41.960 28.570 42.220 28.890 ;
        RECT 40.120 26.530 40.380 26.850 ;
        RECT 39.200 23.470 39.460 23.790 ;
        RECT 40.180 23.110 40.320 26.530 ;
        RECT 41.040 23.130 41.300 23.450 ;
        RECT 40.120 22.790 40.380 23.110 ;
        RECT 39.200 20.925 39.460 21.070 ;
        RECT 39.190 20.555 39.470 20.925 ;
        RECT 40.180 17.670 40.320 22.790 ;
        RECT 41.100 18.010 41.240 23.130 ;
        RECT 42.020 22.770 42.160 28.570 ;
        RECT 41.960 22.450 42.220 22.770 ;
        RECT 42.020 21.410 42.160 22.450 ;
        RECT 41.960 21.090 42.220 21.410 ;
        RECT 41.500 20.070 41.760 20.390 ;
        RECT 41.040 17.690 41.300 18.010 ;
        RECT 40.120 17.350 40.380 17.670 ;
        RECT 40.580 16.670 40.840 16.990 ;
        RECT 40.640 15.290 40.780 16.670 ;
        RECT 41.560 15.970 41.700 20.070 ;
        RECT 41.500 15.650 41.760 15.970 ;
        RECT 40.580 14.970 40.840 15.290 ;
        RECT 38.800 13.730 40.320 13.870 ;
        RECT 40.180 12.910 40.320 13.730 ;
        RECT 40.120 12.590 40.380 12.910 ;
        RECT 41.560 12.230 41.700 15.650 ;
        RECT 36.440 12.140 36.700 12.230 ;
        RECT 36.040 12.000 36.700 12.140 ;
        RECT 36.440 11.910 36.700 12.000 ;
        RECT 37.820 11.910 38.080 12.230 ;
        RECT 41.500 11.910 41.760 12.230 ;
        RECT 42.020 11.890 42.160 21.090 ;
        RECT 42.480 20.050 42.620 53.050 ;
        RECT 42.940 47.250 43.080 94.190 ;
        RECT 43.400 94.170 43.540 120.030 ;
        RECT 46.160 115.250 46.300 158.630 ;
        RECT 46.620 157.410 46.760 158.790 ;
        RECT 47.080 158.770 47.220 164.910 ;
        RECT 47.080 158.630 48.140 158.770 ;
        RECT 47.020 158.110 47.280 158.430 ;
        RECT 47.480 158.110 47.740 158.430 ;
        RECT 46.560 157.090 46.820 157.410 ;
        RECT 46.620 153.670 46.760 157.090 ;
        RECT 47.080 156.390 47.220 158.110 ;
        RECT 47.020 156.070 47.280 156.390 ;
        RECT 47.080 154.690 47.220 156.070 ;
        RECT 47.020 154.370 47.280 154.690 ;
        RECT 46.560 153.350 46.820 153.670 ;
        RECT 47.540 152.990 47.680 158.110 ;
        RECT 46.560 152.670 46.820 152.990 ;
        RECT 47.480 152.670 47.740 152.990 ;
        RECT 46.620 150.610 46.760 152.670 ;
        RECT 47.020 150.970 47.280 151.290 ;
        RECT 46.560 150.290 46.820 150.610 ;
        RECT 47.080 148.910 47.220 150.970 ;
        RECT 48.000 150.610 48.140 158.630 ;
        RECT 49.380 151.290 49.520 165.250 ;
        RECT 49.840 164.890 49.980 167.290 ;
        RECT 49.780 164.570 50.040 164.890 ;
        RECT 49.840 156.730 49.980 164.570 ;
        RECT 50.300 164.550 50.440 170.010 ;
        RECT 51.220 169.900 51.360 174.770 ;
        RECT 52.140 171.010 52.280 174.770 ;
        RECT 52.080 170.690 52.340 171.010 ;
        RECT 52.080 169.900 52.340 169.990 ;
        RECT 51.220 169.760 52.340 169.900 ;
        RECT 52.080 169.670 52.340 169.760 ;
        RECT 50.700 167.630 50.960 167.950 ;
        RECT 50.760 164.890 50.900 167.630 ;
        RECT 52.140 166.930 52.280 169.670 ;
        RECT 52.080 166.610 52.340 166.930 ;
        RECT 52.600 166.590 52.740 175.110 ;
        RECT 53.980 175.030 54.580 175.170 ;
        RECT 53.460 173.070 53.720 173.390 ;
        RECT 52.540 166.270 52.800 166.590 ;
        RECT 53.000 166.270 53.260 166.590 ;
        RECT 50.700 164.570 50.960 164.890 ;
        RECT 50.240 164.230 50.500 164.550 ;
        RECT 50.300 162.510 50.440 164.230 ;
        RECT 50.240 162.190 50.500 162.510 ;
        RECT 50.760 162.170 50.900 164.570 ;
        RECT 53.060 164.550 53.200 166.270 ;
        RECT 53.000 164.230 53.260 164.550 ;
        RECT 51.160 163.890 51.420 164.210 ;
        RECT 51.220 162.170 51.360 163.890 ;
        RECT 53.520 163.610 53.660 173.070 ;
        RECT 53.980 168.290 54.120 175.030 ;
        RECT 55.820 173.730 55.960 177.920 ;
        RECT 56.740 177.810 56.880 180.210 ;
        RECT 57.660 179.170 57.800 180.550 ;
        RECT 57.600 178.850 57.860 179.170 ;
        RECT 57.140 178.510 57.400 178.830 ;
        RECT 56.680 177.490 56.940 177.810 ;
        RECT 57.200 177.210 57.340 178.510 ;
        RECT 56.740 177.070 57.340 177.210 ;
        RECT 56.740 175.430 56.880 177.070 ;
        RECT 57.660 175.430 57.800 178.850 ;
        RECT 60.420 178.490 60.560 181.230 ;
        RECT 60.880 178.830 61.020 181.570 ;
        RECT 61.340 180.190 61.480 189.730 ;
        RECT 61.800 189.370 61.940 190.750 ;
        RECT 63.180 189.710 63.320 196.190 ;
        RECT 63.580 194.490 63.840 194.810 ;
        RECT 63.640 192.770 63.780 194.490 ;
        RECT 69.560 194.150 69.820 194.470 ;
        RECT 63.580 192.450 63.840 192.770 ;
        RECT 69.620 192.090 69.760 194.150 ;
        RECT 69.560 191.770 69.820 192.090 ;
        RECT 65.420 191.090 65.680 191.410 ;
        RECT 65.480 190.050 65.620 191.090 ;
        RECT 65.420 189.730 65.680 190.050 ;
        RECT 63.120 189.390 63.380 189.710 ;
        RECT 61.740 189.050 62.000 189.370 ;
        RECT 64.040 189.050 64.300 189.370 ;
        RECT 66.800 189.050 67.060 189.370 ;
        RECT 61.800 186.650 61.940 189.050 ;
        RECT 63.120 188.710 63.380 189.030 ;
        RECT 61.740 186.330 62.000 186.650 ;
        RECT 63.180 186.310 63.320 188.710 ;
        RECT 64.100 187.330 64.240 189.050 ;
        RECT 64.040 187.010 64.300 187.330 ;
        RECT 66.860 186.310 67.000 189.050 ;
        RECT 63.120 185.990 63.380 186.310 ;
        RECT 66.800 185.990 67.060 186.310 ;
        RECT 64.960 185.650 65.220 185.970 ;
        RECT 64.040 180.210 64.300 180.530 ;
        RECT 61.280 179.870 61.540 180.190 ;
        RECT 62.200 179.870 62.460 180.190 ;
        RECT 60.820 178.510 61.080 178.830 ;
        RECT 60.360 178.170 60.620 178.490 ;
        RECT 56.680 175.110 56.940 175.430 ;
        RECT 57.600 175.110 57.860 175.430 ;
        RECT 58.060 175.110 58.320 175.430 ;
        RECT 55.760 173.410 56.020 173.730 ;
        RECT 55.820 169.990 55.960 173.410 ;
        RECT 56.740 173.390 56.880 175.110 ;
        RECT 56.680 173.070 56.940 173.390 ;
        RECT 55.760 169.670 56.020 169.990 ;
        RECT 56.220 169.670 56.480 169.990 ;
        RECT 53.920 167.970 54.180 168.290 ;
        RECT 53.980 167.610 54.120 167.970 ;
        RECT 53.920 167.290 54.180 167.610 ;
        RECT 53.980 166.590 54.120 167.290 ;
        RECT 53.920 166.270 54.180 166.590 ;
        RECT 55.820 165.480 55.960 169.670 ;
        RECT 56.280 167.270 56.420 169.670 ;
        RECT 58.120 168.290 58.260 175.110 ;
        RECT 60.420 175.090 60.560 178.170 ;
        RECT 61.340 177.470 61.480 179.870 ;
        RECT 61.740 178.510 62.000 178.830 ;
        RECT 62.260 178.740 62.400 179.870 ;
        RECT 62.660 178.740 62.920 178.830 ;
        RECT 62.260 178.600 62.920 178.740 ;
        RECT 62.660 178.510 62.920 178.600 ;
        RECT 61.280 177.150 61.540 177.470 ;
        RECT 61.340 175.770 61.480 177.150 ;
        RECT 61.800 176.450 61.940 178.510 ;
        RECT 62.200 177.830 62.460 178.150 ;
        RECT 63.120 177.830 63.380 178.150 ;
        RECT 61.740 176.130 62.000 176.450 ;
        RECT 61.280 175.450 61.540 175.770 ;
        RECT 60.360 174.770 60.620 175.090 ;
        RECT 60.420 169.310 60.560 174.770 ;
        RECT 62.260 174.750 62.400 177.830 ;
        RECT 62.200 174.430 62.460 174.750 ;
        RECT 61.280 172.730 61.540 173.050 ;
        RECT 61.340 169.990 61.480 172.730 ;
        RECT 62.260 172.710 62.400 174.430 ;
        RECT 62.660 172.730 62.920 173.050 ;
        RECT 62.200 172.390 62.460 172.710 ;
        RECT 61.740 171.710 62.000 172.030 ;
        RECT 61.280 169.670 61.540 169.990 ;
        RECT 60.360 168.990 60.620 169.310 ;
        RECT 58.060 167.970 58.320 168.290 ;
        RECT 58.520 167.970 58.780 168.290 ;
        RECT 56.220 166.950 56.480 167.270 ;
        RECT 55.820 165.340 56.420 165.480 ;
        RECT 54.380 164.570 54.640 164.890 ;
        RECT 55.760 164.570 56.020 164.890 ;
        RECT 52.600 163.470 53.660 163.610 ;
        RECT 52.600 162.850 52.740 163.470 ;
        RECT 52.540 162.530 52.800 162.850 ;
        RECT 50.700 161.850 50.960 162.170 ;
        RECT 51.160 161.850 51.420 162.170 ;
        RECT 51.220 159.110 51.360 161.850 ;
        RECT 51.160 158.790 51.420 159.110 ;
        RECT 49.780 156.410 50.040 156.730 ;
        RECT 51.220 154.090 51.360 158.790 ;
        RECT 51.220 153.950 51.820 154.090 ;
        RECT 49.780 153.350 50.040 153.670 ;
        RECT 51.160 153.350 51.420 153.670 ;
        RECT 49.840 151.970 49.980 153.350 ;
        RECT 49.780 151.650 50.040 151.970 ;
        RECT 49.320 150.970 49.580 151.290 ;
        RECT 47.940 150.290 48.200 150.610 ;
        RECT 47.480 149.950 47.740 150.270 ;
        RECT 47.020 148.590 47.280 148.910 ;
        RECT 47.080 146.530 47.220 148.590 ;
        RECT 47.540 148.230 47.680 149.950 ;
        RECT 47.480 147.910 47.740 148.230 ;
        RECT 51.220 147.890 51.360 153.350 ;
        RECT 51.160 147.570 51.420 147.890 ;
        RECT 47.020 146.210 47.280 146.530 ;
        RECT 51.160 145.530 51.420 145.850 ;
        RECT 51.220 143.810 51.360 145.530 ;
        RECT 51.160 143.490 51.420 143.810 ;
        RECT 51.680 140.750 51.820 153.950 ;
        RECT 52.080 148.930 52.340 149.250 ;
        RECT 52.140 148.570 52.280 148.930 ;
        RECT 52.080 148.250 52.340 148.570 ;
        RECT 51.620 140.430 51.880 140.750 ;
        RECT 52.140 140.410 52.280 148.250 ;
        RECT 52.600 142.790 52.740 162.530 ;
        RECT 54.440 157.070 54.580 164.570 ;
        RECT 55.820 162.170 55.960 164.570 ;
        RECT 56.280 162.170 56.420 165.340 ;
        RECT 58.580 162.850 58.720 167.970 ;
        RECT 59.900 167.520 60.160 167.610 ;
        RECT 60.420 167.520 60.560 168.990 ;
        RECT 61.340 167.610 61.480 169.670 ;
        RECT 61.800 169.650 61.940 171.710 ;
        RECT 62.720 171.010 62.860 172.730 ;
        RECT 62.660 170.690 62.920 171.010 ;
        RECT 62.190 170.155 62.470 170.525 ;
        RECT 62.200 170.010 62.460 170.155 ;
        RECT 61.740 169.330 62.000 169.650 ;
        RECT 63.180 167.950 63.320 177.830 ;
        RECT 64.100 177.470 64.240 180.210 ;
        RECT 64.040 177.150 64.300 177.470 ;
        RECT 65.020 175.430 65.160 185.650 ;
        RECT 69.620 181.210 69.760 191.770 ;
        RECT 69.560 180.890 69.820 181.210 ;
        RECT 65.420 180.550 65.680 180.870 ;
        RECT 65.480 179.170 65.620 180.550 ;
        RECT 65.420 178.850 65.680 179.170 ;
        RECT 64.960 175.110 65.220 175.430 ;
        RECT 63.580 174.430 63.840 174.750 ;
        RECT 63.640 173.050 63.780 174.430 ;
        RECT 63.580 172.730 63.840 173.050 ;
        RECT 64.040 172.730 64.300 173.050 ;
        RECT 64.100 172.370 64.240 172.730 ;
        RECT 64.500 172.390 64.760 172.710 ;
        RECT 64.040 172.050 64.300 172.370 ;
        RECT 63.580 171.710 63.840 172.030 ;
        RECT 63.640 170.670 63.780 171.710 ;
        RECT 63.580 170.350 63.840 170.670 ;
        RECT 64.100 169.990 64.240 172.050 ;
        RECT 64.040 169.670 64.300 169.990 ;
        RECT 63.120 167.630 63.380 167.950 ;
        RECT 59.900 167.380 60.560 167.520 ;
        RECT 59.900 167.290 60.160 167.380 ;
        RECT 61.280 167.290 61.540 167.610 ;
        RECT 64.040 167.290 64.300 167.610 ;
        RECT 60.820 166.950 61.080 167.270 ;
        RECT 60.880 164.890 61.020 166.950 ;
        RECT 63.580 166.270 63.840 166.590 ;
        RECT 60.820 164.570 61.080 164.890 ;
        RECT 58.520 162.530 58.780 162.850 ;
        RECT 55.760 161.850 56.020 162.170 ;
        RECT 56.220 161.850 56.480 162.170 ;
        RECT 57.140 160.830 57.400 161.150 ;
        RECT 57.200 159.110 57.340 160.830 ;
        RECT 57.140 158.790 57.400 159.110 ;
        RECT 57.600 158.790 57.860 159.110 ;
        RECT 55.300 158.110 55.560 158.430 ;
        RECT 54.380 156.750 54.640 157.070 ;
        RECT 53.460 155.390 53.720 155.710 ;
        RECT 53.920 155.390 54.180 155.710 ;
        RECT 53.520 153.670 53.660 155.390 ;
        RECT 53.980 154.350 54.120 155.390 ;
        RECT 55.360 154.690 55.500 158.110 ;
        RECT 57.660 156.730 57.800 158.790 ;
        RECT 57.600 156.410 57.860 156.730 ;
        RECT 55.300 154.370 55.560 154.690 ;
        RECT 53.920 154.030 54.180 154.350 ;
        RECT 53.460 153.350 53.720 153.670 ;
        RECT 54.840 153.580 55.100 153.670 ;
        RECT 55.360 153.580 55.500 154.370 ;
        RECT 58.580 154.010 58.720 162.530 ;
        RECT 59.440 162.190 59.700 162.510 ;
        RECT 55.760 153.690 56.020 154.010 ;
        RECT 58.520 153.690 58.780 154.010 ;
        RECT 54.840 153.440 55.500 153.580 ;
        RECT 54.840 153.350 55.100 153.440 ;
        RECT 53.920 152.670 54.180 152.990 ;
        RECT 53.980 148.230 54.120 152.670 ;
        RECT 55.300 150.970 55.560 151.290 ;
        RECT 53.460 147.910 53.720 148.230 ;
        RECT 53.920 147.910 54.180 148.230 ;
        RECT 53.000 147.230 53.260 147.550 ;
        RECT 53.060 146.530 53.200 147.230 ;
        RECT 53.520 146.530 53.660 147.910 ;
        RECT 54.380 147.800 54.640 147.890 ;
        RECT 55.360 147.800 55.500 150.970 ;
        RECT 55.820 149.330 55.960 153.690 ;
        RECT 56.680 153.350 56.940 153.670 ;
        RECT 56.220 152.670 56.480 152.990 ;
        RECT 56.280 150.270 56.420 152.670 ;
        RECT 56.740 151.290 56.880 153.350 ;
        RECT 56.680 150.970 56.940 151.290 ;
        RECT 56.220 149.950 56.480 150.270 ;
        RECT 57.140 149.950 57.400 150.270 ;
        RECT 55.820 149.250 56.420 149.330 ;
        RECT 55.820 149.190 56.480 149.250 ;
        RECT 56.220 148.930 56.480 149.190 ;
        RECT 54.380 147.660 55.500 147.800 ;
        RECT 54.380 147.570 54.640 147.660 ;
        RECT 53.000 146.210 53.260 146.530 ;
        RECT 53.460 146.210 53.720 146.530 ;
        RECT 53.000 145.530 53.260 145.850 ;
        RECT 53.060 142.790 53.200 145.530 ;
        RECT 55.360 143.810 55.500 147.660 ;
        RECT 57.200 146.190 57.340 149.950 ;
        RECT 58.060 147.570 58.320 147.890 ;
        RECT 57.140 145.870 57.400 146.190 ;
        RECT 55.300 143.490 55.560 143.810 ;
        RECT 52.540 142.470 52.800 142.790 ;
        RECT 53.000 142.470 53.260 142.790 ;
        RECT 57.600 142.470 57.860 142.790 ;
        RECT 52.600 140.410 52.740 142.470 ;
        RECT 53.060 141.090 53.200 142.470 ;
        RECT 53.460 142.130 53.720 142.450 ;
        RECT 57.140 142.130 57.400 142.450 ;
        RECT 53.000 140.770 53.260 141.090 ;
        RECT 53.520 140.410 53.660 142.130 ;
        RECT 49.320 140.090 49.580 140.410 ;
        RECT 52.080 140.090 52.340 140.410 ;
        RECT 52.540 140.090 52.800 140.410 ;
        RECT 53.460 140.090 53.720 140.410 ;
        RECT 47.540 138.370 49.060 138.450 ;
        RECT 49.380 138.370 49.520 140.090 ;
        RECT 50.700 139.750 50.960 140.070 ;
        RECT 47.480 138.310 49.060 138.370 ;
        RECT 47.480 138.050 47.740 138.310 ;
        RECT 48.400 137.710 48.660 138.030 ;
        RECT 46.560 137.205 46.820 137.350 ;
        RECT 46.550 136.835 46.830 137.205 ;
        RECT 47.940 136.690 48.200 137.010 ;
        RECT 46.560 136.350 46.820 136.670 ;
        RECT 46.620 132.930 46.760 136.350 ;
        RECT 48.000 134.630 48.140 136.690 ;
        RECT 48.460 134.970 48.600 137.710 ;
        RECT 48.920 136.670 49.060 138.310 ;
        RECT 49.320 138.050 49.580 138.370 ;
        RECT 50.760 137.690 50.900 139.750 ;
        RECT 52.140 139.130 52.280 140.090 ;
        RECT 51.680 138.990 52.280 139.130 ;
        RECT 50.700 137.370 50.960 137.690 ;
        RECT 48.860 136.350 49.120 136.670 ;
        RECT 48.400 134.650 48.660 134.970 ;
        RECT 47.940 134.310 48.200 134.630 ;
        RECT 48.920 133.950 49.060 136.350 ;
        RECT 50.760 134.970 50.900 137.370 ;
        RECT 51.160 136.690 51.420 137.010 ;
        RECT 51.220 135.310 51.360 136.690 ;
        RECT 51.160 134.990 51.420 135.310 ;
        RECT 50.700 134.650 50.960 134.970 ;
        RECT 48.860 133.630 49.120 133.950 ;
        RECT 46.560 132.610 46.820 132.930 ;
        RECT 46.620 130.210 46.760 132.610 ;
        RECT 46.560 129.890 46.820 130.210 ;
        RECT 46.620 125.790 46.760 129.890 ;
        RECT 50.760 129.610 50.900 134.650 ;
        RECT 50.300 129.530 50.900 129.610 ;
        RECT 50.240 129.470 50.900 129.530 ;
        RECT 50.240 129.210 50.500 129.470 ;
        RECT 47.480 128.190 47.740 128.510 ;
        RECT 47.540 126.130 47.680 128.190 ;
        RECT 50.300 126.470 50.440 129.210 ;
        RECT 50.240 126.150 50.500 126.470 ;
        RECT 47.480 125.810 47.740 126.130 ;
        RECT 46.560 125.470 46.820 125.790 ;
        RECT 48.860 120.030 49.120 120.350 ;
        RECT 48.920 118.650 49.060 120.030 ;
        RECT 50.300 118.990 50.440 126.150 ;
        RECT 50.240 118.670 50.500 118.990 ;
        RECT 48.860 118.330 49.120 118.650 ;
        RECT 50.300 115.590 50.440 118.670 ;
        RECT 50.240 115.270 50.500 115.590 ;
        RECT 46.100 114.930 46.360 115.250 ;
        RECT 49.320 114.590 49.580 114.910 ;
        RECT 43.800 112.890 44.060 113.210 ;
        RECT 43.860 104.030 44.000 112.890 ;
        RECT 49.380 109.810 49.520 114.590 ;
        RECT 49.780 110.850 50.040 111.170 ;
        RECT 49.320 109.490 49.580 109.810 ;
        RECT 48.400 109.150 48.660 109.470 ;
        RECT 48.460 107.770 48.600 109.150 ;
        RECT 49.380 107.770 49.520 109.490 ;
        RECT 49.840 107.770 49.980 110.850 ;
        RECT 50.300 110.490 50.440 115.270 ;
        RECT 50.240 110.170 50.500 110.490 ;
        RECT 48.400 107.450 48.660 107.770 ;
        RECT 49.320 107.450 49.580 107.770 ;
        RECT 49.780 107.450 50.040 107.770 ;
        RECT 43.800 103.710 44.060 104.030 ;
        RECT 43.340 93.850 43.600 94.170 ;
        RECT 43.860 90.340 44.000 103.710 ;
        RECT 48.460 102.670 48.600 107.450 ;
        RECT 48.860 107.110 49.120 107.430 ;
        RECT 48.920 104.370 49.060 107.110 ;
        RECT 51.220 105.730 51.360 134.990 ;
        RECT 51.680 132.250 51.820 138.990 ;
        RECT 53.000 136.410 53.260 136.670 ;
        RECT 53.520 136.410 53.660 140.090 ;
        RECT 53.920 137.370 54.180 137.690 ;
        RECT 53.000 136.350 53.660 136.410 ;
        RECT 53.060 136.270 53.660 136.350 ;
        RECT 52.080 135.330 52.340 135.650 ;
        RECT 52.140 132.250 52.280 135.330 ;
        RECT 51.620 131.930 51.880 132.250 ;
        RECT 52.080 131.930 52.340 132.250 ;
        RECT 53.060 127.490 53.200 136.270 ;
        RECT 53.460 134.990 53.720 135.310 ;
        RECT 53.520 131.910 53.660 134.990 ;
        RECT 53.980 131.910 54.120 137.370 ;
        RECT 55.760 137.030 56.020 137.350 ;
        RECT 55.820 131.910 55.960 137.030 ;
        RECT 57.200 137.010 57.340 142.130 ;
        RECT 57.660 141.090 57.800 142.470 ;
        RECT 57.600 140.770 57.860 141.090 ;
        RECT 57.140 136.690 57.400 137.010 ;
        RECT 58.120 136.670 58.260 147.570 ;
        RECT 58.580 146.190 58.720 153.690 ;
        RECT 58.980 153.350 59.240 153.670 ;
        RECT 59.040 151.290 59.180 153.350 ;
        RECT 58.980 150.970 59.240 151.290 ;
        RECT 58.520 145.870 58.780 146.190 ;
        RECT 59.040 145.850 59.180 150.970 ;
        RECT 58.980 145.530 59.240 145.850 ;
        RECT 59.500 142.450 59.640 162.190 ;
        RECT 60.880 154.010 61.020 164.570 ;
        RECT 62.200 158.790 62.460 159.110 ;
        RECT 63.120 158.790 63.380 159.110 ;
        RECT 62.260 154.090 62.400 158.790 ;
        RECT 63.180 156.050 63.320 158.790 ;
        RECT 63.120 155.730 63.380 156.050 ;
        RECT 60.820 153.690 61.080 154.010 ;
        RECT 62.260 153.950 63.320 154.090 ;
        RECT 60.880 151.290 61.020 153.690 ;
        RECT 62.200 153.350 62.460 153.670 ;
        RECT 62.260 151.290 62.400 153.350 ;
        RECT 63.180 151.630 63.320 153.950 ;
        RECT 63.120 151.310 63.380 151.630 ;
        RECT 60.820 150.970 61.080 151.290 ;
        RECT 62.200 150.970 62.460 151.290 ;
        RECT 62.260 150.610 62.400 150.970 ;
        RECT 62.200 150.290 62.460 150.610 ;
        RECT 63.180 150.270 63.320 151.310 ;
        RECT 61.740 149.950 62.000 150.270 ;
        RECT 63.120 149.950 63.380 150.270 ;
        RECT 61.800 148.230 61.940 149.950 ;
        RECT 59.900 147.910 60.160 148.230 ;
        RECT 61.740 147.910 62.000 148.230 ;
        RECT 59.960 145.850 60.100 147.910 ;
        RECT 60.820 147.570 61.080 147.890 ;
        RECT 60.880 145.850 61.020 147.570 ;
        RECT 59.900 145.530 60.160 145.850 ;
        RECT 60.820 145.530 61.080 145.850 ;
        RECT 60.360 145.190 60.620 145.510 ;
        RECT 59.440 142.130 59.700 142.450 ;
        RECT 60.420 140.410 60.560 145.190 ;
        RECT 61.800 143.210 61.940 147.910 ;
        RECT 63.640 146.190 63.780 166.270 ;
        RECT 64.100 165.570 64.240 167.290 ;
        RECT 64.040 165.250 64.300 165.570 ;
        RECT 64.560 164.210 64.700 172.390 ;
        RECT 65.020 172.030 65.160 175.110 ;
        RECT 65.480 173.050 65.620 178.850 ;
        RECT 65.880 173.070 66.140 173.390 ;
        RECT 65.420 172.730 65.680 173.050 ;
        RECT 64.960 171.710 65.220 172.030 ;
        RECT 65.480 171.010 65.620 172.730 ;
        RECT 65.420 170.690 65.680 171.010 ;
        RECT 64.960 170.350 65.220 170.670 ;
        RECT 65.480 170.525 65.620 170.690 ;
        RECT 65.020 169.310 65.160 170.350 ;
        RECT 65.410 170.155 65.690 170.525 ;
        RECT 65.940 169.990 66.080 173.070 ;
        RECT 66.800 172.730 67.060 173.050 ;
        RECT 66.860 170.670 67.000 172.730 ;
        RECT 68.640 170.690 68.900 171.010 ;
        RECT 66.800 170.350 67.060 170.670 ;
        RECT 65.880 169.670 66.140 169.990 ;
        RECT 66.860 169.310 67.000 170.350 ;
        RECT 68.700 169.650 68.840 170.690 ;
        RECT 69.620 170.330 69.760 180.890 ;
        RECT 69.560 170.010 69.820 170.330 ;
        RECT 68.640 169.330 68.900 169.650 ;
        RECT 64.960 168.990 65.220 169.310 ;
        RECT 65.420 168.990 65.680 169.310 ;
        RECT 65.880 168.990 66.140 169.310 ;
        RECT 66.800 168.990 67.060 169.310 ;
        RECT 65.480 165.570 65.620 168.990 ;
        RECT 65.420 165.250 65.680 165.570 ;
        RECT 65.940 164.210 66.080 168.990 ;
        RECT 69.620 167.610 69.760 170.010 ;
        RECT 69.560 167.290 69.820 167.610 ;
        RECT 69.620 164.550 69.760 167.290 ;
        RECT 69.560 164.230 69.820 164.550 ;
        RECT 64.500 163.890 64.760 164.210 ;
        RECT 65.880 163.890 66.140 164.210 ;
        RECT 69.620 162.510 69.760 164.230 ;
        RECT 69.560 162.190 69.820 162.510 ;
        RECT 64.500 158.790 64.760 159.110 ;
        RECT 64.960 158.790 65.220 159.110 ;
        RECT 64.040 155.730 64.300 156.050 ;
        RECT 64.100 154.690 64.240 155.730 ;
        RECT 64.040 154.370 64.300 154.690 ;
        RECT 64.040 153.350 64.300 153.670 ;
        RECT 64.100 151.970 64.240 153.350 ;
        RECT 64.040 151.650 64.300 151.970 ;
        RECT 64.560 148.910 64.700 158.790 ;
        RECT 65.020 156.390 65.160 158.790 ;
        RECT 69.620 158.770 69.760 162.190 ;
        RECT 69.620 158.630 70.680 158.770 ;
        RECT 66.800 158.110 67.060 158.430 ;
        RECT 66.860 157.070 67.000 158.110 ;
        RECT 65.880 156.750 66.140 157.070 ;
        RECT 66.800 156.750 67.060 157.070 ;
        RECT 67.720 156.750 67.980 157.070 ;
        RECT 64.960 156.070 65.220 156.390 ;
        RECT 64.960 155.390 65.220 155.710 ;
        RECT 65.020 154.350 65.160 155.390 ;
        RECT 64.960 154.030 65.220 154.350 ;
        RECT 64.500 148.590 64.760 148.910 ;
        RECT 64.500 147.230 64.760 147.550 ;
        RECT 63.580 145.870 63.840 146.190 ;
        RECT 64.040 145.530 64.300 145.850 ;
        RECT 63.580 145.190 63.840 145.510 ;
        RECT 61.340 143.070 61.940 143.210 ;
        RECT 58.520 140.090 58.780 140.410 ;
        RECT 60.360 140.090 60.620 140.410 ;
        RECT 58.580 137.350 58.720 140.090 ;
        RECT 58.520 137.030 58.780 137.350 ;
        RECT 58.980 136.690 59.240 137.010 ;
        RECT 58.060 136.350 58.320 136.670 ;
        RECT 58.120 135.560 58.260 136.350 ;
        RECT 58.120 135.420 58.720 135.560 ;
        RECT 58.060 134.650 58.320 134.970 ;
        RECT 58.120 132.930 58.260 134.650 ;
        RECT 58.580 134.290 58.720 135.420 ;
        RECT 58.520 133.970 58.780 134.290 ;
        RECT 58.580 132.930 58.720 133.970 ;
        RECT 58.060 132.610 58.320 132.930 ;
        RECT 58.520 132.610 58.780 132.930 ;
        RECT 57.140 132.270 57.400 132.590 ;
        RECT 53.460 131.590 53.720 131.910 ;
        RECT 53.920 131.590 54.180 131.910 ;
        RECT 55.760 131.590 56.020 131.910 ;
        RECT 53.460 130.910 53.720 131.230 ;
        RECT 53.520 129.870 53.660 130.910 ;
        RECT 55.820 130.210 55.960 131.590 ;
        RECT 55.760 129.890 56.020 130.210 ;
        RECT 53.460 129.550 53.720 129.870 ;
        RECT 53.000 127.170 53.260 127.490 ;
        RECT 57.200 126.470 57.340 132.270 ;
        RECT 59.040 131.570 59.180 136.690 ;
        RECT 60.420 136.670 60.560 140.090 ;
        RECT 61.340 137.010 61.480 143.070 ;
        RECT 61.740 142.130 62.000 142.450 ;
        RECT 63.120 142.130 63.380 142.450 ;
        RECT 61.800 140.070 61.940 142.130 ;
        RECT 61.740 139.750 62.000 140.070 ;
        RECT 61.280 136.690 61.540 137.010 ;
        RECT 60.360 136.580 60.620 136.670 ;
        RECT 59.960 136.440 60.620 136.580 ;
        RECT 59.960 131.570 60.100 136.440 ;
        RECT 60.360 136.350 60.620 136.440 ;
        RECT 60.360 134.650 60.620 134.970 ;
        RECT 60.420 132.930 60.560 134.650 ;
        RECT 60.820 133.630 61.080 133.950 ;
        RECT 60.360 132.610 60.620 132.930 ;
        RECT 58.980 131.250 59.240 131.570 ;
        RECT 59.900 131.250 60.160 131.570 ;
        RECT 59.960 130.210 60.100 131.250 ;
        RECT 59.900 129.890 60.160 130.210 ;
        RECT 59.900 129.210 60.160 129.530 ;
        RECT 59.960 127.490 60.100 129.210 ;
        RECT 59.900 127.170 60.160 127.490 ;
        RECT 60.880 126.810 61.020 133.630 ;
        RECT 61.340 132.930 61.480 136.690 ;
        RECT 61.280 132.610 61.540 132.930 ;
        RECT 61.800 129.870 61.940 139.750 ;
        RECT 63.180 135.650 63.320 142.130 ;
        RECT 63.120 135.330 63.380 135.650 ;
        RECT 63.640 135.310 63.780 145.190 ;
        RECT 64.100 137.205 64.240 145.530 ;
        RECT 64.560 145.510 64.700 147.230 ;
        RECT 65.020 146.530 65.160 154.030 ;
        RECT 65.420 152.670 65.680 152.990 ;
        RECT 64.960 146.210 65.220 146.530 ;
        RECT 65.480 145.850 65.620 152.670 ;
        RECT 65.940 151.630 66.080 156.750 ;
        RECT 66.340 154.370 66.600 154.690 ;
        RECT 66.400 153.670 66.540 154.370 ;
        RECT 67.260 154.030 67.520 154.350 ;
        RECT 67.320 153.670 67.460 154.030 ;
        RECT 66.340 153.350 66.600 153.670 ;
        RECT 67.260 153.350 67.520 153.670 ;
        RECT 65.880 151.310 66.140 151.630 ;
        RECT 65.940 150.950 66.080 151.310 ;
        RECT 65.880 150.630 66.140 150.950 ;
        RECT 65.880 148.590 66.140 148.910 ;
        RECT 65.420 145.530 65.680 145.850 ;
        RECT 64.500 145.190 64.760 145.510 ;
        RECT 65.940 142.790 66.080 148.590 ;
        RECT 66.400 147.970 66.540 153.350 ;
        RECT 66.800 151.650 67.060 151.970 ;
        RECT 66.860 150.690 67.000 151.650 ;
        RECT 66.860 150.550 67.460 150.690 ;
        RECT 67.320 148.230 67.460 150.550 ;
        RECT 66.400 147.830 67.000 147.970 ;
        RECT 67.260 147.910 67.520 148.230 ;
        RECT 66.860 143.470 67.000 147.830 ;
        RECT 67.260 145.190 67.520 145.510 ;
        RECT 66.800 143.150 67.060 143.470 ;
        RECT 67.320 143.130 67.460 145.190 ;
        RECT 67.260 142.810 67.520 143.130 ;
        RECT 65.880 142.470 66.140 142.790 ;
        RECT 67.780 142.450 67.920 156.750 ;
        RECT 70.540 155.710 70.680 158.630 ;
        RECT 70.480 155.390 70.740 155.710 ;
        RECT 72.320 155.390 72.580 155.710 ;
        RECT 70.540 154.010 70.680 155.390 ;
        RECT 70.020 153.690 70.280 154.010 ;
        RECT 70.480 153.690 70.740 154.010 ;
        RECT 68.640 150.630 68.900 150.950 ;
        RECT 68.180 150.290 68.440 150.610 ;
        RECT 68.240 148.230 68.380 150.290 ;
        RECT 68.180 147.910 68.440 148.230 ;
        RECT 68.700 142.450 68.840 150.630 ;
        RECT 70.080 150.610 70.220 153.690 ;
        RECT 70.480 152.670 70.740 152.990 ;
        RECT 70.540 151.630 70.680 152.670 ;
        RECT 70.480 151.310 70.740 151.630 ;
        RECT 72.380 151.290 72.520 155.390 ;
        RECT 72.320 150.970 72.580 151.290 ;
        RECT 70.020 150.290 70.280 150.610 ;
        RECT 74.160 147.910 74.420 148.230 ;
        RECT 74.220 146.530 74.360 147.910 ;
        RECT 74.160 146.210 74.420 146.530 ;
        RECT 69.100 142.470 69.360 142.790 ;
        RECT 67.720 142.130 67.980 142.450 ;
        RECT 68.640 142.130 68.900 142.450 ;
        RECT 64.500 141.790 64.760 142.110 ;
        RECT 64.560 140.750 64.700 141.790 ;
        RECT 68.700 141.090 68.840 142.130 ;
        RECT 68.640 140.770 68.900 141.090 ;
        RECT 64.500 140.430 64.760 140.750 ;
        RECT 64.030 136.835 64.310 137.205 ;
        RECT 62.200 134.990 62.460 135.310 ;
        RECT 63.580 134.990 63.840 135.310 ;
        RECT 62.260 134.630 62.400 134.990 ;
        RECT 62.200 134.310 62.460 134.630 ;
        RECT 63.580 134.370 63.840 134.630 ;
        RECT 64.100 134.370 64.240 136.835 ;
        RECT 69.160 134.970 69.300 142.470 ;
        RECT 69.100 134.650 69.360 134.970 ;
        RECT 69.560 134.650 69.820 134.970 ;
        RECT 63.580 134.310 64.240 134.370 ;
        RECT 65.420 134.310 65.680 134.630 ;
        RECT 61.740 129.550 62.000 129.870 ;
        RECT 62.260 127.150 62.400 134.310 ;
        RECT 63.640 134.230 64.240 134.310 ;
        RECT 65.480 132.930 65.620 134.310 ;
        RECT 65.420 132.610 65.680 132.930 ;
        RECT 69.620 131.480 69.760 134.650 ;
        RECT 68.700 131.340 69.760 131.480 ;
        RECT 68.700 129.870 68.840 131.340 ;
        RECT 66.340 129.550 66.600 129.870 ;
        RECT 68.640 129.550 68.900 129.870 ;
        RECT 62.200 126.830 62.460 127.150 ;
        RECT 60.820 126.490 61.080 126.810 ;
        RECT 57.140 126.150 57.400 126.470 ;
        RECT 52.080 120.710 52.340 121.030 ;
        RECT 59.900 120.710 60.160 121.030 ;
        RECT 60.360 120.710 60.620 121.030 ;
        RECT 61.280 120.940 61.540 121.030 ;
        RECT 60.880 120.800 61.540 120.940 ;
        RECT 52.140 113.890 52.280 120.710 ;
        RECT 58.060 120.370 58.320 120.690 ;
        RECT 53.920 120.030 54.180 120.350 ;
        RECT 53.980 115.590 54.120 120.030 ;
        RECT 53.920 115.270 54.180 115.590 ;
        RECT 52.080 113.570 52.340 113.890 ;
        RECT 58.120 113.210 58.260 120.370 ;
        RECT 59.440 118.330 59.700 118.650 ;
        RECT 59.500 116.610 59.640 118.330 ;
        RECT 59.960 116.610 60.100 120.710 ;
        RECT 59.440 116.290 59.700 116.610 ;
        RECT 59.900 116.290 60.160 116.610 ;
        RECT 58.520 114.930 58.780 115.250 ;
        RECT 58.580 113.890 58.720 114.930 ;
        RECT 60.420 113.890 60.560 120.710 ;
        RECT 60.880 117.630 61.020 120.800 ;
        RECT 61.280 120.710 61.540 120.800 ;
        RECT 66.400 118.650 66.540 129.550 ;
        RECT 65.880 118.330 66.140 118.650 ;
        RECT 66.340 118.330 66.600 118.650 ;
        RECT 69.100 118.330 69.360 118.650 ;
        RECT 60.820 117.310 61.080 117.630 ;
        RECT 60.880 115.590 61.020 117.310 ;
        RECT 65.940 116.610 66.080 118.330 ;
        RECT 65.880 116.290 66.140 116.610 ;
        RECT 60.820 115.270 61.080 115.590 ;
        RECT 64.040 115.270 64.300 115.590 ;
        RECT 65.420 115.270 65.680 115.590 ;
        RECT 58.520 113.570 58.780 113.890 ;
        RECT 60.360 113.570 60.620 113.890 ;
        RECT 58.060 112.890 58.320 113.210 ;
        RECT 60.820 112.890 61.080 113.210 ;
        RECT 62.200 112.890 62.460 113.210 ;
        RECT 58.120 110.470 58.260 112.890 ;
        RECT 57.200 110.330 58.260 110.470 ;
        RECT 56.680 109.830 56.940 110.150 ;
        RECT 56.740 108.450 56.880 109.830 ;
        RECT 57.200 109.470 57.340 110.330 ;
        RECT 60.880 109.470 61.020 112.890 ;
        RECT 62.260 110.830 62.400 112.890 ;
        RECT 64.100 112.870 64.240 115.270 ;
        RECT 64.960 114.930 65.220 115.250 ;
        RECT 64.040 112.550 64.300 112.870 ;
        RECT 62.200 110.510 62.460 110.830 ;
        RECT 57.140 109.150 57.400 109.470 ;
        RECT 58.980 109.150 59.240 109.470 ;
        RECT 60.820 109.150 61.080 109.470 ;
        RECT 61.280 109.150 61.540 109.470 ;
        RECT 57.200 108.450 57.340 109.150 ;
        RECT 56.680 108.130 56.940 108.450 ;
        RECT 57.140 108.130 57.400 108.450 ;
        RECT 55.760 107.450 56.020 107.770 ;
        RECT 55.820 105.730 55.960 107.450 ;
        RECT 59.040 107.430 59.180 109.150 ;
        RECT 58.980 107.110 59.240 107.430 ;
        RECT 59.900 107.110 60.160 107.430 ;
        RECT 56.220 106.770 56.480 107.090 ;
        RECT 51.160 105.410 51.420 105.730 ;
        RECT 55.760 105.410 56.020 105.730 ;
        RECT 49.320 105.070 49.580 105.390 ;
        RECT 48.860 104.050 49.120 104.370 ;
        RECT 48.400 102.350 48.660 102.670 ;
        RECT 46.100 101.670 46.360 101.990 ;
        RECT 47.480 101.670 47.740 101.990 ;
        RECT 44.260 100.990 44.520 101.310 ;
        RECT 44.320 93.830 44.460 100.990 ;
        RECT 46.160 97.570 46.300 101.670 ;
        RECT 47.540 100.290 47.680 101.670 ;
        RECT 47.480 99.970 47.740 100.290 ;
        RECT 46.100 97.250 46.360 97.570 ;
        RECT 44.260 93.510 44.520 93.830 ;
        RECT 47.540 93.490 47.680 99.970 ;
        RECT 47.940 98.610 48.200 98.930 ;
        RECT 48.000 95.870 48.140 98.610 ;
        RECT 48.460 96.890 48.600 102.350 ;
        RECT 48.920 101.310 49.060 104.050 ;
        RECT 49.380 103.010 49.520 105.070 ;
        RECT 49.320 102.690 49.580 103.010 ;
        RECT 48.860 100.990 49.120 101.310 ;
        RECT 48.920 97.230 49.060 100.990 ;
        RECT 49.320 98.950 49.580 99.270 ;
        RECT 48.860 96.910 49.120 97.230 ;
        RECT 48.400 96.570 48.660 96.890 ;
        RECT 49.380 96.210 49.520 98.950 ;
        RECT 49.320 95.890 49.580 96.210 ;
        RECT 47.940 95.550 48.200 95.870 ;
        RECT 48.000 94.170 48.140 95.550 ;
        RECT 47.940 93.850 48.200 94.170 ;
        RECT 47.480 93.170 47.740 93.490 ;
        RECT 48.000 91.110 48.140 93.850 ;
        RECT 47.940 90.790 48.200 91.110 ;
        RECT 49.380 90.430 49.520 95.890 ;
        RECT 50.700 93.850 50.960 94.170 ;
        RECT 43.400 90.200 44.000 90.340 ;
        RECT 43.400 83.630 43.540 90.200 ;
        RECT 49.320 90.110 49.580 90.430 ;
        RECT 44.720 87.730 44.980 88.050 ;
        RECT 44.780 86.690 44.920 87.730 ;
        RECT 44.260 86.370 44.520 86.690 ;
        RECT 44.720 86.370 44.980 86.690 ;
        RECT 44.320 86.010 44.460 86.370 ;
        RECT 48.860 86.030 49.120 86.350 ;
        RECT 44.260 85.690 44.520 86.010 ;
        RECT 43.340 83.310 43.600 83.630 ;
        RECT 43.400 71.810 43.540 83.310 ;
        RECT 44.320 77.170 44.460 85.690 ;
        RECT 45.640 85.010 45.900 85.330 ;
        RECT 45.180 82.290 45.440 82.610 ;
        RECT 44.720 81.950 44.980 82.270 ;
        RECT 44.780 80.910 44.920 81.950 ;
        RECT 44.720 80.590 44.980 80.910 ;
        RECT 45.240 78.530 45.380 82.290 ;
        RECT 45.180 78.210 45.440 78.530 ;
        RECT 44.260 76.850 44.520 77.170 ;
        RECT 43.800 76.510 44.060 76.830 ;
        RECT 43.860 72.410 44.000 76.510 ;
        RECT 44.260 75.150 44.520 75.470 ;
        RECT 44.320 73.090 44.460 75.150 ;
        RECT 45.180 74.810 45.440 75.130 ;
        RECT 44.720 73.790 44.980 74.110 ;
        RECT 44.260 72.770 44.520 73.090 ;
        RECT 43.800 72.090 44.060 72.410 ;
        RECT 43.400 71.670 44.000 71.810 ;
        RECT 43.340 63.590 43.600 63.910 ;
        RECT 43.400 59.490 43.540 63.590 ;
        RECT 43.860 61.190 44.000 71.670 ;
        RECT 44.320 66.970 44.460 72.770 ;
        RECT 44.780 72.070 44.920 73.790 ;
        RECT 45.240 73.090 45.380 74.810 ;
        RECT 45.180 72.770 45.440 73.090 ;
        RECT 44.720 71.750 44.980 72.070 ;
        RECT 44.260 66.650 44.520 66.970 ;
        RECT 44.780 61.530 44.920 71.750 ;
        RECT 45.700 70.030 45.840 85.010 ;
        RECT 47.940 82.970 48.200 83.290 ;
        RECT 46.560 81.950 46.820 82.270 ;
        RECT 46.620 78.530 46.760 81.950 ;
        RECT 46.560 78.210 46.820 78.530 ;
        RECT 47.480 76.510 47.740 76.830 ;
        RECT 46.560 71.070 46.820 71.390 ;
        RECT 45.640 69.710 45.900 70.030 ;
        RECT 45.700 69.350 45.840 69.710 ;
        RECT 45.640 69.030 45.900 69.350 ;
        RECT 46.620 64.930 46.760 71.070 ;
        RECT 47.540 66.970 47.680 76.510 ;
        RECT 48.000 75.470 48.140 82.970 ;
        RECT 48.920 81.250 49.060 86.030 ;
        RECT 49.380 85.670 49.520 90.110 ;
        RECT 49.320 85.350 49.580 85.670 ;
        RECT 49.380 83.290 49.520 85.350 ;
        RECT 49.320 82.970 49.580 83.290 ;
        RECT 48.860 80.930 49.120 81.250 ;
        RECT 47.940 75.150 48.200 75.470 ;
        RECT 48.000 72.410 48.140 75.150 ;
        RECT 47.940 72.090 48.200 72.410 ;
        RECT 48.000 68.920 48.140 72.090 ;
        RECT 49.380 72.070 49.520 82.970 ;
        RECT 49.780 81.950 50.040 82.270 ;
        RECT 49.840 81.250 49.980 81.950 ;
        RECT 49.780 80.930 50.040 81.250 ;
        RECT 50.760 77.850 50.900 93.850 ;
        RECT 50.700 77.530 50.960 77.850 ;
        RECT 50.240 77.190 50.500 77.510 ;
        RECT 50.300 75.810 50.440 77.190 ;
        RECT 50.240 75.490 50.500 75.810 ;
        RECT 49.320 71.750 49.580 72.070 ;
        RECT 49.780 69.370 50.040 69.690 ;
        RECT 48.400 68.920 48.660 69.010 ;
        RECT 48.000 68.780 48.660 68.920 ;
        RECT 48.400 68.690 48.660 68.780 ;
        RECT 47.480 66.650 47.740 66.970 ;
        RECT 49.320 65.970 49.580 66.290 ;
        RECT 49.380 64.930 49.520 65.970 ;
        RECT 46.560 64.610 46.820 64.930 ;
        RECT 49.320 64.610 49.580 64.930 ;
        RECT 45.180 63.250 45.440 63.570 ;
        RECT 44.720 61.210 44.980 61.530 ;
        RECT 43.800 60.870 44.060 61.190 ;
        RECT 44.720 60.190 44.980 60.510 ;
        RECT 43.340 59.170 43.600 59.490 ;
        RECT 43.400 55.750 43.540 59.170 ;
        RECT 44.780 58.470 44.920 60.190 ;
        RECT 45.240 59.490 45.380 63.250 ;
        RECT 47.480 60.530 47.740 60.850 ;
        RECT 47.540 59.490 47.680 60.530 ;
        RECT 45.180 59.170 45.440 59.490 ;
        RECT 47.480 59.170 47.740 59.490 ;
        RECT 44.720 58.150 44.980 58.470 ;
        RECT 47.940 58.150 48.200 58.470 ;
        RECT 43.340 55.430 43.600 55.750 ;
        RECT 47.480 55.090 47.740 55.410 ;
        RECT 47.540 53.710 47.680 55.090 ;
        RECT 47.480 53.390 47.740 53.710 ;
        RECT 45.640 52.710 45.900 53.030 ;
        RECT 47.020 52.710 47.280 53.030 ;
        RECT 44.720 52.030 44.980 52.350 ;
        RECT 43.800 49.990 44.060 50.310 ;
        RECT 42.880 46.930 43.140 47.250 ;
        RECT 42.940 45.210 43.080 46.930 ;
        RECT 42.880 44.890 43.140 45.210 ;
        RECT 43.340 38.770 43.600 39.090 ;
        RECT 43.400 36.710 43.540 38.770 ;
        RECT 43.340 36.390 43.600 36.710 ;
        RECT 42.880 35.710 43.140 36.030 ;
        RECT 42.940 28.290 43.080 35.710 ;
        RECT 43.400 34.330 43.540 36.390 ;
        RECT 43.340 34.010 43.600 34.330 ;
        RECT 43.340 31.970 43.600 32.290 ;
        RECT 43.400 28.970 43.540 31.970 ;
        RECT 43.860 29.570 44.000 49.990 ;
        RECT 44.780 48.270 44.920 52.030 ;
        RECT 44.720 47.950 44.980 48.270 ;
        RECT 45.180 45.570 45.440 45.890 ;
        RECT 45.240 42.490 45.380 45.570 ;
        RECT 44.260 42.170 44.520 42.490 ;
        RECT 45.180 42.170 45.440 42.490 ;
        RECT 44.320 39.430 44.460 42.170 ;
        RECT 45.240 40.450 45.380 42.170 ;
        RECT 45.180 40.130 45.440 40.450 ;
        RECT 44.260 39.110 44.520 39.430 ;
        RECT 44.320 31.610 44.460 39.110 ;
        RECT 45.240 37.730 45.380 40.130 ;
        RECT 45.180 37.410 45.440 37.730 ;
        RECT 45.240 36.030 45.380 37.410 ;
        RECT 44.720 35.710 44.980 36.030 ;
        RECT 45.180 35.710 45.440 36.030 ;
        RECT 44.260 31.290 44.520 31.610 ;
        RECT 44.780 30.930 44.920 35.710 ;
        RECT 45.240 31.610 45.380 35.710 ;
        RECT 45.180 31.290 45.440 31.610 ;
        RECT 44.720 30.610 44.980 30.930 ;
        RECT 43.800 29.250 44.060 29.570 ;
        RECT 43.400 28.830 44.000 28.970 ;
        RECT 43.860 28.550 44.000 28.830 ;
        RECT 44.260 28.570 44.520 28.890 ;
        RECT 42.940 28.210 43.540 28.290 ;
        RECT 43.800 28.230 44.060 28.550 ;
        RECT 42.940 28.150 43.600 28.210 ;
        RECT 43.340 27.890 43.600 28.150 ;
        RECT 43.860 21.070 44.000 28.230 ;
        RECT 44.320 22.430 44.460 28.570 ;
        RECT 44.780 27.870 44.920 30.610 ;
        RECT 44.720 27.550 44.980 27.870 ;
        RECT 44.720 25.850 44.980 26.170 ;
        RECT 44.780 23.790 44.920 25.850 ;
        RECT 44.720 23.470 44.980 23.790 ;
        RECT 44.260 22.110 44.520 22.430 ;
        RECT 43.800 20.750 44.060 21.070 ;
        RECT 42.420 19.730 42.680 20.050 ;
        RECT 42.880 17.350 43.140 17.670 ;
        RECT 42.940 13.250 43.080 17.350 ;
        RECT 45.700 14.270 45.840 52.710 ;
        RECT 47.080 51.330 47.220 52.710 ;
        RECT 47.540 51.330 47.680 53.390 ;
        RECT 48.000 53.030 48.140 58.150 ;
        RECT 49.840 56.770 49.980 69.370 ;
        RECT 50.760 63.230 50.900 77.530 ;
        RECT 51.220 70.370 51.360 105.410 ;
        RECT 56.280 103.010 56.420 106.770 ;
        RECT 58.060 106.430 58.320 106.750 ;
        RECT 57.600 105.410 57.860 105.730 ;
        RECT 56.220 102.690 56.480 103.010 ;
        RECT 57.660 102.330 57.800 105.410 ;
        RECT 57.600 102.010 57.860 102.330 ;
        RECT 58.120 101.730 58.260 106.430 ;
        RECT 59.040 104.710 59.180 107.110 ;
        RECT 58.980 104.390 59.240 104.710 ;
        RECT 59.440 102.690 59.700 103.010 ;
        RECT 58.980 102.350 59.240 102.670 ;
        RECT 57.660 101.590 58.260 101.730 ;
        RECT 57.660 101.310 57.800 101.590 ;
        RECT 53.920 100.990 54.180 101.310 ;
        RECT 57.600 100.990 57.860 101.310 ;
        RECT 53.980 99.610 54.120 100.990 ;
        RECT 53.920 99.290 54.180 99.610 ;
        RECT 57.140 98.950 57.400 99.270 ;
        RECT 57.200 97.570 57.340 98.950 ;
        RECT 57.140 97.250 57.400 97.570 ;
        RECT 53.920 93.510 54.180 93.830 ;
        RECT 53.980 92.130 54.120 93.510 ;
        RECT 53.920 91.810 54.180 92.130 ;
        RECT 57.200 84.990 57.340 97.250 ;
        RECT 57.660 94.170 57.800 100.990 ;
        RECT 59.040 99.270 59.180 102.350 ;
        RECT 59.500 99.270 59.640 102.690 ;
        RECT 59.960 102.670 60.100 107.110 ;
        RECT 60.820 106.770 61.080 107.090 ;
        RECT 60.880 105.390 61.020 106.770 ;
        RECT 61.340 105.730 61.480 109.150 ;
        RECT 61.740 107.450 62.000 107.770 ;
        RECT 61.280 105.410 61.540 105.730 ;
        RECT 60.820 105.070 61.080 105.390 ;
        RECT 60.820 104.390 61.080 104.710 ;
        RECT 61.800 104.450 61.940 107.450 ;
        RECT 62.260 107.170 62.400 110.510 ;
        RECT 62.660 109.830 62.920 110.150 ;
        RECT 62.720 108.450 62.860 109.830 ;
        RECT 63.120 109.490 63.380 109.810 ;
        RECT 62.660 108.130 62.920 108.450 ;
        RECT 63.180 108.110 63.320 109.490 ;
        RECT 63.120 107.790 63.380 108.110 ;
        RECT 62.260 107.090 62.860 107.170 ;
        RECT 62.260 107.030 62.920 107.090 ;
        RECT 62.660 106.770 62.920 107.030 ;
        RECT 64.100 105.390 64.240 112.550 ;
        RECT 65.020 110.150 65.160 114.930 ;
        RECT 64.960 109.830 65.220 110.150 ;
        RECT 65.480 108.110 65.620 115.270 ;
        RECT 69.160 110.150 69.300 118.330 ;
        RECT 80.600 112.890 80.860 113.210 ;
        RECT 71.400 111.870 71.660 112.190 ;
        RECT 69.100 109.830 69.360 110.150 ;
        RECT 66.800 109.490 67.060 109.810 ;
        RECT 66.340 109.150 66.600 109.470 ;
        RECT 65.420 107.790 65.680 108.110 ;
        RECT 66.400 107.430 66.540 109.150 ;
        RECT 66.340 107.110 66.600 107.430 ;
        RECT 64.500 106.770 64.760 107.090 ;
        RECT 64.560 105.730 64.700 106.770 ;
        RECT 66.860 106.750 67.000 109.490 ;
        RECT 67.260 107.450 67.520 107.770 ;
        RECT 66.800 106.430 67.060 106.750 ;
        RECT 67.320 105.730 67.460 107.450 ;
        RECT 70.940 106.770 71.200 107.090 ;
        RECT 64.500 105.410 64.760 105.730 ;
        RECT 65.420 105.410 65.680 105.730 ;
        RECT 67.260 105.410 67.520 105.730 ;
        RECT 64.040 105.070 64.300 105.390 ;
        RECT 59.900 102.350 60.160 102.670 ;
        RECT 59.900 100.990 60.160 101.310 ;
        RECT 58.980 98.950 59.240 99.270 ;
        RECT 59.440 98.950 59.700 99.270 ;
        RECT 58.520 98.270 58.780 98.590 ;
        RECT 58.060 97.250 58.320 97.570 ;
        RECT 57.600 93.850 57.860 94.170 ;
        RECT 58.120 85.670 58.260 97.250 ;
        RECT 58.580 96.890 58.720 98.270 ;
        RECT 59.960 97.570 60.100 100.990 ;
        RECT 60.360 99.630 60.620 99.950 ;
        RECT 59.900 97.250 60.160 97.570 ;
        RECT 58.520 96.570 58.780 96.890 ;
        RECT 58.580 86.010 58.720 96.570 ;
        RECT 60.420 96.550 60.560 99.630 ;
        RECT 60.360 96.230 60.620 96.550 ;
        RECT 60.360 93.510 60.620 93.830 ;
        RECT 59.440 93.060 59.700 93.150 ;
        RECT 59.440 92.920 60.100 93.060 ;
        RECT 59.440 92.830 59.700 92.920 ;
        RECT 58.970 91.955 59.250 92.325 ;
        RECT 59.040 91.790 59.180 91.955 ;
        RECT 58.980 91.470 59.240 91.790 ;
        RECT 59.440 90.110 59.700 90.430 ;
        RECT 59.500 88.050 59.640 90.110 ;
        RECT 59.440 87.730 59.700 88.050 ;
        RECT 58.520 85.690 58.780 86.010 ;
        RECT 58.980 85.690 59.240 86.010 ;
        RECT 58.060 85.350 58.320 85.670 ;
        RECT 57.140 84.670 57.400 84.990 ;
        RECT 58.120 83.370 58.260 85.350 ;
        RECT 57.660 83.230 58.260 83.370 ;
        RECT 57.660 82.950 57.800 83.230 ;
        RECT 57.600 82.630 57.860 82.950 ;
        RECT 58.520 82.630 58.780 82.950 ;
        RECT 58.060 81.950 58.320 82.270 ;
        RECT 51.620 76.510 51.880 76.830 ;
        RECT 51.160 70.050 51.420 70.370 ;
        RECT 51.220 66.630 51.360 70.050 ;
        RECT 51.160 66.310 51.420 66.630 ;
        RECT 51.160 63.930 51.420 64.250 ;
        RECT 50.700 62.910 50.960 63.230 ;
        RECT 50.240 60.870 50.500 61.190 ;
        RECT 50.300 59.490 50.440 60.870 ;
        RECT 50.240 59.170 50.500 59.490 ;
        RECT 49.780 56.450 50.040 56.770 ;
        RECT 50.300 56.090 50.440 59.170 ;
        RECT 50.240 55.770 50.500 56.090 ;
        RECT 51.220 53.030 51.360 63.930 ;
        RECT 51.680 62.210 51.820 76.510 ;
        RECT 56.220 74.810 56.480 75.130 ;
        RECT 56.280 72.070 56.420 74.810 ;
        RECT 58.120 72.070 58.260 81.950 ;
        RECT 58.580 80.570 58.720 82.630 ;
        RECT 59.040 81.250 59.180 85.690 ;
        RECT 58.980 80.930 59.240 81.250 ;
        RECT 58.520 80.250 58.780 80.570 ;
        RECT 58.580 77.170 58.720 80.250 ;
        RECT 58.520 76.850 58.780 77.170 ;
        RECT 59.500 75.130 59.640 87.730 ;
        RECT 59.960 82.950 60.100 92.920 ;
        RECT 60.420 91.450 60.560 93.510 ;
        RECT 60.880 93.490 61.020 104.390 ;
        RECT 61.800 104.310 62.400 104.450 ;
        RECT 62.260 104.030 62.400 104.310 ;
        RECT 61.280 103.710 61.540 104.030 ;
        RECT 62.200 103.710 62.460 104.030 ;
        RECT 61.340 102.330 61.480 103.710 ;
        RECT 61.280 102.010 61.540 102.330 ;
        RECT 61.340 96.890 61.480 102.010 ;
        RECT 61.280 96.570 61.540 96.890 ;
        RECT 61.340 94.850 61.480 96.570 ;
        RECT 62.660 96.230 62.920 96.550 ;
        RECT 65.480 96.405 65.620 105.410 ;
        RECT 67.720 105.070 67.980 105.390 ;
        RECT 67.260 102.010 67.520 102.330 ;
        RECT 65.880 101.670 66.140 101.990 ;
        RECT 65.940 101.310 66.080 101.670 ;
        RECT 67.320 101.310 67.460 102.010 ;
        RECT 65.880 100.990 66.140 101.310 ;
        RECT 67.260 100.990 67.520 101.310 ;
        RECT 61.280 94.530 61.540 94.850 ;
        RECT 61.340 94.110 62.400 94.250 ;
        RECT 60.820 93.170 61.080 93.490 ;
        RECT 60.360 91.130 60.620 91.450 ;
        RECT 61.340 91.110 61.480 94.110 ;
        RECT 61.740 93.510 62.000 93.830 ;
        RECT 61.280 90.790 61.540 91.110 ;
        RECT 61.800 90.430 61.940 93.510 ;
        RECT 62.260 93.150 62.400 94.110 ;
        RECT 62.720 93.830 62.860 96.230 ;
        RECT 64.960 95.890 65.220 96.210 ;
        RECT 65.410 96.035 65.690 96.405 ;
        RECT 65.020 93.830 65.160 95.890 ;
        RECT 62.660 93.510 62.920 93.830 ;
        RECT 64.960 93.510 65.220 93.830 ;
        RECT 62.200 92.830 62.460 93.150 ;
        RECT 62.720 91.450 62.860 93.510 ;
        RECT 64.500 93.170 64.760 93.490 ;
        RECT 62.200 91.130 62.460 91.450 ;
        RECT 62.660 91.130 62.920 91.450 ;
        RECT 64.040 91.130 64.300 91.450 ;
        RECT 61.740 90.110 62.000 90.430 ;
        RECT 60.820 88.410 61.080 88.730 ;
        RECT 60.880 86.690 61.020 88.410 ;
        RECT 62.260 87.710 62.400 91.130 ;
        RECT 62.720 88.050 62.860 91.130 ;
        RECT 64.100 90.430 64.240 91.130 ;
        RECT 64.040 90.110 64.300 90.430 ;
        RECT 62.660 87.960 62.920 88.050 ;
        RECT 62.660 87.820 63.320 87.960 ;
        RECT 62.660 87.730 62.920 87.820 ;
        RECT 62.200 87.390 62.460 87.710 ;
        RECT 60.820 86.370 61.080 86.690 ;
        RECT 60.880 86.010 61.020 86.370 ;
        RECT 61.740 86.030 62.000 86.350 ;
        RECT 60.820 85.690 61.080 86.010 ;
        RECT 60.820 84.670 61.080 84.990 ;
        RECT 60.360 83.650 60.620 83.970 ;
        RECT 59.900 82.630 60.160 82.950 ;
        RECT 59.440 74.810 59.700 75.130 ;
        RECT 59.440 74.130 59.700 74.450 ;
        RECT 59.500 72.750 59.640 74.130 ;
        RECT 59.440 72.430 59.700 72.750 ;
        RECT 56.220 71.750 56.480 72.070 ;
        RECT 58.060 71.750 58.320 72.070 ;
        RECT 56.280 69.690 56.420 71.750 ;
        RECT 59.500 70.370 59.640 72.430 ;
        RECT 59.440 70.050 59.700 70.370 ;
        RECT 58.520 69.710 58.780 70.030 ;
        RECT 56.220 69.370 56.480 69.690 ;
        RECT 56.280 66.970 56.420 69.370 ;
        RECT 56.220 66.650 56.480 66.970 ;
        RECT 57.600 66.310 57.860 66.630 ;
        RECT 56.680 63.590 56.940 63.910 ;
        RECT 52.540 62.910 52.800 63.230 ;
        RECT 51.620 61.890 51.880 62.210 ;
        RECT 52.080 60.190 52.340 60.510 ;
        RECT 52.140 59.150 52.280 60.190 ;
        RECT 52.080 58.830 52.340 59.150 ;
        RECT 52.600 56.090 52.740 62.910 ;
        RECT 56.740 58.810 56.880 63.590 ;
        RECT 57.660 60.850 57.800 66.310 ;
        RECT 58.060 60.870 58.320 61.190 ;
        RECT 57.600 60.530 57.860 60.850 ;
        RECT 58.120 58.810 58.260 60.870 ;
        RECT 56.680 58.490 56.940 58.810 ;
        RECT 58.060 58.490 58.320 58.810 ;
        RECT 58.580 58.720 58.720 69.710 ;
        RECT 58.980 68.350 59.240 68.670 ;
        RECT 59.040 66.290 59.180 68.350 ;
        RECT 58.980 65.970 59.240 66.290 ;
        RECT 59.440 65.630 59.700 65.950 ;
        RECT 59.500 64.930 59.640 65.630 ;
        RECT 59.440 64.610 59.700 64.930 ;
        RECT 59.960 61.530 60.100 82.630 ;
        RECT 60.420 79.550 60.560 83.650 ;
        RECT 60.880 82.950 61.020 84.670 ;
        RECT 61.800 83.970 61.940 86.030 ;
        RECT 62.660 85.690 62.920 86.010 ;
        RECT 61.740 83.650 62.000 83.970 ;
        RECT 62.720 82.950 62.860 85.690 ;
        RECT 60.820 82.630 61.080 82.950 ;
        RECT 62.660 82.860 62.920 82.950 ;
        RECT 62.260 82.720 62.920 82.860 ;
        RECT 61.280 80.930 61.540 81.250 ;
        RECT 60.360 79.230 60.620 79.550 ;
        RECT 60.420 78.530 60.560 79.230 ;
        RECT 60.360 78.210 60.620 78.530 ;
        RECT 61.340 77.170 61.480 80.930 ;
        RECT 62.260 79.890 62.400 82.720 ;
        RECT 62.660 82.630 62.920 82.720 ;
        RECT 62.660 81.950 62.920 82.270 ;
        RECT 62.720 81.250 62.860 81.950 ;
        RECT 62.660 80.930 62.920 81.250 ;
        RECT 62.200 79.570 62.460 79.890 ;
        RECT 62.190 79.290 62.470 79.405 ;
        RECT 61.800 79.150 62.470 79.290 ;
        RECT 61.280 76.850 61.540 77.170 ;
        RECT 61.280 71.750 61.540 72.070 ;
        RECT 60.810 69.515 61.090 69.885 ;
        RECT 60.820 69.370 61.080 69.515 ;
        RECT 61.340 69.205 61.480 71.750 ;
        RECT 61.270 68.835 61.550 69.205 ;
        RECT 60.360 66.650 60.620 66.970 ;
        RECT 59.900 61.210 60.160 61.530 ;
        RECT 60.420 61.190 60.560 66.650 ;
        RECT 60.820 63.930 61.080 64.250 ;
        RECT 60.360 60.870 60.620 61.190 ;
        RECT 59.900 60.530 60.160 60.850 ;
        RECT 58.980 60.190 59.240 60.510 ;
        RECT 59.440 60.190 59.700 60.510 ;
        RECT 59.040 59.490 59.180 60.190 ;
        RECT 58.980 59.170 59.240 59.490 ;
        RECT 59.500 59.150 59.640 60.190 ;
        RECT 59.440 58.830 59.700 59.150 ;
        RECT 58.980 58.720 59.240 58.810 ;
        RECT 58.580 58.580 59.240 58.720 ;
        RECT 58.980 58.490 59.240 58.580 ;
        RECT 57.600 56.110 57.860 56.430 ;
        RECT 52.540 55.770 52.800 56.090 ;
        RECT 56.680 55.430 56.940 55.750 ;
        RECT 52.540 54.750 52.800 55.070 ;
        RECT 52.600 53.030 52.740 54.750 ;
        RECT 47.940 52.710 48.200 53.030 ;
        RECT 51.160 52.710 51.420 53.030 ;
        RECT 52.540 52.710 52.800 53.030 ;
        RECT 47.020 51.010 47.280 51.330 ;
        RECT 47.480 51.010 47.740 51.330 ;
        RECT 46.100 49.650 46.360 49.970 ;
        RECT 46.160 47.930 46.300 49.650 ;
        RECT 46.100 47.610 46.360 47.930 ;
        RECT 46.160 42.490 46.300 47.610 ;
        RECT 48.000 46.910 48.140 52.710 ;
        RECT 50.700 49.650 50.960 49.970 ;
        RECT 50.760 48.610 50.900 49.650 ;
        RECT 50.700 48.290 50.960 48.610 ;
        RECT 51.220 47.250 51.360 52.710 ;
        RECT 52.600 51.330 52.740 52.710 ;
        RECT 53.000 52.030 53.260 52.350 ;
        RECT 52.540 51.010 52.800 51.330 ;
        RECT 53.060 48.610 53.200 52.030 ;
        RECT 56.740 51.330 56.880 55.430 ;
        RECT 56.680 51.010 56.940 51.330 ;
        RECT 53.460 49.990 53.720 50.310 ;
        RECT 53.520 48.610 53.660 49.990 ;
        RECT 54.380 49.310 54.640 49.630 ;
        RECT 53.000 48.290 53.260 48.610 ;
        RECT 53.460 48.290 53.720 48.610 ;
        RECT 53.000 47.270 53.260 47.590 ;
        RECT 51.160 46.930 51.420 47.250 ;
        RECT 47.940 46.590 48.200 46.910 ;
        RECT 47.940 44.890 48.200 45.210 ;
        RECT 48.000 42.830 48.140 44.890 ;
        RECT 48.400 44.210 48.660 44.530 ;
        RECT 47.940 42.510 48.200 42.830 ;
        RECT 46.100 42.170 46.360 42.490 ;
        RECT 47.480 38.770 47.740 39.090 ;
        RECT 46.560 38.430 46.820 38.750 ;
        RECT 46.620 37.390 46.760 38.430 ;
        RECT 47.020 37.410 47.280 37.730 ;
        RECT 46.560 37.070 46.820 37.390 ;
        RECT 47.080 31.610 47.220 37.410 ;
        RECT 47.540 35.010 47.680 38.770 ;
        RECT 48.460 38.750 48.600 44.210 ;
        RECT 49.320 43.870 49.580 44.190 ;
        RECT 48.860 42.170 49.120 42.490 ;
        RECT 48.920 39.430 49.060 42.170 ;
        RECT 49.380 41.810 49.520 43.870 ;
        RECT 52.540 41.830 52.800 42.150 ;
        RECT 49.320 41.490 49.580 41.810 ;
        RECT 48.860 39.110 49.120 39.430 ;
        RECT 48.400 38.430 48.660 38.750 ;
        RECT 49.380 37.050 49.520 41.490 ;
        RECT 50.700 38.770 50.960 39.090 ;
        RECT 49.320 36.730 49.580 37.050 ;
        RECT 50.760 36.710 50.900 38.770 ;
        RECT 50.700 36.390 50.960 36.710 ;
        RECT 47.480 34.690 47.740 35.010 ;
        RECT 50.240 32.990 50.500 33.310 ;
        RECT 47.940 31.630 48.200 31.950 ;
        RECT 47.020 31.290 47.280 31.610 ;
        RECT 48.000 28.550 48.140 31.630 ;
        RECT 49.320 31.290 49.580 31.610 ;
        RECT 49.380 29.570 49.520 31.290 ;
        RECT 49.320 29.250 49.580 29.570 ;
        RECT 46.100 28.230 46.360 28.550 ;
        RECT 47.940 28.230 48.200 28.550 ;
        RECT 46.160 26.170 46.300 28.230 ;
        RECT 46.100 25.850 46.360 26.170 ;
        RECT 48.000 25.570 48.140 28.230 ;
        RECT 49.780 27.890 50.040 28.210 ;
        RECT 46.160 25.430 48.140 25.570 ;
        RECT 48.400 25.510 48.660 25.830 ;
        RECT 46.160 23.110 46.300 25.430 ;
        RECT 47.940 24.890 48.200 25.150 ;
        RECT 47.540 24.830 48.200 24.890 ;
        RECT 47.540 24.750 48.140 24.830 ;
        RECT 46.100 22.790 46.360 23.110 ;
        RECT 47.540 22.430 47.680 24.750 ;
        RECT 48.460 24.210 48.600 25.510 ;
        RECT 48.000 24.070 48.600 24.210 ;
        RECT 48.000 22.430 48.140 24.070 ;
        RECT 48.400 22.450 48.660 22.770 ;
        RECT 47.480 22.110 47.740 22.430 ;
        RECT 47.940 22.110 48.200 22.430 ;
        RECT 45.640 13.950 45.900 14.270 ;
        RECT 42.880 12.930 43.140 13.250 ;
        RECT 47.540 12.570 47.680 22.110 ;
        RECT 48.000 21.070 48.140 22.110 ;
        RECT 48.460 21.410 48.600 22.450 ;
        RECT 48.400 21.090 48.660 21.410 ;
        RECT 47.940 20.750 48.200 21.070 ;
        RECT 48.000 17.670 48.140 20.750 ;
        RECT 48.860 20.070 49.120 20.390 ;
        RECT 48.400 19.730 48.660 20.050 ;
        RECT 48.460 17.670 48.600 19.730 ;
        RECT 48.920 17.670 49.060 20.070 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 48.400 17.350 48.660 17.670 ;
        RECT 48.860 17.350 49.120 17.670 ;
        RECT 49.320 17.350 49.580 17.670 ;
        RECT 47.940 16.670 48.200 16.990 ;
        RECT 48.000 15.290 48.140 16.670 ;
        RECT 49.380 15.970 49.520 17.350 ;
        RECT 49.320 15.650 49.580 15.970 ;
        RECT 47.940 14.970 48.200 15.290 ;
        RECT 47.480 12.250 47.740 12.570 ;
        RECT 49.840 12.230 49.980 27.890 ;
        RECT 50.300 20.730 50.440 32.990 ;
        RECT 50.760 30.590 50.900 36.390 ;
        RECT 52.600 36.030 52.740 41.830 ;
        RECT 53.060 36.370 53.200 47.270 ;
        RECT 54.440 45.890 54.580 49.310 ;
        RECT 54.380 45.570 54.640 45.890 ;
        RECT 55.300 45.570 55.560 45.890 ;
        RECT 55.360 44.870 55.500 45.570 ;
        RECT 55.300 44.550 55.560 44.870 ;
        RECT 57.140 44.550 57.400 44.870 ;
        RECT 54.840 44.210 55.100 44.530 ;
        RECT 54.900 42.490 55.040 44.210 ;
        RECT 53.460 42.170 53.720 42.490 ;
        RECT 54.840 42.170 55.100 42.490 ;
        RECT 53.520 40.450 53.660 42.170 ;
        RECT 53.460 40.130 53.720 40.450 ;
        RECT 53.520 36.710 53.660 40.130 ;
        RECT 54.380 38.430 54.640 38.750 ;
        RECT 54.440 37.050 54.580 38.430 ;
        RECT 54.900 37.050 55.040 42.170 ;
        RECT 56.680 37.410 56.940 37.730 ;
        RECT 54.380 36.730 54.640 37.050 ;
        RECT 54.840 36.730 55.100 37.050 ;
        RECT 53.460 36.390 53.720 36.710 ;
        RECT 53.000 36.050 53.260 36.370 ;
        RECT 52.540 35.710 52.800 36.030 ;
        RECT 50.700 30.270 50.960 30.590 ;
        RECT 51.160 30.270 51.420 30.590 ;
        RECT 50.760 28.890 50.900 30.270 ;
        RECT 50.700 28.570 50.960 28.890 ;
        RECT 50.760 26.510 50.900 28.570 ;
        RECT 51.220 28.210 51.360 30.270 ;
        RECT 51.160 27.890 51.420 28.210 ;
        RECT 52.080 27.890 52.340 28.210 ;
        RECT 50.700 26.190 50.960 26.510 ;
        RECT 50.240 20.410 50.500 20.730 ;
        RECT 50.300 18.690 50.440 20.410 ;
        RECT 50.240 18.370 50.500 18.690 ;
        RECT 50.300 16.990 50.440 18.370 ;
        RECT 50.760 17.670 50.900 26.190 ;
        RECT 52.140 25.490 52.280 27.890 ;
        RECT 52.600 27.870 52.740 35.710 ;
        RECT 54.440 34.330 54.580 36.730 ;
        RECT 54.380 34.010 54.640 34.330 ;
        RECT 52.540 27.550 52.800 27.870 ;
        RECT 52.600 26.080 52.740 27.550 ;
        RECT 53.000 26.080 53.260 26.170 ;
        RECT 52.600 25.940 53.260 26.080 ;
        RECT 53.000 25.850 53.260 25.940 ;
        RECT 52.080 25.170 52.340 25.490 ;
        RECT 53.060 20.730 53.200 25.850 ;
        RECT 54.900 25.490 55.040 36.730 ;
        RECT 55.300 35.710 55.560 36.030 ;
        RECT 55.360 28.550 55.500 35.710 ;
        RECT 55.760 33.330 56.020 33.650 ;
        RECT 55.820 32.290 55.960 33.330 ;
        RECT 56.220 32.990 56.480 33.310 ;
        RECT 55.760 31.970 56.020 32.290 ;
        RECT 56.280 31.610 56.420 32.990 ;
        RECT 56.220 31.290 56.480 31.610 ;
        RECT 55.300 28.230 55.560 28.550 ;
        RECT 56.220 28.230 56.480 28.550 ;
        RECT 55.300 27.550 55.560 27.870 ;
        RECT 55.360 26.170 55.500 27.550 ;
        RECT 56.280 26.170 56.420 28.230 ;
        RECT 56.740 26.850 56.880 37.410 ;
        RECT 57.200 30.590 57.340 44.550 ;
        RECT 57.660 39.850 57.800 56.110 ;
        RECT 58.120 53.030 58.260 58.490 ;
        RECT 59.040 56.770 59.180 58.490 ;
        RECT 59.960 58.210 60.100 60.530 ;
        RECT 60.880 58.810 61.020 63.930 ;
        RECT 61.800 63.910 61.940 79.150 ;
        RECT 62.190 79.035 62.470 79.150 ;
        RECT 63.180 77.930 63.320 87.820 ;
        RECT 64.560 86.690 64.700 93.170 ;
        RECT 65.020 91.450 65.160 93.510 ;
        RECT 64.960 91.130 65.220 91.450 ;
        RECT 65.020 89.410 65.160 91.130 ;
        RECT 65.480 91.110 65.620 96.035 ;
        RECT 65.420 90.790 65.680 91.110 ;
        RECT 64.960 89.090 65.220 89.410 ;
        RECT 64.960 88.070 65.220 88.390 ;
        RECT 64.500 86.600 64.760 86.690 ;
        RECT 64.100 86.460 64.760 86.600 ;
        RECT 63.580 80.930 63.840 81.250 ;
        RECT 62.720 77.790 63.320 77.930 ;
        RECT 62.200 76.510 62.460 76.830 ;
        RECT 62.260 75.470 62.400 76.510 ;
        RECT 62.720 75.810 62.860 77.790 ;
        RECT 63.120 77.190 63.380 77.510 ;
        RECT 62.660 75.490 62.920 75.810 ;
        RECT 62.200 75.150 62.460 75.470 ;
        RECT 63.180 75.130 63.320 77.190 ;
        RECT 63.120 74.810 63.380 75.130 ;
        RECT 63.640 74.790 63.780 80.930 ;
        RECT 64.100 75.130 64.240 86.460 ;
        RECT 64.500 86.370 64.760 86.460 ;
        RECT 65.020 86.010 65.160 88.070 ;
        RECT 64.960 85.690 65.220 86.010 ;
        RECT 65.020 82.950 65.160 85.690 ;
        RECT 65.480 83.290 65.620 90.790 ;
        RECT 65.420 82.970 65.680 83.290 ;
        RECT 64.960 82.630 65.220 82.950 ;
        RECT 65.020 80.910 65.160 82.630 ;
        RECT 64.960 80.590 65.220 80.910 ;
        RECT 64.500 79.910 64.760 80.230 ;
        RECT 64.040 74.810 64.300 75.130 ;
        RECT 62.660 74.700 62.920 74.790 ;
        RECT 62.260 74.560 62.920 74.700 ;
        RECT 62.260 70.370 62.400 74.560 ;
        RECT 62.660 74.470 62.920 74.560 ;
        RECT 63.580 74.470 63.840 74.790 ;
        RECT 64.100 74.020 64.240 74.810 ;
        RECT 63.180 73.880 64.240 74.020 ;
        RECT 62.660 72.090 62.920 72.410 ;
        RECT 62.720 71.730 62.860 72.090 ;
        RECT 62.660 71.410 62.920 71.730 ;
        RECT 62.720 70.370 62.860 71.410 ;
        RECT 63.180 70.370 63.320 73.880 ;
        RECT 63.580 72.090 63.840 72.410 ;
        RECT 62.200 70.050 62.460 70.370 ;
        RECT 62.660 70.050 62.920 70.370 ;
        RECT 63.120 70.050 63.380 70.370 ;
        RECT 62.200 69.600 62.460 69.690 ;
        RECT 62.200 69.460 63.320 69.600 ;
        RECT 62.200 69.370 62.460 69.460 ;
        RECT 62.660 68.690 62.920 69.010 ;
        RECT 62.720 66.630 62.860 68.690 ;
        RECT 63.180 66.630 63.320 69.460 ;
        RECT 62.660 66.310 62.920 66.630 ;
        RECT 63.120 66.310 63.380 66.630 ;
        RECT 63.180 64.250 63.320 66.310 ;
        RECT 63.640 66.290 63.780 72.090 ;
        RECT 64.560 72.070 64.700 79.910 ;
        RECT 64.960 79.405 65.220 79.550 ;
        RECT 64.950 79.035 65.230 79.405 ;
        RECT 65.940 78.190 66.080 100.990 ;
        RECT 67.260 99.290 67.520 99.610 ;
        RECT 66.800 98.610 67.060 98.930 ;
        RECT 66.860 97.570 67.000 98.610 ;
        RECT 67.320 98.590 67.460 99.290 ;
        RECT 67.260 98.270 67.520 98.590 ;
        RECT 66.800 97.250 67.060 97.570 ;
        RECT 66.340 96.570 66.600 96.890 ;
        RECT 66.400 94.510 66.540 96.570 ;
        RECT 66.800 96.230 67.060 96.550 ;
        RECT 66.860 94.850 67.000 96.230 ;
        RECT 67.320 94.850 67.460 98.270 ;
        RECT 67.780 96.890 67.920 105.070 ;
        RECT 71.000 104.710 71.140 106.770 ;
        RECT 70.940 104.390 71.200 104.710 ;
        RECT 69.100 103.710 69.360 104.030 ;
        RECT 68.180 102.690 68.440 103.010 ;
        RECT 68.240 96.890 68.380 102.690 ;
        RECT 69.160 102.330 69.300 103.710 ;
        RECT 68.640 102.010 68.900 102.330 ;
        RECT 69.100 102.010 69.360 102.330 ;
        RECT 68.700 97.570 68.840 102.010 ;
        RECT 69.100 100.990 69.360 101.310 ;
        RECT 69.160 99.610 69.300 100.990 ;
        RECT 69.560 99.630 69.820 99.950 ;
        RECT 69.100 99.290 69.360 99.610 ;
        RECT 68.640 97.250 68.900 97.570 ;
        RECT 67.720 96.570 67.980 96.890 ;
        RECT 68.180 96.570 68.440 96.890 ;
        RECT 67.720 95.890 67.980 96.210 ;
        RECT 68.640 95.890 68.900 96.210 ;
        RECT 66.800 94.530 67.060 94.850 ;
        RECT 67.260 94.530 67.520 94.850 ;
        RECT 66.340 94.190 66.600 94.510 ;
        RECT 66.400 85.670 66.540 94.190 ;
        RECT 66.800 93.510 67.060 93.830 ;
        RECT 66.860 86.690 67.000 93.510 ;
        RECT 67.780 92.325 67.920 95.890 ;
        RECT 68.700 93.150 68.840 95.890 ;
        RECT 68.640 92.830 68.900 93.150 ;
        RECT 67.710 91.955 67.990 92.325 ;
        RECT 66.800 86.370 67.060 86.690 ;
        RECT 66.340 85.350 66.600 85.670 ;
        RECT 66.340 84.670 66.600 84.990 ;
        RECT 66.400 81.250 66.540 84.670 ;
        RECT 66.860 82.950 67.000 86.370 ;
        RECT 67.260 85.350 67.520 85.670 ;
        RECT 66.800 82.630 67.060 82.950 ;
        RECT 66.340 80.930 66.600 81.250 ;
        RECT 66.800 79.570 67.060 79.890 ;
        RECT 65.880 77.870 66.140 78.190 ;
        RECT 65.940 77.510 66.080 77.870 ;
        RECT 65.880 77.190 66.140 77.510 ;
        RECT 65.420 75.490 65.680 75.810 ;
        RECT 65.870 75.635 66.150 76.005 ;
        RECT 64.960 72.770 65.220 73.090 ;
        RECT 64.500 71.980 64.760 72.070 ;
        RECT 64.100 71.840 64.760 71.980 ;
        RECT 63.580 65.970 63.840 66.290 ;
        RECT 63.120 63.930 63.380 64.250 ;
        RECT 61.740 63.590 62.000 63.910 ;
        RECT 64.100 63.570 64.240 71.840 ;
        RECT 64.500 71.750 64.760 71.840 ;
        RECT 64.490 68.835 64.770 69.205 ;
        RECT 64.560 68.670 64.700 68.835 ;
        RECT 64.500 68.350 64.760 68.670 ;
        RECT 64.500 66.990 64.760 67.310 ;
        RECT 64.560 64.250 64.700 66.990 ;
        RECT 64.500 63.930 64.760 64.250 ;
        RECT 64.040 63.250 64.300 63.570 ;
        RECT 62.660 61.210 62.920 61.530 ;
        RECT 60.820 58.490 61.080 58.810 ;
        RECT 59.500 58.070 60.100 58.210 ;
        RECT 58.980 56.450 59.240 56.770 ;
        RECT 59.040 55.750 59.180 56.450 ;
        RECT 58.980 55.430 59.240 55.750 ;
        RECT 58.520 54.750 58.780 55.070 ;
        RECT 58.060 52.710 58.320 53.030 ;
        RECT 58.580 50.310 58.720 54.750 ;
        RECT 58.520 49.990 58.780 50.310 ;
        RECT 58.520 44.210 58.780 44.530 ;
        RECT 58.580 42.490 58.720 44.210 ;
        RECT 59.500 42.830 59.640 58.070 ;
        RECT 59.890 57.275 60.170 57.645 ;
        RECT 62.200 57.470 62.460 57.790 ;
        RECT 59.960 56.090 60.100 57.275 ;
        RECT 59.900 55.770 60.160 56.090 ;
        RECT 60.820 55.430 61.080 55.750 ;
        RECT 61.280 55.490 61.540 55.750 ;
        RECT 62.260 55.490 62.400 57.470 ;
        RECT 62.720 55.750 62.860 61.210 ;
        RECT 63.120 59.170 63.380 59.490 ;
        RECT 63.180 55.750 63.320 59.170 ;
        RECT 61.280 55.430 62.400 55.490 ;
        RECT 62.660 55.430 62.920 55.750 ;
        RECT 63.120 55.430 63.380 55.750 ;
        RECT 63.580 55.430 63.840 55.750 ;
        RECT 59.900 55.090 60.160 55.410 ;
        RECT 59.960 52.690 60.100 55.090 ;
        RECT 60.880 54.050 61.020 55.430 ;
        RECT 61.340 55.350 62.400 55.430 ;
        RECT 61.280 54.750 61.540 55.070 ;
        RECT 60.820 53.730 61.080 54.050 ;
        RECT 61.340 53.370 61.480 54.750 ;
        RECT 61.280 53.050 61.540 53.370 ;
        RECT 59.900 52.370 60.160 52.690 ;
        RECT 62.260 52.350 62.400 55.350 ;
        RECT 63.640 55.070 63.780 55.430 ;
        RECT 63.120 54.750 63.380 55.070 ;
        RECT 63.580 54.750 63.840 55.070 ;
        RECT 63.180 53.030 63.320 54.750 ;
        RECT 63.580 53.390 63.840 53.710 ;
        RECT 63.120 52.710 63.380 53.030 ;
        RECT 62.200 52.030 62.460 52.350 ;
        RECT 63.640 49.970 63.780 53.390 ;
        RECT 64.100 53.370 64.240 63.250 ;
        RECT 65.020 63.230 65.160 72.770 ;
        RECT 65.480 72.410 65.620 75.490 ;
        RECT 65.940 75.470 66.080 75.635 ;
        RECT 65.880 75.150 66.140 75.470 ;
        RECT 66.340 74.810 66.600 75.130 ;
        RECT 66.400 74.450 66.540 74.810 ;
        RECT 66.340 74.130 66.600 74.450 ;
        RECT 65.420 72.090 65.680 72.410 ;
        RECT 66.860 72.070 67.000 79.570 ;
        RECT 67.320 72.070 67.460 85.350 ;
        RECT 67.780 84.990 67.920 91.955 ;
        RECT 68.700 91.450 68.840 92.830 ;
        RECT 68.640 91.130 68.900 91.450 ;
        RECT 69.160 91.110 69.300 99.290 ;
        RECT 69.620 96.210 69.760 99.630 ;
        RECT 71.460 96.800 71.600 111.870 ;
        RECT 80.660 111.170 80.800 112.890 ;
        RECT 81.970 112.355 82.250 112.725 ;
        RECT 81.980 112.210 82.240 112.355 ;
        RECT 80.600 110.850 80.860 111.170 ;
        RECT 71.860 109.830 72.120 110.150 ;
        RECT 79.680 109.830 79.940 110.150 ;
        RECT 80.600 109.830 80.860 110.150 ;
        RECT 71.920 107.770 72.060 109.830 ;
        RECT 71.860 107.450 72.120 107.770 ;
        RECT 73.240 107.450 73.500 107.770 ;
        RECT 73.300 105.730 73.440 107.450 ;
        RECT 79.740 107.430 79.880 109.830 ;
        RECT 79.680 107.110 79.940 107.430 ;
        RECT 79.220 106.430 79.480 106.750 ;
        RECT 73.240 105.410 73.500 105.730 ;
        RECT 76.920 104.730 77.180 105.050 ;
        RECT 75.080 103.710 75.340 104.030 ;
        RECT 72.320 101.330 72.580 101.650 ;
        RECT 71.860 96.800 72.120 96.890 ;
        RECT 71.000 96.660 72.120 96.800 ;
        RECT 70.480 96.230 70.740 96.550 ;
        RECT 69.560 95.890 69.820 96.210 ;
        RECT 70.020 95.550 70.280 95.870 ;
        RECT 70.080 94.510 70.220 95.550 ;
        RECT 70.540 94.850 70.680 96.230 ;
        RECT 70.480 94.530 70.740 94.850 ;
        RECT 70.020 94.190 70.280 94.510 ;
        RECT 70.020 91.130 70.280 91.450 ;
        RECT 69.100 90.790 69.360 91.110 ;
        RECT 70.080 90.770 70.220 91.130 ;
        RECT 70.020 90.450 70.280 90.770 ;
        RECT 70.080 87.710 70.220 90.450 ;
        RECT 71.000 90.430 71.140 96.660 ;
        RECT 71.860 96.570 72.120 96.660 ;
        RECT 71.390 96.035 71.670 96.405 ;
        RECT 71.460 95.870 71.600 96.035 ;
        RECT 71.400 95.550 71.660 95.870 ;
        RECT 72.380 94.170 72.520 101.330 ;
        RECT 72.780 98.950 73.040 99.270 ;
        RECT 72.320 93.850 72.580 94.170 ;
        RECT 72.320 91.130 72.580 91.450 ;
        RECT 71.400 90.790 71.660 91.110 ;
        RECT 70.940 90.110 71.200 90.430 ;
        RECT 71.000 88.390 71.140 90.110 ;
        RECT 71.460 88.390 71.600 90.790 ;
        RECT 72.380 88.730 72.520 91.130 ;
        RECT 72.320 88.410 72.580 88.730 ;
        RECT 70.940 88.070 71.200 88.390 ;
        RECT 71.400 88.070 71.660 88.390 ;
        RECT 70.020 87.390 70.280 87.710 ;
        RECT 67.720 84.670 67.980 84.990 ;
        RECT 67.720 83.650 67.980 83.970 ;
        RECT 67.780 77.930 67.920 83.650 ;
        RECT 70.080 83.630 70.220 87.390 ;
        RECT 71.460 86.600 71.600 88.070 ;
        RECT 71.460 86.460 72.060 86.600 ;
        RECT 70.940 86.030 71.200 86.350 ;
        RECT 70.020 83.310 70.280 83.630 ;
        RECT 69.100 82.970 69.360 83.290 ;
        RECT 68.640 82.290 68.900 82.610 ;
        RECT 68.180 81.950 68.440 82.270 ;
        RECT 68.240 79.550 68.380 81.950 ;
        RECT 68.180 79.230 68.440 79.550 ;
        RECT 67.780 77.790 68.380 77.930 ;
        RECT 68.240 77.510 68.380 77.790 ;
        RECT 67.720 77.190 67.980 77.510 ;
        RECT 68.180 77.190 68.440 77.510 ;
        RECT 67.780 76.005 67.920 77.190 ;
        RECT 67.710 75.635 67.990 76.005 ;
        RECT 67.720 74.130 67.980 74.450 ;
        RECT 66.800 71.750 67.060 72.070 ;
        RECT 67.260 71.750 67.520 72.070 ;
        RECT 65.420 71.410 65.680 71.730 ;
        RECT 65.480 66.630 65.620 71.410 ;
        RECT 65.880 71.070 66.140 71.390 ;
        RECT 66.340 71.070 66.600 71.390 ;
        RECT 65.940 70.370 66.080 71.070 ;
        RECT 65.880 70.050 66.140 70.370 ;
        RECT 65.880 69.370 66.140 69.690 ;
        RECT 65.940 67.650 66.080 69.370 ;
        RECT 66.400 69.350 66.540 71.070 ;
        RECT 66.340 69.030 66.600 69.350 ;
        RECT 65.880 67.330 66.140 67.650 ;
        RECT 66.340 66.990 66.600 67.310 ;
        RECT 65.420 66.310 65.680 66.630 ;
        RECT 65.880 65.970 66.140 66.290 ;
        RECT 65.940 64.250 66.080 65.970 ;
        RECT 65.880 63.930 66.140 64.250 ;
        RECT 64.960 62.910 65.220 63.230 ;
        RECT 65.020 61.190 65.160 62.910 ;
        RECT 65.940 61.530 66.080 63.930 ;
        RECT 65.880 61.210 66.140 61.530 ;
        RECT 64.960 60.870 65.220 61.190 ;
        RECT 65.020 57.645 65.160 60.870 ;
        RECT 65.940 58.470 66.080 61.210 ;
        RECT 65.880 58.150 66.140 58.470 ;
        RECT 64.950 57.275 65.230 57.645 ;
        RECT 65.880 57.470 66.140 57.790 ;
        RECT 64.500 56.450 64.760 56.770 ;
        RECT 64.960 56.450 65.220 56.770 ;
        RECT 64.560 55.750 64.700 56.450 ;
        RECT 65.020 55.750 65.160 56.450 ;
        RECT 65.420 56.110 65.680 56.430 ;
        RECT 64.500 55.430 64.760 55.750 ;
        RECT 64.960 55.430 65.220 55.750 ;
        RECT 64.560 54.050 64.700 55.430 ;
        RECT 65.480 55.410 65.620 56.110 ;
        RECT 65.940 55.750 66.080 57.470 ;
        RECT 66.400 56.090 66.540 66.990 ;
        RECT 66.860 59.150 67.000 71.750 ;
        RECT 67.780 71.390 67.920 74.130 ;
        RECT 67.720 71.300 67.980 71.390 ;
        RECT 67.320 71.160 67.980 71.300 ;
        RECT 67.320 69.885 67.460 71.160 ;
        RECT 67.720 71.070 67.980 71.160 ;
        RECT 68.240 70.450 68.380 77.190 ;
        RECT 68.700 73.090 68.840 82.290 ;
        RECT 69.160 80.910 69.300 82.970 ;
        RECT 69.560 82.290 69.820 82.610 ;
        RECT 69.100 80.590 69.360 80.910 ;
        RECT 69.100 77.930 69.360 78.190 ;
        RECT 69.620 77.930 69.760 82.290 ;
        RECT 69.100 77.870 69.760 77.930 ;
        RECT 69.160 77.790 69.760 77.870 ;
        RECT 68.640 72.770 68.900 73.090 ;
        RECT 69.100 72.090 69.360 72.410 ;
        RECT 69.160 71.130 69.300 72.090 ;
        RECT 67.780 70.310 68.380 70.450 ;
        RECT 68.700 70.990 69.300 71.130 ;
        RECT 67.250 69.515 67.530 69.885 ;
        RECT 67.320 66.970 67.460 69.515 ;
        RECT 67.780 68.670 67.920 70.310 ;
        RECT 68.180 69.770 68.440 70.030 ;
        RECT 68.700 69.770 68.840 70.990 ;
        RECT 69.100 70.050 69.360 70.370 ;
        RECT 68.180 69.710 68.840 69.770 ;
        RECT 68.240 69.630 68.840 69.710 ;
        RECT 68.180 69.260 68.440 69.350 ;
        RECT 69.160 69.260 69.300 70.050 ;
        RECT 69.620 69.690 69.760 77.790 ;
        RECT 70.080 75.210 70.220 83.310 ;
        RECT 71.000 77.510 71.140 86.030 ;
        RECT 71.920 86.010 72.060 86.460 ;
        RECT 72.380 86.350 72.520 88.410 ;
        RECT 72.320 86.030 72.580 86.350 ;
        RECT 72.840 86.010 72.980 98.950 ;
        RECT 74.620 98.610 74.880 98.930 ;
        RECT 74.680 97.570 74.820 98.610 ;
        RECT 74.620 97.250 74.880 97.570 ;
        RECT 73.700 95.890 73.960 96.210 ;
        RECT 73.240 92.830 73.500 93.150 ;
        RECT 73.300 92.130 73.440 92.830 ;
        RECT 73.240 91.810 73.500 92.130 ;
        RECT 71.400 85.690 71.660 86.010 ;
        RECT 71.860 85.690 72.120 86.010 ;
        RECT 72.780 85.690 73.040 86.010 ;
        RECT 71.460 80.570 71.600 85.690 ;
        RECT 71.920 82.520 72.060 85.690 ;
        RECT 71.920 82.380 72.520 82.520 ;
        RECT 71.400 80.250 71.660 80.570 ;
        RECT 72.380 77.510 72.520 82.380 ;
        RECT 72.840 77.850 72.980 85.690 ;
        RECT 73.760 82.950 73.900 95.890 ;
        RECT 75.140 92.130 75.280 103.710 ;
        RECT 76.980 103.010 77.120 104.730 ;
        RECT 79.280 104.710 79.420 106.430 ;
        RECT 80.660 105.730 80.800 109.830 ;
        RECT 81.980 109.325 82.240 109.470 ;
        RECT 81.970 108.955 82.250 109.325 ;
        RECT 80.600 105.410 80.860 105.730 ;
        RECT 79.220 104.390 79.480 104.710 ;
        RECT 79.680 104.390 79.940 104.710 ;
        RECT 76.920 102.690 77.180 103.010 ;
        RECT 79.740 101.990 79.880 104.390 ;
        RECT 79.680 101.670 79.940 101.990 ;
        RECT 76.460 100.990 76.720 101.310 ;
        RECT 76.520 97.570 76.660 100.990 ;
        RECT 79.740 100.290 79.880 101.670 ;
        RECT 79.680 99.970 79.940 100.290 ;
        RECT 77.380 98.270 77.640 98.590 ;
        RECT 76.460 97.250 76.720 97.570 ;
        RECT 77.440 96.550 77.580 98.270 ;
        RECT 76.920 96.230 77.180 96.550 ;
        RECT 77.380 96.230 77.640 96.550 ;
        RECT 76.980 94.850 77.120 96.230 ;
        RECT 76.920 94.530 77.180 94.850 ;
        RECT 75.080 91.810 75.340 92.130 ;
        RECT 74.160 88.070 74.420 88.390 ;
        RECT 81.980 88.070 82.240 88.390 ;
        RECT 73.700 82.630 73.960 82.950 ;
        RECT 72.780 77.530 73.040 77.850 ;
        RECT 70.480 77.190 70.740 77.510 ;
        RECT 70.940 77.190 71.200 77.510 ;
        RECT 72.320 77.190 72.580 77.510 ;
        RECT 70.540 75.810 70.680 77.190 ;
        RECT 70.480 75.490 70.740 75.810 ;
        RECT 70.080 75.130 70.680 75.210 ;
        RECT 70.080 75.070 70.740 75.130 ;
        RECT 70.480 74.810 70.740 75.070 ;
        RECT 69.560 69.370 69.820 69.690 ;
        RECT 70.020 69.370 70.280 69.690 ;
        RECT 68.180 69.120 69.300 69.260 ;
        RECT 68.180 69.030 68.440 69.120 ;
        RECT 67.720 68.350 67.980 68.670 ;
        RECT 67.780 67.650 67.920 68.350 ;
        RECT 67.720 67.330 67.980 67.650 ;
        RECT 69.100 66.990 69.360 67.310 ;
        RECT 67.260 66.650 67.520 66.970 ;
        RECT 69.160 64.250 69.300 66.990 ;
        RECT 69.620 64.590 69.760 69.370 ;
        RECT 70.080 67.650 70.220 69.370 ;
        RECT 70.020 67.330 70.280 67.650 ;
        RECT 70.540 67.050 70.680 74.810 ;
        RECT 71.000 72.410 71.140 77.190 ;
        RECT 71.400 76.510 71.660 76.830 ;
        RECT 70.940 72.090 71.200 72.410 ;
        RECT 70.080 66.910 70.680 67.050 ;
        RECT 69.560 64.270 69.820 64.590 ;
        RECT 68.640 63.930 68.900 64.250 ;
        RECT 69.100 63.930 69.360 64.250 ;
        RECT 68.700 63.570 68.840 63.930 ;
        RECT 68.640 63.250 68.900 63.570 ;
        RECT 69.160 62.170 69.300 63.930 ;
        RECT 69.620 63.570 69.760 64.270 ;
        RECT 69.560 63.250 69.820 63.570 ;
        RECT 68.700 62.030 69.300 62.170 ;
        RECT 66.800 58.830 67.060 59.150 ;
        RECT 66.340 55.770 66.600 56.090 ;
        RECT 66.860 56.000 67.000 58.830 ;
        RECT 67.720 56.000 67.980 56.090 ;
        RECT 66.860 55.860 67.980 56.000 ;
        RECT 67.720 55.770 67.980 55.860 ;
        RECT 65.880 55.430 66.140 55.750 ;
        RECT 65.420 55.090 65.680 55.410 ;
        RECT 64.500 53.730 64.760 54.050 ;
        RECT 64.040 53.050 64.300 53.370 ;
        RECT 64.560 53.280 64.700 53.730 ;
        RECT 66.400 53.710 66.540 55.770 ;
        RECT 68.700 55.750 68.840 62.030 ;
        RECT 69.100 61.210 69.360 61.530 ;
        RECT 69.160 58.810 69.300 61.210 ;
        RECT 70.080 61.190 70.220 66.910 ;
        RECT 71.000 66.290 71.140 72.090 ;
        RECT 71.460 69.690 71.600 76.510 ;
        RECT 71.860 74.470 72.120 74.790 ;
        RECT 71.400 69.370 71.660 69.690 ;
        RECT 71.460 67.310 71.600 69.370 ;
        RECT 71.920 69.350 72.060 74.470 ;
        RECT 72.380 70.370 72.520 77.190 ;
        RECT 72.840 72.410 72.980 77.530 ;
        RECT 73.760 77.170 73.900 82.630 ;
        RECT 73.700 76.850 73.960 77.170 ;
        RECT 72.780 72.090 73.040 72.410 ;
        RECT 73.700 72.090 73.960 72.410 ;
        RECT 73.240 71.410 73.500 71.730 ;
        RECT 72.320 70.050 72.580 70.370 ;
        RECT 71.860 69.030 72.120 69.350 ;
        RECT 71.400 66.990 71.660 67.310 ;
        RECT 72.380 66.970 72.520 70.050 ;
        RECT 72.320 66.650 72.580 66.970 ;
        RECT 71.400 66.310 71.660 66.630 ;
        RECT 70.940 65.970 71.200 66.290 ;
        RECT 71.000 65.690 71.140 65.970 ;
        RECT 70.540 65.550 71.140 65.690 ;
        RECT 70.020 60.870 70.280 61.190 ;
        RECT 69.100 58.490 69.360 58.810 ;
        RECT 70.020 58.490 70.280 58.810 ;
        RECT 69.560 57.810 69.820 58.130 ;
        RECT 69.620 56.770 69.760 57.810 ;
        RECT 69.100 56.450 69.360 56.770 ;
        RECT 69.560 56.450 69.820 56.770 ;
        RECT 68.180 55.430 68.440 55.750 ;
        RECT 68.640 55.430 68.900 55.750 ;
        RECT 68.240 55.070 68.380 55.430 ;
        RECT 68.180 54.750 68.440 55.070 ;
        RECT 66.340 53.390 66.600 53.710 ;
        RECT 64.960 53.280 65.220 53.370 ;
        RECT 64.560 53.140 65.220 53.280 ;
        RECT 64.960 53.050 65.220 53.140 ;
        RECT 67.720 52.030 67.980 52.350 ;
        RECT 67.780 50.310 67.920 52.030 ;
        RECT 68.240 50.990 68.380 54.750 ;
        RECT 68.700 53.370 68.840 55.430 ;
        RECT 69.160 54.130 69.300 56.450 ;
        RECT 69.160 53.990 69.760 54.130 ;
        RECT 70.080 54.050 70.220 58.490 ;
        RECT 70.540 55.660 70.680 65.550 ;
        RECT 70.940 63.930 71.200 64.250 ;
        RECT 71.000 62.210 71.140 63.930 ;
        RECT 70.940 61.890 71.200 62.210 ;
        RECT 71.460 59.490 71.600 66.310 ;
        RECT 71.860 65.970 72.120 66.290 ;
        RECT 71.920 64.590 72.060 65.970 ;
        RECT 71.860 64.270 72.120 64.590 ;
        RECT 72.380 64.160 72.520 66.650 ;
        RECT 72.780 64.160 73.040 64.250 ;
        RECT 72.380 64.020 73.040 64.160 ;
        RECT 71.860 60.870 72.120 61.190 ;
        RECT 71.400 59.170 71.660 59.490 ;
        RECT 70.940 55.660 71.200 55.750 ;
        RECT 70.540 55.520 71.200 55.660 ;
        RECT 70.940 55.430 71.200 55.520 ;
        RECT 69.100 53.390 69.360 53.710 ;
        RECT 68.640 53.050 68.900 53.370 ;
        RECT 68.180 50.670 68.440 50.990 ;
        RECT 69.160 50.310 69.300 53.390 ;
        RECT 67.720 49.990 67.980 50.310 ;
        RECT 69.100 49.990 69.360 50.310 ;
        RECT 63.580 49.650 63.840 49.970 ;
        RECT 69.620 48.270 69.760 53.990 ;
        RECT 70.020 53.730 70.280 54.050 ;
        RECT 71.920 53.710 72.060 60.870 ;
        RECT 72.380 55.750 72.520 64.020 ;
        RECT 72.780 63.930 73.040 64.020 ;
        RECT 72.780 63.250 73.040 63.570 ;
        RECT 72.840 57.790 72.980 63.250 ;
        RECT 73.300 58.810 73.440 71.410 ;
        RECT 73.760 64.250 73.900 72.090 ;
        RECT 74.220 71.390 74.360 88.070 ;
        RECT 79.220 87.390 79.480 87.710 ;
        RECT 75.080 85.690 75.340 86.010 ;
        RECT 75.140 83.970 75.280 85.690 ;
        RECT 76.920 84.670 77.180 84.990 ;
        RECT 75.080 83.650 75.340 83.970 ;
        RECT 76.980 82.610 77.120 84.670 ;
        RECT 79.280 82.950 79.420 87.390 ;
        RECT 82.040 86.690 82.180 88.070 ;
        RECT 79.680 86.370 79.940 86.690 ;
        RECT 81.980 86.370 82.240 86.690 ;
        RECT 79.740 82.950 79.880 86.370 ;
        RECT 81.060 85.690 81.320 86.010 ;
        RECT 81.120 83.970 81.260 85.690 ;
        RECT 81.970 85.155 82.250 85.525 ;
        RECT 81.980 85.010 82.240 85.155 ;
        RECT 81.060 83.650 81.320 83.970 ;
        RECT 79.220 82.630 79.480 82.950 ;
        RECT 79.680 82.630 79.940 82.950 ;
        RECT 76.920 82.290 77.180 82.610 ;
        RECT 80.600 80.250 80.860 80.570 ;
        RECT 78.760 79.230 79.020 79.550 ;
        RECT 79.220 79.230 79.480 79.550 ;
        RECT 78.300 78.210 78.560 78.530 ;
        RECT 75.540 76.850 75.800 77.170 ;
        RECT 75.600 75.810 75.740 76.850 ;
        RECT 77.840 76.510 78.100 76.830 ;
        RECT 75.540 75.490 75.800 75.810 ;
        RECT 77.900 75.470 78.040 76.510 ;
        RECT 77.840 75.150 78.100 75.470 ;
        RECT 78.360 74.790 78.500 78.210 ;
        RECT 78.820 77.510 78.960 79.230 ;
        RECT 78.760 77.190 79.020 77.510 ;
        RECT 79.280 75.810 79.420 79.230 ;
        RECT 80.660 78.530 80.800 80.250 ;
        RECT 80.600 78.210 80.860 78.530 ;
        RECT 81.970 78.355 82.250 78.725 ;
        RECT 81.980 78.210 82.240 78.355 ;
        RECT 79.220 75.490 79.480 75.810 ;
        RECT 80.600 74.810 80.860 75.130 ;
        RECT 78.300 74.470 78.560 74.790 ;
        RECT 80.660 73.090 80.800 74.810 ;
        RECT 81.060 73.790 81.320 74.110 ;
        RECT 80.600 72.770 80.860 73.090 ;
        RECT 80.140 71.750 80.400 72.070 ;
        RECT 75.080 71.410 75.340 71.730 ;
        RECT 74.160 71.070 74.420 71.390 ;
        RECT 75.140 70.370 75.280 71.410 ;
        RECT 75.080 70.050 75.340 70.370 ;
        RECT 79.680 66.310 79.940 66.630 ;
        RECT 75.080 65.970 75.340 66.290 ;
        RECT 73.700 63.930 73.960 64.250 ;
        RECT 74.620 63.930 74.880 64.250 ;
        RECT 73.760 61.530 73.900 63.930 ;
        RECT 73.700 61.210 73.960 61.530 ;
        RECT 73.240 58.490 73.500 58.810 ;
        RECT 72.780 57.470 73.040 57.790 ;
        RECT 72.320 55.430 72.580 55.750 ;
        RECT 71.860 53.390 72.120 53.710 ;
        RECT 72.320 52.940 72.580 53.030 ;
        RECT 72.840 52.940 72.980 57.470 ;
        RECT 73.760 56.090 73.900 61.210 ;
        RECT 73.700 56.000 73.960 56.090 ;
        RECT 73.300 55.860 73.960 56.000 ;
        RECT 73.300 53.370 73.440 55.860 ;
        RECT 73.700 55.770 73.960 55.860 ;
        RECT 73.240 53.050 73.500 53.370 ;
        RECT 74.160 53.050 74.420 53.370 ;
        RECT 72.320 52.800 72.980 52.940 ;
        RECT 72.320 52.710 72.580 52.800 ;
        RECT 73.300 50.990 73.440 53.050 ;
        RECT 74.220 51.330 74.360 53.050 ;
        RECT 74.160 51.010 74.420 51.330 ;
        RECT 73.240 50.670 73.500 50.990 ;
        RECT 70.480 49.310 70.740 49.630 ;
        RECT 70.020 48.290 70.280 48.610 ;
        RECT 69.560 47.950 69.820 48.270 ;
        RECT 64.040 45.570 64.300 45.890 ;
        RECT 64.100 44.870 64.240 45.570 ;
        RECT 66.340 44.890 66.600 45.210 ;
        RECT 60.820 44.550 61.080 44.870 ;
        RECT 62.660 44.780 62.920 44.870 ;
        RECT 64.040 44.780 64.300 44.870 ;
        RECT 62.660 44.640 63.320 44.780 ;
        RECT 62.660 44.550 62.920 44.640 ;
        RECT 60.880 44.190 61.020 44.550 ;
        RECT 60.820 43.870 61.080 44.190 ;
        RECT 59.440 42.510 59.700 42.830 ;
        RECT 58.520 42.170 58.780 42.490 ;
        RECT 59.440 41.830 59.700 42.150 ;
        RECT 57.660 39.710 58.260 39.850 ;
        RECT 57.600 38.770 57.860 39.090 ;
        RECT 57.660 37.730 57.800 38.770 ;
        RECT 57.600 37.410 57.860 37.730 ;
        RECT 57.140 30.270 57.400 30.590 ;
        RECT 56.680 26.530 56.940 26.850 ;
        RECT 55.300 25.850 55.560 26.170 ;
        RECT 56.220 25.850 56.480 26.170 ;
        RECT 54.840 25.170 55.100 25.490 ;
        RECT 53.000 20.410 53.260 20.730 ;
        RECT 51.160 19.390 51.420 19.710 ;
        RECT 51.220 17.670 51.360 19.390 ;
        RECT 50.700 17.350 50.960 17.670 ;
        RECT 51.160 17.350 51.420 17.670 ;
        RECT 50.240 16.670 50.500 16.990 ;
        RECT 50.760 15.630 50.900 17.350 ;
        RECT 54.840 16.670 55.100 16.990 ;
        RECT 50.700 15.310 50.960 15.630 ;
        RECT 54.900 14.610 55.040 16.670 ;
        RECT 54.840 14.290 55.100 14.610 ;
        RECT 49.780 11.910 50.040 12.230 ;
        RECT 55.360 11.890 55.500 25.850 ;
        RECT 56.280 20.730 56.420 25.850 ;
        RECT 58.120 21.410 58.260 39.710 ;
        RECT 59.500 39.430 59.640 41.830 ;
        RECT 60.880 39.430 61.020 43.870 ;
        RECT 61.280 42.170 61.540 42.490 ;
        RECT 59.440 39.110 59.700 39.430 ;
        RECT 60.820 39.110 61.080 39.430 ;
        RECT 60.880 37.050 61.020 39.110 ;
        RECT 61.340 37.390 61.480 42.170 ;
        RECT 62.200 38.770 62.460 39.090 ;
        RECT 61.280 37.070 61.540 37.390 ;
        RECT 58.980 36.730 59.240 37.050 ;
        RECT 60.820 36.730 61.080 37.050 ;
        RECT 61.740 36.730 62.000 37.050 ;
        RECT 59.040 36.030 59.180 36.730 ;
        RECT 58.980 35.710 59.240 36.030 ;
        RECT 59.040 33.990 59.180 35.710 ;
        RECT 58.980 33.670 59.240 33.990 ;
        RECT 59.440 31.970 59.700 32.290 ;
        RECT 59.500 26.170 59.640 31.970 ;
        RECT 59.900 28.230 60.160 28.550 ;
        RECT 59.960 26.510 60.100 28.230 ;
        RECT 59.900 26.190 60.160 26.510 ;
        RECT 59.440 26.080 59.700 26.170 ;
        RECT 58.580 25.940 59.700 26.080 ;
        RECT 58.060 21.090 58.320 21.410 ;
        RECT 56.220 20.410 56.480 20.730 ;
        RECT 56.280 15.630 56.420 20.410 ;
        RECT 58.120 20.390 58.260 21.090 ;
        RECT 58.580 20.730 58.720 25.940 ;
        RECT 59.440 25.850 59.700 25.940 ;
        RECT 60.360 25.850 60.620 26.170 ;
        RECT 60.420 25.570 60.560 25.850 ;
        RECT 59.500 25.490 60.560 25.570 ;
        RECT 59.440 25.430 60.560 25.490 ;
        RECT 59.440 25.170 59.700 25.430 ;
        RECT 59.500 20.730 59.640 25.170 ;
        RECT 60.880 23.110 61.020 36.730 ;
        RECT 61.800 36.370 61.940 36.730 ;
        RECT 61.740 36.050 62.000 36.370 ;
        RECT 61.740 31.630 62.000 31.950 ;
        RECT 61.800 29.650 61.940 31.630 ;
        RECT 62.260 29.650 62.400 38.770 ;
        RECT 63.180 38.750 63.320 44.640 ;
        RECT 63.640 44.640 64.300 44.780 ;
        RECT 63.120 38.430 63.380 38.750 ;
        RECT 63.180 37.050 63.320 38.430 ;
        RECT 63.640 37.390 63.780 44.640 ;
        RECT 64.040 44.550 64.300 44.640 ;
        RECT 66.400 44.530 66.540 44.890 ;
        RECT 64.500 44.210 64.760 44.530 ;
        RECT 66.340 44.210 66.600 44.530 ;
        RECT 67.260 44.210 67.520 44.530 ;
        RECT 64.560 41.210 64.700 44.210 ;
        RECT 65.420 43.870 65.680 44.190 ;
        RECT 64.560 41.070 65.160 41.210 ;
        RECT 64.500 40.130 64.760 40.450 ;
        RECT 64.040 39.110 64.300 39.430 ;
        RECT 64.100 38.750 64.240 39.110 ;
        RECT 64.040 38.430 64.300 38.750 ;
        RECT 63.580 37.070 63.840 37.390 ;
        RECT 64.560 37.050 64.700 40.130 ;
        RECT 65.020 39.430 65.160 41.070 ;
        RECT 65.480 39.770 65.620 43.870 ;
        RECT 66.400 43.170 66.540 44.210 ;
        RECT 66.340 42.850 66.600 43.170 ;
        RECT 65.880 42.170 66.140 42.490 ;
        RECT 65.940 40.450 66.080 42.170 ;
        RECT 65.880 40.130 66.140 40.450 ;
        RECT 65.420 39.450 65.680 39.770 ;
        RECT 64.960 39.110 65.220 39.430 ;
        RECT 65.420 38.430 65.680 38.750 ;
        RECT 66.800 38.660 67.060 38.750 ;
        RECT 67.320 38.660 67.460 44.210 ;
        RECT 66.800 38.520 67.460 38.660 ;
        RECT 66.800 38.430 67.060 38.520 ;
        RECT 63.120 36.730 63.380 37.050 ;
        RECT 64.500 36.960 64.760 37.050 ;
        RECT 64.100 36.820 64.760 36.960 ;
        RECT 61.800 29.510 62.400 29.650 ;
        RECT 62.200 27.550 62.460 27.870 ;
        RECT 61.740 26.530 62.000 26.850 ;
        RECT 61.800 25.490 61.940 26.530 ;
        RECT 62.260 26.170 62.400 27.550 ;
        RECT 62.200 25.850 62.460 26.170 ;
        RECT 61.740 25.170 62.000 25.490 ;
        RECT 60.820 22.790 61.080 23.110 ;
        RECT 58.520 20.410 58.780 20.730 ;
        RECT 59.440 20.640 59.700 20.730 ;
        RECT 59.040 20.500 59.700 20.640 ;
        RECT 57.590 19.875 57.870 20.245 ;
        RECT 58.060 20.070 58.320 20.390 ;
        RECT 57.600 19.730 57.860 19.875 ;
        RECT 56.220 15.310 56.480 15.630 ;
        RECT 58.580 15.290 58.720 20.410 ;
        RECT 59.040 15.540 59.180 20.500 ;
        RECT 59.440 20.410 59.700 20.500 ;
        RECT 59.900 20.410 60.160 20.730 ;
        RECT 59.440 19.390 59.700 19.710 ;
        RECT 59.500 17.330 59.640 19.390 ;
        RECT 59.440 17.010 59.700 17.330 ;
        RECT 59.960 16.990 60.100 20.410 ;
        RECT 61.280 20.070 61.540 20.390 ;
        RECT 59.900 16.670 60.160 16.990 ;
        RECT 59.440 15.540 59.700 15.630 ;
        RECT 59.040 15.400 59.700 15.540 ;
        RECT 59.440 15.310 59.700 15.400 ;
        RECT 58.520 14.970 58.780 15.290 ;
        RECT 57.140 14.630 57.400 14.950 ;
        RECT 57.200 12.230 57.340 14.630 ;
        RECT 59.960 12.230 60.100 16.670 ;
        RECT 61.340 12.570 61.480 20.070 ;
        RECT 62.660 19.960 62.920 20.050 ;
        RECT 61.800 19.820 62.920 19.960 ;
        RECT 61.800 18.690 61.940 19.820 ;
        RECT 62.660 19.730 62.920 19.820 ;
        RECT 61.740 18.370 62.000 18.690 ;
        RECT 62.200 17.350 62.460 17.670 ;
        RECT 62.260 14.950 62.400 17.350 ;
        RECT 62.200 14.630 62.460 14.950 ;
        RECT 61.280 12.250 61.540 12.570 ;
        RECT 63.180 12.230 63.320 36.730 ;
        RECT 64.100 31.270 64.240 36.820 ;
        RECT 64.500 36.730 64.760 36.820 ;
        RECT 65.480 36.710 65.620 38.430 ;
        RECT 65.420 36.390 65.680 36.710 ;
        RECT 64.500 35.940 64.760 36.030 ;
        RECT 65.480 35.940 65.620 36.390 ;
        RECT 67.320 36.030 67.460 38.520 ;
        RECT 67.720 36.730 67.980 37.050 ;
        RECT 64.500 35.800 65.620 35.940 ;
        RECT 64.500 35.710 64.760 35.800 ;
        RECT 67.260 35.710 67.520 36.030 ;
        RECT 64.040 30.950 64.300 31.270 ;
        RECT 64.040 26.420 64.300 26.510 ;
        RECT 64.560 26.420 64.700 35.710 ;
        RECT 66.800 34.350 67.060 34.670 ;
        RECT 66.340 32.990 66.600 33.310 ;
        RECT 66.400 31.270 66.540 32.990 ;
        RECT 66.340 30.950 66.600 31.270 ;
        RECT 65.420 28.230 65.680 28.550 ;
        RECT 64.960 27.890 65.220 28.210 ;
        RECT 65.020 26.850 65.160 27.890 ;
        RECT 64.960 26.530 65.220 26.850 ;
        RECT 65.480 26.510 65.620 28.230 ;
        RECT 64.040 26.280 64.700 26.420 ;
        RECT 64.040 26.190 64.300 26.280 ;
        RECT 65.420 26.190 65.680 26.510 ;
        RECT 64.100 21.410 64.240 26.190 ;
        RECT 66.400 23.450 66.540 30.950 ;
        RECT 66.340 23.130 66.600 23.450 ;
        RECT 64.040 21.090 64.300 21.410 ;
        RECT 65.420 20.410 65.680 20.730 ;
        RECT 65.480 18.690 65.620 20.410 ;
        RECT 65.420 18.600 65.680 18.690 ;
        RECT 65.020 18.460 65.680 18.600 ;
        RECT 65.020 15.970 65.160 18.460 ;
        RECT 65.420 18.370 65.680 18.460 ;
        RECT 66.400 18.010 66.540 23.130 ;
        RECT 66.860 18.690 67.000 34.350 ;
        RECT 67.320 33.650 67.460 35.710 ;
        RECT 67.260 33.330 67.520 33.650 ;
        RECT 67.320 28.210 67.460 33.330 ;
        RECT 67.780 31.950 67.920 36.730 ;
        RECT 67.720 31.630 67.980 31.950 ;
        RECT 67.260 27.890 67.520 28.210 ;
        RECT 67.320 21.070 67.460 27.890 ;
        RECT 67.780 21.070 67.920 31.630 ;
        RECT 69.550 31.435 69.830 31.805 ;
        RECT 69.560 31.290 69.820 31.435 ;
        RECT 70.080 30.930 70.220 48.290 ;
        RECT 70.540 47.930 70.680 49.310 ;
        RECT 70.480 47.610 70.740 47.930 ;
        RECT 71.400 44.550 71.660 44.870 ;
        RECT 71.860 44.550 72.120 44.870 ;
        RECT 72.320 44.550 72.580 44.870 ;
        RECT 70.480 42.510 70.740 42.830 ;
        RECT 70.540 39.430 70.680 42.510 ;
        RECT 71.460 40.450 71.600 44.550 ;
        RECT 71.400 40.130 71.660 40.450 ;
        RECT 70.480 39.110 70.740 39.430 ;
        RECT 71.400 36.730 71.660 37.050 ;
        RECT 71.460 33.990 71.600 36.730 ;
        RECT 71.920 36.710 72.060 44.550 ;
        RECT 71.860 36.390 72.120 36.710 ;
        RECT 72.380 36.370 72.520 44.550 ;
        RECT 73.700 43.870 73.960 44.190 ;
        RECT 73.760 39.090 73.900 43.870 ;
        RECT 73.700 38.770 73.960 39.090 ;
        RECT 74.680 37.050 74.820 63.930 ;
        RECT 73.240 36.730 73.500 37.050 ;
        RECT 74.620 36.730 74.880 37.050 ;
        RECT 72.320 36.050 72.580 36.370 ;
        RECT 73.300 35.010 73.440 36.730 ;
        RECT 73.240 34.690 73.500 35.010 ;
        RECT 74.680 34.330 74.820 36.730 ;
        RECT 74.620 34.010 74.880 34.330 ;
        RECT 71.400 33.670 71.660 33.990 ;
        RECT 72.320 33.670 72.580 33.990 ;
        RECT 69.100 30.610 69.360 30.930 ;
        RECT 70.020 30.610 70.280 30.930 ;
        RECT 69.160 23.020 69.300 30.610 ;
        RECT 71.460 26.250 71.600 33.670 ;
        RECT 71.860 33.330 72.120 33.650 ;
        RECT 71.920 31.950 72.060 33.330 ;
        RECT 72.380 32.290 72.520 33.670 ;
        RECT 72.320 31.970 72.580 32.290 ;
        RECT 71.860 31.630 72.120 31.950 ;
        RECT 72.320 31.290 72.580 31.610 ;
        RECT 73.240 31.290 73.500 31.610 ;
        RECT 74.150 31.435 74.430 31.805 ;
        RECT 74.160 31.290 74.420 31.435 ;
        RECT 72.380 30.930 72.520 31.290 ;
        RECT 72.320 30.610 72.580 30.930 ;
        RECT 73.300 30.590 73.440 31.290 ;
        RECT 74.620 30.610 74.880 30.930 ;
        RECT 73.240 30.270 73.500 30.590 ;
        RECT 71.860 27.890 72.120 28.210 ;
        RECT 71.920 26.850 72.060 27.890 ;
        RECT 72.780 27.550 73.040 27.870 ;
        RECT 71.860 26.530 72.120 26.850 ;
        RECT 70.480 25.850 70.740 26.170 ;
        RECT 70.940 25.850 71.200 26.170 ;
        RECT 71.460 26.110 72.520 26.250 ;
        RECT 70.540 24.130 70.680 25.850 ;
        RECT 70.480 23.810 70.740 24.130 ;
        RECT 70.480 23.130 70.740 23.450 ;
        RECT 69.560 23.020 69.820 23.110 ;
        RECT 69.160 22.880 69.820 23.020 ;
        RECT 69.560 22.790 69.820 22.880 ;
        RECT 67.260 20.750 67.520 21.070 ;
        RECT 67.720 20.750 67.980 21.070 ;
        RECT 66.800 18.370 67.060 18.690 ;
        RECT 66.340 17.690 66.600 18.010 ;
        RECT 66.860 17.670 67.000 18.370 ;
        RECT 66.800 17.350 67.060 17.670 ;
        RECT 65.420 16.670 65.680 16.990 ;
        RECT 64.960 15.650 65.220 15.970 ;
        RECT 65.020 12.230 65.160 15.650 ;
        RECT 65.480 15.290 65.620 16.670 ;
        RECT 65.420 14.970 65.680 15.290 ;
        RECT 67.320 13.870 67.460 20.750 ;
        RECT 69.100 20.410 69.360 20.730 ;
        RECT 69.160 18.010 69.300 20.410 ;
        RECT 69.100 17.690 69.360 18.010 ;
        RECT 67.720 17.350 67.980 17.670 ;
        RECT 67.780 15.970 67.920 17.350 ;
        RECT 67.720 15.650 67.980 15.970 ;
        RECT 69.620 15.290 69.760 22.790 ;
        RECT 70.540 21.410 70.680 23.130 ;
        RECT 70.480 21.090 70.740 21.410 ;
        RECT 70.540 19.710 70.680 21.090 ;
        RECT 71.000 20.730 71.140 25.850 ;
        RECT 71.400 22.790 71.660 23.110 ;
        RECT 71.860 22.790 72.120 23.110 ;
        RECT 71.460 21.410 71.600 22.790 ;
        RECT 71.920 21.410 72.060 22.790 ;
        RECT 71.400 21.090 71.660 21.410 ;
        RECT 71.860 21.090 72.120 21.410 ;
        RECT 72.380 20.730 72.520 26.110 ;
        RECT 72.840 23.110 72.980 27.550 ;
        RECT 73.300 25.830 73.440 30.270 ;
        RECT 74.680 26.170 74.820 30.610 ;
        RECT 74.620 25.850 74.880 26.170 ;
        RECT 73.240 25.510 73.500 25.830 ;
        RECT 75.140 25.570 75.280 65.970 ;
        RECT 76.920 65.630 77.180 65.950 ;
        RECT 77.840 65.630 78.100 65.950 ;
        RECT 79.220 65.630 79.480 65.950 ;
        RECT 76.000 64.270 76.260 64.590 ;
        RECT 76.060 62.210 76.200 64.270 ;
        RECT 76.000 61.890 76.260 62.210 ;
        RECT 75.540 57.470 75.800 57.790 ;
        RECT 75.600 55.750 75.740 57.470 ;
        RECT 75.540 55.430 75.800 55.750 ;
        RECT 76.000 53.050 76.260 53.370 ;
        RECT 76.060 43.170 76.200 53.050 ;
        RECT 76.980 50.650 77.120 65.630 ;
        RECT 77.900 65.125 78.040 65.630 ;
        RECT 77.830 64.755 78.110 65.125 ;
        RECT 78.760 64.610 79.020 64.930 ;
        RECT 77.840 62.910 78.100 63.230 ;
        RECT 77.900 61.530 78.040 62.910 ;
        RECT 78.820 61.530 78.960 64.610 ;
        RECT 77.840 61.210 78.100 61.530 ;
        RECT 78.760 61.210 79.020 61.530 ;
        RECT 79.280 60.850 79.420 65.630 ;
        RECT 79.220 60.530 79.480 60.850 ;
        RECT 77.380 60.190 77.640 60.510 ;
        RECT 77.440 59.490 77.580 60.190 ;
        RECT 79.740 59.490 79.880 66.310 ;
        RECT 80.200 63.570 80.340 71.750 ;
        RECT 80.660 69.690 80.800 72.770 ;
        RECT 81.120 72.070 81.260 73.790 ;
        RECT 81.060 71.750 81.320 72.070 ;
        RECT 81.970 71.555 82.250 71.925 ;
        RECT 82.040 71.390 82.180 71.555 ;
        RECT 81.980 71.070 82.240 71.390 ;
        RECT 80.600 69.370 80.860 69.690 ;
        RECT 82.430 68.155 82.710 68.525 ;
        RECT 81.980 66.310 82.240 66.630 ;
        RECT 82.040 64.930 82.180 66.310 ;
        RECT 80.600 64.610 80.860 64.930 ;
        RECT 81.980 64.610 82.240 64.930 ;
        RECT 80.140 63.250 80.400 63.570 ;
        RECT 80.140 60.870 80.400 61.190 ;
        RECT 77.380 59.170 77.640 59.490 ;
        RECT 79.680 59.170 79.940 59.490 ;
        RECT 77.840 58.150 78.100 58.470 ;
        RECT 77.900 56.770 78.040 58.150 ;
        RECT 80.200 56.770 80.340 60.870 ;
        RECT 80.660 58.810 80.800 64.610 ;
        RECT 82.500 64.250 82.640 68.155 ;
        RECT 82.440 63.930 82.700 64.250 ;
        RECT 81.980 61.725 82.240 61.870 ;
        RECT 81.970 61.355 82.250 61.725 ;
        RECT 81.520 60.870 81.780 61.190 ;
        RECT 80.600 58.490 80.860 58.810 ;
        RECT 81.060 58.490 81.320 58.810 ;
        RECT 77.840 56.450 78.100 56.770 ;
        RECT 80.140 56.450 80.400 56.770 ;
        RECT 77.380 52.030 77.640 52.350 ;
        RECT 79.680 52.030 79.940 52.350 ;
        RECT 77.440 50.650 77.580 52.030 ;
        RECT 79.740 50.650 79.880 52.030 ;
        RECT 76.920 50.330 77.180 50.650 ;
        RECT 77.380 50.330 77.640 50.650 ;
        RECT 79.680 50.330 79.940 50.650 ;
        RECT 81.120 47.250 81.260 58.490 ;
        RECT 81.580 56.770 81.720 60.870 ;
        RECT 81.970 57.955 82.250 58.325 ;
        RECT 81.980 57.810 82.240 57.955 ;
        RECT 81.520 56.450 81.780 56.770 ;
        RECT 81.980 52.030 82.240 52.350 ;
        RECT 82.040 51.525 82.180 52.030 ;
        RECT 81.970 51.155 82.250 51.525 ;
        RECT 82.440 50.330 82.700 50.650 ;
        RECT 82.500 47.930 82.640 50.330 ;
        RECT 82.440 47.610 82.700 47.930 ;
        RECT 81.060 46.930 81.320 47.250 ;
        RECT 76.920 44.210 77.180 44.530 ;
        RECT 76.000 42.850 76.260 43.170 ;
        RECT 75.540 39.110 75.800 39.430 ;
        RECT 75.600 33.990 75.740 39.110 ;
        RECT 76.980 37.050 77.120 44.210 ;
        RECT 81.060 42.170 81.320 42.490 ;
        RECT 81.120 38.750 81.260 42.170 ;
        RECT 82.900 41.490 83.160 41.810 ;
        RECT 82.960 41.325 83.100 41.490 ;
        RECT 82.890 40.955 83.170 41.325 ;
        RECT 81.060 38.430 81.320 38.750 ;
        RECT 76.920 36.730 77.180 37.050 ;
        RECT 76.920 36.050 77.180 36.370 ;
        RECT 75.540 33.670 75.800 33.990 ;
        RECT 75.600 31.270 75.740 33.670 ;
        RECT 76.980 31.950 77.120 36.050 ;
        RECT 79.220 32.990 79.480 33.310 ;
        RECT 76.920 31.630 77.180 31.950 ;
        RECT 79.280 31.610 79.420 32.990 ;
        RECT 81.060 31.970 81.320 32.290 ;
        RECT 79.220 31.290 79.480 31.610 ;
        RECT 75.540 30.950 75.800 31.270 ;
        RECT 75.600 26.510 75.740 30.950 ;
        RECT 76.000 28.910 76.260 29.230 ;
        RECT 75.540 26.190 75.800 26.510 ;
        RECT 74.680 25.430 75.280 25.570 ;
        RECT 73.700 24.830 73.960 25.150 ;
        RECT 73.240 23.130 73.500 23.450 ;
        RECT 72.780 22.790 73.040 23.110 ;
        RECT 72.780 22.110 73.040 22.430 ;
        RECT 72.840 20.730 72.980 22.110 ;
        RECT 70.940 20.410 71.200 20.730 ;
        RECT 71.400 20.410 71.660 20.730 ;
        RECT 72.320 20.640 72.580 20.730 ;
        RECT 71.920 20.500 72.580 20.640 ;
        RECT 70.480 19.390 70.740 19.710 ;
        RECT 70.940 17.350 71.200 17.670 ;
        RECT 71.000 16.990 71.140 17.350 ;
        RECT 70.940 16.670 71.200 16.990 ;
        RECT 71.460 15.290 71.600 20.410 ;
        RECT 71.920 18.350 72.060 20.500 ;
        RECT 72.320 20.410 72.580 20.500 ;
        RECT 72.780 20.410 73.040 20.730 ;
        RECT 72.320 19.390 72.580 19.710 ;
        RECT 71.860 18.030 72.120 18.350 ;
        RECT 72.380 17.670 72.520 19.390 ;
        RECT 71.860 17.350 72.120 17.670 ;
        RECT 72.320 17.350 72.580 17.670 ;
        RECT 72.780 17.350 73.040 17.670 ;
        RECT 69.560 14.970 69.820 15.290 ;
        RECT 71.400 14.970 71.660 15.290 ;
        RECT 69.560 14.290 69.820 14.610 ;
        RECT 66.400 13.730 67.460 13.870 ;
        RECT 57.140 11.910 57.400 12.230 ;
        RECT 59.900 11.910 60.160 12.230 ;
        RECT 63.120 11.910 63.380 12.230 ;
        RECT 64.960 11.910 65.220 12.230 ;
        RECT 66.400 11.890 66.540 13.730 ;
        RECT 69.620 12.230 69.760 14.290 ;
        RECT 71.920 13.250 72.060 17.350 ;
        RECT 72.320 15.650 72.580 15.970 ;
        RECT 71.860 12.930 72.120 13.250 ;
        RECT 72.380 12.570 72.520 15.650 ;
        RECT 72.840 14.270 72.980 17.350 ;
        RECT 73.300 15.630 73.440 23.130 ;
        RECT 73.760 23.110 73.900 24.830 ;
        RECT 73.700 22.790 73.960 23.110 ;
        RECT 73.760 17.670 73.900 22.790 ;
        RECT 74.680 21.070 74.820 25.430 ;
        RECT 75.080 24.830 75.340 25.150 ;
        RECT 75.140 23.790 75.280 24.830 ;
        RECT 75.080 23.470 75.340 23.790 ;
        RECT 75.600 23.450 75.740 26.190 ;
        RECT 75.540 23.130 75.800 23.450 ;
        RECT 75.540 22.450 75.800 22.770 ;
        RECT 74.620 20.750 74.880 21.070 ;
        RECT 75.600 20.390 75.740 22.450 ;
        RECT 75.540 20.070 75.800 20.390 ;
        RECT 73.700 17.350 73.960 17.670 ;
        RECT 73.760 16.990 73.900 17.350 ;
        RECT 73.700 16.670 73.960 16.990 ;
        RECT 74.620 16.670 74.880 16.990 ;
        RECT 75.540 16.670 75.800 16.990 ;
        RECT 73.240 15.310 73.500 15.630 ;
        RECT 73.300 14.950 73.440 15.310 ;
        RECT 74.680 15.290 74.820 16.670 ;
        RECT 74.620 14.970 74.880 15.290 ;
        RECT 73.240 14.630 73.500 14.950 ;
        RECT 72.780 13.950 73.040 14.270 ;
        RECT 73.300 12.570 73.440 14.630 ;
        RECT 75.600 13.250 75.740 16.670 ;
        RECT 76.060 15.290 76.200 28.910 ;
        RECT 78.300 26.190 78.560 26.510 ;
        RECT 77.840 25.850 78.100 26.170 ;
        RECT 77.900 22.430 78.040 25.850 ;
        RECT 77.840 22.110 78.100 22.430 ;
        RECT 77.840 20.410 78.100 20.730 ;
        RECT 77.380 18.030 77.640 18.350 ;
        RECT 76.920 16.670 77.180 16.990 ;
        RECT 76.000 14.970 76.260 15.290 ;
        RECT 75.540 12.930 75.800 13.250 ;
        RECT 72.320 12.250 72.580 12.570 ;
        RECT 73.240 12.250 73.500 12.570 ;
        RECT 76.980 12.230 77.120 16.670 ;
        RECT 69.560 11.910 69.820 12.230 ;
        RECT 76.920 11.910 77.180 12.230 ;
        RECT 32.300 11.570 32.560 11.890 ;
        RECT 41.960 11.570 42.220 11.890 ;
        RECT 55.300 11.570 55.560 11.890 ;
        RECT 66.340 11.570 66.600 11.890 ;
        RECT 32.360 4.000 32.500 11.570 ;
        RECT 35.060 11.230 35.320 11.550 ;
        RECT 38.740 11.230 39.000 11.550 ;
        RECT 41.500 11.230 41.760 11.550 ;
        RECT 45.180 11.230 45.440 11.550 ;
        RECT 48.400 11.230 48.660 11.550 ;
        RECT 51.620 11.230 51.880 11.550 ;
        RECT 54.840 11.230 55.100 11.550 ;
        RECT 58.060 11.230 58.320 11.550 ;
        RECT 61.280 11.230 61.540 11.550 ;
        RECT 64.500 11.230 64.760 11.550 ;
        RECT 67.720 11.230 67.980 11.550 ;
        RECT 35.120 5.170 35.260 11.230 ;
        RECT 35.120 5.030 35.720 5.170 ;
        RECT 35.580 4.000 35.720 5.030 ;
        RECT 38.800 4.000 38.940 11.230 ;
        RECT 41.560 5.850 41.700 11.230 ;
        RECT 41.560 5.710 42.160 5.850 ;
        RECT 42.020 4.000 42.160 5.710 ;
        RECT 45.240 4.000 45.380 11.230 ;
        RECT 48.460 4.000 48.600 11.230 ;
        RECT 51.680 4.000 51.820 11.230 ;
        RECT 54.900 4.000 55.040 11.230 ;
        RECT 58.120 4.000 58.260 11.230 ;
        RECT 61.340 4.000 61.480 11.230 ;
        RECT 64.560 4.000 64.700 11.230 ;
        RECT 67.780 4.000 67.920 11.230 ;
        RECT 70.940 6.470 71.200 6.790 ;
        RECT 71.000 4.000 71.140 6.470 ;
        RECT 74.160 5.450 74.420 5.770 ;
        RECT 74.220 4.000 74.360 5.450 ;
        RECT 77.440 4.000 77.580 18.030 ;
        RECT 77.900 11.890 78.040 20.410 ;
        RECT 78.360 17.670 78.500 26.190 ;
        RECT 79.280 20.730 79.420 31.290 ;
        RECT 81.120 28.550 81.260 31.970 ;
        RECT 81.060 28.230 81.320 28.550 ;
        RECT 82.900 27.725 83.160 27.870 ;
        RECT 82.890 27.355 83.170 27.725 ;
        RECT 82.440 22.110 82.700 22.430 ;
        RECT 82.500 20.730 82.640 22.110 ;
        RECT 79.220 20.410 79.480 20.730 ;
        RECT 82.440 20.410 82.700 20.730 ;
        RECT 87.040 20.070 87.300 20.390 ;
        RECT 83.820 19.730 84.080 20.050 ;
        RECT 80.600 19.390 80.860 19.710 ;
        RECT 78.300 17.350 78.560 17.670 ;
        RECT 80.140 17.350 80.400 17.670 ;
        RECT 79.220 16.670 79.480 16.990 ;
        RECT 77.840 11.570 78.100 11.890 ;
        RECT 79.280 5.770 79.420 16.670 ;
        RECT 80.200 15.970 80.340 17.350 ;
        RECT 80.140 15.650 80.400 15.970 ;
        RECT 79.220 5.450 79.480 5.770 ;
        RECT 80.660 4.000 80.800 19.390 ;
        RECT 81.520 13.950 81.780 14.270 ;
        RECT 81.580 6.790 81.720 13.950 ;
        RECT 81.520 6.470 81.780 6.790 ;
        RECT 83.880 4.000 84.020 19.730 ;
        RECT 87.100 4.000 87.240 20.070 ;
      LAYER met3 ;
        RECT 21.050 198.395 22.630 198.725 ;
        RECT 24.350 195.675 25.930 196.005 ;
        RECT 0.525 195.650 0.855 195.665 ;
        RECT 0.525 195.350 5.210 195.650 ;
        RECT 0.525 195.335 0.855 195.350 ;
        RECT 4.910 194.290 5.210 195.350 ;
        RECT 4.000 193.990 5.210 194.290 ;
        RECT 21.050 192.955 22.630 193.285 ;
        RECT 24.350 190.235 25.930 190.565 ;
        RECT 38.245 189.530 38.575 189.545 ;
        RECT 43.765 189.530 44.095 189.545 ;
        RECT 38.245 189.230 44.095 189.530 ;
        RECT 38.245 189.215 38.575 189.230 ;
        RECT 43.765 189.215 44.095 189.230 ;
        RECT 21.050 187.515 22.630 187.845 ;
        RECT 24.350 184.795 25.930 185.125 ;
        RECT 21.050 182.075 22.630 182.405 ;
        RECT 52.965 180.690 53.295 180.705 ;
        RECT 55.725 180.690 56.055 180.705 ;
        RECT 52.965 180.390 56.055 180.690 ;
        RECT 52.965 180.375 53.295 180.390 ;
        RECT 55.725 180.375 56.055 180.390 ;
        RECT 24.350 179.355 25.930 179.685 ;
        RECT 21.050 176.635 22.630 176.965 ;
        RECT 24.350 173.915 25.930 174.245 ;
        RECT 21.050 171.195 22.630 171.525 ;
        RECT 62.165 170.490 62.495 170.505 ;
        RECT 65.385 170.490 65.715 170.505 ;
        RECT 62.165 170.190 65.715 170.490 ;
        RECT 62.165 170.175 62.495 170.190 ;
        RECT 65.385 170.175 65.715 170.190 ;
        RECT 24.350 168.475 25.930 168.805 ;
        RECT 21.050 165.755 22.630 166.085 ;
        RECT 24.350 163.035 25.930 163.365 ;
        RECT 21.050 160.315 22.630 160.645 ;
        RECT 24.350 157.595 25.930 157.925 ;
        RECT 21.050 154.875 22.630 155.205 ;
        RECT 24.350 152.155 25.930 152.485 ;
        RECT 21.050 149.435 22.630 149.765 ;
        RECT 24.350 146.715 25.930 147.045 ;
        RECT 21.050 143.995 22.630 144.325 ;
        RECT 24.350 141.275 25.930 141.605 ;
        RECT 21.050 138.555 22.630 138.885 ;
        RECT 46.525 137.170 46.855 137.185 ;
        RECT 64.005 137.170 64.335 137.185 ;
        RECT 46.525 136.870 64.335 137.170 ;
        RECT 46.525 136.855 46.855 136.870 ;
        RECT 64.005 136.855 64.335 136.870 ;
        RECT 24.350 135.835 25.930 136.165 ;
        RECT 4.205 133.770 4.535 133.785 ;
        RECT 3.990 133.455 4.535 133.770 ;
        RECT 3.990 133.240 4.290 133.455 ;
        RECT 4.000 132.790 4.290 133.240 ;
        RECT 21.050 133.115 22.630 133.445 ;
        RECT 24.350 130.395 25.930 130.725 ;
        RECT 21.050 127.675 22.630 128.005 ;
        RECT 24.350 124.955 25.930 125.285 ;
        RECT 21.050 122.235 22.630 122.565 ;
        RECT 24.350 119.515 25.930 119.845 ;
        RECT 21.050 116.795 22.630 117.125 ;
        RECT 24.350 114.075 25.930 114.405 ;
        RECT 4.205 113.370 4.535 113.385 ;
        RECT 3.990 113.055 4.535 113.370 ;
        RECT 3.990 112.840 4.290 113.055 ;
        RECT 4.000 112.390 4.290 112.840 ;
        RECT 81.945 112.690 82.275 112.705 ;
        RECT 81.945 112.390 86.000 112.690 ;
        RECT 81.945 112.375 82.275 112.390 ;
        RECT 21.050 111.355 22.630 111.685 ;
        RECT 4.205 109.970 4.535 109.985 ;
        RECT 3.990 109.655 4.535 109.970 ;
        RECT 3.990 109.440 4.290 109.655 ;
        RECT 4.000 108.990 4.290 109.440 ;
        RECT 81.945 109.290 82.275 109.305 ;
        RECT 81.945 108.990 86.000 109.290 ;
        RECT 81.945 108.975 82.275 108.990 ;
        RECT 24.350 108.635 25.930 108.965 ;
        RECT 21.050 105.915 22.630 106.245 ;
        RECT 6.505 105.890 6.835 105.905 ;
        RECT 4.000 105.590 6.835 105.890 ;
        RECT 6.505 105.575 6.835 105.590 ;
        RECT 24.350 103.195 25.930 103.525 ;
        RECT 15.245 102.490 15.575 102.505 ;
        RECT 4.000 102.190 15.575 102.490 ;
        RECT 15.245 102.175 15.575 102.190 ;
        RECT 21.050 100.475 22.630 100.805 ;
        RECT 4.205 99.770 4.535 99.785 ;
        RECT 3.990 99.455 4.535 99.770 ;
        RECT 3.990 99.240 4.290 99.455 ;
        RECT 4.000 98.790 4.290 99.240 ;
        RECT 24.350 97.755 25.930 98.085 ;
        RECT 65.385 96.370 65.715 96.385 ;
        RECT 71.365 96.370 71.695 96.385 ;
        RECT 65.385 96.070 71.695 96.370 ;
        RECT 65.385 96.055 65.715 96.070 ;
        RECT 71.365 96.055 71.695 96.070 ;
        RECT 21.050 95.035 22.630 95.365 ;
        RECT 24.350 92.315 25.930 92.645 ;
        RECT 58.945 92.290 59.275 92.305 ;
        RECT 67.685 92.290 68.015 92.305 ;
        RECT 58.945 91.990 68.015 92.290 ;
        RECT 58.945 91.975 59.275 91.990 ;
        RECT 67.685 91.975 68.015 91.990 ;
        RECT 21.050 89.595 22.630 89.925 ;
        RECT 24.350 86.875 25.930 87.205 ;
        RECT 81.945 85.490 82.275 85.505 ;
        RECT 81.945 85.190 86.000 85.490 ;
        RECT 81.945 85.175 82.275 85.190 ;
        RECT 21.050 84.155 22.630 84.485 ;
        RECT 24.350 81.435 25.930 81.765 ;
        RECT 62.165 79.370 62.495 79.385 ;
        RECT 64.925 79.370 65.255 79.385 ;
        RECT 62.165 79.070 65.255 79.370 ;
        RECT 62.165 79.055 62.495 79.070 ;
        RECT 64.925 79.055 65.255 79.070 ;
        RECT 21.050 78.715 22.630 79.045 ;
        RECT 81.945 78.690 82.275 78.705 ;
        RECT 81.945 78.390 86.000 78.690 ;
        RECT 81.945 78.375 82.275 78.390 ;
        RECT 24.350 75.995 25.930 76.325 ;
        RECT 65.845 75.970 66.175 75.985 ;
        RECT 67.685 75.970 68.015 75.985 ;
        RECT 65.845 75.670 68.015 75.970 ;
        RECT 65.845 75.655 66.175 75.670 ;
        RECT 67.685 75.655 68.015 75.670 ;
        RECT 21.050 73.275 22.630 73.605 ;
        RECT 81.945 71.890 82.275 71.905 ;
        RECT 81.945 71.590 86.000 71.890 ;
        RECT 81.945 71.575 82.275 71.590 ;
        RECT 24.350 70.555 25.930 70.885 ;
        RECT 60.785 69.850 61.115 69.865 ;
        RECT 67.225 69.850 67.555 69.865 ;
        RECT 60.785 69.550 67.555 69.850 ;
        RECT 60.785 69.535 61.115 69.550 ;
        RECT 67.225 69.535 67.555 69.550 ;
        RECT 61.245 69.170 61.575 69.185 ;
        RECT 64.465 69.170 64.795 69.185 ;
        RECT 61.245 68.870 64.795 69.170 ;
        RECT 61.245 68.855 61.575 68.870 ;
        RECT 64.465 68.855 64.795 68.870 ;
        RECT 82.405 68.490 82.735 68.505 ;
        RECT 82.405 68.190 86.000 68.490 ;
        RECT 82.405 68.175 82.735 68.190 ;
        RECT 21.050 67.835 22.630 68.165 ;
        RECT 24.350 65.115 25.930 65.445 ;
        RECT 6.505 65.090 6.835 65.105 ;
        RECT 4.000 64.790 6.835 65.090 ;
        RECT 6.505 64.775 6.835 64.790 ;
        RECT 77.805 65.090 78.135 65.105 ;
        RECT 77.805 64.790 86.000 65.090 ;
        RECT 77.805 64.775 78.135 64.790 ;
        RECT 35.945 63.060 36.275 63.065 ;
        RECT 35.945 63.050 36.530 63.060 ;
        RECT 35.945 62.750 36.730 63.050 ;
        RECT 35.945 62.740 36.530 62.750 ;
        RECT 35.945 62.735 36.275 62.740 ;
        RECT 21.050 62.395 22.630 62.725 ;
        RECT 81.945 61.690 82.275 61.705 ;
        RECT 4.000 61.240 4.290 61.690 ;
        RECT 81.945 61.390 86.000 61.690 ;
        RECT 81.945 61.375 82.275 61.390 ;
        RECT 3.990 61.025 4.290 61.240 ;
        RECT 3.990 60.710 4.535 61.025 ;
        RECT 4.205 60.695 4.535 60.710 ;
        RECT 24.350 59.675 25.930 60.005 ;
        RECT 5.585 58.290 5.915 58.305 ;
        RECT 4.000 57.990 5.915 58.290 ;
        RECT 5.585 57.975 5.915 57.990 ;
        RECT 81.945 58.290 82.275 58.305 ;
        RECT 81.945 57.990 86.000 58.290 ;
        RECT 81.945 57.975 82.275 57.990 ;
        RECT 59.865 57.610 60.195 57.625 ;
        RECT 64.925 57.610 65.255 57.625 ;
        RECT 59.865 57.310 65.255 57.610 ;
        RECT 59.865 57.295 60.195 57.310 ;
        RECT 64.925 57.295 65.255 57.310 ;
        RECT 21.050 56.955 22.630 57.285 ;
        RECT 9.265 54.890 9.595 54.905 ;
        RECT 4.000 54.590 9.595 54.890 ;
        RECT 9.265 54.575 9.595 54.590 ;
        RECT 24.350 54.235 25.930 54.565 ;
        RECT 12.945 53.530 13.275 53.545 ;
        RECT 13.865 53.530 14.195 53.545 ;
        RECT 12.945 53.230 14.195 53.530 ;
        RECT 12.945 53.215 13.275 53.230 ;
        RECT 13.865 53.215 14.195 53.230 ;
        RECT 21.050 51.515 22.630 51.845 ;
        RECT 6.505 51.490 6.835 51.505 ;
        RECT 4.000 51.190 6.835 51.490 ;
        RECT 6.505 51.175 6.835 51.190 ;
        RECT 81.945 51.490 82.275 51.505 ;
        RECT 81.945 51.190 86.000 51.490 ;
        RECT 81.945 51.175 82.275 51.190 ;
        RECT 24.350 48.795 25.930 49.125 ;
        RECT 5.125 48.090 5.455 48.105 ;
        RECT 4.000 47.790 5.455 48.090 ;
        RECT 5.125 47.775 5.455 47.790 ;
        RECT 21.050 46.075 22.630 46.405 ;
        RECT 4.205 45.370 4.535 45.385 ;
        RECT 3.990 45.055 4.535 45.370 ;
        RECT 3.990 44.840 4.290 45.055 ;
        RECT 4.000 44.390 4.290 44.840 ;
        RECT 23.270 44.690 23.650 44.700 ;
        RECT 25.825 44.690 26.155 44.705 ;
        RECT 23.270 44.390 26.155 44.690 ;
        RECT 23.270 44.380 23.650 44.390 ;
        RECT 25.825 44.375 26.155 44.390 ;
        RECT 24.350 43.355 25.930 43.685 ;
        RECT 13.865 41.290 14.195 41.305 ;
        RECT 4.000 40.990 14.195 41.290 ;
        RECT 13.865 40.975 14.195 40.990 ;
        RECT 82.865 41.290 83.195 41.305 ;
        RECT 82.865 40.990 86.000 41.290 ;
        RECT 82.865 40.975 83.195 40.990 ;
        RECT 21.050 40.635 22.630 40.965 ;
        RECT 24.350 37.915 25.930 38.245 ;
        RECT 14.785 37.890 15.115 37.905 ;
        RECT 4.000 37.590 15.115 37.890 ;
        RECT 14.785 37.575 15.115 37.590 ;
        RECT 12.025 36.530 12.355 36.545 ;
        RECT 41.925 36.530 42.255 36.545 ;
        RECT 12.025 36.230 42.255 36.530 ;
        RECT 12.025 36.215 12.355 36.230 ;
        RECT 41.925 36.215 42.255 36.230 ;
        RECT 21.050 35.195 22.630 35.525 ;
        RECT 24.350 32.475 25.930 32.805 ;
        RECT 69.525 31.770 69.855 31.785 ;
        RECT 74.125 31.770 74.455 31.785 ;
        RECT 69.525 31.470 74.455 31.770 ;
        RECT 69.525 31.455 69.855 31.470 ;
        RECT 74.125 31.455 74.455 31.470 ;
        RECT 21.050 29.755 22.630 30.085 ;
        RECT 82.865 27.690 83.195 27.705 ;
        RECT 82.865 27.390 86.000 27.690 ;
        RECT 82.865 27.375 83.195 27.390 ;
        RECT 24.350 27.035 25.930 27.365 ;
        RECT 21.050 24.315 22.630 24.645 ;
        RECT 24.350 21.595 25.930 21.925 ;
        RECT 17.545 20.890 17.875 20.905 ;
        RECT 32.725 20.890 33.055 20.905 ;
        RECT 39.165 20.890 39.495 20.905 ;
        RECT 17.545 20.590 39.495 20.890 ;
        RECT 17.545 20.575 17.875 20.590 ;
        RECT 32.725 20.575 33.055 20.590 ;
        RECT 39.165 20.575 39.495 20.590 ;
        RECT 36.150 20.210 36.530 20.220 ;
        RECT 57.565 20.210 57.895 20.225 ;
        RECT 36.150 19.910 57.895 20.210 ;
        RECT 36.150 19.900 36.530 19.910 ;
        RECT 57.565 19.895 57.895 19.910 ;
        RECT 21.050 18.875 22.630 19.205 ;
        RECT 21.225 18.170 21.555 18.185 ;
        RECT 23.270 18.170 23.650 18.180 ;
        RECT 36.405 18.170 36.735 18.185 ;
        RECT 21.225 17.870 36.735 18.170 ;
        RECT 21.225 17.855 21.555 17.870 ;
        RECT 23.270 17.860 23.650 17.870 ;
        RECT 36.405 17.855 36.735 17.870 ;
        RECT 24.350 16.155 25.930 16.485 ;
        RECT 21.050 13.435 22.630 13.765 ;
        RECT 24.350 10.715 25.930 11.045 ;
      LAYER met4 ;
        RECT 36.175 62.735 36.505 63.065 ;
        RECT 23.295 44.375 23.625 44.705 ;
        RECT 23.310 18.185 23.610 44.375 ;
        RECT 36.190 20.225 36.490 62.735 ;
        RECT 36.175 19.895 36.505 20.225 ;
        RECT 23.295 17.855 23.625 18.185 ;
  END
END main
END LIBRARY

