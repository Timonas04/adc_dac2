MACRO main
  CLASS BLOCK ;
  FOREIGN main ;
  ORIGIN 0.000 0.000 ;
  SIZE 88.945 BY 177.570 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 166.160 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 166.160 ;
    END
  END VPWR
  PIN b0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END b0
  PIN b1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END b1
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END clk
  PIN compr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 84.945 156.440 88.945 157.040 ;
    END
  END compr
  PIN dac[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 17.040 88.945 17.640 ;
    END
  END dac[0]
  PIN dac[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 85.040 88.945 85.640 ;
    END
  END dac[1]
  PIN dac[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 153.040 88.945 153.640 ;
    END
  END dac[2]
  PIN dac[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 91.840 88.945 92.440 ;
    END
  END dac[3]
  PIN dac[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 105.440 88.945 106.040 ;
    END
  END dac[4]
  PIN dac[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 64.640 88.945 65.240 ;
    END
  END dac[5]
  PIN dac[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 68.040 88.945 68.640 ;
    END
  END dac[6]
  PIN dac[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END dac[7]
  PIN dac_coupl
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END dac_coupl
  PIN m0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END m0
  PIN m1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END m1
  PIN reg0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 88.440 88.945 89.040 ;
    END
  END reg0[0]
  PIN reg0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 149.640 88.945 150.240 ;
    END
  END reg0[1]
  PIN reg0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 173.570 74.430 177.570 ;
    END
  END reg0[2]
  PIN reg0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 71.440 88.945 72.040 ;
    END
  END reg0[3]
  PIN reg0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 125.840 88.945 126.440 ;
    END
  END reg0[4]
  PIN reg0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 74.840 88.945 75.440 ;
    END
  END reg0[5]
  PIN reg0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 173.570 77.650 177.570 ;
    END
  END reg0[6]
  PIN reg0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 112.240 88.945 112.840 ;
    END
  END reg0[7]
  PIN reg1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 23.840 88.945 24.440 ;
    END
  END reg1[0]
  PIN reg1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 27.240 88.945 27.840 ;
    END
  END reg1[1]
  PIN reg1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 47.640 88.945 48.240 ;
    END
  END reg1[2]
  PIN reg1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 20.440 88.945 21.040 ;
    END
  END reg1[3]
  PIN reg1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END reg1[4]
  PIN reg1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 61.240 88.945 61.840 ;
    END
  END reg1[5]
  PIN reg1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END reg1[6]
  PIN reg1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END reg1[7]
  PIN reg2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 44.240 88.945 44.840 ;
    END
  END reg2[0]
  PIN reg2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 40.840 88.945 41.440 ;
    END
  END reg2[1]
  PIN reg2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 51.040 88.945 51.640 ;
    END
  END reg2[2]
  PIN reg2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 54.440 88.945 55.040 ;
    END
  END reg2[3]
  PIN reg2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 30.640 88.945 31.240 ;
    END
  END reg2[4]
  PIN reg2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 57.840 88.945 58.440 ;
    END
  END reg2[5]
  PIN reg2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 34.040 88.945 34.640 ;
    END
  END reg2[6]
  PIN reg2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 37.440 88.945 38.040 ;
    END
  END reg2[7]
  PIN reg3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 95.240 88.945 95.840 ;
    END
  END reg3[0]
  PIN reg3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 129.240 88.945 129.840 ;
    END
  END reg3[1]
  PIN reg3[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 142.840 88.945 143.440 ;
    END
  END reg3[2]
  PIN reg3[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 108.840 88.945 109.440 ;
    END
  END reg3[3]
  PIN reg3[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 122.440 88.945 123.040 ;
    END
  END reg3[4]
  PIN reg3[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 78.240 88.945 78.840 ;
    END
  END reg3[5]
  PIN reg3[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 139.440 88.945 140.040 ;
    END
  END reg3[6]
  PIN reg3[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 115.640 88.945 116.240 ;
    END
  END reg3[7]
  PIN reg4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 98.640 88.945 99.240 ;
    END
  END reg4[0]
  PIN reg4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 132.640 88.945 133.240 ;
    END
  END reg4[1]
  PIN reg4[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 173.570 64.770 177.570 ;
    END
  END reg4[2]
  PIN reg4[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 102.040 88.945 102.640 ;
    END
  END reg4[3]
  PIN reg4[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 119.040 88.945 119.640 ;
    END
  END reg4[4]
  PIN reg4[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 81.640 88.945 82.240 ;
    END
  END reg4[5]
  PIN reg4[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 173.570 67.990 177.570 ;
    END
  END reg4[6]
  PIN reg4[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 136.040 88.945 136.640 ;
    END
  END reg4[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 84.945 146.240 88.945 146.840 ;
    END
  END rst
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END rx
  PIN tx
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 173.570 39.010 177.570 ;
    END
  END tx
  OBS
      LAYER nwell ;
        RECT 5.330 164.505 83.450 166.110 ;
      LAYER pwell ;
        RECT 5.525 163.305 6.895 164.115 ;
        RECT 6.905 163.305 12.415 164.115 ;
        RECT 12.425 163.305 17.935 164.115 ;
        RECT 18.415 163.390 18.845 164.175 ;
        RECT 18.865 163.305 24.375 164.115 ;
        RECT 24.385 163.305 29.895 164.115 ;
        RECT 29.905 163.305 31.275 164.115 ;
        RECT 31.295 163.390 31.725 164.175 ;
        RECT 31.745 163.305 37.255 164.115 ;
        RECT 37.265 163.305 39.095 164.115 ;
        RECT 39.105 163.985 40.450 164.215 ;
        RECT 39.105 163.305 40.935 163.985 ;
        RECT 40.945 163.305 43.695 164.115 ;
        RECT 44.175 163.390 44.605 164.175 ;
        RECT 44.625 163.305 50.135 164.115 ;
        RECT 50.145 163.305 51.515 164.115 ;
        RECT 51.525 163.985 52.870 164.215 ;
        RECT 53.365 163.985 54.710 164.215 ;
        RECT 55.205 163.985 56.550 164.215 ;
        RECT 51.525 163.305 53.355 163.985 ;
        RECT 53.365 163.305 55.195 163.985 ;
        RECT 55.205 163.305 57.035 163.985 ;
        RECT 57.055 163.390 57.485 164.175 ;
        RECT 57.990 163.985 59.335 164.215 ;
        RECT 57.505 163.305 59.335 163.985 ;
        RECT 59.345 163.985 60.690 164.215 ;
        RECT 61.495 163.985 62.425 164.215 ;
        RECT 63.795 163.985 64.725 164.215 ;
        RECT 66.095 163.985 67.025 164.215 ;
        RECT 68.085 163.985 69.430 164.215 ;
        RECT 59.345 163.305 61.175 163.985 ;
        RECT 61.495 163.305 63.330 163.985 ;
        RECT 63.795 163.305 65.630 163.985 ;
        RECT 66.095 163.305 67.930 163.985 ;
        RECT 68.085 163.305 69.915 163.985 ;
        RECT 69.935 163.390 70.365 164.175 ;
        RECT 71.435 163.985 72.365 164.215 ;
        RECT 73.735 163.985 74.665 164.215 ;
        RECT 76.035 163.985 76.965 164.215 ;
        RECT 70.530 163.305 72.365 163.985 ;
        RECT 72.830 163.305 74.665 163.985 ;
        RECT 75.130 163.305 76.965 163.985 ;
        RECT 77.745 163.305 80.955 164.215 ;
        RECT 81.885 163.305 83.255 164.115 ;
        RECT 5.665 163.095 5.835 163.305 ;
        RECT 7.045 163.095 7.215 163.305 ;
        RECT 12.565 163.095 12.735 163.305 ;
        RECT 18.085 163.255 18.255 163.285 ;
        RECT 18.080 163.145 18.255 163.255 ;
        RECT 18.085 163.095 18.255 163.145 ;
        RECT 19.005 163.115 19.175 163.305 ;
        RECT 23.605 163.095 23.775 163.285 ;
        RECT 24.525 163.115 24.695 163.305 ;
        RECT 29.125 163.095 29.295 163.285 ;
        RECT 30.045 163.115 30.215 163.305 ;
        RECT 30.960 163.145 31.080 163.255 ;
        RECT 31.885 163.095 32.055 163.305 ;
        RECT 33.720 163.095 33.890 163.285 ;
        RECT 37.405 163.095 37.575 163.305 ;
        RECT 40.625 163.115 40.795 163.305 ;
        RECT 41.085 163.115 41.255 163.305 ;
        RECT 44.765 163.285 44.935 163.305 ;
        RECT 42.925 163.095 43.095 163.285 ;
        RECT 43.840 163.145 43.960 163.255 ;
        RECT 44.760 163.115 44.935 163.285 ;
        RECT 44.760 163.095 44.930 163.115 ;
        RECT 46.145 163.095 46.315 163.285 ;
        RECT 50.285 163.115 50.455 163.305 ;
        RECT 53.045 163.095 53.215 163.305 ;
        RECT 53.505 163.095 53.675 163.285 ;
        RECT 54.885 163.115 55.055 163.305 ;
        RECT 56.725 163.115 56.895 163.305 ;
        RECT 57.645 163.115 57.815 163.305 ;
        RECT 60.865 163.095 61.035 163.305 ;
        RECT 63.165 163.285 63.330 163.305 ;
        RECT 65.465 163.285 65.630 163.305 ;
        RECT 67.765 163.285 67.930 163.305 ;
        RECT 61.335 163.140 61.495 163.250 ;
        RECT 63.165 163.115 63.335 163.285 ;
        RECT 65.465 163.115 65.635 163.285 ;
        RECT 67.765 163.115 67.935 163.285 ;
        RECT 69.145 163.095 69.315 163.285 ;
        RECT 69.605 163.115 69.775 163.305 ;
        RECT 70.530 163.285 70.695 163.305 ;
        RECT 72.830 163.285 72.995 163.305 ;
        RECT 75.130 163.285 75.295 163.305 ;
        RECT 70.525 163.115 70.700 163.285 ;
        RECT 72.825 163.115 72.995 163.285 ;
        RECT 70.530 163.095 70.700 163.115 ;
        RECT 74.210 163.095 74.380 163.285 ;
        RECT 75.125 163.115 75.295 163.285 ;
        RECT 77.420 163.145 77.540 163.255 ;
        RECT 77.885 163.115 78.055 163.305 ;
        RECT 80.645 163.095 80.815 163.285 ;
        RECT 81.115 163.140 81.275 163.260 ;
        RECT 82.945 163.095 83.115 163.305 ;
        RECT 5.525 162.285 6.895 163.095 ;
        RECT 6.905 162.285 12.415 163.095 ;
        RECT 12.425 162.285 17.935 163.095 ;
        RECT 17.945 162.285 23.455 163.095 ;
        RECT 23.465 162.285 28.975 163.095 ;
        RECT 28.985 162.285 30.815 163.095 ;
        RECT 31.295 162.225 31.725 163.010 ;
        RECT 31.745 162.285 33.575 163.095 ;
        RECT 33.595 162.185 37.255 163.095 ;
        RECT 37.265 162.285 42.775 163.095 ;
        RECT 42.785 162.285 44.615 163.095 ;
        RECT 44.645 162.185 45.995 163.095 ;
        RECT 46.005 162.285 51.515 163.095 ;
        RECT 51.525 162.415 53.355 163.095 ;
        RECT 53.475 162.415 56.940 163.095 ;
        RECT 51.525 162.185 52.870 162.415 ;
        RECT 56.020 162.185 56.940 162.415 ;
        RECT 57.055 162.225 57.485 163.010 ;
        RECT 57.600 162.415 61.065 163.095 ;
        RECT 62.145 162.415 69.455 163.095 ;
        RECT 57.600 162.185 58.520 162.415 ;
        RECT 62.145 162.185 63.495 162.415 ;
        RECT 65.030 162.195 65.940 162.415 ;
        RECT 70.385 162.185 73.860 163.095 ;
        RECT 74.065 162.185 77.540 163.095 ;
        RECT 77.745 162.185 80.955 163.095 ;
        RECT 81.885 162.285 83.255 163.095 ;
      LAYER nwell ;
        RECT 5.330 159.065 83.450 161.895 ;
      LAYER pwell ;
        RECT 5.525 157.865 6.895 158.675 ;
        RECT 6.905 157.865 12.415 158.675 ;
        RECT 12.425 157.865 17.935 158.675 ;
        RECT 18.415 157.950 18.845 158.735 ;
        RECT 18.865 157.865 24.375 158.675 ;
        RECT 24.385 157.865 29.895 158.675 ;
        RECT 29.905 157.865 31.735 158.675 ;
        RECT 35.720 158.545 36.630 158.765 ;
        RECT 38.165 158.545 39.515 158.775 ;
        RECT 32.205 157.865 39.515 158.545 ;
        RECT 39.875 158.545 40.805 158.775 ;
        RECT 39.875 157.865 41.710 158.545 ;
        RECT 41.865 157.865 43.695 158.775 ;
        RECT 44.175 157.950 44.605 158.735 ;
        RECT 44.720 158.545 45.640 158.775 ;
        RECT 51.820 158.545 52.730 158.765 ;
        RECT 54.265 158.545 55.615 158.775 ;
        RECT 44.720 157.865 48.185 158.545 ;
        RECT 48.305 157.865 55.615 158.545 ;
        RECT 55.665 158.545 56.595 158.775 ;
        RECT 60.765 158.545 62.115 158.775 ;
        RECT 63.650 158.545 64.560 158.765 ;
        RECT 68.570 158.545 69.915 158.775 ;
        RECT 55.665 157.865 59.565 158.545 ;
        RECT 60.765 157.865 68.075 158.545 ;
        RECT 68.085 157.865 69.915 158.545 ;
        RECT 69.935 157.950 70.365 158.735 ;
        RECT 73.900 158.545 74.810 158.765 ;
        RECT 76.345 158.545 77.695 158.775 ;
        RECT 70.385 157.865 77.695 158.545 ;
        RECT 78.205 157.865 81.415 158.775 ;
        RECT 81.885 157.865 83.255 158.675 ;
        RECT 5.665 157.655 5.835 157.865 ;
        RECT 7.045 157.655 7.215 157.865 ;
        RECT 12.565 157.655 12.735 157.865 ;
        RECT 18.085 157.815 18.255 157.845 ;
        RECT 18.080 157.705 18.255 157.815 ;
        RECT 18.085 157.655 18.255 157.705 ;
        RECT 19.005 157.675 19.175 157.865 ;
        RECT 23.605 157.655 23.775 157.845 ;
        RECT 24.525 157.675 24.695 157.865 ;
        RECT 29.125 157.655 29.295 157.845 ;
        RECT 30.045 157.675 30.215 157.865 ;
        RECT 31.885 157.815 32.055 157.845 ;
        RECT 30.960 157.705 31.080 157.815 ;
        RECT 31.880 157.705 32.055 157.815 ;
        RECT 31.885 157.655 32.055 157.705 ;
        RECT 32.345 157.675 32.515 157.865 ;
        RECT 41.545 157.845 41.710 157.865 ;
        RECT 36.945 157.655 37.115 157.845 ;
        RECT 37.410 157.655 37.580 157.845 ;
        RECT 41.085 157.655 41.255 157.845 ;
        RECT 41.545 157.675 41.715 157.845 ;
        RECT 43.380 157.675 43.550 157.865 ;
        RECT 43.840 157.705 43.960 157.815 ;
        RECT 47.985 157.675 48.155 157.865 ;
        RECT 48.445 157.655 48.615 157.865 ;
        RECT 55.805 157.655 55.975 157.845 ;
        RECT 56.080 157.675 56.250 157.865 ;
        RECT 59.955 157.710 60.115 157.820 ;
        RECT 64.545 157.655 64.715 157.845 ;
        RECT 67.305 157.655 67.475 157.845 ;
        RECT 67.765 157.655 67.935 157.865 ;
        RECT 68.225 157.675 68.395 157.865 ;
        RECT 70.525 157.675 70.695 157.865 ;
        RECT 75.125 157.675 75.295 157.845 ;
        RECT 77.880 157.705 78.000 157.815 ;
        RECT 78.345 157.675 78.515 157.865 ;
        RECT 81.590 157.815 81.760 157.845 ;
        RECT 81.560 157.705 81.760 157.815 ;
        RECT 81.590 157.675 81.760 157.705 ;
        RECT 75.130 157.655 75.295 157.675 ;
        RECT 81.590 157.655 81.700 157.675 ;
        RECT 82.945 157.655 83.115 157.865 ;
        RECT 5.525 156.845 6.895 157.655 ;
        RECT 6.905 156.845 12.415 157.655 ;
        RECT 12.425 156.845 17.935 157.655 ;
        RECT 17.945 156.845 23.455 157.655 ;
        RECT 23.465 156.845 28.975 157.655 ;
        RECT 28.985 156.845 30.815 157.655 ;
        RECT 31.295 156.785 31.725 157.570 ;
        RECT 31.745 156.845 33.575 157.655 ;
        RECT 33.680 156.975 37.145 157.655 ;
        RECT 37.265 156.975 40.850 157.655 ;
        RECT 40.945 156.975 48.255 157.655 ;
        RECT 48.305 156.975 55.615 157.655 ;
        RECT 33.680 156.745 34.600 156.975 ;
        RECT 37.265 156.745 38.185 156.975 ;
        RECT 44.460 156.755 45.370 156.975 ;
        RECT 46.905 156.745 48.255 156.975 ;
        RECT 51.820 156.755 52.730 156.975 ;
        RECT 54.265 156.745 55.615 156.975 ;
        RECT 55.665 156.845 57.035 157.655 ;
        RECT 57.055 156.785 57.485 157.570 ;
        RECT 57.545 156.975 64.855 157.655 ;
        RECT 64.875 156.975 67.615 157.655 ;
        RECT 67.625 156.975 74.935 157.655 ;
        RECT 75.130 156.975 76.965 157.655 ;
        RECT 57.545 156.745 58.895 156.975 ;
        RECT 60.430 156.755 61.340 156.975 ;
        RECT 71.140 156.755 72.050 156.975 ;
        RECT 73.585 156.745 74.935 156.975 ;
        RECT 76.035 156.745 76.965 156.975 ;
        RECT 77.285 156.975 81.700 157.655 ;
        RECT 77.285 156.745 81.215 156.975 ;
        RECT 81.885 156.845 83.255 157.655 ;
      LAYER nwell ;
        RECT 5.330 153.625 83.450 156.455 ;
      LAYER pwell ;
        RECT 5.525 152.425 6.895 153.235 ;
        RECT 6.905 152.425 12.415 153.235 ;
        RECT 12.425 152.425 17.935 153.235 ;
        RECT 18.415 152.510 18.845 153.295 ;
        RECT 18.865 152.425 24.375 153.235 ;
        RECT 24.385 152.425 29.895 153.235 ;
        RECT 30.405 153.105 31.755 153.335 ;
        RECT 33.290 153.105 34.200 153.325 ;
        RECT 38.865 153.245 39.815 153.335 ;
        RECT 30.405 152.425 37.715 153.105 ;
        RECT 37.885 152.425 39.815 153.245 ;
        RECT 40.195 152.425 43.695 153.335 ;
        RECT 44.175 152.510 44.605 153.295 ;
        RECT 44.625 152.425 47.835 153.335 ;
        RECT 47.845 153.135 48.790 153.335 ;
        RECT 47.845 152.455 50.595 153.135 ;
        RECT 50.605 153.105 51.535 153.335 ;
        RECT 58.260 153.105 59.170 153.325 ;
        RECT 60.705 153.105 62.055 153.335 ;
        RECT 47.845 152.425 48.790 152.455 ;
        RECT 5.665 152.215 5.835 152.425 ;
        RECT 7.045 152.215 7.215 152.425 ;
        RECT 12.565 152.215 12.735 152.425 ;
        RECT 18.085 152.375 18.255 152.405 ;
        RECT 18.080 152.265 18.255 152.375 ;
        RECT 18.085 152.215 18.255 152.265 ;
        RECT 19.005 152.235 19.175 152.425 ;
        RECT 23.605 152.215 23.775 152.405 ;
        RECT 24.525 152.235 24.695 152.425 ;
        RECT 27.280 152.215 27.450 152.405 ;
        RECT 28.665 152.215 28.835 152.405 ;
        RECT 30.040 152.265 30.160 152.375 ;
        RECT 31.885 152.215 32.055 152.405 ;
        RECT 37.405 152.235 37.575 152.425 ;
        RECT 37.885 152.405 38.035 152.425 ;
        RECT 40.195 152.405 40.330 152.425 ;
        RECT 37.865 152.235 38.035 152.405 ;
        RECT 39.240 152.265 39.360 152.375 ;
        RECT 39.705 152.215 39.875 152.405 ;
        RECT 40.160 152.235 40.330 152.405 ;
        RECT 43.840 152.265 43.960 152.375 ;
        RECT 44.755 152.235 44.925 152.425 ;
        RECT 5.525 151.405 6.895 152.215 ;
        RECT 6.905 151.405 12.415 152.215 ;
        RECT 12.425 151.405 17.935 152.215 ;
        RECT 17.945 151.405 23.455 152.215 ;
        RECT 23.465 151.405 27.135 152.215 ;
        RECT 27.165 151.305 28.515 152.215 ;
        RECT 28.535 151.305 31.265 152.215 ;
        RECT 31.295 151.345 31.725 152.130 ;
        RECT 31.745 151.535 39.055 152.215 ;
        RECT 39.565 151.535 46.875 152.215 ;
        RECT 47.070 152.185 47.240 152.405 ;
        RECT 50.280 152.235 50.450 152.455 ;
        RECT 50.605 152.425 54.505 153.105 ;
        RECT 54.745 152.425 62.055 153.105 ;
        RECT 62.105 153.105 63.035 153.335 ;
        RECT 66.340 153.105 67.260 153.335 ;
        RECT 62.105 152.425 66.005 153.105 ;
        RECT 66.340 152.425 69.805 153.105 ;
        RECT 69.935 152.510 70.365 153.295 ;
        RECT 70.385 152.425 73.860 153.335 ;
        RECT 78.040 153.105 78.950 153.325 ;
        RECT 80.485 153.105 81.835 153.335 ;
        RECT 74.525 152.425 81.835 153.105 ;
        RECT 81.885 152.425 83.255 153.235 ;
        RECT 51.020 152.235 51.190 152.425 ;
        RECT 49.645 152.185 50.595 152.215 ;
        RECT 35.260 151.315 36.170 151.535 ;
        RECT 37.705 151.305 39.055 151.535 ;
        RECT 43.080 151.315 43.990 151.535 ;
        RECT 45.525 151.305 46.875 151.535 ;
        RECT 46.925 151.505 50.595 152.185 ;
        RECT 49.645 151.305 50.595 151.505 ;
        RECT 50.605 152.185 51.540 152.215 ;
        RECT 53.500 152.185 53.670 152.405 ;
        RECT 54.885 152.235 55.055 152.425 ;
        RECT 56.265 152.215 56.435 152.405 ;
        RECT 56.720 152.265 56.840 152.375 ;
        RECT 57.920 152.215 58.090 152.405 ;
        RECT 62.060 152.215 62.230 152.405 ;
        RECT 62.520 152.235 62.690 152.425 ;
        RECT 69.605 152.405 69.775 152.425 ;
        RECT 69.145 152.215 69.315 152.405 ;
        RECT 69.605 152.235 69.780 152.405 ;
        RECT 70.530 152.235 70.700 152.425 ;
        RECT 74.205 152.375 74.375 152.405 ;
        RECT 74.200 152.265 74.375 152.375 ;
        RECT 69.610 152.215 69.780 152.235 ;
        RECT 74.205 152.215 74.375 152.265 ;
        RECT 74.665 152.215 74.835 152.425 ;
        RECT 82.945 152.215 83.115 152.425 ;
        RECT 50.605 151.985 53.670 152.185 ;
        RECT 50.605 151.505 53.815 151.985 ;
        RECT 50.605 151.305 51.555 151.505 ;
        RECT 52.885 151.305 53.815 151.505 ;
        RECT 53.825 151.535 56.575 152.215 ;
        RECT 53.825 151.305 54.755 151.535 ;
        RECT 57.055 151.345 57.485 152.130 ;
        RECT 57.505 151.535 61.405 152.215 ;
        RECT 61.645 151.535 65.545 152.215 ;
        RECT 65.880 151.535 69.345 152.215 ;
        RECT 57.505 151.305 58.435 151.535 ;
        RECT 61.645 151.305 62.575 151.535 ;
        RECT 65.880 151.305 66.800 151.535 ;
        RECT 69.465 151.305 72.940 152.215 ;
        RECT 73.145 151.435 74.515 152.215 ;
        RECT 74.525 151.535 81.835 152.215 ;
        RECT 78.040 151.315 78.950 151.535 ;
        RECT 80.485 151.305 81.835 151.535 ;
        RECT 81.885 151.405 83.255 152.215 ;
      LAYER nwell ;
        RECT 5.330 148.185 83.450 151.015 ;
      LAYER pwell ;
        RECT 5.525 146.985 6.895 147.795 ;
        RECT 6.905 146.985 12.415 147.795 ;
        RECT 12.425 146.985 17.935 147.795 ;
        RECT 18.415 147.070 18.845 147.855 ;
        RECT 18.865 146.985 24.375 147.795 ;
        RECT 24.385 146.985 28.055 147.795 ;
        RECT 28.525 147.695 29.480 147.895 ;
        RECT 28.525 147.015 30.805 147.695 ;
        RECT 31.875 147.665 32.805 147.895 ;
        RECT 28.525 146.985 29.480 147.015 ;
        RECT 5.665 146.775 5.835 146.985 ;
        RECT 7.045 146.775 7.215 146.985 ;
        RECT 12.565 146.775 12.735 146.985 ;
        RECT 18.085 146.935 18.255 146.965 ;
        RECT 18.080 146.825 18.255 146.935 ;
        RECT 18.085 146.775 18.255 146.825 ;
        RECT 19.005 146.795 19.175 146.985 ;
        RECT 23.605 146.775 23.775 146.965 ;
        RECT 24.525 146.795 24.695 146.985 ;
        RECT 28.200 146.825 28.320 146.935 ;
        RECT 29.125 146.775 29.295 146.965 ;
        RECT 30.510 146.795 30.680 147.015 ;
        RECT 30.970 146.985 32.805 147.665 ;
        RECT 33.125 147.695 34.070 147.895 ;
        RECT 35.405 147.695 36.335 147.895 ;
        RECT 33.125 147.215 36.335 147.695 ;
        RECT 36.440 147.665 37.360 147.895 ;
        RECT 42.680 147.665 43.600 147.895 ;
        RECT 33.125 147.015 36.195 147.215 ;
        RECT 33.125 146.985 34.070 147.015 ;
        RECT 30.970 146.965 31.135 146.985 ;
        RECT 30.965 146.935 31.135 146.965 ;
        RECT 30.960 146.825 31.135 146.935 ;
        RECT 30.965 146.795 31.135 146.825 ;
        RECT 31.895 146.820 32.055 146.930 ;
        RECT 32.810 146.775 32.980 146.965 ;
        RECT 36.025 146.935 36.195 147.015 ;
        RECT 36.440 146.985 39.905 147.665 ;
        RECT 40.135 146.985 43.600 147.665 ;
        RECT 44.175 147.070 44.605 147.855 ;
        RECT 44.625 146.985 45.975 147.895 ;
        RECT 46.005 146.985 49.480 147.895 ;
        RECT 49.685 147.695 50.635 147.895 ;
        RECT 51.965 147.695 52.895 147.895 ;
        RECT 49.685 147.215 52.895 147.695 ;
        RECT 52.905 147.665 53.835 147.895 ;
        RECT 49.685 147.015 52.750 147.215 ;
        RECT 49.685 146.985 50.620 147.015 ;
        RECT 36.020 146.825 36.195 146.935 ;
        RECT 36.025 146.795 36.195 146.825 ;
        RECT 39.705 146.795 39.875 146.985 ;
        RECT 40.165 146.795 40.335 146.985 ;
        RECT 43.385 146.775 43.555 146.965 ;
        RECT 43.845 146.935 44.015 146.965 ;
        RECT 43.840 146.825 44.015 146.935 ;
        RECT 43.845 146.775 44.015 146.825 ;
        RECT 45.690 146.795 45.860 146.985 ;
        RECT 46.150 146.795 46.320 146.985 ;
        RECT 46.615 146.820 46.775 146.930 ;
        RECT 47.525 146.775 47.695 146.965 ;
        RECT 52.580 146.795 52.750 147.015 ;
        RECT 52.905 146.985 55.655 147.665 ;
        RECT 55.665 146.985 58.875 147.895 ;
        RECT 58.885 147.665 59.815 147.895 ;
        RECT 63.025 147.665 63.955 147.895 ;
        RECT 68.675 147.665 69.605 147.895 ;
        RECT 58.885 146.985 62.785 147.665 ;
        RECT 63.025 146.985 66.925 147.665 ;
        RECT 67.770 146.985 69.605 147.665 ;
        RECT 69.935 147.070 70.365 147.855 ;
        RECT 70.480 147.665 71.400 147.895 ;
        RECT 70.480 146.985 73.945 147.665 ;
        RECT 74.065 146.985 77.540 147.895 ;
        RECT 77.745 146.985 81.220 147.895 ;
        RECT 81.885 146.985 83.255 147.795 ;
        RECT 55.345 146.795 55.515 146.985 ;
        RECT 55.795 146.795 55.965 146.985 ;
        RECT 56.725 146.775 56.895 146.965 ;
        RECT 59.300 146.795 59.470 146.985 ;
        RECT 60.865 146.775 61.035 146.965 ;
        RECT 61.325 146.775 61.495 146.965 ;
        RECT 63.440 146.795 63.610 146.985 ;
        RECT 67.770 146.965 67.935 146.985 ;
        RECT 67.300 146.825 67.420 146.935 ;
        RECT 67.765 146.795 67.935 146.965 ;
        RECT 71.905 146.775 72.075 146.965 ;
        RECT 72.355 146.775 72.525 146.965 ;
        RECT 73.745 146.795 73.915 146.985 ;
        RECT 74.210 146.795 74.380 146.985 ;
        RECT 75.585 146.775 75.755 146.965 ;
        RECT 77.415 146.775 77.585 146.965 ;
        RECT 77.890 146.795 78.060 146.985 ;
        RECT 81.555 146.775 81.725 146.965 ;
        RECT 82.945 146.775 83.115 146.985 ;
        RECT 5.525 145.965 6.895 146.775 ;
        RECT 6.905 145.965 12.415 146.775 ;
        RECT 12.425 145.965 17.935 146.775 ;
        RECT 17.945 145.965 23.455 146.775 ;
        RECT 23.465 145.965 28.975 146.775 ;
        RECT 28.985 145.965 30.815 146.775 ;
        RECT 31.295 145.905 31.725 146.690 ;
        RECT 32.665 145.865 35.585 146.775 ;
        RECT 36.385 146.095 43.695 146.775 ;
        RECT 36.385 145.865 37.735 146.095 ;
        RECT 39.270 145.875 40.180 146.095 ;
        RECT 43.715 145.865 46.445 146.775 ;
        RECT 47.385 146.095 54.695 146.775 ;
        RECT 50.900 145.875 51.810 146.095 ;
        RECT 53.345 145.865 54.695 146.095 ;
        RECT 54.745 146.095 57.035 146.775 ;
        RECT 54.745 145.865 55.665 146.095 ;
        RECT 57.055 145.905 57.485 146.690 ;
        RECT 57.600 146.095 61.065 146.775 ;
        RECT 61.185 146.095 68.495 146.775 ;
        RECT 57.600 145.865 58.520 146.095 ;
        RECT 64.700 145.875 65.610 146.095 ;
        RECT 67.145 145.865 68.495 146.095 ;
        RECT 68.640 146.095 72.105 146.775 ;
        RECT 68.640 145.865 69.560 146.095 ;
        RECT 72.225 145.865 75.435 146.775 ;
        RECT 75.445 146.095 77.275 146.775 ;
        RECT 75.930 145.865 77.275 146.095 ;
        RECT 77.285 145.865 80.495 146.775 ;
        RECT 80.505 145.995 81.875 146.775 ;
        RECT 81.885 145.965 83.255 146.775 ;
      LAYER nwell ;
        RECT 5.330 142.745 83.450 145.575 ;
      LAYER pwell ;
        RECT 5.525 141.545 6.895 142.355 ;
        RECT 6.905 141.545 12.415 142.355 ;
        RECT 12.425 141.545 16.095 142.355 ;
        RECT 16.565 141.545 18.395 142.225 ;
        RECT 18.415 141.630 18.845 142.415 ;
        RECT 18.865 141.545 24.375 142.355 ;
        RECT 24.385 141.545 29.895 142.355 ;
        RECT 29.905 141.545 33.575 142.355 ;
        RECT 33.595 141.545 34.945 142.455 ;
        RECT 34.965 141.545 36.315 142.455 ;
        RECT 36.345 141.545 37.715 142.355 ;
        RECT 37.820 142.225 38.740 142.455 ;
        RECT 37.820 141.545 41.285 142.225 ;
        RECT 41.405 141.545 42.775 142.355 ;
        RECT 42.805 141.545 44.155 142.455 ;
        RECT 44.175 141.630 44.605 142.415 ;
        RECT 45.995 142.225 46.915 142.455 ;
        RECT 44.625 141.545 46.915 142.225 ;
        RECT 46.925 141.545 48.755 142.355 ;
        RECT 48.765 142.225 50.110 142.455 ;
        RECT 50.605 142.225 51.535 142.455 ;
        RECT 48.765 141.545 50.595 142.225 ;
        RECT 50.605 141.545 54.505 142.225 ;
        RECT 54.745 141.545 56.835 142.355 ;
        RECT 60.620 142.225 61.540 142.455 ;
        RECT 65.160 142.225 66.070 142.445 ;
        RECT 67.605 142.225 68.955 142.455 ;
        RECT 58.075 141.545 61.540 142.225 ;
        RECT 61.645 141.545 68.955 142.225 ;
        RECT 69.935 141.630 70.365 142.415 ;
        RECT 70.580 141.545 74.055 142.455 ;
        RECT 78.040 142.225 78.950 142.445 ;
        RECT 80.485 142.225 81.835 142.455 ;
        RECT 74.525 141.545 81.835 142.225 ;
        RECT 81.885 141.545 83.255 142.355 ;
        RECT 5.665 141.335 5.835 141.545 ;
        RECT 7.045 141.335 7.215 141.545 ;
        RECT 12.565 141.335 12.735 141.545 ;
        RECT 13.945 141.335 14.115 141.525 ;
        RECT 16.240 141.385 16.360 141.495 ;
        RECT 18.085 141.355 18.255 141.545 ;
        RECT 19.005 141.355 19.175 141.545 ;
        RECT 21.310 141.335 21.480 141.525 ;
        RECT 22.685 141.335 22.855 141.525 ;
        RECT 24.525 141.355 24.695 141.545 ;
        RECT 28.205 141.335 28.375 141.525 ;
        RECT 30.045 141.355 30.215 141.545 ;
        RECT 33.725 141.525 33.895 141.545 ;
        RECT 30.960 141.385 31.080 141.495 ;
        RECT 31.885 141.335 32.055 141.525 ;
        RECT 33.720 141.355 33.895 141.525 ;
        RECT 33.720 141.335 33.890 141.355 ;
        RECT 35.110 141.335 35.280 141.525 ;
        RECT 36.030 141.355 36.200 141.545 ;
        RECT 36.485 141.355 36.655 141.545 ;
        RECT 40.625 141.355 40.795 141.525 ;
        RECT 41.085 141.355 41.255 141.545 ;
        RECT 41.545 141.355 41.715 141.545 ;
        RECT 40.625 141.335 40.790 141.355 ;
        RECT 41.995 141.335 42.165 141.525 ;
        RECT 42.465 141.335 42.635 141.525 ;
        RECT 43.840 141.355 44.010 141.545 ;
        RECT 44.120 141.335 44.290 141.525 ;
        RECT 44.765 141.355 44.935 141.545 ;
        RECT 47.065 141.355 47.235 141.545 ;
        RECT 47.985 141.335 48.155 141.525 ;
        RECT 50.285 141.355 50.455 141.545 ;
        RECT 51.020 141.355 51.190 141.545 ;
        RECT 51.665 141.335 51.835 141.525 ;
        RECT 53.320 141.335 53.490 141.525 ;
        RECT 54.885 141.355 55.055 141.545 ;
        RECT 57.640 141.385 57.760 141.495 ;
        RECT 58.105 141.355 58.275 141.545 ;
        RECT 61.785 141.355 61.955 141.545 ;
        RECT 64.545 141.335 64.715 141.525 ;
        RECT 65.280 141.335 65.450 141.525 ;
        RECT 69.155 141.390 69.315 141.500 ;
        RECT 72.365 141.335 72.535 141.525 ;
        RECT 73.740 141.355 73.910 141.545 ;
        RECT 74.200 141.385 74.320 141.495 ;
        RECT 74.665 141.355 74.835 141.545 ;
        RECT 76.045 141.335 76.215 141.525 ;
        RECT 76.510 141.335 76.680 141.525 ;
        RECT 80.185 141.335 80.355 141.525 ;
        RECT 82.945 141.335 83.115 141.545 ;
        RECT 5.525 140.525 6.895 141.335 ;
        RECT 6.905 140.525 12.415 141.335 ;
        RECT 12.425 140.525 13.795 141.335 ;
        RECT 13.805 140.655 21.115 141.335 ;
        RECT 17.320 140.435 18.230 140.655 ;
        RECT 19.765 140.425 21.115 140.655 ;
        RECT 21.165 140.425 22.515 141.335 ;
        RECT 22.545 140.525 28.055 141.335 ;
        RECT 28.065 140.525 30.815 141.335 ;
        RECT 31.295 140.465 31.725 141.250 ;
        RECT 31.745 140.525 33.575 141.335 ;
        RECT 33.605 140.425 34.955 141.335 ;
        RECT 34.965 140.655 38.550 141.335 ;
        RECT 38.955 140.655 40.790 141.335 ;
        RECT 34.965 140.425 35.885 140.655 ;
        RECT 38.955 140.425 39.885 140.655 ;
        RECT 40.945 140.555 42.315 141.335 ;
        RECT 42.325 140.525 43.695 141.335 ;
        RECT 43.705 140.655 47.605 141.335 ;
        RECT 43.705 140.425 44.635 140.655 ;
        RECT 47.845 140.525 51.515 141.335 ;
        RECT 51.525 140.525 52.895 141.335 ;
        RECT 52.905 140.655 56.805 141.335 ;
        RECT 52.905 140.425 53.835 140.655 ;
        RECT 57.055 140.465 57.485 141.250 ;
        RECT 57.545 140.655 64.855 141.335 ;
        RECT 64.865 140.655 68.765 141.335 ;
        RECT 69.100 140.655 72.565 141.335 ;
        RECT 72.780 140.655 76.245 141.335 ;
        RECT 57.545 140.425 58.895 140.655 ;
        RECT 60.430 140.435 61.340 140.655 ;
        RECT 64.865 140.425 65.795 140.655 ;
        RECT 69.100 140.425 70.020 140.655 ;
        RECT 72.780 140.425 73.700 140.655 ;
        RECT 76.365 140.425 79.840 141.335 ;
        RECT 80.045 140.655 81.875 141.335 ;
        RECT 80.530 140.425 81.875 140.655 ;
        RECT 81.885 140.525 83.255 141.335 ;
      LAYER nwell ;
        RECT 5.330 137.305 83.450 140.135 ;
      LAYER pwell ;
        RECT 5.525 136.105 6.895 136.915 ;
        RECT 6.905 136.105 9.655 136.915 ;
        RECT 13.640 136.785 14.550 137.005 ;
        RECT 16.085 136.785 17.435 137.015 ;
        RECT 10.125 136.105 17.435 136.785 ;
        RECT 18.415 136.190 18.845 136.975 ;
        RECT 18.865 136.105 20.215 137.015 ;
        RECT 23.760 136.785 24.670 137.005 ;
        RECT 26.205 136.785 27.555 137.015 ;
        RECT 31.120 136.785 32.030 137.005 ;
        RECT 33.565 136.785 34.915 137.015 ;
        RECT 20.245 136.105 27.555 136.785 ;
        RECT 27.605 136.105 34.915 136.785 ;
        RECT 35.060 136.785 35.980 137.015 ;
        RECT 35.060 136.105 38.525 136.785 ;
        RECT 38.645 136.105 40.475 136.915 ;
        RECT 40.580 136.785 41.500 137.015 ;
        RECT 40.580 136.105 44.045 136.785 ;
        RECT 44.175 136.190 44.605 136.975 ;
        RECT 44.625 136.105 45.975 137.015 ;
        RECT 46.005 136.105 47.835 136.915 ;
        RECT 51.360 136.785 52.270 137.005 ;
        RECT 53.805 136.785 55.155 137.015 ;
        RECT 47.845 136.105 55.155 136.785 ;
        RECT 55.665 136.785 57.010 137.015 ;
        RECT 60.705 136.785 61.635 137.015 ;
        RECT 55.665 136.105 57.495 136.785 ;
        RECT 57.735 136.105 61.635 136.785 ;
        RECT 61.645 136.785 62.575 137.015 ;
        RECT 65.785 136.785 66.715 137.015 ;
        RECT 61.645 136.105 65.545 136.785 ;
        RECT 65.785 136.105 69.685 136.785 ;
        RECT 69.935 136.190 70.365 136.975 ;
        RECT 73.900 136.785 74.810 137.005 ;
        RECT 76.345 136.785 77.695 137.015 ;
        RECT 70.385 136.105 77.695 136.785 ;
        RECT 77.745 136.105 81.220 137.015 ;
        RECT 81.885 136.105 83.255 136.915 ;
        RECT 5.665 135.895 5.835 136.105 ;
        RECT 7.045 136.055 7.215 136.105 ;
        RECT 7.040 135.945 7.215 136.055 ;
        RECT 7.045 135.915 7.215 135.945 ;
        RECT 8.420 135.895 8.590 136.085 ;
        RECT 8.885 135.895 9.055 136.085 ;
        RECT 9.800 135.945 9.920 136.055 ;
        RECT 10.265 135.915 10.435 136.105 ;
        RECT 12.565 135.895 12.735 136.085 ;
        RECT 16.245 135.895 16.415 136.085 ;
        RECT 17.635 135.950 17.795 136.060 ;
        RECT 19.010 135.915 19.180 136.105 ;
        RECT 20.385 135.915 20.555 136.105 ;
        RECT 23.605 135.895 23.775 136.085 ;
        RECT 27.745 135.915 27.915 136.105 ;
        RECT 31.885 135.895 32.055 136.085 ;
        RECT 38.325 135.915 38.495 136.105 ;
        RECT 38.785 135.915 38.955 136.105 ;
        RECT 39.255 135.940 39.415 136.050 ;
        RECT 40.165 135.895 40.335 136.085 ;
        RECT 43.845 135.915 44.015 136.105 ;
        RECT 44.770 135.915 44.940 136.105 ;
        RECT 46.145 135.915 46.315 136.105 ;
        RECT 47.520 135.945 47.640 136.055 ;
        RECT 47.985 135.915 48.155 136.105 ;
        RECT 48.260 135.895 48.430 136.085 ;
        RECT 55.345 136.055 55.515 136.085 ;
        RECT 55.340 135.945 55.515 136.055 ;
        RECT 55.345 135.895 55.515 135.945 ;
        RECT 55.805 135.895 55.975 136.085 ;
        RECT 57.185 135.915 57.355 136.105 ;
        RECT 61.050 135.915 61.220 136.105 ;
        RECT 62.060 135.915 62.230 136.105 ;
        RECT 62.245 135.895 62.415 136.085 ;
        RECT 62.980 135.895 63.150 136.085 ;
        RECT 66.200 135.915 66.370 136.105 ;
        RECT 66.840 135.945 66.960 136.055 ;
        RECT 70.525 135.915 70.695 136.105 ;
        RECT 74.205 135.895 74.375 136.085 ;
        RECT 74.665 135.895 74.835 136.085 ;
        RECT 77.890 135.915 78.060 136.105 ;
        RECT 81.560 135.945 81.680 136.055 ;
        RECT 82.945 135.895 83.115 136.105 ;
        RECT 5.525 135.085 6.895 135.895 ;
        RECT 7.385 134.985 8.735 135.895 ;
        RECT 8.745 135.215 12.415 135.895 ;
        RECT 12.425 135.215 16.095 135.895 ;
        RECT 16.105 135.215 23.415 135.895 ;
        RECT 23.465 135.215 31.195 135.895 ;
        RECT 11.485 134.985 12.415 135.215 ;
        RECT 15.165 134.985 16.095 135.215 ;
        RECT 19.620 134.995 20.530 135.215 ;
        RECT 22.065 134.985 23.415 135.215 ;
        RECT 26.980 134.995 27.890 135.215 ;
        RECT 29.425 134.985 31.195 135.215 ;
        RECT 31.295 135.025 31.725 135.810 ;
        RECT 31.745 135.215 39.055 135.895 ;
        RECT 40.025 135.215 47.335 135.895 ;
        RECT 35.260 134.995 36.170 135.215 ;
        RECT 37.705 134.985 39.055 135.215 ;
        RECT 43.540 134.995 44.450 135.215 ;
        RECT 45.985 134.985 47.335 135.215 ;
        RECT 47.845 135.215 51.745 135.895 ;
        RECT 52.080 135.215 55.545 135.895 ;
        RECT 47.845 134.985 48.775 135.215 ;
        RECT 52.080 134.985 53.000 135.215 ;
        RECT 55.665 135.085 57.035 135.895 ;
        RECT 57.055 135.025 57.485 135.810 ;
        RECT 57.740 135.215 62.555 135.895 ;
        RECT 62.565 135.215 66.465 135.895 ;
        RECT 67.205 135.215 74.515 135.895 ;
        RECT 74.525 135.215 81.835 135.895 ;
        RECT 62.565 134.985 63.495 135.215 ;
        RECT 67.205 134.985 68.555 135.215 ;
        RECT 70.090 134.995 71.000 135.215 ;
        RECT 78.040 134.995 78.950 135.215 ;
        RECT 80.485 134.985 81.835 135.215 ;
        RECT 81.885 135.085 83.255 135.895 ;
      LAYER nwell ;
        RECT 5.330 131.865 83.450 134.695 ;
      LAYER pwell ;
        RECT 5.525 130.665 6.895 131.475 ;
        RECT 6.905 130.665 9.655 131.475 ;
        RECT 9.665 130.665 12.835 131.575 ;
        RECT 12.885 131.345 13.815 131.575 ;
        RECT 12.885 130.665 16.555 131.345 ;
        RECT 16.565 130.665 18.380 131.575 ;
        RECT 18.415 130.750 18.845 131.535 ;
        RECT 22.525 131.345 23.455 131.575 ;
        RECT 26.205 131.345 27.135 131.575 ;
        RECT 19.785 130.665 23.455 131.345 ;
        RECT 23.465 130.665 27.135 131.345 ;
        RECT 27.145 130.665 28.960 131.575 ;
        RECT 29.000 130.665 30.815 131.575 ;
        RECT 31.305 130.665 32.655 131.575 ;
        RECT 36.180 131.345 37.090 131.565 ;
        RECT 38.625 131.345 39.975 131.575 ;
        RECT 32.665 130.665 39.975 131.345 ;
        RECT 40.025 131.345 40.955 131.575 ;
        RECT 40.025 130.665 43.925 131.345 ;
        RECT 44.175 130.750 44.605 131.535 ;
        RECT 48.140 131.345 49.050 131.565 ;
        RECT 50.585 131.345 51.935 131.575 ;
        RECT 55.500 131.345 56.410 131.565 ;
        RECT 57.945 131.345 59.295 131.575 ;
        RECT 44.625 130.665 51.935 131.345 ;
        RECT 51.985 130.665 59.295 131.345 ;
        RECT 59.385 131.345 60.735 131.575 ;
        RECT 62.270 131.345 63.180 131.565 ;
        RECT 68.675 131.345 69.605 131.575 ;
        RECT 59.385 130.665 66.695 131.345 ;
        RECT 67.770 130.665 69.605 131.345 ;
        RECT 69.935 130.750 70.365 131.535 ;
        RECT 70.480 131.345 71.400 131.575 ;
        RECT 74.160 131.345 75.080 131.575 ;
        RECT 70.480 130.665 73.945 131.345 ;
        RECT 74.160 130.665 77.625 131.345 ;
        RECT 77.745 130.665 81.220 131.575 ;
        RECT 81.885 130.665 83.255 131.475 ;
        RECT 5.665 130.455 5.835 130.665 ;
        RECT 7.045 130.455 7.215 130.665 ;
        RECT 12.565 130.455 12.735 130.665 ;
        RECT 15.320 130.505 15.440 130.615 ;
        RECT 16.245 130.475 16.415 130.665 ;
        RECT 17.625 130.455 17.795 130.645 ;
        RECT 18.085 130.475 18.255 130.665 ;
        RECT 19.015 130.510 19.175 130.620 ;
        RECT 19.925 130.475 20.095 130.665 ;
        RECT 20.845 130.455 21.015 130.645 ;
        RECT 23.605 130.475 23.775 130.665 ;
        RECT 24.065 130.455 24.235 130.645 ;
        RECT 24.525 130.455 24.695 130.645 ;
        RECT 25.905 130.455 26.075 130.645 ;
        RECT 28.210 130.455 28.380 130.645 ;
        RECT 28.665 130.475 28.835 130.665 ;
        RECT 29.125 130.475 29.295 130.665 ;
        RECT 30.965 130.615 31.135 130.645 ;
        RECT 29.580 130.505 29.700 130.615 ;
        RECT 30.960 130.505 31.135 130.615 ;
        RECT 30.965 130.455 31.135 130.505 ;
        RECT 31.420 130.475 31.590 130.665 ;
        RECT 31.880 130.505 32.000 130.615 ;
        RECT 32.345 130.455 32.515 130.645 ;
        RECT 32.805 130.475 32.975 130.665 ;
        RECT 36.025 130.455 36.195 130.645 ;
        RECT 40.440 130.475 40.610 130.665 ;
        RECT 41.085 130.455 41.255 130.645 ;
        RECT 44.765 130.475 44.935 130.665 ;
        RECT 48.720 130.455 48.890 130.645 ;
        RECT 52.125 130.475 52.295 130.665 ;
        RECT 52.580 130.505 52.700 130.615 ;
        RECT 53.320 130.455 53.490 130.645 ;
        RECT 57.645 130.455 57.815 130.645 ;
        RECT 65.925 130.455 66.095 130.645 ;
        RECT 66.385 130.455 66.555 130.665 ;
        RECT 67.770 130.645 67.935 130.665 ;
        RECT 66.855 130.510 67.015 130.620 ;
        RECT 67.765 130.475 67.935 130.645 ;
        RECT 71.720 130.455 71.890 130.645 ;
        RECT 73.745 130.475 73.915 130.665 ;
        RECT 75.575 130.455 75.745 130.645 ;
        RECT 77.425 130.475 77.595 130.665 ;
        RECT 77.890 130.475 78.060 130.665 ;
        RECT 80.645 130.475 80.815 130.645 ;
        RECT 81.115 130.500 81.275 130.610 ;
        RECT 81.560 130.505 81.680 130.615 ;
        RECT 80.645 130.455 80.810 130.475 ;
        RECT 82.945 130.455 83.115 130.665 ;
        RECT 5.525 129.645 6.895 130.455 ;
        RECT 6.905 129.645 12.415 130.455 ;
        RECT 12.425 129.645 15.175 130.455 ;
        RECT 15.645 129.775 17.935 130.455 ;
        RECT 17.945 129.775 21.155 130.455 ;
        RECT 15.645 129.545 16.565 129.775 ;
        RECT 17.945 129.545 19.080 129.775 ;
        RECT 21.165 129.545 24.335 130.455 ;
        RECT 24.385 129.645 25.755 130.455 ;
        RECT 25.765 129.775 28.055 130.455 ;
        RECT 27.135 129.545 28.055 129.775 ;
        RECT 28.065 129.545 29.415 130.455 ;
        RECT 29.915 129.545 31.265 130.455 ;
        RECT 31.295 129.585 31.725 130.370 ;
        RECT 32.315 129.775 35.780 130.455 ;
        RECT 35.885 129.775 40.700 130.455 ;
        RECT 40.945 129.775 48.255 130.455 ;
        RECT 34.860 129.545 35.780 129.775 ;
        RECT 44.460 129.555 45.370 129.775 ;
        RECT 46.905 129.545 48.255 129.775 ;
        RECT 48.305 129.775 52.205 130.455 ;
        RECT 52.905 129.775 56.805 130.455 ;
        RECT 48.305 129.545 49.235 129.775 ;
        RECT 52.905 129.545 53.835 129.775 ;
        RECT 57.055 129.585 57.485 130.370 ;
        RECT 57.505 129.645 58.875 130.455 ;
        RECT 58.925 129.775 66.235 130.455 ;
        RECT 66.245 129.775 71.060 130.455 ;
        RECT 71.305 129.775 75.205 130.455 ;
        RECT 58.925 129.545 60.275 129.775 ;
        RECT 61.810 129.555 62.720 129.775 ;
        RECT 71.305 129.545 72.235 129.775 ;
        RECT 75.445 129.545 78.655 130.455 ;
        RECT 78.975 129.775 80.810 130.455 ;
        RECT 78.975 129.545 79.905 129.775 ;
        RECT 81.885 129.645 83.255 130.455 ;
      LAYER nwell ;
        RECT 5.330 126.425 83.450 129.255 ;
      LAYER pwell ;
        RECT 5.525 125.225 6.895 126.035 ;
        RECT 6.905 125.225 8.275 126.005 ;
        RECT 8.285 125.225 13.795 126.035 ;
        RECT 13.805 125.225 17.475 126.035 ;
        RECT 18.415 125.310 18.845 126.095 ;
        RECT 18.865 125.225 24.375 126.035 ;
        RECT 24.385 125.225 27.135 126.035 ;
        RECT 27.840 125.225 32.655 125.905 ;
        RECT 33.155 125.225 35.875 126.135 ;
        RECT 38.185 125.935 39.140 126.135 ;
        RECT 36.810 125.225 38.175 125.905 ;
        RECT 38.185 125.255 40.465 125.935 ;
        RECT 40.580 125.905 41.500 126.135 ;
        RECT 38.185 125.225 39.140 125.255 ;
        RECT 5.665 125.015 5.835 125.225 ;
        RECT 7.045 125.015 7.215 125.225 ;
        RECT 8.425 125.035 8.595 125.225 ;
        RECT 11.645 125.015 11.815 125.205 ;
        RECT 12.105 125.015 12.275 125.205 ;
        RECT 13.945 125.035 14.115 125.225 ;
        RECT 17.625 125.015 17.795 125.205 ;
        RECT 19.005 125.035 19.175 125.225 ;
        RECT 21.765 125.015 21.935 125.205 ;
        RECT 24.065 125.035 24.235 125.205 ;
        RECT 24.065 125.015 24.215 125.035 ;
        RECT 24.525 125.015 24.695 125.225 ;
        RECT 27.280 125.015 27.450 125.205 ;
        RECT 27.745 125.035 27.915 125.205 ;
        RECT 30.960 125.065 31.080 125.175 ;
        RECT 31.890 125.015 32.060 125.205 ;
        RECT 32.345 125.035 32.515 125.225 ;
        RECT 32.800 125.065 32.920 125.175 ;
        RECT 33.275 125.060 33.435 125.170 ;
        RECT 34.185 125.015 34.355 125.205 ;
        RECT 35.565 125.035 35.735 125.225 ;
        RECT 36.020 125.065 36.140 125.175 ;
        RECT 36.485 125.035 36.655 125.205 ;
        RECT 40.170 125.035 40.340 125.255 ;
        RECT 40.580 125.225 44.045 125.905 ;
        RECT 44.175 125.310 44.605 126.095 ;
        RECT 45.085 125.905 46.015 126.135 ;
        RECT 49.320 125.905 50.240 126.135 ;
        RECT 45.085 125.225 48.985 125.905 ;
        RECT 49.320 125.225 52.785 125.905 ;
        RECT 52.905 125.225 54.735 126.035 ;
        RECT 54.745 125.905 56.090 126.135 ;
        RECT 59.240 125.905 60.160 126.135 ;
        RECT 54.745 125.225 56.575 125.905 ;
        RECT 56.695 125.225 60.160 125.905 ;
        RECT 60.265 125.905 61.610 126.135 ;
        RECT 62.200 125.905 63.120 126.135 ;
        RECT 68.440 125.905 69.360 126.135 ;
        RECT 60.265 125.225 62.095 125.905 ;
        RECT 62.200 125.225 65.665 125.905 ;
        RECT 65.895 125.225 69.360 125.905 ;
        RECT 69.935 125.310 70.365 126.095 ;
        RECT 70.385 125.225 73.595 126.135 ;
        RECT 78.040 125.905 78.950 126.125 ;
        RECT 80.485 125.905 81.835 126.135 ;
        RECT 74.525 125.225 81.835 125.905 ;
        RECT 81.885 125.225 83.255 126.035 ;
        RECT 41.820 125.015 41.990 125.205 ;
        RECT 43.845 125.035 44.015 125.225 ;
        RECT 44.760 125.065 44.880 125.175 ;
        RECT 45.500 125.035 45.670 125.225 ;
        RECT 45.685 125.015 45.855 125.205 ;
        RECT 48.445 125.015 48.615 125.205 ;
        RECT 49.825 125.015 49.995 125.205 ;
        RECT 52.585 125.035 52.755 125.225 ;
        RECT 53.045 125.035 53.215 125.225 ;
        RECT 56.265 125.035 56.435 125.225 ;
        RECT 56.725 125.035 56.895 125.225 ;
        RECT 57.645 125.015 57.815 125.205 ;
        RECT 61.785 125.035 61.955 125.225 ;
        RECT 65.280 125.015 65.450 125.205 ;
        RECT 65.465 125.035 65.635 125.225 ;
        RECT 65.925 125.035 66.095 125.225 ;
        RECT 70.515 125.205 70.685 125.225 ;
        RECT 69.600 125.065 69.720 125.175 ;
        RECT 70.515 125.035 70.695 125.205 ;
        RECT 73.755 125.070 73.915 125.180 ;
        RECT 70.525 125.015 70.695 125.035 ;
        RECT 74.200 125.015 74.370 125.205 ;
        RECT 74.665 125.015 74.835 125.225 ;
        RECT 82.945 125.015 83.115 125.225 ;
        RECT 5.525 124.205 6.895 125.015 ;
        RECT 6.905 124.205 8.275 125.015 ;
        RECT 8.285 124.335 11.955 125.015 ;
        RECT 8.285 124.105 9.215 124.335 ;
        RECT 11.965 124.205 17.475 125.015 ;
        RECT 17.485 124.335 19.315 125.015 ;
        RECT 17.970 124.105 19.315 124.335 ;
        RECT 19.325 124.105 22.075 125.015 ;
        RECT 22.285 124.195 24.215 125.015 ;
        RECT 24.385 124.205 26.215 125.015 ;
        RECT 22.285 124.105 23.235 124.195 ;
        RECT 26.245 124.105 27.595 125.015 ;
        RECT 28.010 124.335 30.435 125.015 ;
        RECT 31.295 124.145 31.725 124.930 ;
        RECT 31.745 124.105 33.095 125.015 ;
        RECT 34.045 124.335 41.355 125.015 ;
        RECT 37.560 124.115 38.470 124.335 ;
        RECT 40.005 124.105 41.355 124.335 ;
        RECT 41.405 124.335 45.305 125.015 ;
        RECT 45.545 124.335 48.285 125.015 ;
        RECT 41.405 124.105 42.335 124.335 ;
        RECT 48.305 124.205 49.675 125.015 ;
        RECT 49.685 124.335 56.995 125.015 ;
        RECT 53.200 124.115 54.110 124.335 ;
        RECT 55.645 124.105 56.995 124.335 ;
        RECT 57.055 124.145 57.485 124.930 ;
        RECT 57.505 124.335 64.815 125.015 ;
        RECT 61.020 124.115 61.930 124.335 ;
        RECT 63.465 124.105 64.815 124.335 ;
        RECT 64.865 124.335 68.765 125.015 ;
        RECT 69.005 124.335 70.835 125.015 ;
        RECT 64.865 124.105 65.795 124.335 ;
        RECT 69.005 124.105 70.350 124.335 ;
        RECT 71.040 124.105 74.515 125.015 ;
        RECT 74.525 124.335 81.835 125.015 ;
        RECT 78.040 124.115 78.950 124.335 ;
        RECT 80.485 124.105 81.835 124.335 ;
        RECT 81.885 124.205 83.255 125.015 ;
      LAYER nwell ;
        RECT 5.330 120.985 83.450 123.815 ;
      LAYER pwell ;
        RECT 5.525 119.785 6.895 120.595 ;
        RECT 10.880 120.465 11.790 120.685 ;
        RECT 13.325 120.465 14.675 120.695 ;
        RECT 7.365 119.785 14.675 120.465 ;
        RECT 14.725 119.785 16.075 120.695 ;
        RECT 16.560 120.015 18.395 120.695 ;
        RECT 16.560 119.785 18.250 120.015 ;
        RECT 18.415 119.870 18.845 120.655 ;
        RECT 18.885 119.785 20.235 120.695 ;
        RECT 25.745 120.465 26.675 120.695 ;
        RECT 29.425 120.465 30.355 120.695 ;
        RECT 32.440 120.465 33.575 120.695 ;
        RECT 20.245 119.785 22.985 120.465 ;
        RECT 23.005 119.785 26.675 120.465 ;
        RECT 26.685 119.785 30.355 120.465 ;
        RECT 30.365 119.785 33.575 120.465 ;
        RECT 33.685 119.785 36.795 120.695 ;
        RECT 36.845 120.465 38.195 120.695 ;
        RECT 39.730 120.465 40.640 120.685 ;
        RECT 36.845 119.785 44.155 120.465 ;
        RECT 44.175 119.870 44.605 120.655 ;
        RECT 44.625 119.785 47.375 120.595 ;
        RECT 47.855 119.785 49.205 120.695 ;
        RECT 49.245 119.785 50.595 120.695 ;
        RECT 50.605 120.465 51.535 120.695 ;
        RECT 54.745 120.465 56.090 120.695 ;
        RECT 50.605 119.785 54.505 120.465 ;
        RECT 54.745 119.785 56.575 120.465 ;
        RECT 56.585 119.785 57.935 120.695 ;
        RECT 57.965 119.785 59.315 120.695 ;
        RECT 59.845 120.465 61.195 120.695 ;
        RECT 62.730 120.465 63.640 120.685 ;
        RECT 68.675 120.465 69.605 120.695 ;
        RECT 59.845 119.785 67.155 120.465 ;
        RECT 67.770 119.785 69.605 120.465 ;
        RECT 69.935 119.870 70.365 120.655 ;
        RECT 70.385 119.785 73.860 120.695 ;
        RECT 74.260 119.785 77.735 120.695 ;
        RECT 77.745 119.785 80.955 120.695 ;
        RECT 81.885 119.785 83.255 120.595 ;
        RECT 5.665 119.575 5.835 119.785 ;
        RECT 7.045 119.735 7.215 119.765 ;
        RECT 7.040 119.625 7.215 119.735 ;
        RECT 7.045 119.575 7.215 119.625 ;
        RECT 7.505 119.595 7.675 119.785 ;
        RECT 14.410 119.575 14.580 119.765 ;
        RECT 14.870 119.595 15.040 119.785 ;
        RECT 18.080 119.595 18.250 119.785 ;
        RECT 19.000 119.575 19.170 119.785 ;
        RECT 19.460 119.625 19.580 119.735 ;
        RECT 19.925 119.575 20.095 119.765 ;
        RECT 20.385 119.595 20.555 119.785 ;
        RECT 23.145 119.595 23.315 119.785 ;
        RECT 24.065 119.575 24.235 119.765 ;
        RECT 26.825 119.595 26.995 119.785 ;
        RECT 30.505 119.595 30.675 119.785 ;
        RECT 31.885 119.575 32.055 119.765 ;
        RECT 33.725 119.595 33.895 119.785 ;
        RECT 37.405 119.575 37.575 119.765 ;
        RECT 42.925 119.575 43.095 119.765 ;
        RECT 43.845 119.595 44.015 119.785 ;
        RECT 44.765 119.595 44.935 119.785 ;
        RECT 45.680 119.625 45.800 119.735 ;
        RECT 46.145 119.575 46.315 119.765 ;
        RECT 47.520 119.625 47.640 119.735 ;
        RECT 48.905 119.595 49.075 119.785 ;
        RECT 49.360 119.595 49.530 119.785 ;
        RECT 51.020 119.595 51.190 119.785 ;
        RECT 53.505 119.575 53.675 119.765 ;
        RECT 56.265 119.595 56.435 119.785 ;
        RECT 57.650 119.595 57.820 119.785 ;
        RECT 59.030 119.595 59.200 119.785 ;
        RECT 59.480 119.625 59.600 119.735 ;
        RECT 60.405 119.575 60.575 119.765 ;
        RECT 62.245 119.575 62.415 119.765 ;
        RECT 62.705 119.575 62.875 119.765 ;
        RECT 65.925 119.575 66.095 119.765 ;
        RECT 66.845 119.595 67.015 119.785 ;
        RECT 67.770 119.765 67.935 119.785 ;
        RECT 67.300 119.625 67.420 119.735 ;
        RECT 67.765 119.595 67.935 119.765 ;
        RECT 70.530 119.595 70.700 119.785 ;
        RECT 73.285 119.595 73.455 119.765 ;
        RECT 73.290 119.575 73.455 119.595 ;
        RECT 75.585 119.575 75.755 119.765 ;
        RECT 77.420 119.595 77.590 119.785 ;
        RECT 80.645 119.595 80.815 119.785 ;
        RECT 81.115 119.620 81.275 119.740 ;
        RECT 80.645 119.575 80.810 119.595 ;
        RECT 82.945 119.575 83.115 119.785 ;
        RECT 5.525 118.765 6.895 119.575 ;
        RECT 6.905 118.895 14.215 119.575 ;
        RECT 10.420 118.675 11.330 118.895 ;
        RECT 12.865 118.665 14.215 118.895 ;
        RECT 14.265 118.665 15.615 119.575 ;
        RECT 15.840 118.665 19.315 119.575 ;
        RECT 19.785 118.665 22.995 119.575 ;
        RECT 23.925 118.895 31.235 119.575 ;
        RECT 27.440 118.675 28.350 118.895 ;
        RECT 29.885 118.665 31.235 118.895 ;
        RECT 31.295 118.705 31.725 119.490 ;
        RECT 31.745 118.765 37.255 119.575 ;
        RECT 37.265 118.765 42.775 119.575 ;
        RECT 42.785 118.765 45.535 119.575 ;
        RECT 46.005 118.895 53.315 119.575 ;
        RECT 53.475 118.895 56.940 119.575 ;
        RECT 49.520 118.675 50.430 118.895 ;
        RECT 51.965 118.665 53.315 118.895 ;
        RECT 56.020 118.665 56.940 118.895 ;
        RECT 57.055 118.705 57.485 119.490 ;
        RECT 57.505 118.665 60.715 119.575 ;
        RECT 60.725 118.895 62.555 119.575 ;
        RECT 60.725 118.665 62.070 118.895 ;
        RECT 62.565 118.665 65.775 119.575 ;
        RECT 65.785 118.895 73.095 119.575 ;
        RECT 73.290 118.895 75.125 119.575 ;
        RECT 69.300 118.675 70.210 118.895 ;
        RECT 71.745 118.665 73.095 118.895 ;
        RECT 74.195 118.665 75.125 118.895 ;
        RECT 75.445 118.665 78.655 119.575 ;
        RECT 78.975 118.895 80.810 119.575 ;
        RECT 78.975 118.665 79.905 118.895 ;
        RECT 81.885 118.765 83.255 119.575 ;
      LAYER nwell ;
        RECT 5.330 115.545 83.450 118.375 ;
      LAYER pwell ;
        RECT 5.525 114.345 6.895 115.155 ;
        RECT 7.825 115.025 8.755 115.255 ;
        RECT 7.825 114.345 11.495 115.025 ;
        RECT 11.505 114.345 12.855 115.255 ;
        RECT 12.885 115.025 14.020 115.255 ;
        RECT 17.440 115.055 18.395 115.255 ;
        RECT 12.885 114.345 16.095 115.025 ;
        RECT 16.115 114.375 18.395 115.055 ;
        RECT 18.415 114.430 18.845 115.215 ;
        RECT 5.665 114.135 5.835 114.345 ;
        RECT 7.045 114.135 7.215 114.325 ;
        RECT 11.185 114.135 11.355 114.345 ;
        RECT 11.650 114.325 11.820 114.345 ;
        RECT 11.645 114.155 11.820 114.325 ;
        RECT 13.940 114.185 14.060 114.295 ;
        RECT 11.645 114.135 11.815 114.155 ;
        RECT 14.405 114.135 14.575 114.325 ;
        RECT 15.785 114.155 15.955 114.345 ;
        RECT 16.240 114.155 16.410 114.375 ;
        RECT 17.440 114.345 18.395 114.375 ;
        RECT 19.060 114.345 22.535 115.255 ;
        RECT 23.595 115.025 24.525 115.255 ;
        RECT 22.690 114.345 24.525 115.025 ;
        RECT 25.345 115.025 26.695 115.255 ;
        RECT 28.230 115.025 29.140 115.245 ;
        RECT 32.705 115.025 34.055 115.255 ;
        RECT 35.590 115.025 36.500 115.245 ;
        RECT 25.345 114.345 32.655 115.025 ;
        RECT 32.705 114.345 40.015 115.025 ;
        RECT 40.025 114.345 41.375 115.255 ;
        RECT 41.405 114.345 44.155 115.155 ;
        RECT 44.175 114.430 44.605 115.215 ;
        RECT 45.545 115.025 46.475 115.255 ;
        RECT 52.340 115.025 53.260 115.255 ;
        RECT 45.545 114.345 49.445 115.025 ;
        RECT 49.795 114.345 53.260 115.025 ;
        RECT 53.365 114.345 56.575 115.255 ;
        RECT 56.585 114.345 58.415 115.255 ;
        RECT 58.425 114.345 60.255 115.255 ;
        RECT 60.265 114.345 63.475 115.255 ;
        RECT 66.140 115.025 67.060 115.255 ;
        RECT 63.595 114.345 67.060 115.025 ;
        RECT 67.165 114.345 69.255 115.155 ;
        RECT 69.935 114.430 70.365 115.215 ;
        RECT 70.580 114.345 74.055 115.255 ;
        RECT 77.580 115.025 78.490 115.245 ;
        RECT 80.025 115.025 81.375 115.255 ;
        RECT 74.065 114.345 81.375 115.025 ;
        RECT 81.885 114.345 83.255 115.155 ;
        RECT 17.625 114.135 17.795 114.325 ;
        RECT 5.525 113.325 6.895 114.135 ;
        RECT 6.905 113.325 9.655 114.135 ;
        RECT 9.665 113.225 11.480 114.135 ;
        RECT 11.505 113.455 13.795 114.135 ;
        RECT 12.875 113.225 13.795 113.455 ;
        RECT 14.365 113.225 17.475 114.135 ;
        RECT 17.485 113.325 19.315 114.135 ;
        RECT 19.465 114.105 19.635 114.325 ;
        RECT 22.220 114.155 22.390 114.345 ;
        RECT 22.690 114.325 22.855 114.345 ;
        RECT 22.680 114.155 22.855 114.325 ;
        RECT 24.985 114.295 25.155 114.325 ;
        RECT 24.980 114.185 25.155 114.295 ;
        RECT 21.590 114.105 22.535 114.135 ;
        RECT 22.680 114.105 22.850 114.155 ;
        RECT 24.985 114.135 25.155 114.185 ;
        RECT 28.210 114.135 28.380 114.325 ;
        RECT 32.345 114.155 32.515 114.345 ;
        RECT 33.265 114.135 33.435 114.325 ;
        RECT 33.735 114.180 33.895 114.290 ;
        RECT 34.645 114.135 34.815 114.325 ;
        RECT 39.705 114.155 39.875 114.345 ;
        RECT 40.170 114.155 40.340 114.345 ;
        RECT 41.545 114.155 41.715 114.345 ;
        RECT 42.005 114.135 42.175 114.325 ;
        RECT 44.775 114.190 44.935 114.300 ;
        RECT 45.960 114.155 46.130 114.345 ;
        RECT 49.825 114.155 49.995 114.345 ;
        RECT 52.585 114.135 52.755 114.325 ;
        RECT 53.045 114.135 53.215 114.325 ;
        RECT 53.505 114.155 53.675 114.345 ;
        RECT 56.275 114.180 56.435 114.290 ;
        RECT 56.730 114.155 56.900 114.345 ;
        RECT 57.645 114.135 57.815 114.325 ;
        RECT 59.940 114.155 60.110 114.345 ;
        RECT 63.165 114.155 63.335 114.345 ;
        RECT 63.625 114.155 63.795 114.345 ;
        RECT 67.305 114.155 67.475 114.345 ;
        RECT 67.765 114.135 67.935 114.325 ;
        RECT 69.150 114.135 69.320 114.325 ;
        RECT 69.605 114.135 69.775 114.325 ;
        RECT 73.740 114.155 73.910 114.345 ;
        RECT 74.205 114.155 74.375 114.345 ;
        RECT 78.805 114.155 78.975 114.325 ;
        RECT 79.265 114.155 79.435 114.325 ;
        RECT 81.560 114.185 81.680 114.295 ;
        RECT 78.805 114.135 78.970 114.155 ;
        RECT 23.880 114.105 24.835 114.135 ;
        RECT 19.465 113.905 22.535 114.105 ;
        RECT 19.325 113.425 22.535 113.905 ;
        RECT 22.555 113.425 24.835 114.105 ;
        RECT 19.325 113.225 20.255 113.425 ;
        RECT 21.590 113.225 22.535 113.425 ;
        RECT 23.880 113.225 24.835 113.425 ;
        RECT 24.885 113.225 28.055 114.135 ;
        RECT 28.065 113.225 30.985 114.135 ;
        RECT 31.295 113.265 31.725 114.050 ;
        RECT 31.745 113.455 33.575 114.135 ;
        RECT 34.505 113.455 41.815 114.135 ;
        RECT 41.865 113.455 49.175 114.135 ;
        RECT 38.020 113.235 38.930 113.455 ;
        RECT 40.465 113.225 41.815 113.455 ;
        RECT 45.380 113.235 46.290 113.455 ;
        RECT 47.825 113.225 49.175 113.455 ;
        RECT 49.320 113.455 52.785 114.135 ;
        RECT 49.320 113.225 50.240 113.455 ;
        RECT 52.905 113.225 56.115 114.135 ;
        RECT 57.055 113.265 57.485 114.050 ;
        RECT 57.555 113.225 60.715 114.135 ;
        RECT 60.765 113.455 68.075 114.135 ;
        RECT 60.765 113.225 62.115 113.455 ;
        RECT 63.650 113.235 64.560 113.455 ;
        RECT 68.085 113.225 69.435 114.135 ;
        RECT 69.465 113.455 76.775 114.135 ;
        RECT 72.980 113.235 73.890 113.455 ;
        RECT 75.425 113.225 76.775 113.455 ;
        RECT 77.135 113.455 78.970 114.135 ;
        RECT 79.270 114.135 79.435 114.155 ;
        RECT 82.945 114.135 83.115 114.345 ;
        RECT 79.270 113.455 81.105 114.135 ;
        RECT 77.135 113.225 78.065 113.455 ;
        RECT 80.175 113.225 81.105 113.455 ;
        RECT 81.885 113.325 83.255 114.135 ;
      LAYER nwell ;
        RECT 5.330 110.105 83.450 112.935 ;
      LAYER pwell ;
        RECT 5.525 108.905 6.895 109.715 ;
        RECT 6.905 108.905 12.415 109.715 ;
        RECT 12.425 108.905 15.175 109.715 ;
        RECT 15.285 108.905 18.395 109.815 ;
        RECT 18.415 108.990 18.845 109.775 ;
        RECT 19.785 108.905 23.440 109.815 ;
        RECT 24.090 108.905 27.960 109.815 ;
        RECT 28.065 108.905 32.880 109.585 ;
        RECT 33.145 108.905 34.495 109.815 ;
        RECT 38.020 109.585 38.930 109.805 ;
        RECT 40.465 109.585 41.815 109.815 ;
        RECT 34.505 108.905 41.815 109.585 ;
        RECT 41.865 108.905 43.695 109.715 ;
        RECT 44.175 108.990 44.605 109.775 ;
        RECT 44.625 109.585 45.555 109.815 ;
        RECT 44.625 108.905 48.525 109.585 ;
        RECT 48.765 108.905 51.975 109.815 ;
        RECT 53.585 109.725 54.535 109.815 ;
        RECT 52.605 108.905 54.535 109.725 ;
        RECT 54.745 108.905 59.560 109.585 ;
        RECT 59.805 108.905 62.725 109.815 ;
        RECT 67.145 109.585 68.075 109.815 ;
        RECT 64.175 108.905 68.075 109.585 ;
        RECT 68.085 109.585 69.430 109.815 ;
        RECT 68.085 108.905 69.915 109.585 ;
        RECT 69.935 108.990 70.365 109.775 ;
        RECT 75.445 109.585 76.790 109.815 ;
        RECT 78.690 109.585 80.035 109.815 ;
        RECT 80.530 109.585 81.875 109.815 ;
        RECT 70.385 108.905 75.200 109.585 ;
        RECT 75.445 108.905 77.275 109.585 ;
        RECT 78.205 108.905 80.035 109.585 ;
        RECT 80.045 108.905 81.875 109.585 ;
        RECT 81.885 108.905 83.255 109.715 ;
        RECT 5.665 108.695 5.835 108.905 ;
        RECT 7.045 108.885 7.215 108.905 ;
        RECT 7.045 108.715 7.225 108.885 ;
        RECT 7.055 108.695 7.225 108.715 ;
        RECT 8.425 108.695 8.595 108.885 ;
        RECT 12.565 108.715 12.735 108.905 ;
        RECT 15.325 108.885 15.495 108.905 ;
        RECT 13.940 108.745 14.060 108.855 ;
        RECT 15.320 108.715 15.495 108.885 ;
        RECT 15.780 108.745 15.900 108.855 ;
        RECT 15.320 108.695 15.490 108.715 ;
        RECT 16.245 108.695 16.415 108.885 ;
        RECT 19.015 108.750 19.175 108.860 ;
        RECT 19.455 108.695 19.625 108.885 ;
        RECT 19.930 108.715 20.100 108.905 ;
        RECT 24.090 108.885 24.235 108.905 ;
        RECT 23.600 108.745 23.720 108.855 ;
        RECT 24.065 108.715 24.235 108.885 ;
        RECT 24.525 108.715 24.695 108.885 ;
        RECT 24.525 108.695 24.690 108.715 ;
        RECT 24.985 108.695 25.155 108.885 ;
        RECT 28.205 108.715 28.375 108.905 ;
        RECT 33.260 108.885 33.430 108.905 ;
        RECT 28.665 108.695 28.835 108.885 ;
        RECT 33.260 108.715 33.435 108.885 ;
        RECT 33.735 108.740 33.895 108.850 ;
        RECT 33.265 108.695 33.435 108.715 ;
        RECT 34.645 108.695 34.815 108.905 ;
        RECT 38.330 108.695 38.500 108.885 ;
        RECT 39.705 108.695 39.875 108.885 ;
        RECT 41.085 108.695 41.255 108.885 ;
        RECT 42.005 108.715 42.175 108.905 ;
        RECT 43.840 108.745 43.960 108.855 ;
        RECT 45.040 108.715 45.210 108.905 ;
        RECT 46.145 108.695 46.315 108.885 ;
        RECT 47.525 108.695 47.695 108.885 ;
        RECT 51.675 108.715 51.845 108.905 ;
        RECT 52.605 108.885 52.755 108.905 ;
        RECT 54.885 108.885 55.055 108.905 ;
        RECT 52.120 108.745 52.240 108.855 ;
        RECT 52.585 108.715 52.755 108.885 ;
        RECT 54.880 108.715 55.055 108.885 ;
        RECT 57.645 108.715 57.815 108.885 ;
        RECT 59.950 108.715 60.120 108.905 ;
        RECT 5.525 107.885 6.895 108.695 ;
        RECT 6.905 107.915 8.275 108.695 ;
        RECT 8.285 107.885 13.795 108.695 ;
        RECT 14.285 107.785 15.635 108.695 ;
        RECT 16.105 107.785 19.315 108.695 ;
        RECT 19.325 107.785 22.535 108.695 ;
        RECT 22.855 108.015 24.690 108.695 ;
        RECT 24.845 108.015 28.515 108.695 ;
        RECT 22.855 107.785 23.785 108.015 ;
        RECT 27.585 107.785 28.515 108.015 ;
        RECT 28.535 107.785 31.265 108.695 ;
        RECT 31.295 107.825 31.725 108.610 ;
        RECT 31.745 108.015 33.575 108.695 ;
        RECT 34.615 108.015 38.080 108.695 ;
        RECT 37.160 107.785 38.080 108.015 ;
        RECT 38.185 107.785 39.535 108.695 ;
        RECT 39.565 107.885 40.935 108.695 ;
        RECT 40.945 108.015 45.760 108.695 ;
        RECT 46.005 107.885 47.375 108.695 ;
        RECT 47.385 108.015 54.695 108.695 ;
        RECT 54.880 108.665 55.050 108.715 ;
        RECT 57.655 108.695 57.815 108.715 ;
        RECT 61.785 108.695 61.955 108.885 ;
        RECT 63.175 108.750 63.335 108.860 ;
        RECT 67.490 108.715 67.660 108.905 ;
        RECT 69.605 108.715 69.775 108.905 ;
        RECT 70.525 108.715 70.695 108.905 ;
        RECT 72.365 108.695 72.535 108.885 ;
        RECT 72.830 108.695 73.000 108.885 ;
        RECT 76.505 108.695 76.675 108.885 ;
        RECT 76.965 108.715 77.135 108.905 ;
        RECT 77.435 108.750 77.595 108.860 ;
        RECT 78.345 108.715 78.515 108.905 ;
        RECT 79.725 108.715 79.895 108.885 ;
        RECT 79.725 108.695 79.890 108.715 ;
        RECT 80.185 108.695 80.355 108.905 ;
        RECT 82.945 108.695 83.115 108.905 ;
        RECT 56.080 108.665 57.035 108.695 ;
        RECT 50.900 107.795 51.810 108.015 ;
        RECT 53.345 107.785 54.695 108.015 ;
        RECT 54.755 107.985 57.035 108.665 ;
        RECT 56.080 107.785 57.035 107.985 ;
        RECT 57.055 107.825 57.485 108.610 ;
        RECT 57.655 107.785 61.310 108.695 ;
        RECT 61.645 108.015 68.955 108.695 ;
        RECT 65.160 107.795 66.070 108.015 ;
        RECT 67.605 107.785 68.955 108.015 ;
        RECT 69.100 108.015 72.565 108.695 ;
        RECT 69.100 107.785 70.020 108.015 ;
        RECT 72.685 107.785 76.160 108.695 ;
        RECT 76.365 107.915 77.735 108.695 ;
        RECT 78.055 108.015 79.890 108.695 ;
        RECT 80.045 108.015 81.875 108.695 ;
        RECT 78.055 107.785 78.985 108.015 ;
        RECT 80.530 107.785 81.875 108.015 ;
        RECT 81.885 107.885 83.255 108.695 ;
      LAYER nwell ;
        RECT 5.330 104.665 83.450 107.495 ;
      LAYER pwell ;
        RECT 5.525 103.465 6.895 104.275 ;
        RECT 7.375 104.145 10.375 104.375 ;
        RECT 11.965 104.145 12.895 104.375 ;
        RECT 7.375 104.055 11.955 104.145 ;
        RECT 7.365 103.695 11.955 104.055 ;
        RECT 7.365 103.505 8.295 103.695 ;
        RECT 7.375 103.465 8.295 103.505 ;
        RECT 10.385 103.465 11.955 103.695 ;
        RECT 11.965 103.465 15.635 104.145 ;
        RECT 15.645 103.695 17.480 104.375 ;
        RECT 15.790 103.465 17.480 103.695 ;
        RECT 18.415 103.550 18.845 104.335 ;
        RECT 18.865 104.145 19.790 104.375 ;
        RECT 23.205 104.145 27.135 104.375 ;
        RECT 30.345 104.145 31.275 104.375 ;
        RECT 18.865 103.465 22.535 104.145 ;
        RECT 22.720 103.465 27.135 104.145 ;
        RECT 27.605 103.465 31.275 104.145 ;
        RECT 31.285 103.465 34.395 104.375 ;
        RECT 38.020 104.145 38.930 104.365 ;
        RECT 40.465 104.145 41.815 104.375 ;
        RECT 34.505 103.465 41.815 104.145 ;
        RECT 41.865 103.465 43.695 104.275 ;
        RECT 44.175 103.550 44.605 104.335 ;
        RECT 44.675 103.465 47.835 104.375 ;
        RECT 48.845 103.465 51.845 104.375 ;
        RECT 51.985 103.465 53.335 104.375 ;
        RECT 53.365 103.465 54.715 104.375 ;
        RECT 57.400 104.145 58.320 104.375 ;
        RECT 54.855 103.465 58.320 104.145 ;
        RECT 58.620 103.465 62.095 104.375 ;
        RECT 62.125 103.465 63.475 104.375 ;
        RECT 63.485 104.145 64.415 104.375 ;
        RECT 63.485 103.465 67.385 104.145 ;
        RECT 67.625 103.465 69.455 104.275 ;
        RECT 69.935 103.550 70.365 104.335 ;
        RECT 71.155 104.145 72.085 104.375 ;
        RECT 71.155 103.465 72.990 104.145 ;
        RECT 73.145 103.465 74.515 104.275 ;
        RECT 78.040 104.145 78.950 104.365 ;
        RECT 80.485 104.145 81.835 104.375 ;
        RECT 74.525 103.465 81.835 104.145 ;
        RECT 81.885 103.465 83.255 104.275 ;
        RECT 5.665 103.255 5.835 103.465 ;
        RECT 7.040 103.305 7.160 103.415 ;
        RECT 7.505 103.255 7.675 103.445 ;
        RECT 11.645 103.275 11.815 103.465 ;
        RECT 15.325 103.275 15.495 103.465 ;
        RECT 15.790 103.275 15.960 103.465 ;
        RECT 17.625 103.255 17.795 103.445 ;
        RECT 18.080 103.410 18.200 103.415 ;
        RECT 18.080 103.305 18.255 103.410 ;
        RECT 18.095 103.300 18.255 103.305 ;
        RECT 5.525 102.445 6.895 103.255 ;
        RECT 7.365 102.575 14.675 103.255 ;
        RECT 10.880 102.355 11.790 102.575 ;
        RECT 13.325 102.345 14.675 102.575 ;
        RECT 14.725 102.345 17.895 103.255 ;
        RECT 19.010 103.225 19.180 103.465 ;
        RECT 22.720 103.445 22.830 103.465 ;
        RECT 22.660 103.410 22.830 103.445 ;
        RECT 22.660 103.300 22.855 103.410 ;
        RECT 27.280 103.305 27.400 103.415 ;
        RECT 22.660 103.275 22.830 103.300 ;
        RECT 27.745 103.275 27.915 103.465 ;
        RECT 30.960 103.255 31.130 103.445 ;
        RECT 34.185 103.275 34.355 103.465 ;
        RECT 34.645 103.275 34.815 103.465 ;
        RECT 38.785 103.255 38.955 103.445 ;
        RECT 39.245 103.255 39.415 103.445 ;
        RECT 42.005 103.275 42.175 103.465 ;
        RECT 43.845 103.415 44.015 103.445 ;
        RECT 43.840 103.305 44.015 103.415 ;
        RECT 43.845 103.255 44.015 103.305 ;
        RECT 44.765 103.275 44.935 103.465 ;
        RECT 47.525 103.255 47.695 103.445 ;
        RECT 47.985 103.255 48.155 103.445 ;
        RECT 48.905 103.275 49.075 103.465 ;
        RECT 51.665 103.255 51.835 103.445 ;
        RECT 52.130 103.275 52.300 103.465 ;
        RECT 53.050 103.255 53.220 103.445 ;
        RECT 54.430 103.275 54.600 103.465 ;
        RECT 54.885 103.275 55.055 103.465 ;
        RECT 56.275 103.300 56.435 103.410 ;
        RECT 57.645 103.255 57.815 103.445 ;
        RECT 59.025 103.255 59.195 103.445 ;
        RECT 61.780 103.275 61.950 103.465 ;
        RECT 62.240 103.275 62.410 103.465 ;
        RECT 62.715 103.300 62.875 103.410 ;
        RECT 63.900 103.275 64.070 103.465 ;
        RECT 66.840 103.255 67.010 103.445 ;
        RECT 67.305 103.255 67.475 103.445 ;
        RECT 67.765 103.275 67.935 103.465 ;
        RECT 72.825 103.445 72.990 103.465 ;
        RECT 69.600 103.305 69.720 103.415 ;
        RECT 70.520 103.305 70.640 103.415 ;
        RECT 72.825 103.275 72.995 103.445 ;
        RECT 73.285 103.275 73.455 103.465 ;
        RECT 74.665 103.445 74.835 103.465 ;
        RECT 74.665 103.275 74.840 103.445 ;
        RECT 74.670 103.255 74.840 103.275 ;
        RECT 78.335 103.255 78.505 103.445 ;
        RECT 81.560 103.305 81.680 103.415 ;
        RECT 82.945 103.255 83.115 103.465 ;
        RECT 21.585 103.225 22.535 103.255 ;
        RECT 18.865 102.545 22.535 103.225 ;
        RECT 21.585 102.345 22.535 102.545 ;
        RECT 23.715 102.345 31.275 103.255 ;
        RECT 31.295 102.385 31.725 103.170 ;
        RECT 31.785 102.575 39.095 103.255 ;
        RECT 31.785 102.345 33.135 102.575 ;
        RECT 34.670 102.355 35.580 102.575 ;
        RECT 39.105 102.445 40.475 103.255 ;
        RECT 40.580 102.575 44.045 103.255 ;
        RECT 44.260 102.575 47.725 103.255 ;
        RECT 40.580 102.345 41.500 102.575 ;
        RECT 44.260 102.345 45.180 102.575 ;
        RECT 47.845 102.445 51.515 103.255 ;
        RECT 51.525 102.445 52.895 103.255 ;
        RECT 52.905 102.345 55.825 103.255 ;
        RECT 57.055 102.385 57.485 103.170 ;
        RECT 57.515 102.345 58.865 103.255 ;
        RECT 58.885 102.445 62.555 103.255 ;
        RECT 63.680 102.345 67.155 103.255 ;
        RECT 67.165 102.575 74.475 103.255 ;
        RECT 70.680 102.355 71.590 102.575 ;
        RECT 73.125 102.345 74.475 102.575 ;
        RECT 74.525 102.345 78.000 103.255 ;
        RECT 78.205 102.345 81.415 103.255 ;
        RECT 81.885 102.445 83.255 103.255 ;
      LAYER nwell ;
        RECT 5.330 99.225 83.450 102.055 ;
      LAYER pwell ;
        RECT 5.525 98.025 6.895 98.835 ;
        RECT 10.420 98.705 11.330 98.925 ;
        RECT 12.865 98.705 14.215 98.935 ;
        RECT 6.905 98.025 14.215 98.705 ;
        RECT 14.265 98.025 15.635 98.835 ;
        RECT 15.645 98.025 18.395 98.935 ;
        RECT 18.415 98.110 18.845 98.895 ;
        RECT 18.865 98.025 20.695 98.835 ;
        RECT 20.705 98.735 21.650 98.935 ;
        RECT 20.705 98.055 23.455 98.735 ;
        RECT 20.705 98.025 21.650 98.055 ;
        RECT 5.665 97.815 5.835 98.025 ;
        RECT 7.045 97.815 7.215 98.025 ;
        RECT 8.885 97.815 9.055 98.005 ;
        RECT 12.105 97.815 12.275 98.005 ;
        RECT 14.405 97.835 14.575 98.025 ;
        RECT 14.860 97.865 14.980 97.975 ;
        RECT 17.160 97.815 17.330 98.005 ;
        RECT 17.620 97.865 17.740 97.975 ;
        RECT 18.085 97.815 18.255 98.025 ;
        RECT 19.005 97.835 19.175 98.025 ;
        RECT 20.845 97.815 21.015 98.005 ;
        RECT 22.225 97.815 22.395 98.005 ;
        RECT 23.140 97.835 23.310 98.055 ;
        RECT 23.565 98.025 26.675 98.935 ;
        RECT 30.200 98.705 31.110 98.925 ;
        RECT 32.645 98.705 33.995 98.935 ;
        RECT 26.685 98.025 33.995 98.705 ;
        RECT 34.045 98.025 37.715 98.835 ;
        RECT 37.920 98.025 41.395 98.935 ;
        RECT 41.405 98.025 43.695 98.935 ;
        RECT 44.175 98.110 44.605 98.895 ;
        RECT 44.625 98.025 46.455 98.935 ;
        RECT 47.385 98.025 50.595 98.935 ;
        RECT 50.605 98.025 54.275 98.835 ;
        RECT 57.955 98.705 58.875 98.935 ;
        RECT 55.290 98.025 58.875 98.705 ;
        RECT 58.895 98.705 60.855 98.935 ;
        RECT 58.895 98.025 61.345 98.705 ;
        RECT 61.645 98.025 67.155 98.835 ;
        RECT 68.085 98.705 69.430 98.935 ;
        RECT 68.085 98.025 69.915 98.705 ;
        RECT 69.935 98.110 70.365 98.895 ;
        RECT 73.900 98.705 74.810 98.925 ;
        RECT 76.345 98.705 77.695 98.935 ;
        RECT 70.385 98.025 77.695 98.705 ;
        RECT 78.205 98.025 81.415 98.935 ;
        RECT 81.885 98.025 83.255 98.835 ;
        RECT 23.605 97.835 23.775 98.025 ;
        RECT 26.825 97.815 26.995 98.025 ;
        RECT 5.525 97.005 6.895 97.815 ;
        RECT 6.905 97.005 8.735 97.815 ;
        RECT 8.785 96.905 11.955 97.815 ;
        RECT 11.965 97.135 14.705 97.815 ;
        RECT 15.640 97.585 17.330 97.815 ;
        RECT 15.640 96.905 17.475 97.585 ;
        RECT 17.945 97.135 20.695 97.815 ;
        RECT 19.765 96.905 20.695 97.135 ;
        RECT 20.715 96.905 22.065 97.815 ;
        RECT 22.085 97.005 23.915 97.815 ;
        RECT 24.055 96.905 27.055 97.815 ;
        RECT 27.145 97.785 28.090 97.815 ;
        RECT 29.580 97.785 29.750 98.005 ;
        RECT 30.045 97.815 30.215 98.005 ;
        RECT 31.885 97.815 32.055 98.005 ;
        RECT 34.185 97.835 34.355 98.025 ;
        RECT 34.645 97.815 34.815 98.005 ;
        RECT 41.080 97.835 41.250 98.025 ;
        RECT 41.545 97.835 41.715 98.025 ;
        RECT 27.145 97.105 29.895 97.785 ;
        RECT 27.145 96.905 28.090 97.105 ;
        RECT 29.905 97.005 31.275 97.815 ;
        RECT 31.295 96.945 31.725 97.730 ;
        RECT 31.745 97.005 34.495 97.815 ;
        RECT 34.505 97.135 41.815 97.815 ;
        RECT 42.010 97.785 42.180 98.005 ;
        RECT 43.840 97.865 43.960 97.975 ;
        RECT 44.770 97.835 44.940 98.025 ;
        RECT 45.225 97.815 45.395 98.005 ;
        RECT 46.615 97.870 46.775 97.980 ;
        RECT 47.515 97.835 47.685 98.025 ;
        RECT 50.745 97.835 50.915 98.025 ;
        RECT 58.560 98.005 58.730 98.025 ;
        RECT 61.325 98.005 61.345 98.025 ;
        RECT 52.580 97.865 52.700 97.975 ;
        RECT 53.960 97.815 54.130 98.005 ;
        RECT 54.425 97.815 54.595 98.005 ;
        RECT 58.560 97.835 58.740 98.005 ;
        RECT 59.020 97.865 59.140 97.975 ;
        RECT 58.570 97.815 58.740 97.835 ;
        RECT 59.485 97.815 59.655 98.005 ;
        RECT 61.325 97.835 61.495 98.005 ;
        RECT 61.785 97.835 61.955 98.025 ;
        RECT 62.980 97.815 63.150 98.005 ;
        RECT 67.315 97.870 67.475 97.980 ;
        RECT 69.605 97.835 69.775 98.025 ;
        RECT 70.525 98.005 70.695 98.025 ;
        RECT 70.065 97.815 70.235 98.005 ;
        RECT 70.525 97.835 70.700 98.005 ;
        RECT 74.200 97.865 74.320 97.975 ;
        RECT 70.530 97.815 70.700 97.835 ;
        RECT 74.665 97.815 74.835 98.005 ;
        RECT 77.880 97.865 78.000 97.975 ;
        RECT 78.345 97.835 78.515 98.025 ;
        RECT 81.560 97.865 81.680 97.975 ;
        RECT 82.945 97.815 83.115 98.025 ;
        RECT 44.140 97.785 45.075 97.815 ;
        RECT 42.010 97.585 45.075 97.785 ;
        RECT 38.020 96.915 38.930 97.135 ;
        RECT 40.465 96.905 41.815 97.135 ;
        RECT 41.865 97.105 45.075 97.585 ;
        RECT 45.085 97.135 52.395 97.815 ;
        RECT 41.865 96.905 42.795 97.105 ;
        RECT 44.125 96.905 45.075 97.105 ;
        RECT 48.600 96.915 49.510 97.135 ;
        RECT 51.045 96.905 52.395 97.135 ;
        RECT 52.925 96.905 54.275 97.815 ;
        RECT 54.295 96.905 57.025 97.815 ;
        RECT 57.055 96.945 57.485 97.730 ;
        RECT 57.505 96.905 58.855 97.815 ;
        RECT 59.345 96.905 62.555 97.815 ;
        RECT 62.565 97.135 66.465 97.815 ;
        RECT 66.800 97.135 70.265 97.815 ;
        RECT 62.565 96.905 63.495 97.135 ;
        RECT 66.800 96.905 67.720 97.135 ;
        RECT 70.385 96.905 73.860 97.815 ;
        RECT 74.525 97.135 81.835 97.815 ;
        RECT 78.040 96.915 78.950 97.135 ;
        RECT 80.485 96.905 81.835 97.135 ;
        RECT 81.885 97.005 83.255 97.815 ;
      LAYER nwell ;
        RECT 5.330 93.785 83.450 96.615 ;
      LAYER pwell ;
        RECT 5.525 92.585 6.895 93.395 ;
        RECT 6.905 92.585 12.415 93.395 ;
        RECT 12.425 92.585 17.935 93.395 ;
        RECT 18.415 92.670 18.845 93.455 ;
        RECT 18.865 92.585 24.375 93.395 ;
        RECT 24.385 92.585 28.055 93.395 ;
        RECT 28.065 92.585 29.435 93.395 ;
        RECT 29.465 92.585 30.815 93.495 ;
        RECT 33.480 93.265 34.400 93.495 ;
        RECT 30.935 92.585 34.400 93.265 ;
        RECT 34.545 93.265 35.895 93.495 ;
        RECT 37.430 93.265 38.340 93.485 ;
        RECT 34.545 92.585 41.855 93.265 ;
        RECT 41.965 92.585 44.155 93.495 ;
        RECT 44.175 92.670 44.605 93.455 ;
        RECT 44.625 93.265 45.555 93.495 ;
        RECT 50.125 93.265 51.055 93.495 ;
        RECT 52.885 93.265 53.815 93.495 ;
        RECT 44.625 92.585 48.295 93.265 ;
        RECT 48.305 92.585 51.055 93.265 ;
        RECT 51.065 92.585 53.815 93.265 ;
        RECT 54.895 92.585 58.550 93.495 ;
        RECT 58.905 92.585 60.255 93.495 ;
        RECT 64.700 93.265 65.610 93.485 ;
        RECT 67.145 93.265 68.495 93.495 ;
        RECT 61.185 92.585 68.495 93.265 ;
        RECT 68.545 92.585 69.915 93.365 ;
        RECT 69.935 92.670 70.365 93.455 ;
        RECT 71.305 92.585 74.515 93.495 ;
        RECT 74.525 92.585 78.000 93.495 ;
        RECT 78.205 92.585 81.415 93.495 ;
        RECT 81.885 92.585 83.255 93.395 ;
        RECT 5.665 92.375 5.835 92.585 ;
        RECT 7.045 92.375 7.215 92.585 ;
        RECT 10.735 92.420 10.895 92.530 ;
        RECT 11.650 92.375 11.820 92.565 ;
        RECT 12.565 92.395 12.735 92.585 ;
        RECT 13.025 92.375 13.195 92.565 ;
        RECT 18.080 92.425 18.200 92.535 ;
        RECT 18.555 92.420 18.715 92.530 ;
        RECT 19.005 92.395 19.175 92.585 ;
        RECT 24.525 92.395 24.695 92.585 ;
        RECT 28.205 92.395 28.375 92.585 ;
        RECT 29.125 92.375 29.295 92.565 ;
        RECT 29.585 92.375 29.755 92.565 ;
        RECT 30.500 92.395 30.670 92.585 ;
        RECT 30.965 92.395 31.135 92.585 ;
        RECT 31.880 92.375 32.050 92.565 ;
        RECT 34.185 92.375 34.355 92.565 ;
        RECT 34.655 92.420 34.815 92.530 ;
        RECT 35.565 92.375 35.735 92.565 ;
        RECT 41.545 92.395 41.715 92.585 ;
        RECT 42.925 92.375 43.095 92.565 ;
        RECT 43.840 92.395 44.010 92.585 ;
        RECT 45.695 92.420 45.855 92.530 ;
        RECT 46.610 92.375 46.780 92.565 ;
        RECT 47.985 92.395 48.155 92.585 ;
        RECT 48.445 92.395 48.615 92.585 ;
        RECT 51.205 92.565 51.375 92.585 ;
        RECT 54.895 92.565 55.055 92.585 ;
        RECT 48.905 92.375 49.075 92.565 ;
        RECT 51.205 92.395 51.380 92.565 ;
        RECT 53.515 92.420 53.675 92.530 ;
        RECT 53.975 92.430 54.135 92.540 ;
        RECT 54.885 92.395 55.055 92.565 ;
        RECT 51.210 92.375 51.380 92.395 ;
        RECT 56.725 92.375 56.895 92.565 ;
        RECT 57.645 92.375 57.815 92.565 ;
        RECT 59.020 92.395 59.190 92.585 ;
        RECT 59.485 92.375 59.655 92.565 ;
        RECT 60.415 92.430 60.575 92.540 ;
        RECT 61.325 92.395 61.495 92.585 ;
        RECT 69.605 92.395 69.775 92.585 ;
        RECT 70.065 92.375 70.235 92.565 ;
        RECT 70.535 92.430 70.695 92.540 ;
        RECT 71.435 92.395 71.605 92.585 ;
        RECT 71.905 92.375 72.075 92.565 ;
        RECT 72.365 92.375 72.535 92.565 ;
        RECT 74.670 92.395 74.840 92.585 ;
        RECT 79.725 92.395 79.895 92.565 ;
        RECT 81.105 92.395 81.275 92.585 ;
        RECT 81.560 92.425 81.680 92.535 ;
        RECT 79.730 92.375 79.895 92.395 ;
        RECT 82.945 92.375 83.115 92.585 ;
        RECT 5.525 91.565 6.895 92.375 ;
        RECT 6.905 91.565 10.575 92.375 ;
        RECT 11.505 91.465 12.855 92.375 ;
        RECT 12.885 91.565 18.395 92.375 ;
        RECT 19.360 91.465 29.380 92.375 ;
        RECT 29.445 91.565 31.275 92.375 ;
        RECT 31.295 91.505 31.725 92.290 ;
        RECT 31.765 91.465 33.115 92.375 ;
        RECT 33.135 91.465 34.485 92.375 ;
        RECT 35.425 91.695 42.735 92.375 ;
        RECT 42.785 91.695 45.535 92.375 ;
        RECT 38.940 91.475 39.850 91.695 ;
        RECT 41.385 91.465 42.735 91.695 ;
        RECT 44.605 91.465 45.535 91.695 ;
        RECT 46.465 91.465 48.655 92.375 ;
        RECT 48.765 91.695 51.055 92.375 ;
        RECT 51.065 91.695 53.340 92.375 ;
        RECT 50.135 91.465 51.055 91.695 ;
        RECT 51.970 91.465 53.340 91.695 ;
        RECT 54.295 91.465 57.025 92.375 ;
        RECT 57.055 91.505 57.485 92.290 ;
        RECT 57.505 91.565 59.335 92.375 ;
        RECT 59.345 91.695 66.655 92.375 ;
        RECT 62.860 91.475 63.770 91.695 ;
        RECT 65.305 91.465 66.655 91.695 ;
        RECT 66.800 91.695 70.265 92.375 ;
        RECT 70.385 91.695 72.215 92.375 ;
        RECT 72.225 91.695 79.535 92.375 ;
        RECT 79.730 91.695 81.565 92.375 ;
        RECT 66.800 91.465 67.720 91.695 ;
        RECT 70.385 91.465 71.730 91.695 ;
        RECT 75.740 91.475 76.650 91.695 ;
        RECT 78.185 91.465 79.535 91.695 ;
        RECT 80.635 91.465 81.565 91.695 ;
        RECT 81.885 91.565 83.255 92.375 ;
      LAYER nwell ;
        RECT 5.330 88.345 83.450 91.175 ;
      LAYER pwell ;
        RECT 5.525 87.145 6.895 87.955 ;
        RECT 6.905 87.825 7.825 88.055 ;
        RECT 9.205 87.825 10.125 88.055 ;
        RECT 6.905 87.145 9.195 87.825 ;
        RECT 9.205 87.145 11.495 87.825 ;
        RECT 11.985 87.145 13.335 88.055 ;
        RECT 16.090 87.825 17.015 88.055 ;
        RECT 13.345 87.145 17.015 87.825 ;
        RECT 17.025 87.145 18.375 88.055 ;
        RECT 18.415 87.230 18.845 88.015 ;
        RECT 18.875 87.145 20.225 88.055 ;
        RECT 20.245 87.145 22.075 87.955 ;
        RECT 22.855 87.825 23.785 88.055 ;
        RECT 22.855 87.145 24.690 87.825 ;
        RECT 25.765 87.375 27.600 88.055 ;
        RECT 5.665 86.935 5.835 87.145 ;
        RECT 7.055 86.980 7.215 87.090 ;
        RECT 7.965 86.935 8.135 87.125 ;
        RECT 8.885 86.955 9.055 87.145 ;
        RECT 11.185 86.955 11.355 87.145 ;
        RECT 11.640 86.985 11.760 87.095 ;
        RECT 13.020 86.955 13.190 87.145 ;
        RECT 15.320 86.985 15.440 87.095 ;
        RECT 16.700 86.935 16.870 87.145 ;
        RECT 17.165 86.935 17.335 87.125 ;
        RECT 18.090 86.955 18.260 87.145 ;
        RECT 19.005 86.955 19.175 87.145 ;
        RECT 20.385 86.955 20.555 87.145 ;
        RECT 24.525 87.125 24.690 87.145 ;
        RECT 25.910 87.145 27.600 87.375 ;
        RECT 28.065 87.145 33.575 87.955 ;
        RECT 33.585 87.145 36.335 87.955 ;
        RECT 36.345 87.145 37.695 88.055 ;
        RECT 37.725 87.145 40.935 88.055 ;
        RECT 40.945 87.145 43.695 88.055 ;
        RECT 44.175 87.230 44.605 88.015 ;
        RECT 44.625 87.145 53.730 87.825 ;
        RECT 53.825 87.145 59.335 87.955 ;
        RECT 59.345 87.145 61.175 87.955 ;
        RECT 61.185 87.825 62.115 88.055 ;
        RECT 61.185 87.145 65.085 87.825 ;
        RECT 65.325 87.145 66.695 87.955 ;
        RECT 66.705 87.145 69.915 88.055 ;
        RECT 69.935 87.230 70.365 88.015 ;
        RECT 70.385 87.145 71.755 87.925 ;
        RECT 71.765 87.145 75.240 88.055 ;
        RECT 75.755 87.825 76.685 88.055 ;
        RECT 78.795 87.825 79.725 88.055 ;
        RECT 75.755 87.145 77.590 87.825 ;
        RECT 25.910 87.125 26.080 87.145 ;
        RECT 22.220 86.985 22.340 87.095 ;
        RECT 24.525 86.935 24.695 87.125 ;
        RECT 24.995 86.990 25.155 87.100 ;
        RECT 25.905 86.955 26.080 87.125 ;
        RECT 28.205 86.955 28.375 87.145 ;
        RECT 25.905 86.935 26.075 86.955 ;
        RECT 30.505 86.935 30.675 87.125 ;
        RECT 30.960 86.985 31.080 87.095 ;
        RECT 31.885 86.935 32.055 87.125 ;
        RECT 33.725 86.955 33.895 87.145 ;
        RECT 36.490 86.955 36.660 87.145 ;
        RECT 37.405 86.935 37.575 87.125 ;
        RECT 40.625 86.955 40.795 87.145 ;
        RECT 41.085 86.935 41.255 87.145 ;
        RECT 5.525 86.125 6.895 86.935 ;
        RECT 7.825 86.255 15.135 86.935 ;
        RECT 11.340 86.035 12.250 86.255 ;
        RECT 13.785 86.025 15.135 86.255 ;
        RECT 15.665 86.025 17.015 86.935 ;
        RECT 17.025 86.255 24.335 86.935 ;
        RECT 20.540 86.035 21.450 86.255 ;
        RECT 22.985 86.025 24.335 86.255 ;
        RECT 24.385 86.125 25.755 86.935 ;
        RECT 25.765 86.255 28.055 86.935 ;
        RECT 27.135 86.025 28.055 86.255 ;
        RECT 28.075 86.025 30.805 86.935 ;
        RECT 31.295 86.065 31.725 86.850 ;
        RECT 31.745 86.125 37.255 86.935 ;
        RECT 37.265 86.125 40.935 86.935 ;
        RECT 40.945 86.125 42.315 86.935 ;
        RECT 42.460 86.905 42.630 87.125 ;
        RECT 43.840 86.985 43.960 87.095 ;
        RECT 44.765 86.955 44.935 87.145 ;
        RECT 45.685 86.935 45.855 87.125 ;
        RECT 47.980 86.935 48.150 87.125 ;
        RECT 48.445 86.935 48.615 87.125 ;
        RECT 49.830 86.935 50.000 87.125 ;
        RECT 52.130 86.935 52.300 87.125 ;
        RECT 53.965 86.955 54.135 87.145 ;
        RECT 54.430 86.935 54.600 87.125 ;
        RECT 56.720 86.985 56.840 87.095 ;
        RECT 57.645 86.935 57.815 87.125 ;
        RECT 59.485 86.955 59.655 87.145 ;
        RECT 61.600 86.955 61.770 87.145 ;
        RECT 63.165 86.935 63.335 87.125 ;
        RECT 65.465 86.955 65.635 87.145 ;
        RECT 66.385 86.935 66.555 87.125 ;
        RECT 68.225 86.935 68.395 87.125 ;
        RECT 69.605 86.955 69.775 87.145 ;
        RECT 70.065 86.935 70.235 87.125 ;
        RECT 70.525 86.955 70.695 87.145 ;
        RECT 71.910 86.955 72.080 87.145 ;
        RECT 77.425 87.125 77.590 87.145 ;
        RECT 77.890 87.145 79.725 87.825 ;
        RECT 80.045 87.825 81.390 88.055 ;
        RECT 80.045 87.145 81.875 87.825 ;
        RECT 81.885 87.145 83.255 87.955 ;
        RECT 77.890 87.125 78.055 87.145 ;
        RECT 70.530 86.935 70.695 86.955 ;
        RECT 74.660 86.935 74.830 87.125 ;
        RECT 75.125 86.935 75.295 87.125 ;
        RECT 76.960 86.985 77.080 87.095 ;
        RECT 77.425 86.955 77.595 87.125 ;
        RECT 77.885 86.955 78.055 87.125 ;
        RECT 80.185 86.935 80.355 87.125 ;
        RECT 80.645 86.935 80.815 87.125 ;
        RECT 81.565 86.955 81.735 87.145 ;
        RECT 82.945 86.935 83.115 87.145 ;
        RECT 43.660 86.905 44.615 86.935 ;
        RECT 42.335 86.225 44.615 86.905 ;
        RECT 43.660 86.025 44.615 86.225 ;
        RECT 44.635 86.025 45.985 86.935 ;
        RECT 46.460 86.705 48.150 86.935 ;
        RECT 46.460 86.025 48.295 86.705 ;
        RECT 48.305 86.125 49.675 86.935 ;
        RECT 49.685 86.255 51.960 86.935 ;
        RECT 50.590 86.025 51.960 86.255 ;
        RECT 51.985 86.025 54.195 86.935 ;
        RECT 54.285 86.025 56.495 86.935 ;
        RECT 57.055 86.065 57.485 86.850 ;
        RECT 57.505 86.125 63.015 86.935 ;
        RECT 63.025 86.125 64.855 86.935 ;
        RECT 64.865 86.255 66.695 86.935 ;
        RECT 66.705 86.255 68.535 86.935 ;
        RECT 68.545 86.255 70.375 86.935 ;
        RECT 70.530 86.255 72.365 86.935 ;
        RECT 64.865 86.025 66.210 86.255 ;
        RECT 66.705 86.025 68.050 86.255 ;
        RECT 68.545 86.025 69.890 86.255 ;
        RECT 71.435 86.025 72.365 86.255 ;
        RECT 72.785 86.025 74.975 86.935 ;
        RECT 74.985 86.255 76.815 86.935 ;
        RECT 75.470 86.025 76.815 86.255 ;
        RECT 77.285 86.025 80.495 86.935 ;
        RECT 80.505 86.125 81.875 86.935 ;
        RECT 81.885 86.125 83.255 86.935 ;
      LAYER nwell ;
        RECT 5.330 82.905 83.450 85.735 ;
      LAYER pwell ;
        RECT 5.525 81.705 6.895 82.515 ;
        RECT 10.420 82.385 11.330 82.605 ;
        RECT 12.865 82.385 14.215 82.615 ;
        RECT 17.260 82.385 18.395 82.615 ;
        RECT 6.905 81.705 14.215 82.385 ;
        RECT 15.185 81.705 18.395 82.385 ;
        RECT 18.415 81.790 18.845 82.575 ;
        RECT 18.865 81.705 22.075 82.615 ;
        RECT 22.095 81.705 24.835 82.385 ;
        RECT 24.865 81.705 26.215 82.615 ;
        RECT 29.740 82.385 30.650 82.605 ;
        RECT 32.185 82.385 33.535 82.615 ;
        RECT 26.225 81.705 33.535 82.385 ;
        RECT 33.625 82.385 34.975 82.615 ;
        RECT 36.510 82.385 37.420 82.605 ;
        RECT 33.625 81.705 40.935 82.385 ;
        RECT 40.945 81.705 43.695 82.515 ;
        RECT 44.175 81.790 44.605 82.575 ;
        RECT 44.625 81.705 46.455 82.515 ;
        RECT 46.485 81.705 47.835 82.615 ;
        RECT 49.215 82.385 50.135 82.615 ;
        RECT 47.845 81.705 50.135 82.385 ;
        RECT 50.605 82.415 51.560 82.615 ;
        RECT 50.605 81.735 52.885 82.415 ;
        RECT 50.605 81.705 51.560 81.735 ;
        RECT 5.665 81.495 5.835 81.705 ;
        RECT 7.045 81.495 7.215 81.705 ;
        RECT 14.415 81.550 14.575 81.660 ;
        RECT 15.325 81.515 15.495 81.705 ;
        RECT 17.165 81.495 17.335 81.685 ;
        RECT 19.005 81.515 19.175 81.705 ;
        RECT 19.465 81.515 19.635 81.685 ;
        RECT 19.465 81.495 19.630 81.515 ;
        RECT 21.760 81.495 21.930 81.685 ;
        RECT 24.065 81.515 24.235 81.685 ;
        RECT 24.525 81.655 24.695 81.705 ;
        RECT 24.520 81.545 24.695 81.655 ;
        RECT 24.525 81.515 24.695 81.545 ;
        RECT 24.980 81.685 25.150 81.705 ;
        RECT 24.980 81.515 25.155 81.685 ;
        RECT 26.365 81.515 26.535 81.705 ;
        RECT 24.065 81.495 24.215 81.515 ;
        RECT 24.985 81.495 25.155 81.515 ;
        RECT 5.525 80.685 6.895 81.495 ;
        RECT 6.905 80.815 14.215 81.495 ;
        RECT 10.420 80.595 11.330 80.815 ;
        RECT 12.865 80.585 14.215 80.815 ;
        RECT 14.265 80.815 17.475 81.495 ;
        RECT 17.795 80.815 19.630 81.495 ;
        RECT 20.240 81.265 21.930 81.495 ;
        RECT 14.265 80.585 15.400 80.815 ;
        RECT 17.795 80.585 18.725 80.815 ;
        RECT 20.240 80.585 22.075 81.265 ;
        RECT 22.285 80.675 24.215 81.495 ;
        RECT 24.845 80.815 27.135 81.495 ;
        RECT 27.290 81.465 27.460 81.685 ;
        RECT 30.515 81.540 30.675 81.650 ;
        RECT 31.885 81.495 32.055 81.685 ;
        RECT 29.420 81.465 30.355 81.495 ;
        RECT 27.290 81.265 30.355 81.465 ;
        RECT 22.285 80.585 23.235 80.675 ;
        RECT 26.215 80.585 27.135 80.815 ;
        RECT 27.145 80.785 30.355 81.265 ;
        RECT 27.145 80.585 28.075 80.785 ;
        RECT 29.405 80.585 30.355 80.785 ;
        RECT 31.295 80.625 31.725 81.410 ;
        RECT 31.745 80.685 33.115 81.495 ;
        RECT 33.270 81.465 33.440 81.685 ;
        RECT 36.485 81.515 36.655 81.685 ;
        RECT 36.490 81.495 36.655 81.515 ;
        RECT 38.785 81.495 38.955 81.685 ;
        RECT 40.625 81.515 40.795 81.705 ;
        RECT 41.085 81.515 41.255 81.705 ;
        RECT 44.765 81.685 44.935 81.705 ;
        RECT 42.465 81.495 42.635 81.685 ;
        RECT 43.840 81.545 43.960 81.655 ;
        RECT 44.760 81.515 44.935 81.685 ;
        RECT 46.600 81.685 46.770 81.705 ;
        RECT 46.600 81.515 46.775 81.685 ;
        RECT 44.760 81.495 44.930 81.515 ;
        RECT 46.605 81.495 46.775 81.515 ;
        RECT 47.065 81.495 47.235 81.685 ;
        RECT 47.985 81.515 48.155 81.705 ;
        RECT 52.590 81.685 52.760 81.735 ;
        RECT 52.905 81.705 54.735 82.615 ;
        RECT 55.795 82.385 56.725 82.615 ;
        RECT 54.890 81.705 56.725 82.385 ;
        RECT 57.045 81.705 62.555 82.515 ;
        RECT 62.565 81.705 64.395 82.515 ;
        RECT 64.875 81.705 66.225 82.615 ;
        RECT 66.440 81.705 69.915 82.615 ;
        RECT 69.935 81.790 70.365 82.575 ;
        RECT 73.900 82.385 74.810 82.605 ;
        RECT 76.345 82.385 77.695 82.615 ;
        RECT 70.385 81.705 77.695 82.385 ;
        RECT 77.745 81.705 81.220 82.615 ;
        RECT 81.885 81.705 83.255 82.515 ;
        RECT 50.280 81.545 50.400 81.655 ;
        RECT 35.400 81.465 36.335 81.495 ;
        RECT 33.270 81.265 36.335 81.465 ;
        RECT 33.125 80.785 36.335 81.265 ;
        RECT 36.490 80.815 38.325 81.495 ;
        RECT 33.125 80.585 34.055 80.785 ;
        RECT 35.385 80.585 36.335 80.785 ;
        RECT 37.395 80.585 38.325 80.815 ;
        RECT 38.645 80.685 42.315 81.495 ;
        RECT 42.325 80.685 43.695 81.495 ;
        RECT 43.725 80.585 45.075 81.495 ;
        RECT 45.085 80.815 46.915 81.495 ;
        RECT 45.085 80.585 46.430 80.815 ;
        RECT 47.005 80.585 50.005 81.495 ;
        RECT 50.145 81.465 51.100 81.495 ;
        RECT 52.130 81.465 52.300 81.685 ;
        RECT 52.580 81.515 52.760 81.685 ;
        RECT 53.050 81.515 53.220 81.705 ;
        RECT 54.890 81.685 55.055 81.705 ;
        RECT 52.580 81.465 52.750 81.515 ;
        RECT 54.885 81.495 55.055 81.685 ;
        RECT 57.185 81.515 57.355 81.705 ;
        RECT 59.485 81.495 59.655 81.685 ;
        RECT 59.945 81.495 60.115 81.685 ;
        RECT 61.325 81.495 61.495 81.685 ;
        RECT 62.705 81.515 62.875 81.705 ;
        RECT 64.085 81.495 64.255 81.685 ;
        RECT 64.550 81.655 64.720 81.685 ;
        RECT 64.540 81.545 64.720 81.655 ;
        RECT 64.550 81.495 64.720 81.545 ;
        RECT 65.925 81.515 66.095 81.705 ;
        RECT 66.850 81.495 67.020 81.685 ;
        RECT 69.155 81.540 69.315 81.650 ;
        RECT 69.600 81.515 69.770 81.705 ;
        RECT 70.525 81.515 70.695 81.705 ;
        RECT 71.905 81.515 72.075 81.685 ;
        RECT 74.205 81.515 74.375 81.685 ;
        RECT 71.905 81.495 72.070 81.515 ;
        RECT 74.205 81.495 74.355 81.515 ;
        RECT 74.665 81.495 74.835 81.685 ;
        RECT 77.890 81.515 78.060 81.705 ;
        RECT 81.560 81.545 81.680 81.655 ;
        RECT 82.945 81.495 83.115 81.705 ;
        RECT 53.780 81.465 54.735 81.495 ;
        RECT 50.145 80.785 52.425 81.465 ;
        RECT 52.455 80.785 54.735 81.465 ;
        RECT 54.745 80.815 57.035 81.495 ;
        RECT 50.145 80.585 51.100 80.785 ;
        RECT 53.780 80.585 54.735 80.785 ;
        RECT 56.115 80.585 57.035 80.815 ;
        RECT 57.055 80.625 57.485 81.410 ;
        RECT 57.505 80.815 59.795 81.495 ;
        RECT 57.505 80.585 58.425 80.815 ;
        RECT 59.805 80.685 61.175 81.495 ;
        RECT 61.195 80.585 62.545 81.495 ;
        RECT 62.565 80.815 64.395 81.495 ;
        RECT 64.405 80.815 66.680 81.495 ;
        RECT 62.565 80.585 63.910 80.815 ;
        RECT 65.310 80.585 66.680 80.815 ;
        RECT 66.705 80.585 68.915 81.495 ;
        RECT 70.235 80.815 72.070 81.495 ;
        RECT 70.235 80.585 71.165 80.815 ;
        RECT 72.425 80.675 74.355 81.495 ;
        RECT 74.525 80.815 81.835 81.495 ;
        RECT 72.425 80.585 73.375 80.675 ;
        RECT 78.040 80.595 78.950 80.815 ;
        RECT 80.485 80.585 81.835 80.815 ;
        RECT 81.885 80.685 83.255 81.495 ;
      LAYER nwell ;
        RECT 5.330 77.465 83.450 80.295 ;
      LAYER pwell ;
        RECT 5.525 76.265 6.895 77.075 ;
        RECT 7.825 76.975 8.775 77.175 ;
        RECT 10.105 76.975 11.035 77.175 ;
        RECT 7.825 76.495 11.035 76.975 ;
        RECT 11.965 76.975 12.895 77.175 ;
        RECT 14.230 76.975 15.175 77.175 ;
        RECT 11.965 76.495 15.175 76.975 ;
        RECT 15.185 76.975 16.115 77.175 ;
        RECT 17.445 76.975 18.395 77.175 ;
        RECT 15.185 76.495 18.395 76.975 ;
        RECT 7.825 76.295 10.890 76.495 ;
        RECT 7.825 76.265 8.760 76.295 ;
        RECT 5.665 76.055 5.835 76.265 ;
        RECT 7.045 76.055 7.215 76.245 ;
        RECT 10.720 76.055 10.890 76.295 ;
        RECT 12.105 76.295 15.175 76.495 ;
        RECT 11.185 76.055 11.355 76.245 ;
        RECT 12.105 76.075 12.275 76.295 ;
        RECT 14.230 76.265 15.175 76.295 ;
        RECT 15.330 76.295 18.395 76.495 ;
        RECT 18.415 76.350 18.845 77.135 ;
        RECT 13.480 76.055 13.650 76.245 ;
        RECT 13.945 76.055 14.115 76.245 ;
        RECT 15.330 76.075 15.500 76.295 ;
        RECT 17.460 76.265 18.395 76.295 ;
        RECT 19.060 76.265 22.535 77.175 ;
        RECT 22.545 76.265 24.835 77.175 ;
        RECT 24.865 76.265 26.215 77.175 ;
        RECT 27.455 76.945 28.385 77.175 ;
        RECT 27.455 76.265 29.290 76.945 ;
        RECT 29.445 76.265 33.100 77.175 ;
        RECT 33.165 76.945 34.515 77.175 ;
        RECT 36.050 76.945 36.960 77.165 ;
        RECT 40.485 76.975 41.435 77.175 ;
        RECT 42.765 76.975 43.695 77.175 ;
        RECT 33.165 76.265 40.475 76.945 ;
        RECT 40.485 76.495 43.695 76.975 ;
        RECT 40.485 76.295 43.550 76.495 ;
        RECT 44.175 76.350 44.605 77.135 ;
        RECT 40.485 76.265 41.420 76.295 ;
        RECT 19.465 76.055 19.635 76.245 ;
        RECT 22.220 76.075 22.390 76.265 ;
        RECT 22.685 76.075 22.855 76.265 ;
        RECT 23.145 76.055 23.315 76.245 ;
        RECT 24.980 76.075 25.150 76.265 ;
        RECT 29.125 76.245 29.290 76.265 ;
        RECT 26.365 76.075 26.535 76.245 ;
        RECT 26.825 76.075 26.995 76.245 ;
        RECT 29.125 76.075 29.295 76.245 ;
        RECT 29.590 76.075 29.760 76.265 ;
        RECT 31.880 76.105 32.000 76.215 ;
        RECT 26.365 76.055 26.530 76.075 ;
        RECT 5.525 75.245 6.895 76.055 ;
        RECT 6.905 75.245 9.655 76.055 ;
        RECT 9.685 75.145 11.035 76.055 ;
        RECT 11.045 75.245 12.415 76.055 ;
        RECT 12.445 75.145 13.795 76.055 ;
        RECT 13.805 75.245 19.315 76.055 ;
        RECT 19.325 75.245 22.995 76.055 ;
        RECT 23.005 75.245 24.375 76.055 ;
        RECT 24.695 75.375 26.530 76.055 ;
        RECT 26.845 76.055 26.995 76.075 ;
        RECT 29.130 76.055 29.295 76.075 ;
        RECT 32.345 76.055 32.515 76.245 ;
        RECT 39.705 76.055 39.875 76.245 ;
        RECT 40.165 76.075 40.335 76.265 ;
        RECT 41.085 76.055 41.255 76.245 ;
        RECT 43.380 76.075 43.550 76.295 ;
        RECT 44.625 76.265 46.455 77.175 ;
        RECT 46.465 76.265 49.675 77.175 ;
        RECT 49.695 76.265 51.045 77.175 ;
        RECT 51.260 76.265 54.735 77.175 ;
        RECT 55.815 76.265 59.470 77.175 ;
        RECT 59.805 76.265 63.015 77.175 ;
        RECT 64.075 76.945 65.005 77.175 ;
        RECT 67.585 76.975 68.995 77.175 ;
        RECT 63.170 76.265 65.005 76.945 ;
        RECT 66.260 76.295 68.995 76.975 ;
        RECT 69.935 76.350 70.365 77.135 ;
        RECT 71.725 76.975 73.135 77.175 ;
        RECT 70.400 76.295 73.135 76.975 ;
        RECT 43.840 76.105 43.960 76.215 ;
        RECT 44.770 76.075 44.940 76.265 ;
        RECT 46.605 76.075 46.775 76.265 ;
        RECT 48.450 76.055 48.620 76.245 ;
        RECT 49.825 76.075 49.995 76.265 ;
        RECT 52.120 76.055 52.290 76.245 ;
        RECT 54.420 76.075 54.590 76.265 ;
        RECT 55.815 76.245 55.975 76.265 ;
        RECT 54.895 76.110 55.055 76.220 ;
        RECT 55.805 76.075 55.975 76.245 ;
        RECT 56.720 76.055 56.890 76.245 ;
        RECT 57.645 76.055 57.815 76.245 ;
        RECT 59.945 76.075 60.115 76.265 ;
        RECT 63.170 76.245 63.335 76.265 ;
        RECT 61.140 76.055 61.310 76.245 ;
        RECT 63.165 76.075 63.335 76.245 ;
        RECT 65.475 76.110 65.635 76.220 ;
        RECT 66.385 76.075 66.555 76.295 ;
        RECT 67.600 76.265 68.995 76.295 ;
        RECT 68.225 76.055 68.395 76.245 ;
        RECT 68.680 76.105 68.800 76.215 ;
        RECT 69.145 76.075 69.315 76.245 ;
        RECT 70.525 76.075 70.695 76.295 ;
        RECT 71.740 76.265 73.135 76.295 ;
        RECT 73.145 76.265 75.335 77.175 ;
        RECT 75.445 76.265 78.655 77.175 ;
        RECT 78.665 76.265 81.875 77.175 ;
        RECT 81.885 76.265 83.255 77.075 ;
        RECT 69.175 76.055 69.315 76.075 ;
        RECT 71.910 76.055 72.080 76.245 ;
        RECT 73.290 76.075 73.460 76.265 ;
        RECT 75.575 76.245 75.745 76.265 ;
        RECT 75.575 76.075 75.760 76.245 ;
        RECT 75.590 76.055 75.760 76.075 ;
        RECT 81.105 76.075 81.275 76.245 ;
        RECT 81.565 76.215 81.735 76.265 ;
        RECT 81.560 76.105 81.735 76.215 ;
        RECT 81.565 76.075 81.735 76.105 ;
        RECT 81.105 76.055 81.270 76.075 ;
        RECT 82.945 76.055 83.115 76.265 ;
        RECT 24.695 75.145 25.625 75.375 ;
        RECT 26.845 75.235 28.775 76.055 ;
        RECT 29.130 75.375 30.965 76.055 ;
        RECT 27.825 75.145 28.775 75.235 ;
        RECT 30.035 75.145 30.965 75.375 ;
        RECT 31.295 75.185 31.725 75.970 ;
        RECT 32.205 75.375 39.515 76.055 ;
        RECT 35.720 75.155 36.630 75.375 ;
        RECT 38.165 75.145 39.515 75.375 ;
        RECT 39.565 75.245 40.935 76.055 ;
        RECT 40.945 75.375 48.255 76.055 ;
        RECT 44.460 75.155 45.370 75.375 ;
        RECT 46.905 75.145 48.255 75.375 ;
        RECT 48.305 75.145 51.975 76.055 ;
        RECT 52.005 75.145 53.355 76.055 ;
        RECT 53.560 75.145 57.035 76.055 ;
        RECT 57.055 75.185 57.485 75.970 ;
        RECT 57.505 75.145 60.715 76.055 ;
        RECT 60.725 75.375 64.625 76.055 ;
        RECT 64.960 75.375 68.425 76.055 ;
        RECT 60.725 75.145 61.655 75.375 ;
        RECT 64.960 75.145 65.880 75.375 ;
        RECT 69.175 75.235 71.745 76.055 ;
        RECT 70.155 75.145 71.745 75.235 ;
        RECT 71.765 75.145 75.240 76.055 ;
        RECT 75.445 75.145 78.920 76.055 ;
        RECT 79.435 75.375 81.270 76.055 ;
        RECT 79.435 75.145 80.365 75.375 ;
        RECT 81.885 75.245 83.255 76.055 ;
      LAYER nwell ;
        RECT 5.330 72.025 83.450 74.855 ;
      LAYER pwell ;
        RECT 5.525 70.825 6.895 71.635 ;
        RECT 6.905 70.825 12.415 71.635 ;
        RECT 12.425 70.825 16.095 71.635 ;
        RECT 16.575 70.825 17.925 71.735 ;
        RECT 18.415 70.910 18.845 71.695 ;
        RECT 18.865 70.825 20.695 71.635 ;
        RECT 21.225 70.825 22.995 71.735 ;
        RECT 23.055 70.825 26.215 71.735 ;
        RECT 26.225 70.825 28.975 71.735 ;
        RECT 28.985 70.825 31.735 71.735 ;
        RECT 32.215 70.825 34.945 71.735 ;
        RECT 34.965 70.825 36.795 71.635 ;
        RECT 40.510 71.505 44.120 71.735 ;
        RECT 37.210 70.825 39.635 71.505 ;
        RECT 40.025 70.825 44.120 71.505 ;
        RECT 44.175 70.910 44.605 71.695 ;
        RECT 44.625 71.505 45.555 71.735 ;
        RECT 44.625 70.825 48.525 71.505 ;
        RECT 48.765 70.825 50.135 71.635 ;
        RECT 50.145 71.535 51.075 71.735 ;
        RECT 52.405 71.535 53.355 71.735 ;
        RECT 54.700 71.535 55.655 71.735 ;
        RECT 50.145 71.055 53.355 71.535 ;
        RECT 50.290 70.855 53.355 71.055 ;
        RECT 53.375 70.855 55.655 71.535 ;
        RECT 5.665 70.615 5.835 70.825 ;
        RECT 7.045 70.615 7.215 70.825 ;
        RECT 8.880 70.665 9.000 70.775 ;
        RECT 10.270 70.615 10.440 70.805 ;
        RECT 10.725 70.615 10.895 70.805 ;
        RECT 12.565 70.635 12.735 70.825 ;
        RECT 16.240 70.770 16.360 70.775 ;
        RECT 16.240 70.665 16.415 70.770 ;
        RECT 16.255 70.660 16.415 70.665 ;
        RECT 16.705 70.635 16.875 70.825 ;
        RECT 17.160 70.615 17.330 70.805 ;
        RECT 18.080 70.665 18.200 70.775 ;
        RECT 18.545 70.615 18.715 70.805 ;
        RECT 19.005 70.635 19.175 70.825 ;
        RECT 20.845 70.775 21.015 70.805 ;
        RECT 20.840 70.665 21.015 70.775 ;
        RECT 20.845 70.635 21.015 70.665 ;
        RECT 22.680 70.635 22.850 70.825 ;
        RECT 23.145 70.635 23.315 70.825 ;
        RECT 26.365 70.635 26.535 70.825 ;
        RECT 29.125 70.635 29.295 70.825 ;
        RECT 34.645 70.805 34.815 70.825 ;
        RECT 20.865 70.615 21.015 70.635 ;
        RECT 30.045 70.615 30.215 70.805 ;
        RECT 30.515 70.660 30.675 70.770 ;
        RECT 31.880 70.665 32.000 70.775 ;
        RECT 34.640 70.635 34.815 70.805 ;
        RECT 34.640 70.615 34.810 70.635 ;
        RECT 35.105 70.615 35.275 70.825 ;
        RECT 40.170 70.805 40.340 70.825 ;
        RECT 36.945 70.635 37.115 70.805 ;
        RECT 40.165 70.635 40.340 70.805 ;
        RECT 45.040 70.635 45.210 70.825 ;
        RECT 40.165 70.615 40.335 70.635 ;
        RECT 47.525 70.615 47.695 70.805 ;
        RECT 48.905 70.635 49.075 70.825 ;
        RECT 50.290 70.635 50.460 70.855 ;
        RECT 52.420 70.825 53.355 70.855 ;
        RECT 50.745 70.635 50.915 70.805 ;
        RECT 51.215 70.660 51.375 70.770 ;
        RECT 52.125 70.635 52.295 70.805 ;
        RECT 53.500 70.635 53.670 70.855 ;
        RECT 54.700 70.825 55.655 70.855 ;
        RECT 55.665 70.825 58.875 71.735 ;
        RECT 62.400 71.505 63.310 71.725 ;
        RECT 64.845 71.505 66.195 71.735 ;
        RECT 67.295 71.505 68.225 71.735 ;
        RECT 58.885 70.825 66.195 71.505 ;
        RECT 66.390 70.825 68.225 71.505 ;
        RECT 68.555 70.825 69.905 71.735 ;
        RECT 69.935 70.910 70.365 71.695 ;
        RECT 70.385 70.825 72.155 71.735 ;
        RECT 75.740 71.505 76.650 71.725 ;
        RECT 78.185 71.505 79.535 71.735 ;
        RECT 80.635 71.505 81.565 71.735 ;
        RECT 72.225 70.825 79.535 71.505 ;
        RECT 79.730 70.825 81.565 71.505 ;
        RECT 81.885 70.825 83.255 71.635 ;
        RECT 50.745 70.615 50.910 70.635 ;
        RECT 5.525 69.805 6.895 70.615 ;
        RECT 6.905 69.805 8.735 70.615 ;
        RECT 9.205 69.705 10.555 70.615 ;
        RECT 10.585 69.805 16.095 70.615 ;
        RECT 17.045 69.705 18.395 70.615 ;
        RECT 18.405 69.935 20.695 70.615 ;
        RECT 19.775 69.705 20.695 69.935 ;
        RECT 20.865 69.795 22.795 70.615 ;
        RECT 21.845 69.705 22.795 69.795 ;
        RECT 23.045 69.935 30.355 70.615 ;
        RECT 23.045 69.705 24.395 69.935 ;
        RECT 25.930 69.715 26.840 69.935 ;
        RECT 31.295 69.745 31.725 70.530 ;
        RECT 31.890 69.705 34.955 70.615 ;
        RECT 34.965 69.935 39.780 70.615 ;
        RECT 40.025 69.935 47.335 70.615 ;
        RECT 43.540 69.715 44.450 69.935 ;
        RECT 45.985 69.705 47.335 69.935 ;
        RECT 47.385 69.805 48.755 70.615 ;
        RECT 49.075 69.935 50.910 70.615 ;
        RECT 52.145 70.615 52.295 70.635 ;
        RECT 54.425 70.615 54.595 70.805 ;
        RECT 55.805 70.635 55.975 70.825 ;
        RECT 57.645 70.615 57.815 70.805 ;
        RECT 59.025 70.635 59.195 70.825 ;
        RECT 66.390 70.805 66.555 70.825 ;
        RECT 61.320 70.665 61.440 70.775 ;
        RECT 62.060 70.615 62.230 70.805 ;
        RECT 66.385 70.635 66.555 70.805 ;
        RECT 68.685 70.635 68.855 70.825 ;
        RECT 69.145 70.615 69.315 70.805 ;
        RECT 70.530 70.635 70.700 70.825 ;
        RECT 70.980 70.615 71.150 70.805 ;
        RECT 71.445 70.615 71.615 70.805 ;
        RECT 72.365 70.635 72.535 70.825 ;
        RECT 79.730 70.805 79.895 70.825 ;
        RECT 72.825 70.615 72.995 70.805 ;
        RECT 79.725 70.635 79.895 70.805 ;
        RECT 80.185 70.615 80.355 70.805 ;
        RECT 82.945 70.615 83.115 70.825 ;
        RECT 49.075 69.705 50.005 69.935 ;
        RECT 52.145 69.795 54.075 70.615 ;
        RECT 54.285 69.935 57.025 70.615 ;
        RECT 53.125 69.705 54.075 69.795 ;
        RECT 57.055 69.745 57.485 70.530 ;
        RECT 57.615 69.935 61.080 70.615 ;
        RECT 60.160 69.705 61.080 69.935 ;
        RECT 61.645 69.935 65.545 70.615 ;
        RECT 65.880 69.935 69.345 70.615 ;
        RECT 61.645 69.705 62.575 69.935 ;
        RECT 65.880 69.705 66.800 69.935 ;
        RECT 69.525 69.705 71.295 70.615 ;
        RECT 71.305 69.835 72.675 70.615 ;
        RECT 72.685 69.935 79.995 70.615 ;
        RECT 80.045 69.935 81.875 70.615 ;
        RECT 76.200 69.715 77.110 69.935 ;
        RECT 78.645 69.705 79.995 69.935 ;
        RECT 80.530 69.705 81.875 69.935 ;
        RECT 81.885 69.805 83.255 70.615 ;
      LAYER nwell ;
        RECT 5.330 66.585 83.450 69.415 ;
      LAYER pwell ;
        RECT 5.525 65.385 6.895 66.195 ;
        RECT 10.420 66.065 11.330 66.285 ;
        RECT 12.865 66.065 14.215 66.295 ;
        RECT 6.905 65.385 14.215 66.065 ;
        RECT 14.725 65.385 16.540 66.295 ;
        RECT 16.565 65.385 18.395 66.295 ;
        RECT 18.415 65.470 18.845 66.255 ;
        RECT 18.865 65.385 22.525 66.295 ;
        RECT 23.005 65.385 27.820 66.065 ;
        RECT 28.065 65.385 29.895 66.195 ;
        RECT 33.020 66.065 33.940 66.295 ;
        RECT 36.765 66.095 37.715 66.295 ;
        RECT 30.475 65.385 33.940 66.065 ;
        RECT 34.045 65.415 37.715 66.095 ;
        RECT 5.665 65.175 5.835 65.385 ;
        RECT 7.045 65.195 7.215 65.385 ;
        RECT 10.725 65.175 10.895 65.365 ;
        RECT 13.025 65.195 13.195 65.365 ;
        RECT 14.400 65.225 14.520 65.335 ;
        RECT 13.025 65.175 13.190 65.195 ;
        RECT 14.865 65.175 15.035 65.365 ;
        RECT 15.325 65.195 15.495 65.365 ;
        RECT 16.245 65.195 16.415 65.385 ;
        RECT 15.345 65.175 15.495 65.195 ;
        RECT 17.625 65.175 17.795 65.365 ;
        RECT 18.080 65.195 18.250 65.385 ;
        RECT 21.315 65.220 21.475 65.330 ;
        RECT 5.525 64.365 6.895 65.175 ;
        RECT 7.825 64.495 11.035 65.175 ;
        RECT 11.355 64.495 13.190 65.175 ;
        RECT 7.825 64.265 8.960 64.495 ;
        RECT 11.355 64.265 12.285 64.495 ;
        RECT 13.345 64.265 15.160 65.175 ;
        RECT 15.345 64.355 17.275 65.175 ;
        RECT 16.325 64.265 17.275 64.355 ;
        RECT 17.485 64.265 21.155 65.175 ;
        RECT 22.230 65.145 22.400 65.385 ;
        RECT 22.680 65.225 22.800 65.335 ;
        RECT 23.145 65.195 23.315 65.385 ;
        RECT 25.445 65.195 25.615 65.365 ;
        RECT 28.205 65.195 28.375 65.385 ;
        RECT 29.580 65.225 29.700 65.335 ;
        RECT 25.455 65.175 25.615 65.195 ;
        RECT 30.040 65.175 30.210 65.365 ;
        RECT 30.505 65.195 30.675 65.385 ;
        RECT 32.805 65.175 32.975 65.365 ;
        RECT 34.190 65.195 34.360 65.415 ;
        RECT 36.765 65.385 37.715 65.415 ;
        RECT 37.725 65.385 39.095 66.195 ;
        RECT 39.200 66.065 40.120 66.295 ;
        RECT 39.200 65.385 42.665 66.065 ;
        RECT 42.785 65.385 44.155 66.195 ;
        RECT 44.175 65.470 44.605 66.255 ;
        RECT 44.625 65.385 48.295 66.195 ;
        RECT 49.710 66.065 51.055 66.295 ;
        RECT 49.225 65.385 51.055 66.065 ;
        RECT 51.065 65.385 52.895 66.295 ;
        RECT 55.560 66.065 56.480 66.295 ;
        RECT 53.015 65.385 56.480 66.065 ;
        RECT 56.585 65.385 59.795 66.295 ;
        RECT 63.320 66.065 64.230 66.285 ;
        RECT 65.765 66.065 67.115 66.295 ;
        RECT 59.805 65.385 67.115 66.065 ;
        RECT 68.085 66.065 69.430 66.295 ;
        RECT 68.085 65.385 69.915 66.065 ;
        RECT 69.935 65.470 70.365 66.255 ;
        RECT 70.480 66.065 71.400 66.295 ;
        RECT 76.390 66.065 77.735 66.295 ;
        RECT 70.480 65.385 73.945 66.065 ;
        RECT 74.065 65.385 75.895 66.065 ;
        RECT 75.905 65.385 77.735 66.065 ;
        RECT 77.745 65.385 80.955 66.295 ;
        RECT 81.885 65.385 83.255 66.195 ;
        RECT 37.865 65.195 38.035 65.385 ;
        RECT 40.165 65.175 40.335 65.365 ;
        RECT 42.465 65.195 42.635 65.385 ;
        RECT 42.925 65.195 43.095 65.385 ;
        RECT 42.925 65.175 42.945 65.195 ;
        RECT 43.660 65.175 43.830 65.365 ;
        RECT 44.765 65.195 44.935 65.385 ;
        RECT 48.455 65.230 48.615 65.340 ;
        RECT 49.365 65.195 49.535 65.385 ;
        RECT 50.745 65.175 50.915 65.365 ;
        RECT 51.215 65.220 51.375 65.330 ;
        RECT 52.400 65.175 52.570 65.365 ;
        RECT 52.580 65.195 52.750 65.385 ;
        RECT 53.045 65.195 53.215 65.385 ;
        RECT 56.275 65.220 56.435 65.330 ;
        RECT 56.725 65.195 56.895 65.385 ;
        RECT 57.920 65.175 58.090 65.365 ;
        RECT 59.945 65.195 60.115 65.385 ;
        RECT 61.780 65.225 61.900 65.335 ;
        RECT 62.520 65.175 62.690 65.365 ;
        RECT 66.660 65.175 66.830 65.365 ;
        RECT 67.315 65.230 67.475 65.340 ;
        RECT 69.605 65.195 69.775 65.385 ;
        RECT 73.745 65.175 73.915 65.385 ;
        RECT 75.585 65.195 75.755 65.385 ;
        RECT 76.045 65.365 76.215 65.385 ;
        RECT 76.040 65.195 76.215 65.365 ;
        RECT 76.040 65.175 76.210 65.195 ;
        RECT 76.505 65.175 76.675 65.365 ;
        RECT 77.885 65.175 78.055 65.365 ;
        RECT 80.645 65.195 80.815 65.385 ;
        RECT 81.115 65.220 81.275 65.340 ;
        RECT 82.945 65.175 83.115 65.385 ;
        RECT 24.360 65.145 25.295 65.175 ;
        RECT 22.230 64.945 25.295 65.145 ;
        RECT 22.085 64.465 25.295 64.945 ;
        RECT 22.085 64.265 23.015 64.465 ;
        RECT 24.345 64.265 25.295 64.465 ;
        RECT 25.455 64.265 29.110 65.175 ;
        RECT 29.925 64.265 31.275 65.175 ;
        RECT 31.295 64.305 31.725 65.090 ;
        RECT 31.755 64.265 33.105 65.175 ;
        RECT 33.165 64.495 40.475 65.175 ;
        RECT 40.495 64.495 42.945 65.175 ;
        RECT 43.245 64.495 47.145 65.175 ;
        RECT 47.480 64.495 50.945 65.175 ;
        RECT 51.985 64.495 55.885 65.175 ;
        RECT 33.165 64.265 34.515 64.495 ;
        RECT 36.050 64.275 36.960 64.495 ;
        RECT 40.495 64.265 42.455 64.495 ;
        RECT 43.245 64.265 44.175 64.495 ;
        RECT 47.480 64.265 48.400 64.495 ;
        RECT 51.985 64.265 52.915 64.495 ;
        RECT 57.055 64.305 57.485 65.090 ;
        RECT 57.505 64.495 61.405 65.175 ;
        RECT 62.105 64.495 66.005 65.175 ;
        RECT 66.245 64.495 70.145 65.175 ;
        RECT 70.480 64.495 73.945 65.175 ;
        RECT 57.505 64.265 58.435 64.495 ;
        RECT 62.105 64.265 63.035 64.495 ;
        RECT 66.245 64.265 67.175 64.495 ;
        RECT 70.480 64.265 71.400 64.495 ;
        RECT 74.165 64.265 76.355 65.175 ;
        RECT 76.365 64.395 77.735 65.175 ;
        RECT 77.745 64.265 80.955 65.175 ;
        RECT 81.885 64.365 83.255 65.175 ;
      LAYER nwell ;
        RECT 5.330 61.145 83.450 63.975 ;
      LAYER pwell ;
        RECT 5.525 59.945 6.895 60.755 ;
        RECT 7.380 59.945 9.195 60.855 ;
        RECT 10.575 60.625 11.495 60.855 ;
        RECT 9.205 59.945 11.495 60.625 ;
        RECT 11.505 60.625 12.640 60.855 ;
        RECT 11.505 59.945 14.715 60.625 ;
        RECT 15.645 59.945 18.395 60.855 ;
        RECT 18.415 60.030 18.845 60.815 ;
        RECT 18.865 59.945 20.695 60.755 ;
        RECT 22.780 60.625 23.915 60.855 ;
        RECT 27.440 60.625 28.350 60.845 ;
        RECT 29.885 60.625 31.235 60.855 ;
        RECT 20.705 59.945 23.915 60.625 ;
        RECT 23.925 59.945 31.235 60.625 ;
        RECT 31.295 59.945 34.025 60.855 ;
        RECT 37.560 60.625 38.470 60.845 ;
        RECT 40.005 60.625 41.355 60.855 ;
        RECT 42.455 60.625 43.385 60.855 ;
        RECT 34.045 59.945 41.355 60.625 ;
        RECT 41.550 59.945 43.385 60.625 ;
        RECT 44.175 60.030 44.605 60.815 ;
        RECT 44.635 59.945 45.985 60.855 ;
        RECT 46.005 60.625 46.935 60.855 ;
        RECT 50.185 60.625 51.535 60.855 ;
        RECT 53.070 60.625 53.980 60.845 ;
        RECT 57.965 60.625 59.310 60.855 ;
        RECT 63.320 60.625 64.230 60.845 ;
        RECT 65.765 60.625 67.115 60.855 ;
        RECT 46.005 59.945 49.905 60.625 ;
        RECT 50.185 59.945 57.495 60.625 ;
        RECT 57.965 59.945 59.795 60.625 ;
        RECT 59.805 59.945 67.115 60.625 ;
        RECT 67.165 59.945 69.255 60.755 ;
        RECT 69.935 60.030 70.365 60.815 ;
        RECT 70.385 59.945 75.200 60.625 ;
        RECT 75.445 59.945 78.920 60.855 ;
        RECT 80.175 60.625 81.105 60.855 ;
        RECT 79.270 59.945 81.105 60.625 ;
        RECT 81.885 59.945 83.255 60.755 ;
        RECT 5.665 59.735 5.835 59.945 ;
        RECT 7.040 59.785 7.160 59.895 ;
        RECT 7.505 59.755 7.675 59.945 ;
        RECT 9.345 59.755 9.515 59.945 ;
        RECT 13.945 59.735 14.115 59.925 ;
        RECT 14.405 59.755 14.575 59.945 ;
        RECT 14.875 59.790 15.035 59.900 ;
        RECT 15.785 59.755 15.955 59.945 ;
        RECT 16.245 59.735 16.415 59.925 ;
        RECT 16.705 59.735 16.875 59.925 ;
        RECT 18.540 59.785 18.660 59.895 ;
        RECT 19.005 59.755 19.175 59.945 ;
        RECT 20.845 59.755 21.015 59.945 ;
        RECT 21.765 59.735 21.935 59.925 ;
        RECT 22.230 59.735 22.400 59.925 ;
        RECT 23.605 59.735 23.775 59.925 ;
        RECT 24.065 59.755 24.235 59.945 ;
        RECT 5.525 58.925 6.895 59.735 ;
        RECT 6.945 59.055 14.255 59.735 ;
        RECT 14.265 59.055 16.555 59.735 ;
        RECT 16.565 59.055 18.395 59.735 ;
        RECT 6.945 58.825 8.295 59.055 ;
        RECT 9.830 58.835 10.740 59.055 ;
        RECT 14.265 58.825 15.185 59.055 ;
        RECT 18.865 58.825 22.075 59.735 ;
        RECT 22.085 58.825 23.435 59.735 ;
        RECT 23.465 58.925 24.835 59.735 ;
        RECT 24.845 59.705 25.780 59.735 ;
        RECT 27.740 59.705 27.910 59.925 ;
        RECT 28.205 59.735 28.375 59.925 ;
        RECT 30.960 59.785 31.080 59.895 ;
        RECT 31.425 59.755 31.595 59.945 ;
        RECT 31.885 59.735 32.055 59.925 ;
        RECT 33.265 59.735 33.435 59.925 ;
        RECT 34.185 59.755 34.355 59.945 ;
        RECT 41.550 59.925 41.715 59.945 ;
        RECT 34.645 59.735 34.815 59.925 ;
        RECT 36.945 59.735 37.115 59.925 ;
        RECT 38.780 59.785 38.900 59.895 ;
        RECT 39.245 59.735 39.415 59.925 ;
        RECT 41.545 59.755 41.715 59.925 ;
        RECT 43.840 59.785 43.960 59.895 ;
        RECT 45.685 59.755 45.855 59.945 ;
        RECT 46.420 59.755 46.590 59.945 ;
        RECT 46.610 59.735 46.780 59.925 ;
        RECT 56.725 59.735 56.895 59.925 ;
        RECT 57.185 59.755 57.355 59.945 ;
        RECT 57.645 59.895 57.815 59.925 ;
        RECT 57.640 59.785 57.815 59.895 ;
        RECT 57.645 59.735 57.815 59.785 ;
        RECT 59.485 59.755 59.655 59.945 ;
        RECT 59.945 59.755 60.115 59.945 ;
        RECT 60.405 59.735 60.575 59.925 ;
        RECT 67.305 59.755 67.475 59.945 ;
        RECT 69.145 59.735 69.315 59.925 ;
        RECT 69.605 59.755 69.775 59.925 ;
        RECT 70.525 59.755 70.695 59.945 ;
        RECT 71.905 59.755 72.075 59.925 ;
        RECT 74.200 59.785 74.320 59.895 ;
        RECT 69.625 59.735 69.775 59.755 ;
        RECT 71.910 59.735 72.075 59.755 ;
        RECT 74.665 59.735 74.835 59.925 ;
        RECT 75.590 59.755 75.760 59.945 ;
        RECT 79.270 59.925 79.435 59.945 ;
        RECT 79.265 59.755 79.435 59.925 ;
        RECT 81.560 59.785 81.680 59.895 ;
        RECT 82.945 59.735 83.115 59.945 ;
        RECT 24.845 59.505 27.910 59.705 ;
        RECT 24.845 59.025 28.055 59.505 ;
        RECT 24.845 58.825 25.795 59.025 ;
        RECT 27.125 58.825 28.055 59.025 ;
        RECT 28.075 58.825 30.805 59.735 ;
        RECT 31.295 58.865 31.725 59.650 ;
        RECT 31.745 58.925 33.115 59.735 ;
        RECT 33.125 58.955 34.495 59.735 ;
        RECT 34.505 59.055 36.795 59.735 ;
        RECT 35.875 58.825 36.795 59.055 ;
        RECT 36.805 58.925 38.635 59.735 ;
        RECT 39.105 59.055 46.415 59.735 ;
        RECT 42.620 58.835 43.530 59.055 ;
        RECT 45.065 58.825 46.415 59.055 ;
        RECT 46.465 58.825 49.580 59.735 ;
        RECT 49.725 59.055 57.035 59.735 ;
        RECT 49.725 58.825 51.075 59.055 ;
        RECT 52.610 58.835 53.520 59.055 ;
        RECT 57.055 58.865 57.485 59.650 ;
        RECT 57.505 58.925 60.255 59.735 ;
        RECT 60.265 59.055 67.575 59.735 ;
        RECT 63.780 58.835 64.690 59.055 ;
        RECT 66.225 58.825 67.575 59.055 ;
        RECT 67.625 59.055 69.455 59.735 ;
        RECT 67.625 58.825 68.970 59.055 ;
        RECT 69.625 58.915 71.555 59.735 ;
        RECT 71.910 59.055 73.745 59.735 ;
        RECT 74.525 59.055 81.835 59.735 ;
        RECT 70.605 58.825 71.555 58.915 ;
        RECT 72.815 58.825 73.745 59.055 ;
        RECT 78.040 58.835 78.950 59.055 ;
        RECT 80.485 58.825 81.835 59.055 ;
        RECT 81.885 58.925 83.255 59.735 ;
      LAYER nwell ;
        RECT 5.330 55.705 83.450 58.535 ;
      LAYER pwell ;
        RECT 5.525 54.505 6.895 55.315 ;
        RECT 10.420 55.185 11.330 55.405 ;
        RECT 12.865 55.185 14.215 55.415 ;
        RECT 6.905 54.505 14.215 55.185 ;
        RECT 14.265 54.505 15.615 55.415 ;
        RECT 15.645 54.505 18.395 55.315 ;
        RECT 18.415 54.590 18.845 55.375 ;
        RECT 18.865 54.505 21.615 55.315 ;
        RECT 21.625 54.505 22.975 55.415 ;
        RECT 23.025 54.505 24.375 55.415 ;
        RECT 24.385 54.505 26.215 55.315 ;
        RECT 26.225 55.185 27.145 55.415 ;
        RECT 26.225 54.505 28.515 55.185 ;
        RECT 28.525 54.505 34.035 55.315 ;
        RECT 34.045 54.505 39.555 55.315 ;
        RECT 39.565 54.505 41.395 55.315 ;
        RECT 43.235 55.185 44.155 55.415 ;
        RECT 41.865 54.505 44.155 55.185 ;
        RECT 44.175 54.590 44.605 55.375 ;
        RECT 45.995 55.215 47.350 55.415 ;
        RECT 44.670 55.185 47.350 55.215 ;
        RECT 49.215 55.185 50.135 55.415 ;
        RECT 44.670 54.535 47.835 55.185 ;
        RECT 45.995 54.505 47.835 54.535 ;
        RECT 47.845 54.505 50.135 55.185 ;
        RECT 50.145 54.505 55.655 55.315 ;
        RECT 55.665 54.505 58.415 55.315 ;
        RECT 58.425 54.505 63.240 55.185 ;
        RECT 63.485 54.505 65.315 55.315 ;
        RECT 65.425 54.505 67.615 55.415 ;
        RECT 67.825 55.325 68.775 55.415 ;
        RECT 67.825 54.505 69.755 55.325 ;
        RECT 69.935 54.590 70.365 55.375 ;
        RECT 71.040 54.505 74.515 55.415 ;
        RECT 78.040 55.185 78.950 55.405 ;
        RECT 80.485 55.185 81.835 55.415 ;
        RECT 74.525 54.505 81.835 55.185 ;
        RECT 81.885 54.505 83.255 55.315 ;
        RECT 5.665 54.295 5.835 54.505 ;
        RECT 7.045 54.295 7.215 54.505 ;
        RECT 10.265 54.295 10.435 54.485 ;
        RECT 10.725 54.295 10.895 54.485 ;
        RECT 13.480 54.295 13.650 54.485 ;
        RECT 13.945 54.295 14.115 54.485 ;
        RECT 14.410 54.315 14.580 54.505 ;
        RECT 15.785 54.315 15.955 54.505 ;
        RECT 19.005 54.315 19.175 54.505 ;
        RECT 19.460 54.345 19.580 54.455 ;
        RECT 19.930 54.295 20.100 54.485 ;
        RECT 22.690 54.315 22.860 54.505 ;
        RECT 23.140 54.315 23.310 54.505 ;
        RECT 24.525 54.315 24.695 54.505 ;
        RECT 27.745 54.315 27.915 54.485 ;
        RECT 28.205 54.315 28.375 54.505 ;
        RECT 28.665 54.315 28.835 54.505 ;
        RECT 27.750 54.295 27.915 54.315 ;
        RECT 30.045 54.295 30.215 54.485 ;
        RECT 31.885 54.295 32.055 54.485 ;
        RECT 34.185 54.315 34.355 54.505 ;
        RECT 35.565 54.295 35.735 54.485 ;
        RECT 38.325 54.295 38.495 54.485 ;
        RECT 38.785 54.295 38.955 54.485 ;
        RECT 39.705 54.315 39.875 54.505 ;
        RECT 41.540 54.345 41.660 54.455 ;
        RECT 42.005 54.315 42.175 54.505 ;
        RECT 42.460 54.295 42.630 54.485 ;
        RECT 42.925 54.295 43.095 54.485 ;
        RECT 46.605 54.315 46.775 54.485 ;
        RECT 47.525 54.315 47.695 54.505 ;
        RECT 47.985 54.315 48.155 54.505 ;
        RECT 46.605 54.295 46.770 54.315 ;
        RECT 48.440 54.295 48.610 54.485 ;
        RECT 48.905 54.295 49.075 54.485 ;
        RECT 50.285 54.315 50.455 54.505 ;
        RECT 54.425 54.295 54.595 54.485 ;
        RECT 55.805 54.315 55.975 54.505 ;
        RECT 57.655 54.340 57.815 54.450 ;
        RECT 58.565 54.295 58.735 54.505 ;
        RECT 61.785 54.295 61.955 54.485 ;
        RECT 63.625 54.315 63.795 54.505 ;
        RECT 67.300 54.485 67.470 54.505 ;
        RECT 69.605 54.485 69.755 54.505 ;
        RECT 65.460 54.345 65.580 54.455 ;
        RECT 67.300 54.315 67.475 54.485 ;
        RECT 67.305 54.295 67.475 54.315 ;
        RECT 69.145 54.295 69.315 54.485 ;
        RECT 69.605 54.315 69.775 54.485 ;
        RECT 70.515 54.295 70.685 54.485 ;
        RECT 74.200 54.295 74.370 54.505 ;
        RECT 74.665 54.295 74.835 54.505 ;
        RECT 82.945 54.295 83.115 54.505 ;
        RECT 5.525 53.485 6.895 54.295 ;
        RECT 6.905 53.485 8.275 54.295 ;
        RECT 8.285 53.615 10.575 54.295 ;
        RECT 10.585 53.615 12.415 54.295 ;
        RECT 8.285 53.385 9.205 53.615 ;
        RECT 12.445 53.385 13.795 54.295 ;
        RECT 13.805 53.485 19.315 54.295 ;
        RECT 19.785 53.385 27.535 54.295 ;
        RECT 27.750 53.615 29.585 54.295 ;
        RECT 28.655 53.385 29.585 53.615 ;
        RECT 29.905 53.485 31.275 54.295 ;
        RECT 31.295 53.425 31.725 54.210 ;
        RECT 31.745 53.485 35.415 54.295 ;
        RECT 35.425 53.485 36.795 54.295 ;
        RECT 36.805 53.385 38.620 54.295 ;
        RECT 38.645 53.485 41.395 54.295 ;
        RECT 41.425 53.385 42.775 54.295 ;
        RECT 42.785 53.485 44.615 54.295 ;
        RECT 44.935 53.615 46.770 54.295 ;
        RECT 44.935 53.385 45.865 53.615 ;
        RECT 46.925 53.385 48.755 54.295 ;
        RECT 48.765 53.485 54.275 54.295 ;
        RECT 54.285 53.485 57.035 54.295 ;
        RECT 57.055 53.425 57.485 54.210 ;
        RECT 58.475 53.385 61.635 54.295 ;
        RECT 61.645 53.485 65.315 54.295 ;
        RECT 65.785 53.615 67.615 54.295 ;
        RECT 67.625 53.615 69.455 54.295 ;
        RECT 65.785 53.385 67.130 53.615 ;
        RECT 67.625 53.385 68.970 53.615 ;
        RECT 69.465 53.515 70.835 54.295 ;
        RECT 71.040 53.385 74.515 54.295 ;
        RECT 74.525 53.615 81.835 54.295 ;
        RECT 78.040 53.395 78.950 53.615 ;
        RECT 80.485 53.385 81.835 53.615 ;
        RECT 81.885 53.485 83.255 54.295 ;
      LAYER nwell ;
        RECT 5.330 50.265 83.450 53.095 ;
      LAYER pwell ;
        RECT 5.525 49.065 6.895 49.875 ;
        RECT 6.905 49.065 12.415 49.875 ;
        RECT 12.425 49.065 15.175 49.875 ;
        RECT 15.655 49.065 18.385 49.975 ;
        RECT 18.415 49.150 18.845 49.935 ;
        RECT 26.265 49.745 27.615 49.975 ;
        RECT 29.150 49.745 30.060 49.965 ;
        RECT 33.585 49.775 34.515 49.975 ;
        RECT 35.845 49.775 36.795 49.975 ;
        RECT 19.325 49.065 21.155 49.745 ;
        RECT 21.400 49.065 26.215 49.745 ;
        RECT 26.265 49.065 33.575 49.745 ;
        RECT 33.585 49.295 36.795 49.775 ;
        RECT 39.460 49.745 40.380 49.975 ;
        RECT 33.730 49.095 36.795 49.295 ;
        RECT 5.665 48.855 5.835 49.065 ;
        RECT 7.045 48.855 7.215 49.065 ;
        RECT 12.565 48.855 12.735 49.065 ;
        RECT 13.950 48.855 14.120 49.045 ;
        RECT 15.320 48.905 15.440 49.015 ;
        RECT 15.785 48.855 15.955 49.065 ;
        RECT 19.005 49.015 19.175 49.045 ;
        RECT 19.000 48.905 19.175 49.015 ;
        RECT 19.005 48.855 19.175 48.905 ;
        RECT 19.465 48.875 19.635 49.065 ;
        RECT 22.695 48.900 22.855 49.010 ;
        RECT 25.905 48.875 26.075 49.065 ;
        RECT 27.285 48.875 27.455 49.045 ;
        RECT 27.285 48.855 27.430 48.875 ;
        RECT 30.045 48.855 30.215 49.045 ;
        RECT 30.515 48.900 30.675 49.010 ;
        RECT 33.265 48.875 33.435 49.065 ;
        RECT 33.730 49.045 33.900 49.095 ;
        RECT 35.860 49.065 36.795 49.095 ;
        RECT 36.915 49.065 40.380 49.745 ;
        RECT 40.500 49.065 42.315 49.975 ;
        RECT 42.805 49.065 44.155 49.975 ;
        RECT 44.175 49.150 44.605 49.935 ;
        RECT 44.720 49.745 45.640 49.975 ;
        RECT 49.320 49.745 50.240 49.975 ;
        RECT 44.720 49.065 48.185 49.745 ;
        RECT 49.320 49.065 52.785 49.745 ;
        RECT 52.905 49.065 55.655 49.875 ;
        RECT 59.180 49.745 60.090 49.965 ;
        RECT 61.625 49.745 62.975 49.975 ;
        RECT 55.665 49.065 62.975 49.745 ;
        RECT 63.025 49.065 64.395 49.875 ;
        RECT 64.405 49.745 65.750 49.975 ;
        RECT 64.405 49.065 66.235 49.745 ;
        RECT 66.245 49.065 69.720 49.975 ;
        RECT 69.935 49.150 70.365 49.935 ;
        RECT 73.900 49.745 74.810 49.965 ;
        RECT 76.345 49.745 77.695 49.975 ;
        RECT 70.385 49.065 77.695 49.745 ;
        RECT 78.055 49.745 78.985 49.975 ;
        RECT 80.530 49.745 81.875 49.975 ;
        RECT 78.055 49.065 79.890 49.745 ;
        RECT 80.045 49.065 81.875 49.745 ;
        RECT 81.885 49.065 83.255 49.875 ;
        RECT 33.725 48.875 33.900 49.045 ;
        RECT 34.180 48.905 34.300 49.015 ;
        RECT 36.945 48.875 37.115 49.065 ;
        RECT 40.625 48.875 40.795 49.065 ;
        RECT 33.725 48.855 33.895 48.875 ;
        RECT 41.545 48.855 41.715 49.045 ;
        RECT 42.005 48.855 42.175 49.045 ;
        RECT 42.460 48.905 42.580 49.015 ;
        RECT 43.840 48.875 44.010 49.065 ;
        RECT 45.685 48.855 45.855 49.045 ;
        RECT 47.985 48.875 48.155 49.065 ;
        RECT 48.455 49.015 48.615 49.020 ;
        RECT 48.440 48.910 48.615 49.015 ;
        RECT 48.440 48.905 48.560 48.910 ;
        RECT 48.905 48.855 49.075 49.045 ;
        RECT 52.585 48.875 52.755 49.065 ;
        RECT 53.045 48.875 53.215 49.065 ;
        RECT 55.805 48.875 55.975 49.065 ;
        RECT 56.720 48.905 56.840 49.015 ;
        RECT 57.645 48.855 57.815 49.045 ;
        RECT 63.165 48.875 63.335 49.065 ;
        RECT 65.465 48.855 65.635 49.045 ;
        RECT 65.925 48.875 66.095 49.065 ;
        RECT 66.390 48.875 66.560 49.065 ;
        RECT 70.525 48.875 70.695 49.065 ;
        RECT 79.725 49.045 79.890 49.065 ;
        RECT 75.585 48.855 75.755 49.045 ;
        RECT 76.055 48.900 76.215 49.010 ;
        RECT 76.965 48.875 77.135 49.045 ;
        RECT 79.265 48.875 79.435 49.045 ;
        RECT 79.725 48.875 79.895 49.045 ;
        RECT 80.185 48.875 80.355 49.065 ;
        RECT 81.560 48.905 81.680 49.015 ;
        RECT 76.970 48.855 77.135 48.875 ;
        RECT 79.270 48.855 79.435 48.875 ;
        RECT 82.945 48.855 83.115 49.065 ;
        RECT 5.525 48.045 6.895 48.855 ;
        RECT 6.905 48.045 12.415 48.855 ;
        RECT 12.425 48.045 13.795 48.855 ;
        RECT 13.805 47.945 15.635 48.855 ;
        RECT 15.745 47.945 18.855 48.855 ;
        RECT 18.865 48.175 22.535 48.855 ;
        RECT 21.605 47.945 22.535 48.175 ;
        RECT 23.560 47.945 27.430 48.855 ;
        RECT 27.605 48.175 30.355 48.855 ;
        RECT 27.605 47.945 28.535 48.175 ;
        RECT 31.295 47.985 31.725 48.770 ;
        RECT 31.745 48.175 34.035 48.855 ;
        RECT 34.545 48.175 41.855 48.855 ;
        RECT 41.975 48.175 45.440 48.855 ;
        RECT 31.745 47.945 32.665 48.175 ;
        RECT 34.545 47.945 35.895 48.175 ;
        RECT 37.430 47.955 38.340 48.175 ;
        RECT 44.520 47.945 45.440 48.175 ;
        RECT 45.545 47.945 48.295 48.855 ;
        RECT 48.765 48.175 56.495 48.855 ;
        RECT 52.280 47.955 53.190 48.175 ;
        RECT 54.725 47.945 56.495 48.175 ;
        RECT 57.055 47.985 57.485 48.770 ;
        RECT 57.505 48.175 65.235 48.855 ;
        RECT 65.325 48.175 72.635 48.855 ;
        RECT 61.020 47.955 61.930 48.175 ;
        RECT 63.465 47.945 65.235 48.175 ;
        RECT 68.840 47.955 69.750 48.175 ;
        RECT 71.285 47.945 72.635 48.175 ;
        RECT 72.685 47.945 75.895 48.855 ;
        RECT 76.970 48.175 78.805 48.855 ;
        RECT 79.270 48.175 81.105 48.855 ;
        RECT 77.875 47.945 78.805 48.175 ;
        RECT 80.175 47.945 81.105 48.175 ;
        RECT 81.885 48.045 83.255 48.855 ;
      LAYER nwell ;
        RECT 5.330 44.825 83.450 47.655 ;
      LAYER pwell ;
        RECT 5.525 43.625 6.895 44.435 ;
        RECT 6.905 43.625 8.735 44.435 ;
        RECT 8.745 44.305 9.665 44.535 ;
        RECT 8.745 43.625 11.035 44.305 ;
        RECT 11.045 43.625 12.860 44.535 ;
        RECT 12.885 43.625 15.635 44.435 ;
        RECT 17.155 44.305 18.085 44.535 ;
        RECT 16.250 43.625 18.085 44.305 ;
        RECT 18.415 43.710 18.845 44.495 ;
        RECT 20.670 44.335 21.615 44.535 ;
        RECT 18.865 43.655 21.615 44.335 ;
        RECT 5.665 43.415 5.835 43.625 ;
        RECT 7.045 43.435 7.215 43.625 ;
        RECT 10.725 43.435 10.895 43.625 ;
        RECT 12.565 43.435 12.735 43.625 ;
        RECT 13.025 43.435 13.195 43.625 ;
        RECT 16.250 43.605 16.415 43.625 ;
        RECT 13.945 43.415 14.115 43.605 ;
        RECT 14.405 43.415 14.575 43.605 ;
        RECT 15.780 43.465 15.900 43.575 ;
        RECT 16.245 43.435 16.415 43.605 ;
        RECT 16.710 43.415 16.880 43.605 ;
        RECT 18.085 43.415 18.255 43.605 ;
        RECT 19.010 43.435 19.180 43.655 ;
        RECT 20.670 43.625 21.615 43.655 ;
        RECT 22.545 43.625 25.755 44.535 ;
        RECT 38.020 44.305 38.930 44.525 ;
        RECT 40.465 44.305 41.815 44.535 ;
        RECT 43.235 44.305 44.155 44.535 ;
        RECT 26.630 43.625 29.055 44.305 ;
        RECT 29.680 43.625 34.495 44.305 ;
        RECT 34.505 43.625 41.815 44.305 ;
        RECT 41.865 43.625 44.155 44.305 ;
        RECT 44.175 43.710 44.605 44.495 ;
        RECT 48.140 44.305 49.050 44.525 ;
        RECT 50.585 44.305 51.935 44.535 ;
        RECT 57.045 44.305 57.975 44.535 ;
        RECT 68.500 44.335 69.455 44.535 ;
        RECT 44.625 43.625 51.935 44.305 ;
        RECT 52.220 43.625 57.035 44.305 ;
        RECT 57.045 43.625 60.945 44.305 ;
        RECT 62.340 43.625 67.155 44.305 ;
        RECT 67.175 43.655 69.455 44.335 ;
        RECT 69.935 43.710 70.365 44.495 ;
        RECT 70.695 44.305 71.625 44.535 ;
        RECT 21.775 43.470 21.935 43.580 ;
        RECT 22.685 43.435 22.855 43.625 ;
        RECT 23.605 43.435 23.775 43.605 ;
        RECT 23.605 43.415 23.770 43.435 ;
        RECT 24.065 43.415 24.235 43.605 ;
        RECT 25.900 43.465 26.020 43.575 ;
        RECT 26.365 43.415 26.535 43.605 ;
        RECT 29.585 43.415 29.755 43.605 ;
        RECT 33.725 43.435 33.895 43.605 ;
        RECT 34.185 43.575 34.355 43.625 ;
        RECT 34.180 43.465 34.355 43.575 ;
        RECT 34.185 43.435 34.355 43.465 ;
        RECT 33.725 43.415 33.875 43.435 ;
        RECT 34.645 43.415 34.815 43.625 ;
        RECT 42.005 43.415 42.175 43.625 ;
        RECT 44.765 43.435 44.935 43.625 ;
        RECT 49.365 43.415 49.535 43.605 ;
        RECT 52.400 43.415 52.570 43.605 ;
        RECT 56.275 43.460 56.435 43.570 ;
        RECT 56.725 43.435 56.895 43.625 ;
        RECT 57.460 43.435 57.630 43.625 ;
        RECT 66.845 43.605 67.015 43.625 ;
        RECT 57.655 43.460 57.815 43.570 ;
        RECT 58.840 43.415 59.010 43.605 ;
        RECT 61.335 43.470 61.495 43.580 ;
        RECT 62.980 43.415 63.150 43.605 ;
        RECT 66.845 43.435 67.020 43.605 ;
        RECT 67.300 43.435 67.470 43.655 ;
        RECT 68.500 43.625 69.455 43.655 ;
        RECT 70.695 43.625 72.530 44.305 ;
        RECT 72.685 43.625 74.055 44.435 ;
        RECT 74.065 43.625 77.540 44.535 ;
        RECT 78.055 44.305 78.985 44.535 ;
        RECT 80.530 44.305 81.875 44.535 ;
        RECT 78.055 43.625 79.890 44.305 ;
        RECT 80.045 43.625 81.875 44.305 ;
        RECT 81.885 43.625 83.255 44.435 ;
        RECT 72.365 43.605 72.530 43.625 ;
        RECT 69.600 43.465 69.720 43.575 ;
        RECT 70.520 43.465 70.640 43.575 ;
        RECT 72.365 43.435 72.535 43.605 ;
        RECT 72.825 43.435 72.995 43.625 ;
        RECT 74.210 43.605 74.380 43.625 ;
        RECT 79.725 43.605 79.890 43.625 ;
        RECT 74.200 43.435 74.380 43.605 ;
        RECT 66.850 43.415 67.020 43.435 ;
        RECT 74.200 43.415 74.370 43.435 ;
        RECT 74.665 43.415 74.835 43.605 ;
        RECT 79.725 43.435 79.895 43.605 ;
        RECT 80.185 43.435 80.355 43.625 ;
        RECT 82.945 43.415 83.115 43.625 ;
        RECT 5.525 42.605 6.895 43.415 ;
        RECT 6.945 42.735 14.255 43.415 ;
        RECT 14.265 42.735 16.555 43.415 ;
        RECT 6.945 42.505 8.295 42.735 ;
        RECT 9.830 42.515 10.740 42.735 ;
        RECT 15.635 42.505 16.555 42.735 ;
        RECT 16.565 42.505 17.915 43.415 ;
        RECT 17.945 42.605 21.615 43.415 ;
        RECT 21.935 42.735 23.770 43.415 ;
        RECT 23.925 42.735 26.215 43.415 ;
        RECT 21.935 42.505 22.865 42.735 ;
        RECT 25.295 42.505 26.215 42.735 ;
        RECT 26.305 42.505 29.305 43.415 ;
        RECT 29.445 42.605 31.275 43.415 ;
        RECT 31.295 42.545 31.725 43.330 ;
        RECT 31.945 42.595 33.875 43.415 ;
        RECT 34.505 42.735 41.815 43.415 ;
        RECT 41.865 42.735 49.175 43.415 ;
        RECT 31.945 42.505 32.895 42.595 ;
        RECT 38.020 42.515 38.930 42.735 ;
        RECT 40.465 42.505 41.815 42.735 ;
        RECT 45.380 42.515 46.290 42.735 ;
        RECT 47.825 42.505 49.175 42.735 ;
        RECT 49.225 42.605 51.315 43.415 ;
        RECT 51.985 42.735 55.885 43.415 ;
        RECT 51.985 42.505 52.915 42.735 ;
        RECT 57.055 42.545 57.485 43.330 ;
        RECT 58.425 42.735 62.325 43.415 ;
        RECT 62.565 42.735 66.465 43.415 ;
        RECT 58.425 42.505 59.355 42.735 ;
        RECT 62.565 42.505 63.495 42.735 ;
        RECT 66.705 42.505 70.180 43.415 ;
        RECT 71.040 42.505 74.515 43.415 ;
        RECT 74.525 42.735 81.835 43.415 ;
        RECT 78.040 42.515 78.950 42.735 ;
        RECT 80.485 42.505 81.835 42.735 ;
        RECT 81.885 42.605 83.255 43.415 ;
      LAYER nwell ;
        RECT 5.330 39.385 83.450 42.215 ;
      LAYER pwell ;
        RECT 5.525 38.185 6.895 38.995 ;
        RECT 11.340 38.865 12.250 39.085 ;
        RECT 13.785 38.865 15.135 39.095 ;
        RECT 7.825 38.185 15.135 38.865 ;
        RECT 15.185 38.865 16.320 39.095 ;
        RECT 15.185 38.185 18.395 38.865 ;
        RECT 18.415 38.270 18.845 39.055 ;
        RECT 18.865 38.185 20.680 39.095 ;
        RECT 20.705 38.185 22.055 39.095 ;
        RECT 22.085 38.185 25.755 38.995 ;
        RECT 25.765 38.895 26.715 39.095 ;
        RECT 28.045 38.895 28.975 39.095 ;
        RECT 25.765 38.415 28.975 38.895 ;
        RECT 28.985 38.865 30.120 39.095 ;
        RECT 25.765 38.215 28.830 38.415 ;
        RECT 25.765 38.185 26.700 38.215 ;
        RECT 5.665 37.975 5.835 38.185 ;
        RECT 7.965 38.165 8.135 38.185 ;
        RECT 7.055 38.030 7.215 38.140 ;
        RECT 7.960 37.995 8.135 38.165 ;
        RECT 7.960 37.975 8.130 37.995 ;
        RECT 8.425 37.975 8.595 38.165 ;
        RECT 17.625 37.975 17.795 38.165 ;
        RECT 18.085 38.135 18.255 38.185 ;
        RECT 18.080 38.025 18.255 38.135 ;
        RECT 18.085 37.995 18.255 38.025 ;
        RECT 20.385 37.995 20.555 38.185 ;
        RECT 20.850 37.995 21.020 38.185 ;
        RECT 22.225 38.165 22.395 38.185 ;
        RECT 21.760 37.975 21.930 38.165 ;
        RECT 22.225 37.995 22.400 38.165 ;
        RECT 22.230 37.975 22.400 37.995 ;
        RECT 24.065 37.975 24.235 38.165 ;
        RECT 28.660 37.995 28.830 38.215 ;
        RECT 28.985 38.185 32.195 38.865 ;
        RECT 32.205 38.185 35.125 39.095 ;
        RECT 35.735 38.865 36.665 39.095 ;
        RECT 35.735 38.185 37.570 38.865 ;
        RECT 37.725 38.185 39.095 38.995 ;
        RECT 39.125 38.185 40.475 39.095 ;
        RECT 40.580 38.865 41.500 39.095 ;
        RECT 40.580 38.185 44.045 38.865 ;
        RECT 44.175 38.270 44.605 39.055 ;
        RECT 44.625 38.895 45.580 39.095 ;
        RECT 44.625 38.215 46.905 38.895 ;
        RECT 47.425 38.865 48.775 39.095 ;
        RECT 50.310 38.865 51.220 39.085 ;
        RECT 56.085 38.895 57.465 39.095 ;
        RECT 44.625 38.185 45.580 38.215 ;
        RECT 31.885 37.975 32.055 38.185 ;
        RECT 32.350 37.995 32.520 38.185 ;
        RECT 37.405 38.165 37.570 38.185 ;
        RECT 37.405 37.995 37.575 38.165 ;
        RECT 37.865 37.995 38.035 38.185 ;
        RECT 39.240 38.165 39.410 38.185 ;
        RECT 39.240 37.995 39.420 38.165 ;
        RECT 39.250 37.975 39.420 37.995 ;
        RECT 41.085 37.975 41.255 38.165 ;
        RECT 43.845 37.995 44.015 38.185 ;
        RECT 44.315 38.020 44.475 38.130 ;
        RECT 45.225 37.975 45.395 38.165 ;
        RECT 46.610 37.995 46.780 38.215 ;
        RECT 47.425 38.185 54.735 38.865 ;
        RECT 54.760 38.215 57.465 38.895 ;
        RECT 61.020 38.865 61.930 39.085 ;
        RECT 63.465 38.865 65.235 39.095 ;
        RECT 47.060 38.025 47.180 38.135 ;
        RECT 54.425 37.995 54.595 38.185 ;
        RECT 54.885 37.995 55.055 38.215 ;
        RECT 56.085 38.185 57.465 38.215 ;
        RECT 57.505 38.185 65.235 38.865 ;
        RECT 65.325 38.895 66.270 39.095 ;
        RECT 67.605 38.895 68.535 39.095 ;
        RECT 65.325 38.415 68.535 38.895 ;
        RECT 65.325 38.215 68.395 38.415 ;
        RECT 65.325 38.185 66.270 38.215 ;
        RECT 55.805 37.975 55.975 38.165 ;
        RECT 56.275 38.020 56.435 38.130 ;
        RECT 57.645 37.975 57.815 38.185 ;
        RECT 65.465 37.975 65.635 38.165 ;
        RECT 68.225 37.995 68.395 38.215 ;
        RECT 68.545 38.185 69.915 38.995 ;
        RECT 69.935 38.270 70.365 39.055 ;
        RECT 70.580 38.185 74.055 39.095 ;
        RECT 78.040 38.865 78.950 39.085 ;
        RECT 80.485 38.865 81.835 39.095 ;
        RECT 74.525 38.185 81.835 38.865 ;
        RECT 81.885 38.185 83.255 38.995 ;
        RECT 68.685 37.995 68.855 38.185 ;
        RECT 73.740 37.995 73.910 38.185 ;
        RECT 74.200 38.025 74.320 38.135 ;
        RECT 74.665 37.995 74.835 38.185 ;
        RECT 79.725 37.975 79.895 38.165 ;
        RECT 80.185 37.975 80.355 38.165 ;
        RECT 82.945 37.975 83.115 38.185 ;
        RECT 5.525 37.165 6.895 37.975 ;
        RECT 6.925 37.065 8.275 37.975 ;
        RECT 8.285 37.295 15.595 37.975 ;
        RECT 11.800 37.075 12.710 37.295 ;
        RECT 14.245 37.065 15.595 37.295 ;
        RECT 15.645 37.295 17.935 37.975 ;
        RECT 15.645 37.065 16.565 37.295 ;
        RECT 18.600 37.065 22.075 37.975 ;
        RECT 22.085 37.065 23.915 37.975 ;
        RECT 23.925 37.295 31.235 37.975 ;
        RECT 27.440 37.075 28.350 37.295 ;
        RECT 29.885 37.065 31.235 37.295 ;
        RECT 31.295 37.105 31.725 37.890 ;
        RECT 31.745 37.295 39.055 37.975 ;
        RECT 35.260 37.075 36.170 37.295 ;
        RECT 37.705 37.065 39.055 37.295 ;
        RECT 39.105 37.065 40.935 37.975 ;
        RECT 41.045 37.065 44.155 37.975 ;
        RECT 45.085 37.295 52.395 37.975 ;
        RECT 48.600 37.075 49.510 37.295 ;
        RECT 51.045 37.065 52.395 37.295 ;
        RECT 52.540 37.295 56.005 37.975 ;
        RECT 52.540 37.065 53.460 37.295 ;
        RECT 57.055 37.105 57.485 37.890 ;
        RECT 57.505 37.295 65.235 37.975 ;
        RECT 65.325 37.295 72.635 37.975 ;
        RECT 61.020 37.075 61.930 37.295 ;
        RECT 63.465 37.065 65.235 37.295 ;
        RECT 68.840 37.075 69.750 37.295 ;
        RECT 71.285 37.065 72.635 37.295 ;
        RECT 72.725 37.295 80.035 37.975 ;
        RECT 80.045 37.295 81.875 37.975 ;
        RECT 72.725 37.065 74.075 37.295 ;
        RECT 75.610 37.075 76.520 37.295 ;
        RECT 80.530 37.065 81.875 37.295 ;
        RECT 81.885 37.165 83.255 37.975 ;
      LAYER nwell ;
        RECT 5.330 33.945 83.450 36.775 ;
      LAYER pwell ;
        RECT 5.525 32.745 6.895 33.555 ;
        RECT 7.405 32.745 10.575 33.655 ;
        RECT 11.955 33.425 12.875 33.655 ;
        RECT 15.175 33.425 16.095 33.655 ;
        RECT 17.475 33.425 18.395 33.655 ;
        RECT 10.585 32.745 12.875 33.425 ;
        RECT 13.805 32.745 16.095 33.425 ;
        RECT 16.105 32.745 18.395 33.425 ;
        RECT 18.415 32.830 18.845 33.615 ;
        RECT 22.380 33.425 23.290 33.645 ;
        RECT 24.825 33.425 26.175 33.655 ;
        RECT 18.865 32.745 26.175 33.425 ;
        RECT 26.225 32.745 27.575 33.655 ;
        RECT 31.120 33.425 32.030 33.645 ;
        RECT 33.565 33.425 34.915 33.655 ;
        RECT 27.605 32.745 34.915 33.425 ;
        RECT 34.965 33.425 35.885 33.655 ;
        RECT 34.965 32.745 37.255 33.425 ;
        RECT 37.265 32.745 39.095 33.555 ;
        RECT 39.105 32.745 40.455 33.655 ;
        RECT 40.485 32.745 44.155 33.555 ;
        RECT 44.175 32.830 44.605 33.615 ;
        RECT 44.625 32.745 45.995 33.555 ;
        RECT 46.100 33.425 47.020 33.655 ;
        RECT 49.780 33.425 50.700 33.655 ;
        RECT 56.105 33.425 57.035 33.655 ;
        RECT 46.100 32.745 49.565 33.425 ;
        RECT 49.780 32.745 53.245 33.425 ;
        RECT 53.365 32.745 57.035 33.425 ;
        RECT 57.505 33.425 58.435 33.655 ;
        RECT 57.505 32.745 61.405 33.425 ;
        RECT 61.645 32.745 63.015 33.555 ;
        RECT 63.025 33.425 64.370 33.655 ;
        RECT 63.025 32.745 64.855 33.425 ;
        RECT 64.865 32.745 68.340 33.655 ;
        RECT 68.545 32.745 69.915 33.555 ;
        RECT 69.935 32.830 70.365 33.615 ;
        RECT 70.385 32.745 73.595 33.655 ;
        RECT 78.040 33.425 78.950 33.645 ;
        RECT 80.485 33.425 81.835 33.655 ;
        RECT 74.525 32.745 81.835 33.425 ;
        RECT 81.885 32.745 83.255 33.555 ;
        RECT 5.665 32.535 5.835 32.745 ;
        RECT 7.045 32.695 7.215 32.725 ;
        RECT 7.040 32.585 7.215 32.695 ;
        RECT 7.045 32.535 7.215 32.585 ;
        RECT 7.505 32.555 7.675 32.745 ;
        RECT 10.725 32.555 10.895 32.745 ;
        RECT 12.560 32.585 12.680 32.695 ;
        RECT 13.025 32.535 13.195 32.725 ;
        RECT 13.945 32.555 14.115 32.745 ;
        RECT 16.245 32.535 16.415 32.745 ;
        RECT 19.005 32.555 19.175 32.745 ;
        RECT 25.445 32.535 25.615 32.725 ;
        RECT 25.905 32.535 26.075 32.725 ;
        RECT 26.370 32.555 26.540 32.745 ;
        RECT 27.745 32.555 27.915 32.745 ;
        RECT 29.585 32.535 29.755 32.725 ;
        RECT 30.045 32.535 30.215 32.725 ;
        RECT 31.885 32.535 32.055 32.725 ;
        RECT 34.645 32.535 34.815 32.725 ;
        RECT 36.945 32.555 37.115 32.745 ;
        RECT 37.405 32.555 37.575 32.745 ;
        RECT 40.170 32.725 40.340 32.745 ;
        RECT 40.165 32.555 40.340 32.725 ;
        RECT 40.625 32.555 40.795 32.745 ;
        RECT 44.765 32.555 44.935 32.745 ;
        RECT 40.165 32.535 40.335 32.555 ;
        RECT 45.685 32.535 45.855 32.725 ;
        RECT 48.450 32.535 48.620 32.725 ;
        RECT 48.910 32.535 49.080 32.725 ;
        RECT 49.365 32.555 49.535 32.745 ;
        RECT 50.755 32.580 50.915 32.690 ;
        RECT 53.045 32.555 53.215 32.745 ;
        RECT 53.505 32.535 53.675 32.745 ;
        RECT 5.525 31.725 6.895 32.535 ;
        RECT 6.905 31.725 12.415 32.535 ;
        RECT 12.925 31.625 16.095 32.535 ;
        RECT 16.105 31.855 23.415 32.535 ;
        RECT 19.620 31.635 20.530 31.855 ;
        RECT 22.065 31.625 23.415 31.855 ;
        RECT 23.465 31.855 25.755 32.535 ;
        RECT 23.465 31.625 24.385 31.855 ;
        RECT 25.765 31.725 27.135 32.535 ;
        RECT 27.145 31.855 29.895 32.535 ;
        RECT 27.145 31.625 28.075 31.855 ;
        RECT 29.905 31.725 31.275 32.535 ;
        RECT 31.295 31.665 31.725 32.450 ;
        RECT 31.755 31.625 34.485 32.535 ;
        RECT 34.505 31.725 40.015 32.535 ;
        RECT 40.025 31.725 45.535 32.535 ;
        RECT 45.545 31.725 47.375 32.535 ;
        RECT 47.385 31.625 48.735 32.535 ;
        RECT 48.765 31.625 50.595 32.535 ;
        RECT 51.525 31.855 53.815 32.535 ;
        RECT 53.970 32.505 54.140 32.725 ;
        RECT 57.180 32.585 57.300 32.695 ;
        RECT 56.100 32.505 57.035 32.535 ;
        RECT 53.970 32.305 57.035 32.505 ;
        RECT 57.645 32.505 57.815 32.725 ;
        RECT 57.920 32.555 58.090 32.745 ;
        RECT 60.875 32.580 61.035 32.690 ;
        RECT 61.785 32.555 61.955 32.745 ;
        RECT 63.165 32.535 63.335 32.725 ;
        RECT 64.545 32.555 64.715 32.745 ;
        RECT 65.010 32.725 65.180 32.745 ;
        RECT 65.005 32.555 65.180 32.725 ;
        RECT 67.305 32.555 67.475 32.725 ;
        RECT 68.685 32.555 68.855 32.745 ;
        RECT 69.605 32.555 69.775 32.725 ;
        RECT 70.060 32.585 70.180 32.695 ;
        RECT 70.525 32.555 70.695 32.745 ;
        RECT 72.365 32.555 72.535 32.725 ;
        RECT 65.005 32.535 65.175 32.555 ;
        RECT 67.305 32.535 67.470 32.555 ;
        RECT 69.605 32.535 69.770 32.555 ;
        RECT 72.365 32.535 72.530 32.555 ;
        RECT 72.825 32.535 72.995 32.725 ;
        RECT 73.755 32.590 73.915 32.700 ;
        RECT 74.665 32.555 74.835 32.745 ;
        RECT 77.880 32.535 78.050 32.725 ;
        RECT 81.105 32.535 81.275 32.725 ;
        RECT 81.560 32.585 81.680 32.695 ;
        RECT 82.945 32.535 83.115 32.745 ;
        RECT 59.770 32.505 60.715 32.535 ;
        RECT 51.525 31.625 52.445 31.855 ;
        RECT 53.825 31.825 57.035 32.305 ;
        RECT 53.825 31.625 54.755 31.825 ;
        RECT 56.085 31.625 57.035 31.825 ;
        RECT 57.055 31.665 57.485 32.450 ;
        RECT 57.645 32.305 60.715 32.505 ;
        RECT 57.505 31.825 60.715 32.305 ;
        RECT 57.505 31.625 58.435 31.825 ;
        RECT 59.770 31.625 60.715 31.825 ;
        RECT 61.645 31.855 63.475 32.535 ;
        RECT 63.485 31.855 65.315 32.535 ;
        RECT 65.635 31.855 67.470 32.535 ;
        RECT 67.935 31.855 69.770 32.535 ;
        RECT 70.695 31.855 72.530 32.535 ;
        RECT 72.685 31.855 74.515 32.535 ;
        RECT 61.645 31.625 62.990 31.855 ;
        RECT 63.485 31.625 64.830 31.855 ;
        RECT 65.635 31.625 66.565 31.855 ;
        RECT 67.935 31.625 68.865 31.855 ;
        RECT 70.695 31.625 71.625 31.855 ;
        RECT 73.170 31.625 74.515 31.855 ;
        RECT 74.720 31.625 78.195 32.535 ;
        RECT 78.205 31.625 81.415 32.535 ;
        RECT 81.885 31.725 83.255 32.535 ;
      LAYER nwell ;
        RECT 5.330 28.505 83.450 31.335 ;
      LAYER pwell ;
        RECT 5.525 27.305 6.895 28.115 ;
        RECT 6.905 27.305 12.415 28.115 ;
        RECT 12.425 27.305 17.935 28.115 ;
        RECT 18.415 27.390 18.845 28.175 ;
        RECT 18.905 27.985 20.255 28.215 ;
        RECT 21.790 27.985 22.700 28.205 ;
        RECT 29.740 27.985 30.650 28.205 ;
        RECT 32.185 27.985 33.535 28.215 ;
        RECT 18.905 27.305 26.215 27.985 ;
        RECT 26.225 27.305 33.535 27.985 ;
        RECT 33.585 27.305 39.095 28.115 ;
        RECT 39.105 27.305 42.775 28.115 ;
        RECT 42.785 27.305 44.155 28.115 ;
        RECT 44.175 27.390 44.605 28.175 ;
        RECT 44.625 27.305 50.135 28.115 ;
        RECT 50.145 27.305 51.975 28.115 ;
        RECT 52.465 27.305 53.815 28.215 ;
        RECT 53.825 27.305 55.175 28.215 ;
        RECT 55.205 27.305 56.575 28.115 ;
        RECT 56.595 27.305 57.945 28.215 ;
        RECT 57.965 27.305 59.335 28.115 ;
        RECT 59.345 27.985 60.690 28.215 ;
        RECT 61.185 27.985 62.530 28.215 ;
        RECT 63.335 27.985 64.265 28.215 ;
        RECT 66.375 27.985 67.305 28.215 ;
        RECT 68.675 27.985 69.605 28.215 ;
        RECT 59.345 27.305 61.175 27.985 ;
        RECT 61.185 27.305 63.015 27.985 ;
        RECT 63.335 27.305 65.170 27.985 ;
        RECT 5.665 27.095 5.835 27.305 ;
        RECT 7.045 27.095 7.215 27.305 ;
        RECT 12.565 27.095 12.735 27.305 ;
        RECT 18.085 27.255 18.255 27.285 ;
        RECT 18.080 27.145 18.255 27.255 ;
        RECT 18.085 27.095 18.255 27.145 ;
        RECT 23.605 27.095 23.775 27.285 ;
        RECT 25.905 27.115 26.075 27.305 ;
        RECT 26.365 27.115 26.535 27.305 ;
        RECT 29.125 27.095 29.295 27.285 ;
        RECT 30.960 27.145 31.080 27.255 ;
        RECT 31.885 27.095 32.055 27.285 ;
        RECT 33.725 27.115 33.895 27.305 ;
        RECT 37.405 27.095 37.575 27.285 ;
        RECT 39.245 27.115 39.415 27.305 ;
        RECT 42.925 27.095 43.095 27.305 ;
        RECT 44.765 27.115 44.935 27.305 ;
        RECT 48.445 27.095 48.615 27.285 ;
        RECT 50.285 27.115 50.455 27.305 ;
        RECT 50.750 27.095 50.920 27.285 ;
        RECT 52.120 27.145 52.240 27.255 ;
        RECT 52.580 27.115 52.750 27.305 ;
        RECT 53.970 27.285 54.140 27.305 ;
        RECT 53.045 27.115 53.215 27.285 ;
        RECT 53.500 27.145 53.620 27.255 ;
        RECT 53.965 27.115 54.140 27.285 ;
        RECT 55.345 27.115 55.515 27.305 ;
        RECT 56.725 27.115 56.895 27.305 ;
        RECT 57.640 27.145 57.760 27.255 ;
        RECT 58.105 27.115 58.275 27.305 ;
        RECT 53.045 27.095 53.210 27.115 ;
        RECT 5.525 26.285 6.895 27.095 ;
        RECT 6.905 26.285 12.415 27.095 ;
        RECT 12.425 26.285 17.935 27.095 ;
        RECT 17.945 26.285 23.455 27.095 ;
        RECT 23.465 26.285 28.975 27.095 ;
        RECT 28.985 26.285 30.815 27.095 ;
        RECT 31.295 26.225 31.725 27.010 ;
        RECT 31.745 26.285 37.255 27.095 ;
        RECT 37.265 26.285 42.775 27.095 ;
        RECT 42.785 26.285 48.295 27.095 ;
        RECT 48.305 26.285 49.675 27.095 ;
        RECT 49.685 26.185 51.035 27.095 ;
        RECT 51.375 26.415 53.210 27.095 ;
        RECT 53.965 27.065 54.135 27.115 ;
        RECT 58.380 27.095 58.550 27.285 ;
        RECT 60.865 27.115 61.035 27.305 ;
        RECT 62.520 27.095 62.690 27.285 ;
        RECT 62.705 27.115 62.875 27.305 ;
        RECT 65.005 27.285 65.170 27.305 ;
        RECT 65.470 27.305 67.305 27.985 ;
        RECT 67.770 27.305 69.605 27.985 ;
        RECT 69.935 27.390 70.365 28.175 ;
        RECT 70.385 27.305 73.595 28.215 ;
        RECT 73.605 27.305 76.815 28.215 ;
        RECT 77.285 27.305 80.760 28.215 ;
        RECT 81.885 27.305 83.255 28.115 ;
        RECT 65.470 27.285 65.635 27.305 ;
        RECT 67.770 27.285 67.935 27.305 ;
        RECT 65.005 27.115 65.175 27.285 ;
        RECT 65.465 27.115 65.635 27.285 ;
        RECT 66.390 27.095 66.560 27.285 ;
        RECT 67.765 27.115 67.935 27.285 ;
        RECT 70.525 27.115 70.695 27.305 ;
        RECT 73.285 27.095 73.455 27.285 ;
        RECT 73.750 27.095 73.920 27.285 ;
        RECT 76.505 27.115 76.675 27.305 ;
        RECT 76.960 27.145 77.080 27.255 ;
        RECT 77.430 27.095 77.600 27.305 ;
        RECT 81.115 27.140 81.275 27.260 ;
        RECT 82.945 27.095 83.115 27.305 ;
        RECT 56.090 27.065 57.035 27.095 ;
        RECT 53.965 26.865 57.035 27.065 ;
        RECT 51.375 26.185 52.305 26.415 ;
        RECT 53.825 26.385 57.035 26.865 ;
        RECT 53.825 26.185 54.755 26.385 ;
        RECT 56.090 26.185 57.035 26.385 ;
        RECT 57.055 26.225 57.485 27.010 ;
        RECT 57.965 26.415 61.865 27.095 ;
        RECT 62.105 26.415 66.005 27.095 ;
        RECT 57.965 26.185 58.895 26.415 ;
        RECT 62.105 26.185 63.035 26.415 ;
        RECT 66.245 26.185 69.720 27.095 ;
        RECT 70.020 26.415 73.485 27.095 ;
        RECT 70.020 26.185 70.940 26.415 ;
        RECT 73.605 26.185 77.080 27.095 ;
        RECT 77.285 26.185 80.760 27.095 ;
        RECT 81.885 26.285 83.255 27.095 ;
      LAYER nwell ;
        RECT 5.330 23.065 83.450 25.895 ;
      LAYER pwell ;
        RECT 5.525 21.865 6.895 22.675 ;
        RECT 6.905 21.865 12.415 22.675 ;
        RECT 12.425 21.865 17.935 22.675 ;
        RECT 18.415 21.950 18.845 22.735 ;
        RECT 18.865 21.865 24.375 22.675 ;
        RECT 24.385 21.865 29.895 22.675 ;
        RECT 29.905 21.865 35.415 22.675 ;
        RECT 35.425 21.865 40.935 22.675 ;
        RECT 40.945 21.865 43.695 22.675 ;
        RECT 44.175 21.950 44.605 22.735 ;
        RECT 44.625 21.865 46.455 22.775 ;
        RECT 47.605 22.685 48.555 22.775 ;
        RECT 46.625 21.865 48.555 22.685 ;
        RECT 52.280 22.545 53.190 22.765 ;
        RECT 54.725 22.545 56.075 22.775 ;
        RECT 60.560 22.545 61.470 22.765 ;
        RECT 63.005 22.545 64.775 22.775 ;
        RECT 48.765 21.865 56.075 22.545 ;
        RECT 57.045 21.865 64.775 22.545 ;
        RECT 64.865 22.545 65.795 22.775 ;
        RECT 64.865 21.865 68.765 22.545 ;
        RECT 69.935 21.950 70.365 22.735 ;
        RECT 70.425 22.545 71.775 22.775 ;
        RECT 73.310 22.545 74.220 22.765 ;
        RECT 70.425 21.865 77.735 22.545 ;
        RECT 77.745 21.865 81.220 22.775 ;
        RECT 81.885 21.865 83.255 22.675 ;
        RECT 5.665 21.655 5.835 21.865 ;
        RECT 7.045 21.655 7.215 21.865 ;
        RECT 12.565 21.655 12.735 21.865 ;
        RECT 18.085 21.815 18.255 21.845 ;
        RECT 18.080 21.705 18.255 21.815 ;
        RECT 18.085 21.655 18.255 21.705 ;
        RECT 19.005 21.675 19.175 21.865 ;
        RECT 23.605 21.655 23.775 21.845 ;
        RECT 24.525 21.675 24.695 21.865 ;
        RECT 29.125 21.655 29.295 21.845 ;
        RECT 30.045 21.675 30.215 21.865 ;
        RECT 30.960 21.705 31.080 21.815 ;
        RECT 31.885 21.655 32.055 21.845 ;
        RECT 35.565 21.675 35.735 21.865 ;
        RECT 37.405 21.655 37.575 21.845 ;
        RECT 41.085 21.675 41.255 21.865 ;
        RECT 42.005 21.675 42.175 21.845 ;
        RECT 43.840 21.705 43.960 21.815 ;
        RECT 44.305 21.675 44.475 21.845 ;
        RECT 42.005 21.655 42.170 21.675 ;
        RECT 44.305 21.655 44.455 21.675 ;
        RECT 44.770 21.655 44.940 21.865 ;
        RECT 46.625 21.845 46.775 21.865 ;
        RECT 46.605 21.675 46.775 21.845 ;
        RECT 48.455 21.700 48.615 21.810 ;
        RECT 48.905 21.675 49.075 21.865 ;
        RECT 49.365 21.655 49.535 21.845 ;
        RECT 56.275 21.710 56.435 21.820 ;
        RECT 57.185 21.675 57.355 21.865 ;
        RECT 65.005 21.655 65.175 21.845 ;
        RECT 65.280 21.675 65.450 21.865 ;
        RECT 65.465 21.655 65.635 21.845 ;
        RECT 69.155 21.710 69.315 21.820 ;
        RECT 72.820 21.705 72.940 21.815 ;
        RECT 77.425 21.675 77.595 21.865 ;
        RECT 77.890 21.675 78.060 21.865 ;
        RECT 80.185 21.655 80.355 21.845 ;
        RECT 80.645 21.655 80.815 21.845 ;
        RECT 81.560 21.705 81.680 21.815 ;
        RECT 82.945 21.655 83.115 21.865 ;
        RECT 5.525 20.845 6.895 21.655 ;
        RECT 6.905 20.845 12.415 21.655 ;
        RECT 12.425 20.845 17.935 21.655 ;
        RECT 17.945 20.845 23.455 21.655 ;
        RECT 23.465 20.845 28.975 21.655 ;
        RECT 28.985 20.845 30.815 21.655 ;
        RECT 31.295 20.785 31.725 21.570 ;
        RECT 31.745 20.845 37.255 21.655 ;
        RECT 37.265 20.845 40.015 21.655 ;
        RECT 40.335 20.975 42.170 21.655 ;
        RECT 40.335 20.745 41.265 20.975 ;
        RECT 42.525 20.835 44.455 21.655 ;
        RECT 42.525 20.745 43.475 20.835 ;
        RECT 44.625 20.745 48.295 21.655 ;
        RECT 49.225 20.975 56.955 21.655 ;
        RECT 52.740 20.755 53.650 20.975 ;
        RECT 55.185 20.745 56.955 20.975 ;
        RECT 57.055 20.785 57.485 21.570 ;
        RECT 57.585 20.975 65.315 21.655 ;
        RECT 65.325 20.975 72.635 21.655 ;
        RECT 57.585 20.745 59.355 20.975 ;
        RECT 60.890 20.755 61.800 20.975 ;
        RECT 68.840 20.755 69.750 20.975 ;
        RECT 71.285 20.745 72.635 20.975 ;
        RECT 73.185 20.975 80.495 21.655 ;
        RECT 73.185 20.745 74.535 20.975 ;
        RECT 76.070 20.755 76.980 20.975 ;
        RECT 80.505 20.845 81.875 21.655 ;
        RECT 81.885 20.845 83.255 21.655 ;
      LAYER nwell ;
        RECT 5.330 17.625 83.450 20.455 ;
      LAYER pwell ;
        RECT 5.525 16.425 6.895 17.235 ;
        RECT 6.905 16.425 12.415 17.235 ;
        RECT 12.425 16.425 17.935 17.235 ;
        RECT 18.415 16.510 18.845 17.295 ;
        RECT 18.865 16.425 24.375 17.235 ;
        RECT 24.385 16.425 29.895 17.235 ;
        RECT 29.905 16.425 35.415 17.235 ;
        RECT 35.425 16.425 40.935 17.235 ;
        RECT 40.945 16.425 42.775 17.235 ;
        RECT 42.785 16.425 44.155 17.205 ;
        RECT 44.175 16.510 44.605 17.295 ;
        RECT 48.200 17.105 49.120 17.335 ;
        RECT 52.740 17.105 53.650 17.325 ;
        RECT 55.185 17.105 56.535 17.335 ;
        RECT 57.955 17.105 58.875 17.335 ;
        RECT 63.320 17.105 64.230 17.325 ;
        RECT 65.765 17.105 67.115 17.335 ;
        RECT 68.215 17.105 69.145 17.335 ;
        RECT 45.655 16.425 49.120 17.105 ;
        RECT 49.225 16.425 56.535 17.105 ;
        RECT 56.585 16.425 58.875 17.105 ;
        RECT 59.805 16.425 67.115 17.105 ;
        RECT 67.310 16.425 69.145 17.105 ;
        RECT 69.935 16.510 70.365 17.295 ;
        RECT 70.385 16.425 73.860 17.335 ;
        RECT 78.040 17.105 78.950 17.325 ;
        RECT 80.485 17.105 81.835 17.335 ;
        RECT 74.525 16.425 81.835 17.105 ;
        RECT 81.885 16.425 83.255 17.235 ;
        RECT 5.665 16.215 5.835 16.425 ;
        RECT 7.045 16.215 7.215 16.425 ;
        RECT 12.565 16.215 12.735 16.425 ;
        RECT 18.085 16.375 18.255 16.405 ;
        RECT 18.080 16.265 18.255 16.375 ;
        RECT 18.085 16.215 18.255 16.265 ;
        RECT 19.005 16.235 19.175 16.425 ;
        RECT 23.605 16.215 23.775 16.405 ;
        RECT 24.525 16.235 24.695 16.425 ;
        RECT 29.125 16.215 29.295 16.405 ;
        RECT 30.045 16.235 30.215 16.425 ;
        RECT 30.960 16.265 31.080 16.375 ;
        RECT 31.885 16.215 32.055 16.405 ;
        RECT 35.565 16.235 35.735 16.425 ;
        RECT 37.405 16.215 37.575 16.405 ;
        RECT 40.165 16.215 40.335 16.405 ;
        RECT 41.085 16.235 41.255 16.425 ;
        RECT 43.845 16.235 44.015 16.425 ;
        RECT 44.775 16.270 44.935 16.380 ;
        RECT 45.685 16.235 45.855 16.425 ;
        RECT 47.525 16.215 47.695 16.405 ;
        RECT 49.365 16.235 49.535 16.425 ;
        RECT 51.215 16.260 51.375 16.370 ;
        RECT 52.400 16.215 52.570 16.405 ;
        RECT 56.275 16.260 56.435 16.370 ;
        RECT 56.725 16.235 56.895 16.425 ;
        RECT 57.645 16.215 57.815 16.405 ;
        RECT 59.035 16.270 59.195 16.380 ;
        RECT 59.945 16.235 60.115 16.425 ;
        RECT 67.310 16.405 67.475 16.425 ;
        RECT 63.160 16.265 63.280 16.375 ;
        RECT 63.625 16.215 63.795 16.405 ;
        RECT 67.305 16.235 67.475 16.405 ;
        RECT 69.600 16.265 69.720 16.375 ;
        RECT 70.530 16.235 70.700 16.425 ;
        RECT 70.985 16.215 71.155 16.405 ;
        RECT 72.365 16.235 72.535 16.405 ;
        RECT 74.200 16.265 74.320 16.375 ;
        RECT 72.370 16.215 72.535 16.235 ;
        RECT 74.665 16.215 74.835 16.425 ;
        RECT 82.945 16.215 83.115 16.425 ;
        RECT 5.525 15.405 6.895 16.215 ;
        RECT 6.905 15.405 12.415 16.215 ;
        RECT 12.425 15.405 17.935 16.215 ;
        RECT 17.945 15.405 23.455 16.215 ;
        RECT 23.465 15.405 28.975 16.215 ;
        RECT 28.985 15.405 30.815 16.215 ;
        RECT 31.295 15.345 31.725 16.130 ;
        RECT 31.745 15.405 37.255 16.215 ;
        RECT 37.265 15.405 40.015 16.215 ;
        RECT 40.025 15.535 47.335 16.215 ;
        RECT 43.540 15.315 44.450 15.535 ;
        RECT 45.985 15.305 47.335 15.535 ;
        RECT 47.385 15.405 51.055 16.215 ;
        RECT 51.985 15.535 55.885 16.215 ;
        RECT 51.985 15.305 52.915 15.535 ;
        RECT 57.055 15.345 57.485 16.130 ;
        RECT 57.505 15.405 63.015 16.215 ;
        RECT 63.485 15.535 70.795 16.215 ;
        RECT 67.000 15.315 67.910 15.535 ;
        RECT 69.445 15.305 70.795 15.535 ;
        RECT 70.845 15.435 72.215 16.215 ;
        RECT 72.370 15.535 74.205 16.215 ;
        RECT 74.525 15.535 81.835 16.215 ;
        RECT 73.275 15.305 74.205 15.535 ;
        RECT 78.040 15.315 78.950 15.535 ;
        RECT 80.485 15.305 81.835 15.535 ;
        RECT 81.885 15.405 83.255 16.215 ;
      LAYER nwell ;
        RECT 5.330 12.185 83.450 15.015 ;
      LAYER pwell ;
        RECT 5.525 10.985 6.895 11.795 ;
        RECT 6.905 10.985 12.415 11.795 ;
        RECT 12.425 10.985 17.935 11.795 ;
        RECT 18.415 11.070 18.845 11.855 ;
        RECT 18.865 10.985 24.375 11.795 ;
        RECT 24.385 10.985 29.895 11.795 ;
        RECT 29.905 10.985 31.275 11.795 ;
        RECT 31.295 11.070 31.725 11.855 ;
        RECT 31.745 10.985 35.415 11.795 ;
        RECT 36.545 11.665 40.475 11.895 ;
        RECT 42.325 11.665 43.670 11.895 ;
        RECT 36.060 10.985 40.475 11.665 ;
        RECT 40.485 10.985 42.315 11.665 ;
        RECT 42.325 10.985 44.155 11.665 ;
        RECT 44.175 11.070 44.605 11.855 ;
        RECT 45.545 11.665 46.890 11.895 ;
        RECT 45.545 10.985 47.375 11.665 ;
        RECT 47.385 10.985 48.755 11.795 ;
        RECT 48.765 10.985 50.595 11.665 ;
        RECT 50.605 10.985 56.115 11.795 ;
        RECT 57.055 11.070 57.485 11.855 ;
        RECT 57.505 10.985 63.015 11.795 ;
        RECT 63.025 10.985 64.855 11.795 ;
        RECT 64.865 11.665 66.210 11.895 ;
        RECT 64.865 10.985 66.695 11.665 ;
        RECT 66.705 10.985 68.075 11.795 ;
        RECT 68.085 11.665 69.430 11.895 ;
        RECT 68.085 10.985 69.915 11.665 ;
        RECT 69.935 11.070 70.365 11.855 ;
        RECT 71.305 11.665 72.650 11.895 ;
        RECT 73.630 11.665 74.975 11.895 ;
        RECT 75.470 11.665 76.815 11.895 ;
        RECT 77.875 11.665 78.805 11.895 ;
        RECT 80.530 11.665 81.875 11.895 ;
        RECT 71.305 10.985 73.135 11.665 ;
        RECT 73.145 10.985 74.975 11.665 ;
        RECT 74.985 10.985 76.815 11.665 ;
        RECT 76.970 10.985 78.805 11.665 ;
        RECT 80.045 10.985 81.875 11.665 ;
        RECT 81.885 10.985 83.255 11.795 ;
        RECT 5.665 10.795 5.835 10.985 ;
        RECT 7.045 10.795 7.215 10.985 ;
        RECT 12.565 10.795 12.735 10.985 ;
        RECT 18.080 10.825 18.200 10.935 ;
        RECT 19.005 10.795 19.175 10.985 ;
        RECT 24.525 10.795 24.695 10.985 ;
        RECT 30.045 10.795 30.215 10.985 ;
        RECT 31.885 10.795 32.055 10.985 ;
        RECT 36.060 10.965 36.170 10.985 ;
        RECT 35.560 10.825 35.680 10.935 ;
        RECT 36.000 10.795 36.170 10.965 ;
        RECT 40.625 10.795 40.795 10.985 ;
        RECT 43.845 10.795 44.015 10.985 ;
        RECT 44.775 10.830 44.935 10.940 ;
        RECT 47.065 10.795 47.235 10.985 ;
        RECT 47.525 10.795 47.695 10.985 ;
        RECT 48.905 10.795 49.075 10.985 ;
        RECT 50.745 10.795 50.915 10.985 ;
        RECT 56.275 10.830 56.435 10.940 ;
        RECT 57.645 10.795 57.815 10.985 ;
        RECT 63.165 10.795 63.335 10.985 ;
        RECT 66.385 10.795 66.555 10.985 ;
        RECT 66.845 10.795 67.015 10.985 ;
        RECT 69.605 10.795 69.775 10.985 ;
        RECT 70.535 10.830 70.695 10.940 ;
        RECT 72.825 10.795 72.995 10.985 ;
        RECT 73.285 10.795 73.455 10.985 ;
        RECT 75.125 10.795 75.295 10.985 ;
        RECT 76.970 10.965 77.135 10.985 ;
        RECT 76.965 10.795 77.135 10.965 ;
        RECT 79.275 10.830 79.435 10.940 ;
        RECT 80.185 10.795 80.355 10.985 ;
        RECT 82.945 10.795 83.115 10.985 ;
      LAYER li1 ;
        RECT 5.520 165.835 83.260 166.005 ;
        RECT 5.605 164.745 6.815 165.835 ;
        RECT 6.985 165.400 12.330 165.835 ;
        RECT 12.505 165.400 17.850 165.835 ;
        RECT 5.605 164.035 6.125 164.575 ;
        RECT 6.295 164.205 6.815 164.745 ;
        RECT 5.605 163.285 6.815 164.035 ;
        RECT 8.570 163.830 8.910 164.660 ;
        RECT 10.390 164.150 10.740 165.400 ;
        RECT 14.090 163.830 14.430 164.660 ;
        RECT 15.910 164.150 16.260 165.400 ;
        RECT 18.485 164.670 18.775 165.835 ;
        RECT 18.945 165.400 24.290 165.835 ;
        RECT 24.465 165.400 29.810 165.835 ;
        RECT 6.985 163.285 12.330 163.830 ;
        RECT 12.505 163.285 17.850 163.830 ;
        RECT 18.485 163.285 18.775 164.010 ;
        RECT 20.530 163.830 20.870 164.660 ;
        RECT 22.350 164.150 22.700 165.400 ;
        RECT 26.050 163.830 26.390 164.660 ;
        RECT 27.870 164.150 28.220 165.400 ;
        RECT 29.985 164.745 31.195 165.835 ;
        RECT 29.985 164.035 30.505 164.575 ;
        RECT 30.675 164.205 31.195 164.745 ;
        RECT 31.365 164.670 31.655 165.835 ;
        RECT 31.825 165.400 37.170 165.835 ;
        RECT 18.945 163.285 24.290 163.830 ;
        RECT 24.465 163.285 29.810 163.830 ;
        RECT 29.985 163.285 31.195 164.035 ;
        RECT 31.365 163.285 31.655 164.010 ;
        RECT 33.410 163.830 33.750 164.660 ;
        RECT 35.230 164.150 35.580 165.400 ;
        RECT 37.345 164.745 39.015 165.835 ;
        RECT 37.345 164.055 38.095 164.575 ;
        RECT 38.265 164.225 39.015 164.745 ;
        RECT 39.190 164.685 39.450 165.835 ;
        RECT 39.625 164.760 39.880 165.665 ;
        RECT 40.050 165.075 40.380 165.835 ;
        RECT 40.595 164.905 40.765 165.665 ;
        RECT 31.825 163.285 37.170 163.830 ;
        RECT 37.345 163.285 39.015 164.055 ;
        RECT 39.190 163.285 39.450 164.125 ;
        RECT 39.625 164.030 39.795 164.760 ;
        RECT 40.050 164.735 40.765 164.905 ;
        RECT 41.025 164.745 43.615 165.835 ;
        RECT 40.050 164.525 40.220 164.735 ;
        RECT 39.965 164.195 40.220 164.525 ;
        RECT 39.625 163.455 39.880 164.030 ;
        RECT 40.050 164.005 40.220 164.195 ;
        RECT 40.500 164.185 40.855 164.555 ;
        RECT 41.025 164.055 42.235 164.575 ;
        RECT 42.405 164.225 43.615 164.745 ;
        RECT 44.245 164.670 44.535 165.835 ;
        RECT 44.705 165.400 50.050 165.835 ;
        RECT 40.050 163.835 40.765 164.005 ;
        RECT 40.050 163.285 40.380 163.665 ;
        RECT 40.595 163.455 40.765 163.835 ;
        RECT 41.025 163.285 43.615 164.055 ;
        RECT 44.245 163.285 44.535 164.010 ;
        RECT 46.290 163.830 46.630 164.660 ;
        RECT 48.110 164.150 48.460 165.400 ;
        RECT 50.225 164.745 51.435 165.835 ;
        RECT 50.225 164.035 50.745 164.575 ;
        RECT 50.915 164.205 51.435 164.745 ;
        RECT 51.610 164.685 51.870 165.835 ;
        RECT 52.045 164.760 52.300 165.665 ;
        RECT 52.470 165.075 52.800 165.835 ;
        RECT 53.015 164.905 53.185 165.665 ;
        RECT 44.705 163.285 50.050 163.830 ;
        RECT 50.225 163.285 51.435 164.035 ;
        RECT 51.610 163.285 51.870 164.125 ;
        RECT 52.045 164.030 52.215 164.760 ;
        RECT 52.470 164.735 53.185 164.905 ;
        RECT 52.470 164.525 52.640 164.735 ;
        RECT 53.450 164.685 53.710 165.835 ;
        RECT 53.885 164.760 54.140 165.665 ;
        RECT 54.310 165.075 54.640 165.835 ;
        RECT 54.855 164.905 55.025 165.665 ;
        RECT 52.385 164.195 52.640 164.525 ;
        RECT 52.045 163.455 52.300 164.030 ;
        RECT 52.470 164.005 52.640 164.195 ;
        RECT 52.920 164.185 53.275 164.555 ;
        RECT 52.470 163.835 53.185 164.005 ;
        RECT 52.470 163.285 52.800 163.665 ;
        RECT 53.015 163.455 53.185 163.835 ;
        RECT 53.450 163.285 53.710 164.125 ;
        RECT 53.885 164.030 54.055 164.760 ;
        RECT 54.310 164.735 55.025 164.905 ;
        RECT 54.310 164.525 54.480 164.735 ;
        RECT 55.290 164.685 55.550 165.835 ;
        RECT 55.725 164.760 55.980 165.665 ;
        RECT 56.150 165.075 56.480 165.835 ;
        RECT 56.695 164.905 56.865 165.665 ;
        RECT 54.225 164.195 54.480 164.525 ;
        RECT 53.885 163.455 54.140 164.030 ;
        RECT 54.310 164.005 54.480 164.195 ;
        RECT 54.760 164.185 55.115 164.555 ;
        RECT 54.310 163.835 55.025 164.005 ;
        RECT 54.310 163.285 54.640 163.665 ;
        RECT 54.855 163.455 55.025 163.835 ;
        RECT 55.290 163.285 55.550 164.125 ;
        RECT 55.725 164.030 55.895 164.760 ;
        RECT 56.150 164.735 56.865 164.905 ;
        RECT 56.150 164.525 56.320 164.735 ;
        RECT 57.125 164.670 57.415 165.835 ;
        RECT 57.675 164.905 57.845 165.665 ;
        RECT 58.060 165.075 58.390 165.835 ;
        RECT 57.675 164.735 58.390 164.905 ;
        RECT 58.560 164.760 58.815 165.665 ;
        RECT 56.065 164.195 56.320 164.525 ;
        RECT 55.725 163.455 55.980 164.030 ;
        RECT 56.150 164.005 56.320 164.195 ;
        RECT 56.600 164.185 56.955 164.555 ;
        RECT 57.585 164.185 57.940 164.555 ;
        RECT 58.220 164.525 58.390 164.735 ;
        RECT 58.220 164.195 58.475 164.525 ;
        RECT 56.150 163.835 56.865 164.005 ;
        RECT 56.150 163.285 56.480 163.665 ;
        RECT 56.695 163.455 56.865 163.835 ;
        RECT 57.125 163.285 57.415 164.010 ;
        RECT 58.220 164.005 58.390 164.195 ;
        RECT 58.645 164.030 58.815 164.760 ;
        RECT 58.990 164.685 59.250 165.835 ;
        RECT 59.430 164.685 59.690 165.835 ;
        RECT 59.865 164.760 60.120 165.665 ;
        RECT 60.290 165.075 60.620 165.835 ;
        RECT 60.835 164.905 61.005 165.665 ;
        RECT 57.675 163.835 58.390 164.005 ;
        RECT 57.675 163.455 57.845 163.835 ;
        RECT 58.060 163.285 58.390 163.665 ;
        RECT 58.560 163.455 58.815 164.030 ;
        RECT 58.990 163.285 59.250 164.125 ;
        RECT 59.430 163.285 59.690 164.125 ;
        RECT 59.865 164.030 60.035 164.760 ;
        RECT 60.290 164.735 61.005 164.905 ;
        RECT 61.300 165.045 61.835 165.665 ;
        RECT 60.290 164.525 60.460 164.735 ;
        RECT 60.205 164.195 60.460 164.525 ;
        RECT 59.865 163.455 60.120 164.030 ;
        RECT 60.290 164.005 60.460 164.195 ;
        RECT 60.740 164.185 61.095 164.555 ;
        RECT 61.300 164.025 61.615 165.045 ;
        RECT 62.005 165.035 62.335 165.835 ;
        RECT 63.600 165.045 64.135 165.665 ;
        RECT 62.820 164.865 63.210 165.040 ;
        RECT 61.785 164.695 63.210 164.865 ;
        RECT 61.785 164.195 61.955 164.695 ;
        RECT 60.290 163.835 61.005 164.005 ;
        RECT 60.290 163.285 60.620 163.665 ;
        RECT 60.835 163.455 61.005 163.835 ;
        RECT 61.300 163.455 61.915 164.025 ;
        RECT 62.205 163.965 62.470 164.525 ;
        RECT 62.640 163.795 62.810 164.695 ;
        RECT 62.980 163.965 63.335 164.525 ;
        RECT 63.600 164.025 63.915 165.045 ;
        RECT 64.305 165.035 64.635 165.835 ;
        RECT 65.900 165.045 66.435 165.665 ;
        RECT 65.120 164.865 65.510 165.040 ;
        RECT 64.085 164.695 65.510 164.865 ;
        RECT 64.085 164.195 64.255 164.695 ;
        RECT 62.085 163.285 62.300 163.795 ;
        RECT 62.530 163.465 62.810 163.795 ;
        RECT 62.990 163.285 63.230 163.795 ;
        RECT 63.600 163.455 64.215 164.025 ;
        RECT 64.505 163.965 64.770 164.525 ;
        RECT 64.940 163.795 65.110 164.695 ;
        RECT 65.280 163.965 65.635 164.525 ;
        RECT 65.900 164.025 66.215 165.045 ;
        RECT 66.605 165.035 66.935 165.835 ;
        RECT 67.420 164.865 67.810 165.040 ;
        RECT 66.385 164.695 67.810 164.865 ;
        RECT 66.385 164.195 66.555 164.695 ;
        RECT 64.385 163.285 64.600 163.795 ;
        RECT 64.830 163.465 65.110 163.795 ;
        RECT 65.290 163.285 65.530 163.795 ;
        RECT 65.900 163.455 66.515 164.025 ;
        RECT 66.805 163.965 67.070 164.525 ;
        RECT 67.240 163.795 67.410 164.695 ;
        RECT 68.170 164.685 68.430 165.835 ;
        RECT 68.605 164.760 68.860 165.665 ;
        RECT 69.030 165.075 69.360 165.835 ;
        RECT 69.575 164.905 69.745 165.665 ;
        RECT 67.580 163.965 67.935 164.525 ;
        RECT 66.685 163.285 66.900 163.795 ;
        RECT 67.130 163.465 67.410 163.795 ;
        RECT 67.590 163.285 67.830 163.795 ;
        RECT 68.170 163.285 68.430 164.125 ;
        RECT 68.605 164.030 68.775 164.760 ;
        RECT 69.030 164.735 69.745 164.905 ;
        RECT 69.030 164.525 69.200 164.735 ;
        RECT 70.005 164.670 70.295 165.835 ;
        RECT 70.650 164.865 71.040 165.040 ;
        RECT 71.525 165.035 71.855 165.835 ;
        RECT 72.025 165.045 72.560 165.665 ;
        RECT 70.650 164.695 72.075 164.865 ;
        RECT 68.945 164.195 69.200 164.525 ;
        RECT 68.605 163.455 68.860 164.030 ;
        RECT 69.030 164.005 69.200 164.195 ;
        RECT 69.480 164.185 69.835 164.555 ;
        RECT 69.030 163.835 69.745 164.005 ;
        RECT 69.030 163.285 69.360 163.665 ;
        RECT 69.575 163.455 69.745 163.835 ;
        RECT 70.005 163.285 70.295 164.010 ;
        RECT 70.525 163.965 70.880 164.525 ;
        RECT 71.050 163.795 71.220 164.695 ;
        RECT 71.390 163.965 71.655 164.525 ;
        RECT 71.905 164.195 72.075 164.695 ;
        RECT 72.245 164.025 72.560 165.045 ;
        RECT 72.950 164.865 73.340 165.040 ;
        RECT 73.825 165.035 74.155 165.835 ;
        RECT 74.325 165.045 74.860 165.665 ;
        RECT 72.950 164.695 74.375 164.865 ;
        RECT 70.630 163.285 70.870 163.795 ;
        RECT 71.050 163.465 71.330 163.795 ;
        RECT 71.560 163.285 71.775 163.795 ;
        RECT 71.945 163.455 72.560 164.025 ;
        RECT 72.825 163.965 73.180 164.525 ;
        RECT 73.350 163.795 73.520 164.695 ;
        RECT 73.690 163.965 73.955 164.525 ;
        RECT 74.205 164.195 74.375 164.695 ;
        RECT 74.545 164.025 74.860 165.045 ;
        RECT 75.250 164.865 75.640 165.040 ;
        RECT 76.125 165.035 76.455 165.835 ;
        RECT 76.625 165.045 77.160 165.665 ;
        RECT 75.250 164.695 76.675 164.865 ;
        RECT 72.930 163.285 73.170 163.795 ;
        RECT 73.350 163.465 73.630 163.795 ;
        RECT 73.860 163.285 74.075 163.795 ;
        RECT 74.245 163.455 74.860 164.025 ;
        RECT 75.125 163.965 75.480 164.525 ;
        RECT 75.650 163.795 75.820 164.695 ;
        RECT 75.990 163.965 76.255 164.525 ;
        RECT 76.505 164.195 76.675 164.695 ;
        RECT 76.845 164.025 77.160 165.045 ;
        RECT 77.830 165.445 78.165 165.665 ;
        RECT 79.170 165.455 79.525 165.835 ;
        RECT 77.830 164.825 78.085 165.445 ;
        RECT 78.335 165.285 78.565 165.325 ;
        RECT 79.695 165.285 79.945 165.665 ;
        RECT 78.335 165.085 79.945 165.285 ;
        RECT 78.335 164.995 78.520 165.085 ;
        RECT 79.110 165.075 79.945 165.085 ;
        RECT 80.195 165.055 80.445 165.835 ;
        RECT 80.615 164.985 80.875 165.665 ;
        RECT 78.675 164.885 79.005 164.915 ;
        RECT 78.675 164.825 80.475 164.885 ;
        RECT 77.830 164.715 80.535 164.825 ;
        RECT 77.830 164.655 79.005 164.715 ;
        RECT 80.335 164.680 80.535 164.715 ;
        RECT 77.825 164.275 78.315 164.475 ;
        RECT 78.505 164.275 78.980 164.485 ;
        RECT 75.230 163.285 75.470 163.795 ;
        RECT 75.650 163.465 75.930 163.795 ;
        RECT 76.160 163.285 76.375 163.795 ;
        RECT 76.545 163.455 77.160 164.025 ;
        RECT 77.830 163.285 78.285 164.050 ;
        RECT 78.760 163.875 78.980 164.275 ;
        RECT 79.225 164.275 79.555 164.485 ;
        RECT 79.225 163.875 79.435 164.275 ;
        RECT 79.725 164.240 80.135 164.545 ;
        RECT 80.365 164.105 80.535 164.680 ;
        RECT 80.265 163.985 80.535 164.105 ;
        RECT 79.690 163.940 80.535 163.985 ;
        RECT 79.690 163.815 80.445 163.940 ;
        RECT 79.690 163.665 79.860 163.815 ;
        RECT 80.705 163.795 80.875 164.985 ;
        RECT 81.965 164.745 83.175 165.835 ;
        RECT 81.965 164.205 82.485 164.745 ;
        RECT 82.655 164.035 83.175 164.575 ;
        RECT 80.645 163.785 80.875 163.795 ;
        RECT 78.560 163.455 79.860 163.665 ;
        RECT 80.115 163.285 80.445 163.645 ;
        RECT 80.615 163.455 80.875 163.785 ;
        RECT 81.965 163.285 83.175 164.035 ;
        RECT 5.520 163.115 83.260 163.285 ;
        RECT 5.605 162.365 6.815 163.115 ;
        RECT 6.985 162.570 12.330 163.115 ;
        RECT 12.505 162.570 17.850 163.115 ;
        RECT 18.025 162.570 23.370 163.115 ;
        RECT 23.545 162.570 28.890 163.115 ;
        RECT 5.605 161.825 6.125 162.365 ;
        RECT 6.295 161.655 6.815 162.195 ;
        RECT 8.570 161.740 8.910 162.570 ;
        RECT 5.605 160.565 6.815 161.655 ;
        RECT 10.390 161.000 10.740 162.250 ;
        RECT 14.090 161.740 14.430 162.570 ;
        RECT 15.910 161.000 16.260 162.250 ;
        RECT 19.610 161.740 19.950 162.570 ;
        RECT 21.430 161.000 21.780 162.250 ;
        RECT 25.130 161.740 25.470 162.570 ;
        RECT 29.065 162.345 30.735 163.115 ;
        RECT 31.365 162.390 31.655 163.115 ;
        RECT 31.825 162.345 33.495 163.115 ;
        RECT 26.950 161.000 27.300 162.250 ;
        RECT 29.065 161.825 29.815 162.345 ;
        RECT 29.985 161.655 30.735 162.175 ;
        RECT 31.825 161.825 32.575 162.345 ;
        RECT 6.985 160.565 12.330 161.000 ;
        RECT 12.505 160.565 17.850 161.000 ;
        RECT 18.025 160.565 23.370 161.000 ;
        RECT 23.545 160.565 28.890 161.000 ;
        RECT 29.065 160.565 30.735 161.655 ;
        RECT 31.365 160.565 31.655 161.730 ;
        RECT 32.745 161.655 33.495 162.175 ;
        RECT 31.825 160.565 33.495 161.655 ;
        RECT 33.665 162.130 33.935 162.945 ;
        RECT 34.105 162.375 34.775 163.115 ;
        RECT 34.945 162.545 35.240 162.890 ;
        RECT 35.420 162.715 35.795 163.115 ;
        RECT 36.010 162.545 36.340 162.890 ;
        RECT 34.945 162.375 36.340 162.545 ;
        RECT 36.590 162.375 37.175 162.945 ;
        RECT 37.345 162.570 42.690 163.115 ;
        RECT 33.665 160.735 34.015 162.130 ;
        RECT 34.185 161.705 34.355 162.205 ;
        RECT 34.525 161.875 34.860 162.205 ;
        RECT 35.030 161.875 35.370 162.205 ;
        RECT 34.185 161.535 34.930 161.705 ;
        RECT 34.185 160.565 34.590 161.365 ;
        RECT 34.760 160.905 34.930 161.535 ;
        RECT 35.100 161.130 35.370 161.875 ;
        RECT 35.560 161.875 35.850 162.205 ;
        RECT 36.020 161.875 36.420 162.205 ;
        RECT 35.560 161.130 35.795 161.875 ;
        RECT 36.590 161.705 36.760 162.375 ;
        RECT 36.930 161.875 37.175 162.205 ;
        RECT 38.930 161.740 39.270 162.570 ;
        RECT 42.865 162.345 44.535 163.115 ;
        RECT 35.965 161.535 37.175 161.705 ;
        RECT 35.965 160.905 36.295 161.535 ;
        RECT 34.760 160.735 36.295 160.905 ;
        RECT 36.480 160.565 36.715 161.365 ;
        RECT 36.885 160.735 37.175 161.535 ;
        RECT 40.750 161.000 41.100 162.250 ;
        RECT 42.865 161.825 43.615 162.345 ;
        RECT 44.705 162.315 45.015 163.115 ;
        RECT 45.220 162.315 45.915 162.945 ;
        RECT 46.085 162.570 51.430 163.115 ;
        RECT 43.785 161.655 44.535 162.175 ;
        RECT 44.715 161.875 45.050 162.145 ;
        RECT 45.220 161.715 45.390 162.315 ;
        RECT 45.560 161.875 45.895 162.125 ;
        RECT 47.670 161.740 48.010 162.570 ;
        RECT 51.610 162.275 51.870 163.115 ;
        RECT 52.045 162.370 52.300 162.945 ;
        RECT 52.470 162.735 52.800 163.115 ;
        RECT 53.015 162.565 53.185 162.945 ;
        RECT 52.470 162.395 53.185 162.565 ;
        RECT 53.560 162.485 53.845 162.945 ;
        RECT 54.015 162.655 54.285 163.115 ;
        RECT 37.345 160.565 42.690 161.000 ;
        RECT 42.865 160.565 44.535 161.655 ;
        RECT 44.705 160.565 44.985 161.705 ;
        RECT 45.155 160.735 45.485 161.715 ;
        RECT 45.655 160.565 45.915 161.705 ;
        RECT 49.490 161.000 49.840 162.250 ;
        RECT 46.085 160.565 51.430 161.000 ;
        RECT 51.610 160.565 51.870 161.715 ;
        RECT 52.045 161.640 52.215 162.370 ;
        RECT 52.470 162.205 52.640 162.395 ;
        RECT 53.560 162.315 54.515 162.485 ;
        RECT 52.385 161.875 52.640 162.205 ;
        RECT 52.470 161.665 52.640 161.875 ;
        RECT 52.920 161.845 53.275 162.215 ;
        RECT 52.045 160.735 52.300 161.640 ;
        RECT 52.470 161.495 53.185 161.665 ;
        RECT 53.445 161.585 54.135 162.145 ;
        RECT 52.470 160.565 52.800 161.325 ;
        RECT 53.015 160.735 53.185 161.495 ;
        RECT 54.305 161.415 54.515 162.315 ;
        RECT 53.560 161.195 54.515 161.415 ;
        RECT 54.685 162.145 55.085 162.945 ;
        RECT 55.275 162.485 55.555 162.945 ;
        RECT 56.075 162.655 56.400 163.115 ;
        RECT 55.275 162.315 56.400 162.485 ;
        RECT 56.570 162.375 56.955 162.945 ;
        RECT 57.125 162.390 57.415 163.115 ;
        RECT 55.950 162.205 56.400 162.315 ;
        RECT 54.685 161.585 55.780 162.145 ;
        RECT 55.950 161.875 56.505 162.205 ;
        RECT 53.560 160.735 53.845 161.195 ;
        RECT 54.015 160.565 54.285 161.025 ;
        RECT 54.685 160.735 55.085 161.585 ;
        RECT 55.950 161.415 56.400 161.875 ;
        RECT 56.675 161.705 56.955 162.375 ;
        RECT 57.585 162.375 57.970 162.945 ;
        RECT 58.140 162.655 58.465 163.115 ;
        RECT 58.985 162.485 59.265 162.945 ;
        RECT 55.275 161.195 56.400 161.415 ;
        RECT 55.275 160.735 55.555 161.195 ;
        RECT 56.075 160.565 56.400 161.025 ;
        RECT 56.570 160.735 56.955 161.705 ;
        RECT 57.125 160.565 57.415 161.730 ;
        RECT 57.585 161.705 57.865 162.375 ;
        RECT 58.140 162.315 59.265 162.485 ;
        RECT 58.140 162.205 58.590 162.315 ;
        RECT 58.035 161.875 58.590 162.205 ;
        RECT 59.455 162.145 59.855 162.945 ;
        RECT 60.255 162.655 60.525 163.115 ;
        RECT 60.695 162.485 60.980 162.945 ;
        RECT 57.585 160.735 57.970 161.705 ;
        RECT 58.140 161.415 58.590 161.875 ;
        RECT 58.760 161.585 59.855 162.145 ;
        RECT 58.140 161.195 59.265 161.415 ;
        RECT 58.140 160.565 58.465 161.025 ;
        RECT 58.985 160.735 59.265 161.195 ;
        RECT 59.455 160.735 59.855 161.585 ;
        RECT 60.025 162.315 60.980 162.485 ;
        RECT 62.235 162.460 62.565 162.895 ;
        RECT 62.735 162.505 62.905 163.115 ;
        RECT 62.185 162.375 62.565 162.460 ;
        RECT 63.075 162.375 63.405 162.900 ;
        RECT 63.665 162.585 63.875 163.115 ;
        RECT 64.150 162.665 64.935 162.835 ;
        RECT 65.105 162.665 65.510 162.835 ;
        RECT 62.185 162.335 62.410 162.375 ;
        RECT 60.025 161.415 60.235 162.315 ;
        RECT 60.405 161.585 61.095 162.145 ;
        RECT 62.185 161.755 62.355 162.335 ;
        RECT 63.075 162.205 63.275 162.375 ;
        RECT 64.150 162.205 64.320 162.665 ;
        RECT 62.525 161.875 63.275 162.205 ;
        RECT 63.445 161.875 64.320 162.205 ;
        RECT 62.185 161.705 62.400 161.755 ;
        RECT 62.185 161.625 62.575 161.705 ;
        RECT 60.025 161.195 60.980 161.415 ;
        RECT 60.255 160.565 60.525 161.025 ;
        RECT 60.695 160.735 60.980 161.195 ;
        RECT 62.245 160.780 62.575 161.625 ;
        RECT 63.085 161.670 63.275 161.875 ;
        RECT 62.745 160.565 62.915 161.575 ;
        RECT 63.085 161.295 63.980 161.670 ;
        RECT 63.085 160.735 63.425 161.295 ;
        RECT 63.655 160.565 63.970 161.065 ;
        RECT 64.150 161.035 64.320 161.875 ;
        RECT 64.490 162.165 64.955 162.495 ;
        RECT 65.340 162.435 65.510 162.665 ;
        RECT 65.690 162.615 66.060 163.115 ;
        RECT 66.380 162.665 67.055 162.835 ;
        RECT 67.250 162.665 67.585 162.835 ;
        RECT 64.490 161.205 64.810 162.165 ;
        RECT 65.340 162.135 66.170 162.435 ;
        RECT 64.980 161.235 65.170 161.955 ;
        RECT 65.340 161.065 65.510 162.135 ;
        RECT 65.970 162.105 66.170 162.135 ;
        RECT 65.680 161.885 65.850 161.955 ;
        RECT 66.380 161.885 66.550 162.665 ;
        RECT 67.415 162.525 67.585 162.665 ;
        RECT 67.755 162.655 68.005 163.115 ;
        RECT 65.680 161.715 66.550 161.885 ;
        RECT 66.720 162.245 67.245 162.465 ;
        RECT 67.415 162.395 67.640 162.525 ;
        RECT 65.680 161.625 66.190 161.715 ;
        RECT 64.150 160.865 65.035 161.035 ;
        RECT 65.260 160.735 65.510 161.065 ;
        RECT 65.680 160.565 65.850 161.365 ;
        RECT 66.020 161.010 66.190 161.625 ;
        RECT 66.720 161.545 66.890 162.245 ;
        RECT 66.360 161.180 66.890 161.545 ;
        RECT 67.060 161.480 67.300 162.075 ;
        RECT 67.470 161.290 67.640 162.395 ;
        RECT 67.810 161.535 68.090 162.485 ;
        RECT 67.335 161.160 67.640 161.290 ;
        RECT 66.020 160.840 67.125 161.010 ;
        RECT 67.335 160.735 67.585 161.160 ;
        RECT 67.755 160.565 68.020 161.025 ;
        RECT 68.260 160.735 68.445 162.855 ;
        RECT 68.615 162.735 68.945 163.115 ;
        RECT 69.115 162.565 69.285 162.855 ;
        RECT 68.620 162.395 69.285 162.565 ;
        RECT 68.620 161.405 68.850 162.395 ;
        RECT 70.465 162.315 70.805 162.945 ;
        RECT 70.975 162.315 71.225 163.115 ;
        RECT 71.415 162.465 71.745 162.945 ;
        RECT 71.915 162.655 72.140 163.115 ;
        RECT 72.310 162.465 72.640 162.945 ;
        RECT 69.020 161.575 69.370 162.225 ;
        RECT 70.465 161.705 70.640 162.315 ;
        RECT 71.415 162.295 72.640 162.465 ;
        RECT 73.270 162.335 73.770 162.945 ;
        RECT 70.810 161.955 71.505 162.125 ;
        RECT 71.335 161.705 71.505 161.955 ;
        RECT 71.680 161.925 72.100 162.125 ;
        RECT 72.270 161.925 72.600 162.125 ;
        RECT 72.770 161.925 73.100 162.125 ;
        RECT 73.270 161.705 73.440 162.335 ;
        RECT 74.145 162.315 74.485 162.945 ;
        RECT 74.655 162.315 74.905 163.115 ;
        RECT 75.095 162.465 75.425 162.945 ;
        RECT 75.595 162.655 75.820 163.115 ;
        RECT 75.990 162.465 76.320 162.945 ;
        RECT 73.625 161.875 73.975 162.125 ;
        RECT 74.145 161.705 74.320 162.315 ;
        RECT 75.095 162.295 76.320 162.465 ;
        RECT 76.950 162.335 77.450 162.945 ;
        RECT 77.825 162.615 78.085 162.945 ;
        RECT 78.255 162.755 78.585 163.115 ;
        RECT 78.840 162.735 80.140 162.945 ;
        RECT 74.490 161.955 75.185 162.125 ;
        RECT 75.015 161.705 75.185 161.955 ;
        RECT 75.360 161.925 75.780 162.125 ;
        RECT 75.950 161.925 76.280 162.125 ;
        RECT 76.450 161.925 76.780 162.125 ;
        RECT 76.950 161.705 77.120 162.335 ;
        RECT 77.305 161.875 77.655 162.125 ;
        RECT 68.620 161.235 69.285 161.405 ;
        RECT 68.615 160.565 68.945 161.065 ;
        RECT 69.115 160.735 69.285 161.235 ;
        RECT 70.465 160.735 70.805 161.705 ;
        RECT 70.975 160.565 71.145 161.705 ;
        RECT 71.335 161.535 73.770 161.705 ;
        RECT 71.415 160.565 71.665 161.365 ;
        RECT 72.310 160.735 72.640 161.535 ;
        RECT 72.940 160.565 73.270 161.365 ;
        RECT 73.440 160.735 73.770 161.535 ;
        RECT 74.145 160.735 74.485 161.705 ;
        RECT 74.655 160.565 74.825 161.705 ;
        RECT 75.015 161.535 77.450 161.705 ;
        RECT 75.095 160.565 75.345 161.365 ;
        RECT 75.990 160.735 76.320 161.535 ;
        RECT 76.620 160.565 76.950 161.365 ;
        RECT 77.120 160.735 77.450 161.535 ;
        RECT 77.825 161.415 77.995 162.615 ;
        RECT 78.840 162.585 79.010 162.735 ;
        RECT 78.255 162.460 79.010 162.585 ;
        RECT 78.165 162.415 79.010 162.460 ;
        RECT 78.165 162.295 78.435 162.415 ;
        RECT 78.165 161.720 78.335 162.295 ;
        RECT 78.565 161.855 78.975 162.160 ;
        RECT 79.265 162.125 79.475 162.525 ;
        RECT 79.145 161.915 79.475 162.125 ;
        RECT 79.720 162.125 79.940 162.525 ;
        RECT 80.415 162.350 80.870 163.115 ;
        RECT 81.965 162.365 83.175 163.115 ;
        RECT 79.720 161.915 80.195 162.125 ;
        RECT 80.385 161.925 80.875 162.125 ;
        RECT 78.165 161.685 78.365 161.720 ;
        RECT 79.695 161.685 80.870 161.745 ;
        RECT 78.165 161.575 80.870 161.685 ;
        RECT 78.225 161.515 80.025 161.575 ;
        RECT 79.695 161.485 80.025 161.515 ;
        RECT 77.825 160.735 78.085 161.415 ;
        RECT 78.255 160.565 78.505 161.345 ;
        RECT 78.755 161.315 79.590 161.325 ;
        RECT 80.180 161.315 80.365 161.405 ;
        RECT 78.755 161.115 80.365 161.315 ;
        RECT 78.755 160.735 79.005 161.115 ;
        RECT 80.135 161.075 80.365 161.115 ;
        RECT 80.615 160.955 80.870 161.575 ;
        RECT 79.175 160.565 79.530 160.945 ;
        RECT 80.535 160.735 80.870 160.955 ;
        RECT 81.965 161.655 82.485 162.195 ;
        RECT 82.655 161.825 83.175 162.365 ;
        RECT 81.965 160.565 83.175 161.655 ;
        RECT 5.520 160.395 83.260 160.565 ;
        RECT 5.605 159.305 6.815 160.395 ;
        RECT 6.985 159.960 12.330 160.395 ;
        RECT 12.505 159.960 17.850 160.395 ;
        RECT 5.605 158.595 6.125 159.135 ;
        RECT 6.295 158.765 6.815 159.305 ;
        RECT 5.605 157.845 6.815 158.595 ;
        RECT 8.570 158.390 8.910 159.220 ;
        RECT 10.390 158.710 10.740 159.960 ;
        RECT 14.090 158.390 14.430 159.220 ;
        RECT 15.910 158.710 16.260 159.960 ;
        RECT 18.485 159.230 18.775 160.395 ;
        RECT 18.945 159.960 24.290 160.395 ;
        RECT 24.465 159.960 29.810 160.395 ;
        RECT 6.985 157.845 12.330 158.390 ;
        RECT 12.505 157.845 17.850 158.390 ;
        RECT 18.485 157.845 18.775 158.570 ;
        RECT 20.530 158.390 20.870 159.220 ;
        RECT 22.350 158.710 22.700 159.960 ;
        RECT 26.050 158.390 26.390 159.220 ;
        RECT 27.870 158.710 28.220 159.960 ;
        RECT 29.985 159.305 31.655 160.395 ;
        RECT 32.375 159.725 32.545 160.225 ;
        RECT 32.715 159.895 33.045 160.395 ;
        RECT 32.375 159.555 33.040 159.725 ;
        RECT 29.985 158.615 30.735 159.135 ;
        RECT 30.905 158.785 31.655 159.305 ;
        RECT 32.290 158.735 32.640 159.385 ;
        RECT 18.945 157.845 24.290 158.390 ;
        RECT 24.465 157.845 29.810 158.390 ;
        RECT 29.985 157.845 31.655 158.615 ;
        RECT 32.810 158.565 33.040 159.555 ;
        RECT 32.375 158.395 33.040 158.565 ;
        RECT 32.375 158.105 32.545 158.395 ;
        RECT 32.715 157.845 33.045 158.225 ;
        RECT 33.215 158.105 33.400 160.225 ;
        RECT 33.640 159.935 33.905 160.395 ;
        RECT 34.075 159.800 34.325 160.225 ;
        RECT 34.535 159.950 35.640 160.120 ;
        RECT 34.020 159.670 34.325 159.800 ;
        RECT 33.570 158.475 33.850 159.425 ;
        RECT 34.020 158.565 34.190 159.670 ;
        RECT 34.360 158.885 34.600 159.480 ;
        RECT 34.770 159.415 35.300 159.780 ;
        RECT 34.770 158.715 34.940 159.415 ;
        RECT 35.470 159.335 35.640 159.950 ;
        RECT 35.810 159.595 35.980 160.395 ;
        RECT 36.150 159.895 36.400 160.225 ;
        RECT 36.625 159.925 37.510 160.095 ;
        RECT 35.470 159.245 35.980 159.335 ;
        RECT 34.020 158.435 34.245 158.565 ;
        RECT 34.415 158.495 34.940 158.715 ;
        RECT 35.110 159.075 35.980 159.245 ;
        RECT 33.655 157.845 33.905 158.305 ;
        RECT 34.075 158.295 34.245 158.435 ;
        RECT 35.110 158.295 35.280 159.075 ;
        RECT 35.810 159.005 35.980 159.075 ;
        RECT 35.490 158.825 35.690 158.855 ;
        RECT 36.150 158.825 36.320 159.895 ;
        RECT 36.490 159.005 36.680 159.725 ;
        RECT 35.490 158.525 36.320 158.825 ;
        RECT 36.850 158.795 37.170 159.755 ;
        RECT 34.075 158.125 34.410 158.295 ;
        RECT 34.605 158.125 35.280 158.295 ;
        RECT 35.600 157.845 35.970 158.345 ;
        RECT 36.150 158.295 36.320 158.525 ;
        RECT 36.705 158.465 37.170 158.795 ;
        RECT 37.340 159.085 37.510 159.925 ;
        RECT 37.690 159.895 38.005 160.395 ;
        RECT 38.235 159.665 38.575 160.225 ;
        RECT 37.680 159.290 38.575 159.665 ;
        RECT 38.745 159.385 38.915 160.395 ;
        RECT 38.385 159.085 38.575 159.290 ;
        RECT 39.085 159.335 39.415 160.180 ;
        RECT 39.680 159.605 40.215 160.225 ;
        RECT 39.085 159.255 39.475 159.335 ;
        RECT 39.260 159.205 39.475 159.255 ;
        RECT 37.340 158.755 38.215 159.085 ;
        RECT 38.385 158.755 39.135 159.085 ;
        RECT 37.340 158.295 37.510 158.755 ;
        RECT 38.385 158.585 38.585 158.755 ;
        RECT 39.305 158.625 39.475 159.205 ;
        RECT 39.250 158.585 39.475 158.625 ;
        RECT 36.150 158.125 36.555 158.295 ;
        RECT 36.725 158.125 37.510 158.295 ;
        RECT 37.785 157.845 37.995 158.375 ;
        RECT 38.255 158.060 38.585 158.585 ;
        RECT 39.095 158.500 39.475 158.585 ;
        RECT 39.680 158.585 39.995 159.605 ;
        RECT 40.385 159.595 40.715 160.395 ;
        RECT 41.200 159.425 41.590 159.600 ;
        RECT 41.950 159.595 42.205 160.395 ;
        RECT 42.405 159.545 42.735 160.225 ;
        RECT 40.165 159.255 41.590 159.425 ;
        RECT 40.165 158.755 40.335 159.255 ;
        RECT 38.755 157.845 38.925 158.455 ;
        RECT 39.095 158.065 39.425 158.500 ;
        RECT 39.680 158.015 40.295 158.585 ;
        RECT 40.585 158.525 40.850 159.085 ;
        RECT 41.020 158.355 41.190 159.255 ;
        RECT 41.360 158.525 41.715 159.085 ;
        RECT 41.950 159.055 42.195 159.415 ;
        RECT 42.385 159.265 42.735 159.545 ;
        RECT 42.385 158.885 42.555 159.265 ;
        RECT 42.915 159.085 43.110 160.135 ;
        RECT 43.290 159.255 43.610 160.395 ;
        RECT 44.245 159.230 44.535 160.395 ;
        RECT 44.705 159.255 45.090 160.225 ;
        RECT 45.260 159.935 45.585 160.395 ;
        RECT 46.105 159.765 46.385 160.225 ;
        RECT 45.260 159.545 46.385 159.765 ;
        RECT 42.035 158.715 42.555 158.885 ;
        RECT 42.725 158.755 43.110 159.085 ;
        RECT 43.290 159.035 43.550 159.085 ;
        RECT 43.290 158.865 43.555 159.035 ;
        RECT 43.290 158.755 43.550 158.865 ;
        RECT 42.035 158.355 42.205 158.715 ;
        RECT 44.705 158.585 44.985 159.255 ;
        RECT 45.260 159.085 45.710 159.545 ;
        RECT 46.575 159.375 46.975 160.225 ;
        RECT 47.375 159.935 47.645 160.395 ;
        RECT 47.815 159.765 48.100 160.225 ;
        RECT 45.155 158.755 45.710 159.085 ;
        RECT 45.880 158.815 46.975 159.375 ;
        RECT 45.260 158.645 45.710 158.755 ;
        RECT 40.465 157.845 40.680 158.355 ;
        RECT 40.910 158.025 41.190 158.355 ;
        RECT 41.370 157.845 41.610 158.355 ;
        RECT 42.005 158.185 42.205 158.355 ;
        RECT 42.035 158.150 42.205 158.185 ;
        RECT 42.395 158.375 43.610 158.545 ;
        RECT 42.395 158.070 42.625 158.375 ;
        RECT 42.795 157.845 43.125 158.205 ;
        RECT 43.320 158.025 43.610 158.375 ;
        RECT 44.245 157.845 44.535 158.570 ;
        RECT 44.705 158.015 45.090 158.585 ;
        RECT 45.260 158.475 46.385 158.645 ;
        RECT 45.260 157.845 45.585 158.305 ;
        RECT 46.105 158.015 46.385 158.475 ;
        RECT 46.575 158.015 46.975 158.815 ;
        RECT 47.145 159.545 48.100 159.765 ;
        RECT 48.475 159.725 48.645 160.225 ;
        RECT 48.815 159.895 49.145 160.395 ;
        RECT 48.475 159.555 49.140 159.725 ;
        RECT 47.145 158.645 47.355 159.545 ;
        RECT 47.525 158.815 48.215 159.375 ;
        RECT 48.390 158.735 48.740 159.385 ;
        RECT 47.145 158.475 48.100 158.645 ;
        RECT 48.910 158.565 49.140 159.555 ;
        RECT 47.375 157.845 47.645 158.305 ;
        RECT 47.815 158.015 48.100 158.475 ;
        RECT 48.475 158.395 49.140 158.565 ;
        RECT 48.475 158.105 48.645 158.395 ;
        RECT 48.815 157.845 49.145 158.225 ;
        RECT 49.315 158.105 49.500 160.225 ;
        RECT 49.740 159.935 50.005 160.395 ;
        RECT 50.175 159.800 50.425 160.225 ;
        RECT 50.635 159.950 51.740 160.120 ;
        RECT 50.120 159.670 50.425 159.800 ;
        RECT 49.670 158.475 49.950 159.425 ;
        RECT 50.120 158.565 50.290 159.670 ;
        RECT 50.460 158.885 50.700 159.480 ;
        RECT 50.870 159.415 51.400 159.780 ;
        RECT 50.870 158.715 51.040 159.415 ;
        RECT 51.570 159.335 51.740 159.950 ;
        RECT 51.910 159.595 52.080 160.395 ;
        RECT 52.250 159.895 52.500 160.225 ;
        RECT 52.725 159.925 53.610 160.095 ;
        RECT 51.570 159.245 52.080 159.335 ;
        RECT 50.120 158.435 50.345 158.565 ;
        RECT 50.515 158.495 51.040 158.715 ;
        RECT 51.210 159.075 52.080 159.245 ;
        RECT 49.755 157.845 50.005 158.305 ;
        RECT 50.175 158.295 50.345 158.435 ;
        RECT 51.210 158.295 51.380 159.075 ;
        RECT 51.910 159.005 52.080 159.075 ;
        RECT 51.590 158.825 51.790 158.855 ;
        RECT 52.250 158.825 52.420 159.895 ;
        RECT 52.590 159.005 52.780 159.725 ;
        RECT 51.590 158.525 52.420 158.825 ;
        RECT 52.950 158.795 53.270 159.755 ;
        RECT 50.175 158.125 50.510 158.295 ;
        RECT 50.705 158.125 51.380 158.295 ;
        RECT 51.700 157.845 52.070 158.345 ;
        RECT 52.250 158.295 52.420 158.525 ;
        RECT 52.805 158.465 53.270 158.795 ;
        RECT 53.440 159.085 53.610 159.925 ;
        RECT 53.790 159.895 54.105 160.395 ;
        RECT 54.335 159.665 54.675 160.225 ;
        RECT 53.780 159.290 54.675 159.665 ;
        RECT 54.845 159.385 55.015 160.395 ;
        RECT 54.485 159.085 54.675 159.290 ;
        RECT 55.185 159.335 55.515 160.180 ;
        RECT 55.185 159.255 55.575 159.335 ;
        RECT 55.360 159.205 55.575 159.255 ;
        RECT 53.440 158.755 54.315 159.085 ;
        RECT 54.485 158.755 55.235 159.085 ;
        RECT 53.440 158.295 53.610 158.755 ;
        RECT 54.485 158.585 54.685 158.755 ;
        RECT 55.405 158.625 55.575 159.205 ;
        RECT 55.350 158.585 55.575 158.625 ;
        RECT 52.250 158.125 52.655 158.295 ;
        RECT 52.825 158.125 53.610 158.295 ;
        RECT 53.885 157.845 54.095 158.375 ;
        RECT 54.355 158.060 54.685 158.585 ;
        RECT 55.195 158.500 55.575 158.585 ;
        RECT 55.750 159.255 56.085 160.225 ;
        RECT 56.255 159.255 56.425 160.395 ;
        RECT 56.595 160.055 58.625 160.225 ;
        RECT 55.750 158.585 55.920 159.255 ;
        RECT 56.595 159.085 56.765 160.055 ;
        RECT 56.090 158.755 56.345 159.085 ;
        RECT 56.570 158.755 56.765 159.085 ;
        RECT 56.935 159.715 58.060 159.885 ;
        RECT 56.175 158.585 56.345 158.755 ;
        RECT 56.935 158.585 57.105 159.715 ;
        RECT 54.855 157.845 55.025 158.455 ;
        RECT 55.195 158.065 55.525 158.500 ;
        RECT 55.750 158.015 56.005 158.585 ;
        RECT 56.175 158.415 57.105 158.585 ;
        RECT 57.275 159.375 58.285 159.545 ;
        RECT 57.275 158.575 57.445 159.375 ;
        RECT 56.930 158.380 57.105 158.415 ;
        RECT 56.175 157.845 56.505 158.245 ;
        RECT 56.930 158.015 57.460 158.380 ;
        RECT 57.650 158.355 57.925 159.175 ;
        RECT 57.645 158.185 57.925 158.355 ;
        RECT 57.650 158.015 57.925 158.185 ;
        RECT 58.095 158.015 58.285 159.375 ;
        RECT 58.455 159.390 58.625 160.055 ;
        RECT 58.795 159.635 58.965 160.395 ;
        RECT 59.200 159.635 59.715 160.045 ;
        RECT 58.455 159.200 59.205 159.390 ;
        RECT 59.375 158.825 59.715 159.635 ;
        RECT 60.865 159.335 61.195 160.180 ;
        RECT 61.365 159.385 61.535 160.395 ;
        RECT 61.705 159.665 62.045 160.225 ;
        RECT 62.275 159.895 62.590 160.395 ;
        RECT 62.770 159.925 63.655 160.095 ;
        RECT 58.485 158.655 59.715 158.825 ;
        RECT 60.805 159.255 61.195 159.335 ;
        RECT 61.705 159.290 62.600 159.665 ;
        RECT 60.805 159.205 61.020 159.255 ;
        RECT 58.465 157.845 58.975 158.380 ;
        RECT 59.195 158.050 59.440 158.655 ;
        RECT 60.805 158.625 60.975 159.205 ;
        RECT 61.705 159.085 61.895 159.290 ;
        RECT 62.770 159.085 62.940 159.925 ;
        RECT 63.880 159.895 64.130 160.225 ;
        RECT 61.145 158.755 61.895 159.085 ;
        RECT 62.065 158.755 62.940 159.085 ;
        RECT 60.805 158.585 61.030 158.625 ;
        RECT 61.695 158.585 61.895 158.755 ;
        RECT 60.805 158.500 61.185 158.585 ;
        RECT 60.855 158.065 61.185 158.500 ;
        RECT 61.355 157.845 61.525 158.455 ;
        RECT 61.695 158.060 62.025 158.585 ;
        RECT 62.285 157.845 62.495 158.375 ;
        RECT 62.770 158.295 62.940 158.755 ;
        RECT 63.110 158.795 63.430 159.755 ;
        RECT 63.600 159.005 63.790 159.725 ;
        RECT 63.960 158.825 64.130 159.895 ;
        RECT 64.300 159.595 64.470 160.395 ;
        RECT 64.640 159.950 65.745 160.120 ;
        RECT 64.640 159.335 64.810 159.950 ;
        RECT 65.955 159.800 66.205 160.225 ;
        RECT 66.375 159.935 66.640 160.395 ;
        RECT 64.980 159.415 65.510 159.780 ;
        RECT 65.955 159.670 66.260 159.800 ;
        RECT 64.300 159.245 64.810 159.335 ;
        RECT 64.300 159.075 65.170 159.245 ;
        RECT 64.300 159.005 64.470 159.075 ;
        RECT 64.590 158.825 64.790 158.855 ;
        RECT 63.110 158.465 63.575 158.795 ;
        RECT 63.960 158.525 64.790 158.825 ;
        RECT 63.960 158.295 64.130 158.525 ;
        RECT 62.770 158.125 63.555 158.295 ;
        RECT 63.725 158.125 64.130 158.295 ;
        RECT 64.310 157.845 64.680 158.345 ;
        RECT 65.000 158.295 65.170 159.075 ;
        RECT 65.340 158.715 65.510 159.415 ;
        RECT 65.680 158.885 65.920 159.480 ;
        RECT 65.340 158.495 65.865 158.715 ;
        RECT 66.090 158.565 66.260 159.670 ;
        RECT 66.035 158.435 66.260 158.565 ;
        RECT 66.430 158.475 66.710 159.425 ;
        RECT 66.035 158.295 66.205 158.435 ;
        RECT 65.000 158.125 65.675 158.295 ;
        RECT 65.870 158.125 66.205 158.295 ;
        RECT 66.375 157.845 66.625 158.305 ;
        RECT 66.880 158.105 67.065 160.225 ;
        RECT 67.235 159.895 67.565 160.395 ;
        RECT 67.735 159.725 67.905 160.225 ;
        RECT 67.240 159.555 67.905 159.725 ;
        RECT 67.240 158.565 67.470 159.555 ;
        RECT 68.255 159.465 68.425 160.225 ;
        RECT 68.640 159.635 68.970 160.395 ;
        RECT 67.640 158.735 67.990 159.385 ;
        RECT 68.255 159.295 68.970 159.465 ;
        RECT 69.140 159.320 69.395 160.225 ;
        RECT 68.165 158.745 68.520 159.115 ;
        RECT 68.800 159.085 68.970 159.295 ;
        RECT 68.800 158.755 69.055 159.085 ;
        RECT 68.800 158.565 68.970 158.755 ;
        RECT 69.225 158.590 69.395 159.320 ;
        RECT 69.570 159.245 69.830 160.395 ;
        RECT 70.005 159.230 70.295 160.395 ;
        RECT 70.555 159.725 70.725 160.225 ;
        RECT 70.895 159.895 71.225 160.395 ;
        RECT 70.555 159.555 71.220 159.725 ;
        RECT 70.470 158.735 70.820 159.385 ;
        RECT 67.240 158.395 67.905 158.565 ;
        RECT 67.235 157.845 67.565 158.225 ;
        RECT 67.735 158.105 67.905 158.395 ;
        RECT 68.255 158.395 68.970 158.565 ;
        RECT 68.255 158.015 68.425 158.395 ;
        RECT 68.640 157.845 68.970 158.225 ;
        RECT 69.140 158.015 69.395 158.590 ;
        RECT 69.570 157.845 69.830 158.685 ;
        RECT 70.005 157.845 70.295 158.570 ;
        RECT 70.990 158.565 71.220 159.555 ;
        RECT 70.555 158.395 71.220 158.565 ;
        RECT 70.555 158.105 70.725 158.395 ;
        RECT 70.895 157.845 71.225 158.225 ;
        RECT 71.395 158.105 71.580 160.225 ;
        RECT 71.820 159.935 72.085 160.395 ;
        RECT 72.255 159.800 72.505 160.225 ;
        RECT 72.715 159.950 73.820 160.120 ;
        RECT 72.200 159.670 72.505 159.800 ;
        RECT 71.750 158.475 72.030 159.425 ;
        RECT 72.200 158.565 72.370 159.670 ;
        RECT 72.540 158.885 72.780 159.480 ;
        RECT 72.950 159.415 73.480 159.780 ;
        RECT 72.950 158.715 73.120 159.415 ;
        RECT 73.650 159.335 73.820 159.950 ;
        RECT 73.990 159.595 74.160 160.395 ;
        RECT 74.330 159.895 74.580 160.225 ;
        RECT 74.805 159.925 75.690 160.095 ;
        RECT 73.650 159.245 74.160 159.335 ;
        RECT 72.200 158.435 72.425 158.565 ;
        RECT 72.595 158.495 73.120 158.715 ;
        RECT 73.290 159.075 74.160 159.245 ;
        RECT 71.835 157.845 72.085 158.305 ;
        RECT 72.255 158.295 72.425 158.435 ;
        RECT 73.290 158.295 73.460 159.075 ;
        RECT 73.990 159.005 74.160 159.075 ;
        RECT 73.670 158.825 73.870 158.855 ;
        RECT 74.330 158.825 74.500 159.895 ;
        RECT 74.670 159.005 74.860 159.725 ;
        RECT 73.670 158.525 74.500 158.825 ;
        RECT 75.030 158.795 75.350 159.755 ;
        RECT 72.255 158.125 72.590 158.295 ;
        RECT 72.785 158.125 73.460 158.295 ;
        RECT 73.780 157.845 74.150 158.345 ;
        RECT 74.330 158.295 74.500 158.525 ;
        RECT 74.885 158.465 75.350 158.795 ;
        RECT 75.520 159.085 75.690 159.925 ;
        RECT 75.870 159.895 76.185 160.395 ;
        RECT 76.415 159.665 76.755 160.225 ;
        RECT 75.860 159.290 76.755 159.665 ;
        RECT 76.925 159.385 77.095 160.395 ;
        RECT 76.565 159.085 76.755 159.290 ;
        RECT 77.265 159.335 77.595 160.180 ;
        RECT 78.290 160.005 78.625 160.225 ;
        RECT 79.630 160.015 79.985 160.395 ;
        RECT 78.290 159.385 78.545 160.005 ;
        RECT 78.795 159.845 79.025 159.885 ;
        RECT 80.155 159.845 80.405 160.225 ;
        RECT 78.795 159.645 80.405 159.845 ;
        RECT 78.795 159.555 78.980 159.645 ;
        RECT 79.570 159.635 80.405 159.645 ;
        RECT 80.655 159.615 80.905 160.395 ;
        RECT 81.075 159.545 81.335 160.225 ;
        RECT 79.135 159.445 79.465 159.475 ;
        RECT 79.135 159.385 80.935 159.445 ;
        RECT 77.265 159.255 77.655 159.335 ;
        RECT 77.440 159.205 77.655 159.255 ;
        RECT 78.290 159.275 80.995 159.385 ;
        RECT 78.290 159.215 79.465 159.275 ;
        RECT 80.795 159.240 80.995 159.275 ;
        RECT 75.520 158.755 76.395 159.085 ;
        RECT 76.565 158.755 77.315 159.085 ;
        RECT 75.520 158.295 75.690 158.755 ;
        RECT 76.565 158.585 76.765 158.755 ;
        RECT 77.485 158.625 77.655 159.205 ;
        RECT 78.285 158.835 78.775 159.035 ;
        RECT 78.965 158.835 79.440 159.045 ;
        RECT 77.430 158.585 77.655 158.625 ;
        RECT 74.330 158.125 74.735 158.295 ;
        RECT 74.905 158.125 75.690 158.295 ;
        RECT 75.965 157.845 76.175 158.375 ;
        RECT 76.435 158.060 76.765 158.585 ;
        RECT 77.275 158.500 77.655 158.585 ;
        RECT 76.935 157.845 77.105 158.455 ;
        RECT 77.275 158.065 77.605 158.500 ;
        RECT 78.290 157.845 78.745 158.610 ;
        RECT 79.220 158.435 79.440 158.835 ;
        RECT 79.685 158.835 80.015 159.045 ;
        RECT 79.685 158.435 79.895 158.835 ;
        RECT 80.185 158.800 80.595 159.105 ;
        RECT 80.825 158.665 80.995 159.240 ;
        RECT 80.725 158.545 80.995 158.665 ;
        RECT 80.150 158.500 80.995 158.545 ;
        RECT 80.150 158.375 80.905 158.500 ;
        RECT 80.150 158.225 80.320 158.375 ;
        RECT 81.165 158.345 81.335 159.545 ;
        RECT 81.965 159.305 83.175 160.395 ;
        RECT 81.965 158.765 82.485 159.305 ;
        RECT 82.655 158.595 83.175 159.135 ;
        RECT 79.020 158.015 80.320 158.225 ;
        RECT 80.575 157.845 80.905 158.205 ;
        RECT 81.075 158.015 81.335 158.345 ;
        RECT 81.965 157.845 83.175 158.595 ;
        RECT 5.520 157.675 83.260 157.845 ;
        RECT 5.605 156.925 6.815 157.675 ;
        RECT 6.985 157.130 12.330 157.675 ;
        RECT 12.505 157.130 17.850 157.675 ;
        RECT 18.025 157.130 23.370 157.675 ;
        RECT 23.545 157.130 28.890 157.675 ;
        RECT 5.605 156.385 6.125 156.925 ;
        RECT 6.295 156.215 6.815 156.755 ;
        RECT 8.570 156.300 8.910 157.130 ;
        RECT 5.605 155.125 6.815 156.215 ;
        RECT 10.390 155.560 10.740 156.810 ;
        RECT 14.090 156.300 14.430 157.130 ;
        RECT 15.910 155.560 16.260 156.810 ;
        RECT 19.610 156.300 19.950 157.130 ;
        RECT 21.430 155.560 21.780 156.810 ;
        RECT 25.130 156.300 25.470 157.130 ;
        RECT 29.065 156.905 30.735 157.675 ;
        RECT 31.365 156.950 31.655 157.675 ;
        RECT 31.825 156.905 33.495 157.675 ;
        RECT 33.665 156.935 34.050 157.505 ;
        RECT 34.220 157.215 34.545 157.675 ;
        RECT 35.065 157.045 35.345 157.505 ;
        RECT 26.950 155.560 27.300 156.810 ;
        RECT 29.065 156.385 29.815 156.905 ;
        RECT 29.985 156.215 30.735 156.735 ;
        RECT 31.825 156.385 32.575 156.905 ;
        RECT 6.985 155.125 12.330 155.560 ;
        RECT 12.505 155.125 17.850 155.560 ;
        RECT 18.025 155.125 23.370 155.560 ;
        RECT 23.545 155.125 28.890 155.560 ;
        RECT 29.065 155.125 30.735 156.215 ;
        RECT 31.365 155.125 31.655 156.290 ;
        RECT 32.745 156.215 33.495 156.735 ;
        RECT 31.825 155.125 33.495 156.215 ;
        RECT 33.665 156.265 33.945 156.935 ;
        RECT 34.220 156.875 35.345 157.045 ;
        RECT 34.220 156.765 34.670 156.875 ;
        RECT 34.115 156.435 34.670 156.765 ;
        RECT 35.535 156.705 35.935 157.505 ;
        RECT 36.335 157.215 36.605 157.675 ;
        RECT 36.775 157.045 37.060 157.505 ;
        RECT 33.665 155.295 34.050 156.265 ;
        RECT 34.220 155.975 34.670 156.435 ;
        RECT 34.840 156.145 35.935 156.705 ;
        RECT 34.220 155.755 35.345 155.975 ;
        RECT 34.220 155.125 34.545 155.585 ;
        RECT 35.065 155.295 35.345 155.755 ;
        RECT 35.535 155.295 35.935 156.145 ;
        RECT 36.105 156.875 37.060 157.045 ;
        RECT 37.345 156.950 37.605 157.505 ;
        RECT 37.775 157.230 38.205 157.675 ;
        RECT 38.440 157.105 38.610 157.505 ;
        RECT 38.780 157.275 39.500 157.675 ;
        RECT 36.105 155.975 36.315 156.875 ;
        RECT 36.485 156.145 37.175 156.705 ;
        RECT 37.345 156.235 37.520 156.950 ;
        RECT 38.440 156.935 39.320 157.105 ;
        RECT 39.670 157.060 39.840 157.505 ;
        RECT 40.415 157.165 40.815 157.675 ;
        RECT 37.690 156.435 37.945 156.765 ;
        RECT 36.105 155.755 37.060 155.975 ;
        RECT 36.335 155.125 36.605 155.585 ;
        RECT 36.775 155.295 37.060 155.755 ;
        RECT 37.345 155.295 37.605 156.235 ;
        RECT 37.775 155.955 37.945 156.435 ;
        RECT 38.170 156.145 38.500 156.765 ;
        RECT 38.670 156.385 38.960 156.765 ;
        RECT 39.150 156.215 39.320 156.935 ;
        RECT 38.800 156.045 39.320 156.215 ;
        RECT 39.490 156.890 39.840 157.060 ;
        RECT 41.115 157.125 41.285 157.415 ;
        RECT 41.455 157.295 41.785 157.675 ;
        RECT 37.775 155.785 38.535 155.955 ;
        RECT 38.800 155.855 38.970 156.045 ;
        RECT 39.490 155.865 39.660 156.890 ;
        RECT 40.080 156.405 40.340 156.995 ;
        RECT 39.860 156.105 40.340 156.405 ;
        RECT 40.540 156.105 40.800 156.995 ;
        RECT 41.115 156.955 41.780 157.125 ;
        RECT 41.030 156.135 41.380 156.785 ;
        RECT 41.550 155.965 41.780 156.955 ;
        RECT 38.365 155.560 38.535 155.785 ;
        RECT 39.250 155.695 39.660 155.865 ;
        RECT 39.835 155.755 40.775 155.925 ;
        RECT 39.250 155.560 39.505 155.695 ;
        RECT 37.775 155.125 38.105 155.525 ;
        RECT 38.365 155.390 39.505 155.560 ;
        RECT 39.835 155.505 40.005 155.755 ;
        RECT 39.250 155.295 39.505 155.390 ;
        RECT 39.675 155.335 40.005 155.505 ;
        RECT 40.175 155.125 40.425 155.585 ;
        RECT 40.595 155.295 40.775 155.755 ;
        RECT 41.115 155.795 41.780 155.965 ;
        RECT 41.115 155.295 41.285 155.795 ;
        RECT 41.455 155.125 41.785 155.625 ;
        RECT 41.955 155.295 42.140 157.415 ;
        RECT 42.395 157.215 42.645 157.675 ;
        RECT 42.815 157.225 43.150 157.395 ;
        RECT 43.345 157.225 44.020 157.395 ;
        RECT 42.815 157.085 42.985 157.225 ;
        RECT 42.310 156.095 42.590 157.045 ;
        RECT 42.760 156.955 42.985 157.085 ;
        RECT 42.760 155.850 42.930 156.955 ;
        RECT 43.155 156.805 43.680 157.025 ;
        RECT 43.100 156.040 43.340 156.635 ;
        RECT 43.510 156.105 43.680 156.805 ;
        RECT 43.850 156.445 44.020 157.225 ;
        RECT 44.340 157.175 44.710 157.675 ;
        RECT 44.890 157.225 45.295 157.395 ;
        RECT 45.465 157.225 46.250 157.395 ;
        RECT 44.890 156.995 45.060 157.225 ;
        RECT 44.230 156.695 45.060 156.995 ;
        RECT 45.445 156.725 45.910 157.055 ;
        RECT 44.230 156.665 44.430 156.695 ;
        RECT 44.550 156.445 44.720 156.515 ;
        RECT 43.850 156.275 44.720 156.445 ;
        RECT 44.210 156.185 44.720 156.275 ;
        RECT 42.760 155.720 43.065 155.850 ;
        RECT 43.510 155.740 44.040 156.105 ;
        RECT 42.380 155.125 42.645 155.585 ;
        RECT 42.815 155.295 43.065 155.720 ;
        RECT 44.210 155.570 44.380 156.185 ;
        RECT 43.275 155.400 44.380 155.570 ;
        RECT 44.550 155.125 44.720 155.925 ;
        RECT 44.890 155.625 45.060 156.695 ;
        RECT 45.230 155.795 45.420 156.515 ;
        RECT 45.590 155.765 45.910 156.725 ;
        RECT 46.080 156.765 46.250 157.225 ;
        RECT 46.525 157.145 46.735 157.675 ;
        RECT 46.995 156.935 47.325 157.460 ;
        RECT 47.495 157.065 47.665 157.675 ;
        RECT 47.835 157.020 48.165 157.455 ;
        RECT 48.475 157.125 48.645 157.415 ;
        RECT 48.815 157.295 49.145 157.675 ;
        RECT 47.835 156.935 48.215 157.020 ;
        RECT 48.475 156.955 49.140 157.125 ;
        RECT 47.125 156.765 47.325 156.935 ;
        RECT 47.990 156.895 48.215 156.935 ;
        RECT 46.080 156.435 46.955 156.765 ;
        RECT 47.125 156.435 47.875 156.765 ;
        RECT 44.890 155.295 45.140 155.625 ;
        RECT 46.080 155.595 46.250 156.435 ;
        RECT 47.125 156.230 47.315 156.435 ;
        RECT 48.045 156.315 48.215 156.895 ;
        RECT 48.000 156.265 48.215 156.315 ;
        RECT 46.420 155.855 47.315 156.230 ;
        RECT 47.825 156.185 48.215 156.265 ;
        RECT 45.365 155.425 46.250 155.595 ;
        RECT 46.430 155.125 46.745 155.625 ;
        RECT 46.975 155.295 47.315 155.855 ;
        RECT 47.485 155.125 47.655 156.135 ;
        RECT 47.825 155.340 48.155 156.185 ;
        RECT 48.390 156.135 48.740 156.785 ;
        RECT 48.910 155.965 49.140 156.955 ;
        RECT 48.475 155.795 49.140 155.965 ;
        RECT 48.475 155.295 48.645 155.795 ;
        RECT 48.815 155.125 49.145 155.625 ;
        RECT 49.315 155.295 49.500 157.415 ;
        RECT 49.755 157.215 50.005 157.675 ;
        RECT 50.175 157.225 50.510 157.395 ;
        RECT 50.705 157.225 51.380 157.395 ;
        RECT 50.175 157.085 50.345 157.225 ;
        RECT 49.670 156.095 49.950 157.045 ;
        RECT 50.120 156.955 50.345 157.085 ;
        RECT 50.120 155.850 50.290 156.955 ;
        RECT 50.515 156.805 51.040 157.025 ;
        RECT 50.460 156.040 50.700 156.635 ;
        RECT 50.870 156.105 51.040 156.805 ;
        RECT 51.210 156.445 51.380 157.225 ;
        RECT 51.700 157.175 52.070 157.675 ;
        RECT 52.250 157.225 52.655 157.395 ;
        RECT 52.825 157.225 53.610 157.395 ;
        RECT 52.250 156.995 52.420 157.225 ;
        RECT 51.590 156.695 52.420 156.995 ;
        RECT 52.805 156.725 53.270 157.055 ;
        RECT 51.590 156.665 51.790 156.695 ;
        RECT 51.910 156.445 52.080 156.515 ;
        RECT 51.210 156.275 52.080 156.445 ;
        RECT 51.570 156.185 52.080 156.275 ;
        RECT 50.120 155.720 50.425 155.850 ;
        RECT 50.870 155.740 51.400 156.105 ;
        RECT 49.740 155.125 50.005 155.585 ;
        RECT 50.175 155.295 50.425 155.720 ;
        RECT 51.570 155.570 51.740 156.185 ;
        RECT 50.635 155.400 51.740 155.570 ;
        RECT 51.910 155.125 52.080 155.925 ;
        RECT 52.250 155.625 52.420 156.695 ;
        RECT 52.590 155.795 52.780 156.515 ;
        RECT 52.950 155.765 53.270 156.725 ;
        RECT 53.440 156.765 53.610 157.225 ;
        RECT 53.885 157.145 54.095 157.675 ;
        RECT 54.355 156.935 54.685 157.460 ;
        RECT 54.855 157.065 55.025 157.675 ;
        RECT 55.195 157.020 55.525 157.455 ;
        RECT 55.195 156.935 55.575 157.020 ;
        RECT 54.485 156.765 54.685 156.935 ;
        RECT 55.350 156.895 55.575 156.935 ;
        RECT 53.440 156.435 54.315 156.765 ;
        RECT 54.485 156.435 55.235 156.765 ;
        RECT 52.250 155.295 52.500 155.625 ;
        RECT 53.440 155.595 53.610 156.435 ;
        RECT 54.485 156.230 54.675 156.435 ;
        RECT 55.405 156.315 55.575 156.895 ;
        RECT 55.745 156.925 56.955 157.675 ;
        RECT 57.125 156.950 57.415 157.675 ;
        RECT 57.635 157.020 57.965 157.455 ;
        RECT 58.135 157.065 58.305 157.675 ;
        RECT 57.585 156.935 57.965 157.020 ;
        RECT 58.475 156.935 58.805 157.460 ;
        RECT 59.065 157.145 59.275 157.675 ;
        RECT 59.550 157.225 60.335 157.395 ;
        RECT 60.505 157.225 60.910 157.395 ;
        RECT 55.745 156.385 56.265 156.925 ;
        RECT 57.585 156.895 57.810 156.935 ;
        RECT 55.360 156.265 55.575 156.315 ;
        RECT 53.780 155.855 54.675 156.230 ;
        RECT 55.185 156.185 55.575 156.265 ;
        RECT 56.435 156.215 56.955 156.755 ;
        RECT 57.585 156.315 57.755 156.895 ;
        RECT 58.475 156.765 58.675 156.935 ;
        RECT 59.550 156.765 59.720 157.225 ;
        RECT 57.925 156.435 58.675 156.765 ;
        RECT 58.845 156.435 59.720 156.765 ;
        RECT 52.725 155.425 53.610 155.595 ;
        RECT 53.790 155.125 54.105 155.625 ;
        RECT 54.335 155.295 54.675 155.855 ;
        RECT 54.845 155.125 55.015 156.135 ;
        RECT 55.185 155.340 55.515 156.185 ;
        RECT 55.745 155.125 56.955 156.215 ;
        RECT 57.125 155.125 57.415 156.290 ;
        RECT 57.585 156.265 57.800 156.315 ;
        RECT 57.585 156.185 57.975 156.265 ;
        RECT 57.645 155.340 57.975 156.185 ;
        RECT 58.485 156.230 58.675 156.435 ;
        RECT 58.145 155.125 58.315 156.135 ;
        RECT 58.485 155.855 59.380 156.230 ;
        RECT 58.485 155.295 58.825 155.855 ;
        RECT 59.055 155.125 59.370 155.625 ;
        RECT 59.550 155.595 59.720 156.435 ;
        RECT 59.890 156.725 60.355 157.055 ;
        RECT 60.740 156.995 60.910 157.225 ;
        RECT 61.090 157.175 61.460 157.675 ;
        RECT 61.780 157.225 62.455 157.395 ;
        RECT 62.650 157.225 62.985 157.395 ;
        RECT 59.890 155.765 60.210 156.725 ;
        RECT 60.740 156.695 61.570 156.995 ;
        RECT 60.380 155.795 60.570 156.515 ;
        RECT 60.740 155.625 60.910 156.695 ;
        RECT 61.370 156.665 61.570 156.695 ;
        RECT 61.080 156.445 61.250 156.515 ;
        RECT 61.780 156.445 61.950 157.225 ;
        RECT 62.815 157.085 62.985 157.225 ;
        RECT 63.155 157.215 63.405 157.675 ;
        RECT 61.080 156.275 61.950 156.445 ;
        RECT 62.120 156.805 62.645 157.025 ;
        RECT 62.815 156.955 63.040 157.085 ;
        RECT 61.080 156.185 61.590 156.275 ;
        RECT 59.550 155.425 60.435 155.595 ;
        RECT 60.660 155.295 60.910 155.625 ;
        RECT 61.080 155.125 61.250 155.925 ;
        RECT 61.420 155.570 61.590 156.185 ;
        RECT 62.120 156.105 62.290 156.805 ;
        RECT 61.760 155.740 62.290 156.105 ;
        RECT 62.460 156.040 62.700 156.635 ;
        RECT 62.870 155.850 63.040 156.955 ;
        RECT 63.210 156.095 63.490 157.045 ;
        RECT 62.735 155.720 63.040 155.850 ;
        RECT 61.420 155.400 62.525 155.570 ;
        RECT 62.735 155.295 62.985 155.720 ;
        RECT 63.155 155.125 63.420 155.585 ;
        RECT 63.660 155.295 63.845 157.415 ;
        RECT 64.015 157.295 64.345 157.675 ;
        RECT 64.515 157.125 64.685 157.415 ;
        RECT 65.005 157.195 65.285 157.675 ;
        RECT 64.020 156.955 64.685 157.125 ;
        RECT 65.455 157.025 65.715 157.415 ;
        RECT 65.890 157.195 66.145 157.675 ;
        RECT 66.315 157.025 66.610 157.415 ;
        RECT 66.790 157.195 67.065 157.675 ;
        RECT 67.235 157.175 67.535 157.505 ;
        RECT 64.020 155.965 64.250 156.955 ;
        RECT 64.960 156.855 66.610 157.025 ;
        RECT 64.420 156.135 64.770 156.785 ;
        RECT 64.960 156.345 65.365 156.855 ;
        RECT 65.535 156.515 66.675 156.685 ;
        RECT 64.960 156.175 65.715 156.345 ;
        RECT 64.020 155.795 64.685 155.965 ;
        RECT 64.015 155.125 64.345 155.625 ;
        RECT 64.515 155.295 64.685 155.795 ;
        RECT 65.000 155.125 65.285 155.995 ;
        RECT 65.455 155.925 65.715 156.175 ;
        RECT 66.505 156.265 66.675 156.515 ;
        RECT 66.845 156.435 67.195 157.005 ;
        RECT 67.365 156.265 67.535 157.175 ;
        RECT 67.795 157.125 67.965 157.415 ;
        RECT 68.135 157.295 68.465 157.675 ;
        RECT 67.795 156.955 68.460 157.125 ;
        RECT 66.505 156.095 67.535 156.265 ;
        RECT 67.710 156.135 68.060 156.785 ;
        RECT 65.455 155.755 66.575 155.925 ;
        RECT 65.455 155.295 65.715 155.755 ;
        RECT 65.890 155.125 66.145 155.585 ;
        RECT 66.315 155.295 66.575 155.755 ;
        RECT 66.745 155.125 67.055 155.925 ;
        RECT 67.225 155.295 67.535 156.095 ;
        RECT 68.230 155.965 68.460 156.955 ;
        RECT 67.795 155.795 68.460 155.965 ;
        RECT 67.795 155.295 67.965 155.795 ;
        RECT 68.135 155.125 68.465 155.625 ;
        RECT 68.635 155.295 68.820 157.415 ;
        RECT 69.075 157.215 69.325 157.675 ;
        RECT 69.495 157.225 69.830 157.395 ;
        RECT 70.025 157.225 70.700 157.395 ;
        RECT 69.495 157.085 69.665 157.225 ;
        RECT 68.990 156.095 69.270 157.045 ;
        RECT 69.440 156.955 69.665 157.085 ;
        RECT 69.440 155.850 69.610 156.955 ;
        RECT 69.835 156.805 70.360 157.025 ;
        RECT 69.780 156.040 70.020 156.635 ;
        RECT 70.190 156.105 70.360 156.805 ;
        RECT 70.530 156.445 70.700 157.225 ;
        RECT 71.020 157.175 71.390 157.675 ;
        RECT 71.570 157.225 71.975 157.395 ;
        RECT 72.145 157.225 72.930 157.395 ;
        RECT 71.570 156.995 71.740 157.225 ;
        RECT 70.910 156.695 71.740 156.995 ;
        RECT 72.125 156.725 72.590 157.055 ;
        RECT 70.910 156.665 71.110 156.695 ;
        RECT 71.230 156.445 71.400 156.515 ;
        RECT 70.530 156.275 71.400 156.445 ;
        RECT 70.890 156.185 71.400 156.275 ;
        RECT 69.440 155.720 69.745 155.850 ;
        RECT 70.190 155.740 70.720 156.105 ;
        RECT 69.060 155.125 69.325 155.585 ;
        RECT 69.495 155.295 69.745 155.720 ;
        RECT 70.890 155.570 71.060 156.185 ;
        RECT 69.955 155.400 71.060 155.570 ;
        RECT 71.230 155.125 71.400 155.925 ;
        RECT 71.570 155.625 71.740 156.695 ;
        RECT 71.910 155.795 72.100 156.515 ;
        RECT 72.270 155.765 72.590 156.725 ;
        RECT 72.760 156.765 72.930 157.225 ;
        RECT 73.205 157.145 73.415 157.675 ;
        RECT 73.675 156.935 74.005 157.460 ;
        RECT 74.175 157.065 74.345 157.675 ;
        RECT 74.515 157.020 74.845 157.455 ;
        RECT 75.230 157.165 75.470 157.675 ;
        RECT 75.650 157.165 75.930 157.495 ;
        RECT 76.160 157.165 76.375 157.675 ;
        RECT 74.515 156.935 74.895 157.020 ;
        RECT 73.805 156.765 74.005 156.935 ;
        RECT 74.670 156.895 74.895 156.935 ;
        RECT 72.760 156.435 73.635 156.765 ;
        RECT 73.805 156.435 74.555 156.765 ;
        RECT 71.570 155.295 71.820 155.625 ;
        RECT 72.760 155.595 72.930 156.435 ;
        RECT 73.805 156.230 73.995 156.435 ;
        RECT 74.725 156.315 74.895 156.895 ;
        RECT 75.125 156.435 75.480 156.995 ;
        RECT 74.680 156.265 74.895 156.315 ;
        RECT 75.650 156.265 75.820 157.165 ;
        RECT 75.990 156.435 76.255 156.995 ;
        RECT 76.545 156.935 77.160 157.505 ;
        RECT 76.505 156.265 76.675 156.765 ;
        RECT 73.100 155.855 73.995 156.230 ;
        RECT 74.505 156.185 74.895 156.265 ;
        RECT 72.045 155.425 72.930 155.595 ;
        RECT 73.110 155.125 73.425 155.625 ;
        RECT 73.655 155.295 73.995 155.855 ;
        RECT 74.165 155.125 74.335 156.135 ;
        RECT 74.505 155.340 74.835 156.185 ;
        RECT 75.250 156.095 76.675 156.265 ;
        RECT 75.250 155.920 75.640 156.095 ;
        RECT 76.125 155.125 76.455 155.925 ;
        RECT 76.845 155.915 77.160 156.935 ;
        RECT 76.625 155.295 77.160 155.915 ;
        RECT 77.365 156.935 77.625 157.505 ;
        RECT 77.795 157.275 78.180 157.675 ;
        RECT 78.350 157.105 78.605 157.505 ;
        RECT 77.795 156.935 78.605 157.105 ;
        RECT 78.795 156.935 79.040 157.505 ;
        RECT 79.210 157.275 79.595 157.675 ;
        RECT 79.765 157.105 80.020 157.505 ;
        RECT 79.210 156.935 80.020 157.105 ;
        RECT 80.210 156.935 80.635 157.505 ;
        RECT 80.805 157.275 81.190 157.675 ;
        RECT 81.360 157.105 81.795 157.505 ;
        RECT 80.805 156.935 81.795 157.105 ;
        RECT 77.365 156.265 77.550 156.935 ;
        RECT 77.795 156.765 78.145 156.935 ;
        RECT 78.795 156.765 78.965 156.935 ;
        RECT 79.210 156.765 79.560 156.935 ;
        RECT 80.210 156.765 80.560 156.935 ;
        RECT 80.805 156.765 81.140 156.935 ;
        RECT 81.965 156.925 83.175 157.675 ;
        RECT 77.720 156.435 78.145 156.765 ;
        RECT 77.365 155.295 77.625 156.265 ;
        RECT 77.795 155.915 78.145 156.435 ;
        RECT 78.315 156.265 78.965 156.765 ;
        RECT 79.135 156.435 79.560 156.765 ;
        RECT 78.315 156.085 79.040 156.265 ;
        RECT 77.795 155.720 78.605 155.915 ;
        RECT 77.795 155.125 78.180 155.550 ;
        RECT 78.350 155.295 78.605 155.720 ;
        RECT 78.795 155.295 79.040 156.085 ;
        RECT 79.210 155.915 79.560 156.435 ;
        RECT 79.730 156.265 80.560 156.765 ;
        RECT 80.730 156.435 81.140 156.765 ;
        RECT 79.730 156.085 80.635 156.265 ;
        RECT 79.210 155.720 80.040 155.915 ;
        RECT 79.210 155.125 79.595 155.550 ;
        RECT 79.765 155.295 80.040 155.720 ;
        RECT 80.210 155.295 80.635 156.085 ;
        RECT 80.805 155.890 81.140 156.435 ;
        RECT 81.310 156.060 81.795 156.765 ;
        RECT 81.965 156.215 82.485 156.755 ;
        RECT 82.655 156.385 83.175 156.925 ;
        RECT 80.805 155.720 81.795 155.890 ;
        RECT 80.805 155.125 81.190 155.550 ;
        RECT 81.360 155.295 81.795 155.720 ;
        RECT 81.965 155.125 83.175 156.215 ;
        RECT 5.520 154.955 83.260 155.125 ;
        RECT 5.605 153.865 6.815 154.955 ;
        RECT 6.985 154.520 12.330 154.955 ;
        RECT 12.505 154.520 17.850 154.955 ;
        RECT 5.605 153.155 6.125 153.695 ;
        RECT 6.295 153.325 6.815 153.865 ;
        RECT 5.605 152.405 6.815 153.155 ;
        RECT 8.570 152.950 8.910 153.780 ;
        RECT 10.390 153.270 10.740 154.520 ;
        RECT 14.090 152.950 14.430 153.780 ;
        RECT 15.910 153.270 16.260 154.520 ;
        RECT 18.485 153.790 18.775 154.955 ;
        RECT 18.945 154.520 24.290 154.955 ;
        RECT 24.465 154.520 29.810 154.955 ;
        RECT 6.985 152.405 12.330 152.950 ;
        RECT 12.505 152.405 17.850 152.950 ;
        RECT 18.485 152.405 18.775 153.130 ;
        RECT 20.530 152.950 20.870 153.780 ;
        RECT 22.350 153.270 22.700 154.520 ;
        RECT 26.050 152.950 26.390 153.780 ;
        RECT 27.870 153.270 28.220 154.520 ;
        RECT 30.505 153.895 30.835 154.740 ;
        RECT 31.005 153.945 31.175 154.955 ;
        RECT 31.345 154.225 31.685 154.785 ;
        RECT 31.915 154.455 32.230 154.955 ;
        RECT 32.410 154.485 33.295 154.655 ;
        RECT 30.445 153.815 30.835 153.895 ;
        RECT 31.345 153.850 32.240 154.225 ;
        RECT 30.445 153.765 30.660 153.815 ;
        RECT 30.445 153.185 30.615 153.765 ;
        RECT 31.345 153.645 31.535 153.850 ;
        RECT 32.410 153.645 32.580 154.485 ;
        RECT 33.520 154.455 33.770 154.785 ;
        RECT 30.785 153.315 31.535 153.645 ;
        RECT 31.705 153.315 32.580 153.645 ;
        RECT 30.445 153.145 30.670 153.185 ;
        RECT 31.335 153.145 31.535 153.315 ;
        RECT 30.445 153.060 30.825 153.145 ;
        RECT 18.945 152.405 24.290 152.950 ;
        RECT 24.465 152.405 29.810 152.950 ;
        RECT 30.495 152.625 30.825 153.060 ;
        RECT 30.995 152.405 31.165 153.015 ;
        RECT 31.335 152.620 31.665 153.145 ;
        RECT 31.925 152.405 32.135 152.935 ;
        RECT 32.410 152.855 32.580 153.315 ;
        RECT 32.750 153.355 33.070 154.315 ;
        RECT 33.240 153.565 33.430 154.285 ;
        RECT 33.600 153.385 33.770 154.455 ;
        RECT 33.940 154.155 34.110 154.955 ;
        RECT 34.280 154.510 35.385 154.680 ;
        RECT 34.280 153.895 34.450 154.510 ;
        RECT 35.595 154.360 35.845 154.785 ;
        RECT 36.015 154.495 36.280 154.955 ;
        RECT 34.620 153.975 35.150 154.340 ;
        RECT 35.595 154.230 35.900 154.360 ;
        RECT 33.940 153.805 34.450 153.895 ;
        RECT 33.940 153.635 34.810 153.805 ;
        RECT 33.940 153.565 34.110 153.635 ;
        RECT 34.230 153.385 34.430 153.415 ;
        RECT 32.750 153.025 33.215 153.355 ;
        RECT 33.600 153.085 34.430 153.385 ;
        RECT 33.600 152.855 33.770 153.085 ;
        RECT 32.410 152.685 33.195 152.855 ;
        RECT 33.365 152.685 33.770 152.855 ;
        RECT 33.950 152.405 34.320 152.905 ;
        RECT 34.640 152.855 34.810 153.635 ;
        RECT 34.980 153.275 35.150 153.975 ;
        RECT 35.320 153.445 35.560 154.040 ;
        RECT 34.980 153.055 35.505 153.275 ;
        RECT 35.730 153.125 35.900 154.230 ;
        RECT 35.675 152.995 35.900 153.125 ;
        RECT 36.070 153.035 36.350 153.985 ;
        RECT 35.675 152.855 35.845 152.995 ;
        RECT 34.640 152.685 35.315 152.855 ;
        RECT 35.510 152.685 35.845 152.855 ;
        RECT 36.015 152.405 36.265 152.865 ;
        RECT 36.520 152.665 36.705 154.785 ;
        RECT 36.875 154.455 37.205 154.955 ;
        RECT 37.375 154.285 37.545 154.785 ;
        RECT 38.005 154.285 38.285 154.955 ;
        RECT 36.880 154.115 37.545 154.285 ;
        RECT 36.880 153.125 37.110 154.115 ;
        RECT 38.455 154.065 38.755 154.615 ;
        RECT 38.955 154.235 39.285 154.955 ;
        RECT 39.475 154.235 39.935 154.785 ;
        RECT 37.280 153.295 37.630 153.945 ;
        RECT 37.820 153.645 38.085 154.005 ;
        RECT 38.455 153.895 39.395 154.065 ;
        RECT 39.225 153.645 39.395 153.895 ;
        RECT 37.820 153.395 38.495 153.645 ;
        RECT 38.715 153.395 39.055 153.645 ;
        RECT 39.225 153.315 39.515 153.645 ;
        RECT 39.225 153.225 39.395 153.315 ;
        RECT 36.880 152.955 37.545 153.125 ;
        RECT 36.875 152.405 37.205 152.785 ;
        RECT 37.375 152.665 37.545 152.955 ;
        RECT 38.005 153.035 39.395 153.225 ;
        RECT 38.005 152.675 38.335 153.035 ;
        RECT 39.685 152.865 39.935 154.235 ;
        RECT 38.955 152.405 39.205 152.865 ;
        RECT 39.375 152.575 39.935 152.865 ;
        RECT 40.105 153.815 40.490 154.775 ;
        RECT 40.705 154.155 40.995 154.955 ;
        RECT 41.165 154.615 42.530 154.785 ;
        RECT 41.165 153.985 41.335 154.615 ;
        RECT 40.660 153.815 41.335 153.985 ;
        RECT 40.105 153.145 40.280 153.815 ;
        RECT 40.660 153.645 40.830 153.815 ;
        RECT 41.505 153.645 41.830 154.445 ;
        RECT 42.200 154.405 42.530 154.615 ;
        RECT 42.200 154.155 43.155 154.405 ;
        RECT 40.465 153.395 40.830 153.645 ;
        RECT 41.025 153.395 41.275 153.645 ;
        RECT 40.465 153.315 40.655 153.395 ;
        RECT 41.025 153.315 41.195 153.395 ;
        RECT 41.485 153.315 41.830 153.645 ;
        RECT 42.000 153.315 42.275 153.980 ;
        RECT 42.460 153.315 42.815 153.980 ;
        RECT 42.985 153.145 43.155 154.155 ;
        RECT 43.325 153.815 43.615 154.955 ;
        RECT 44.245 153.790 44.535 154.955 ;
        RECT 44.710 154.005 44.975 154.775 ;
        RECT 45.145 154.235 45.475 154.955 ;
        RECT 45.665 154.415 45.925 154.775 ;
        RECT 46.095 154.585 46.425 154.955 ;
        RECT 46.595 154.415 46.855 154.775 ;
        RECT 45.665 154.185 46.855 154.415 ;
        RECT 47.425 154.005 47.715 154.775 ;
        RECT 43.340 153.315 43.615 153.645 ;
        RECT 40.105 152.575 40.615 153.145 ;
        RECT 41.160 152.975 42.560 153.145 ;
        RECT 40.785 152.405 40.955 152.965 ;
        RECT 41.160 152.575 41.490 152.975 ;
        RECT 41.665 152.405 41.995 152.805 ;
        RECT 42.230 152.785 42.560 152.975 ;
        RECT 42.730 152.955 43.155 153.145 ;
        RECT 43.325 152.785 43.615 153.055 ;
        RECT 42.230 152.575 43.615 152.785 ;
        RECT 44.245 152.405 44.535 153.130 ;
        RECT 44.710 152.585 45.045 154.005 ;
        RECT 45.220 153.825 47.715 154.005 ;
        RECT 45.220 153.135 45.445 153.825 ;
        RECT 47.925 153.815 48.195 154.785 ;
        RECT 48.405 154.155 48.685 154.955 ;
        RECT 48.855 154.445 50.510 154.735 ;
        RECT 48.920 154.105 50.510 154.275 ;
        RECT 48.920 153.985 49.090 154.105 ;
        RECT 48.365 153.815 49.090 153.985 ;
        RECT 45.645 153.315 45.925 153.645 ;
        RECT 46.105 153.315 46.680 153.645 ;
        RECT 46.860 153.315 47.295 153.645 ;
        RECT 47.475 153.315 47.745 153.645 ;
        RECT 45.220 152.945 47.705 153.135 ;
        RECT 45.225 152.405 45.970 152.775 ;
        RECT 46.535 152.585 46.790 152.945 ;
        RECT 46.970 152.405 47.300 152.775 ;
        RECT 47.480 152.585 47.705 152.945 ;
        RECT 47.925 153.080 48.095 153.815 ;
        RECT 48.365 153.645 48.535 153.815 ;
        RECT 49.280 153.765 49.995 153.935 ;
        RECT 50.190 153.815 50.510 154.105 ;
        RECT 50.690 153.815 51.025 154.785 ;
        RECT 51.195 153.815 51.365 154.955 ;
        RECT 51.535 154.615 53.565 154.785 ;
        RECT 48.265 153.315 48.535 153.645 ;
        RECT 48.705 153.315 49.110 153.645 ;
        RECT 49.280 153.315 49.990 153.765 ;
        RECT 48.365 153.145 48.535 153.315 ;
        RECT 47.925 152.735 48.195 153.080 ;
        RECT 48.365 152.975 49.975 153.145 ;
        RECT 50.160 153.075 50.510 153.645 ;
        RECT 50.690 153.145 50.860 153.815 ;
        RECT 51.535 153.645 51.705 154.615 ;
        RECT 51.030 153.315 51.285 153.645 ;
        RECT 51.510 153.315 51.705 153.645 ;
        RECT 51.875 154.275 53.000 154.445 ;
        RECT 51.115 153.145 51.285 153.315 ;
        RECT 51.875 153.145 52.045 154.275 ;
        RECT 48.385 152.405 48.765 152.805 ;
        RECT 48.935 152.625 49.105 152.975 ;
        RECT 49.275 152.405 49.605 152.805 ;
        RECT 49.805 152.625 49.975 152.975 ;
        RECT 50.175 152.405 50.505 152.905 ;
        RECT 50.690 152.575 50.945 153.145 ;
        RECT 51.115 152.975 52.045 153.145 ;
        RECT 52.215 153.935 53.225 154.105 ;
        RECT 52.215 153.135 52.385 153.935 ;
        RECT 52.590 153.595 52.865 153.735 ;
        RECT 52.585 153.425 52.865 153.595 ;
        RECT 51.870 152.940 52.045 152.975 ;
        RECT 51.115 152.405 51.445 152.805 ;
        RECT 51.870 152.575 52.400 152.940 ;
        RECT 52.590 152.575 52.865 153.425 ;
        RECT 53.035 152.575 53.225 153.935 ;
        RECT 53.395 153.950 53.565 154.615 ;
        RECT 53.735 154.195 53.905 154.955 ;
        RECT 54.140 154.195 54.655 154.605 ;
        RECT 53.395 153.760 54.145 153.950 ;
        RECT 54.315 153.385 54.655 154.195 ;
        RECT 54.915 154.285 55.085 154.785 ;
        RECT 55.255 154.455 55.585 154.955 ;
        RECT 54.915 154.115 55.580 154.285 ;
        RECT 53.425 153.215 54.655 153.385 ;
        RECT 54.830 153.295 55.180 153.945 ;
        RECT 53.405 152.405 53.915 152.940 ;
        RECT 54.135 152.610 54.380 153.215 ;
        RECT 55.350 153.125 55.580 154.115 ;
        RECT 54.915 152.955 55.580 153.125 ;
        RECT 54.915 152.665 55.085 152.955 ;
        RECT 55.255 152.405 55.585 152.785 ;
        RECT 55.755 152.665 55.940 154.785 ;
        RECT 56.180 154.495 56.445 154.955 ;
        RECT 56.615 154.360 56.865 154.785 ;
        RECT 57.075 154.510 58.180 154.680 ;
        RECT 56.560 154.230 56.865 154.360 ;
        RECT 56.110 153.035 56.390 153.985 ;
        RECT 56.560 153.125 56.730 154.230 ;
        RECT 56.900 153.445 57.140 154.040 ;
        RECT 57.310 153.975 57.840 154.340 ;
        RECT 57.310 153.275 57.480 153.975 ;
        RECT 58.010 153.895 58.180 154.510 ;
        RECT 58.350 154.155 58.520 154.955 ;
        RECT 58.690 154.455 58.940 154.785 ;
        RECT 59.165 154.485 60.050 154.655 ;
        RECT 58.010 153.805 58.520 153.895 ;
        RECT 56.560 152.995 56.785 153.125 ;
        RECT 56.955 153.055 57.480 153.275 ;
        RECT 57.650 153.635 58.520 153.805 ;
        RECT 56.195 152.405 56.445 152.865 ;
        RECT 56.615 152.855 56.785 152.995 ;
        RECT 57.650 152.855 57.820 153.635 ;
        RECT 58.350 153.565 58.520 153.635 ;
        RECT 58.030 153.385 58.230 153.415 ;
        RECT 58.690 153.385 58.860 154.455 ;
        RECT 59.030 153.565 59.220 154.285 ;
        RECT 58.030 153.085 58.860 153.385 ;
        RECT 59.390 153.355 59.710 154.315 ;
        RECT 56.615 152.685 56.950 152.855 ;
        RECT 57.145 152.685 57.820 152.855 ;
        RECT 58.140 152.405 58.510 152.905 ;
        RECT 58.690 152.855 58.860 153.085 ;
        RECT 59.245 153.025 59.710 153.355 ;
        RECT 59.880 153.645 60.050 154.485 ;
        RECT 60.230 154.455 60.545 154.955 ;
        RECT 60.775 154.225 61.115 154.785 ;
        RECT 60.220 153.850 61.115 154.225 ;
        RECT 61.285 153.945 61.455 154.955 ;
        RECT 60.925 153.645 61.115 153.850 ;
        RECT 61.625 153.895 61.955 154.740 ;
        RECT 61.625 153.815 62.015 153.895 ;
        RECT 61.800 153.765 62.015 153.815 ;
        RECT 59.880 153.315 60.755 153.645 ;
        RECT 60.925 153.315 61.675 153.645 ;
        RECT 59.880 152.855 60.050 153.315 ;
        RECT 60.925 153.145 61.125 153.315 ;
        RECT 61.845 153.185 62.015 153.765 ;
        RECT 61.790 153.145 62.015 153.185 ;
        RECT 58.690 152.685 59.095 152.855 ;
        RECT 59.265 152.685 60.050 152.855 ;
        RECT 60.325 152.405 60.535 152.935 ;
        RECT 60.795 152.620 61.125 153.145 ;
        RECT 61.635 153.060 62.015 153.145 ;
        RECT 62.190 153.815 62.525 154.785 ;
        RECT 62.695 153.815 62.865 154.955 ;
        RECT 63.035 154.615 65.065 154.785 ;
        RECT 62.190 153.145 62.360 153.815 ;
        RECT 63.035 153.645 63.205 154.615 ;
        RECT 62.530 153.315 62.785 153.645 ;
        RECT 63.010 153.315 63.205 153.645 ;
        RECT 63.375 154.275 64.500 154.445 ;
        RECT 62.615 153.145 62.785 153.315 ;
        RECT 63.375 153.145 63.545 154.275 ;
        RECT 61.295 152.405 61.465 153.015 ;
        RECT 61.635 152.625 61.965 153.060 ;
        RECT 62.190 152.575 62.445 153.145 ;
        RECT 62.615 152.975 63.545 153.145 ;
        RECT 63.715 153.935 64.725 154.105 ;
        RECT 63.715 153.135 63.885 153.935 ;
        RECT 64.090 153.255 64.365 153.735 ;
        RECT 64.085 153.085 64.365 153.255 ;
        RECT 63.370 152.940 63.545 152.975 ;
        RECT 62.615 152.405 62.945 152.805 ;
        RECT 63.370 152.575 63.900 152.940 ;
        RECT 64.090 152.575 64.365 153.085 ;
        RECT 64.535 152.575 64.725 153.935 ;
        RECT 64.895 153.950 65.065 154.615 ;
        RECT 65.235 154.195 65.405 154.955 ;
        RECT 65.640 154.195 66.155 154.605 ;
        RECT 64.895 153.760 65.645 153.950 ;
        RECT 65.815 153.385 66.155 154.195 ;
        RECT 64.925 153.215 66.155 153.385 ;
        RECT 66.325 153.815 66.710 154.785 ;
        RECT 66.880 154.495 67.205 154.955 ;
        RECT 67.725 154.325 68.005 154.785 ;
        RECT 66.880 154.105 68.005 154.325 ;
        RECT 64.905 152.405 65.415 152.940 ;
        RECT 65.635 152.610 65.880 153.215 ;
        RECT 66.325 153.145 66.605 153.815 ;
        RECT 66.880 153.645 67.330 154.105 ;
        RECT 68.195 153.935 68.595 154.785 ;
        RECT 68.995 154.495 69.265 154.955 ;
        RECT 69.435 154.325 69.720 154.785 ;
        RECT 66.775 153.315 67.330 153.645 ;
        RECT 67.500 153.375 68.595 153.935 ;
        RECT 66.880 153.205 67.330 153.315 ;
        RECT 66.325 152.575 66.710 153.145 ;
        RECT 66.880 153.035 68.005 153.205 ;
        RECT 66.880 152.405 67.205 152.865 ;
        RECT 67.725 152.575 68.005 153.035 ;
        RECT 68.195 152.575 68.595 153.375 ;
        RECT 68.765 154.105 69.720 154.325 ;
        RECT 68.765 153.205 68.975 154.105 ;
        RECT 69.145 153.375 69.835 153.935 ;
        RECT 70.005 153.790 70.295 154.955 ;
        RECT 70.465 153.815 70.805 154.785 ;
        RECT 70.975 153.815 71.145 154.955 ;
        RECT 71.415 154.155 71.665 154.955 ;
        RECT 72.310 153.985 72.640 154.785 ;
        RECT 72.940 154.155 73.270 154.955 ;
        RECT 73.440 153.985 73.770 154.785 ;
        RECT 74.695 154.285 74.865 154.785 ;
        RECT 75.035 154.455 75.365 154.955 ;
        RECT 74.695 154.115 75.360 154.285 ;
        RECT 71.335 153.815 73.770 153.985 ;
        RECT 70.465 153.255 70.640 153.815 ;
        RECT 71.335 153.565 71.505 153.815 ;
        RECT 70.810 153.395 71.505 153.565 ;
        RECT 71.680 153.395 72.100 153.595 ;
        RECT 72.270 153.395 72.600 153.595 ;
        RECT 72.770 153.395 73.100 153.595 ;
        RECT 70.465 153.205 70.695 153.255 ;
        RECT 68.765 153.035 69.720 153.205 ;
        RECT 68.995 152.405 69.265 152.865 ;
        RECT 69.435 152.575 69.720 153.035 ;
        RECT 70.005 152.405 70.295 153.130 ;
        RECT 70.465 152.575 70.805 153.205 ;
        RECT 70.975 152.405 71.225 153.205 ;
        RECT 71.415 153.055 72.640 153.225 ;
        RECT 71.415 152.575 71.745 153.055 ;
        RECT 71.915 152.405 72.140 152.865 ;
        RECT 72.310 152.575 72.640 153.055 ;
        RECT 73.270 153.185 73.440 153.815 ;
        RECT 73.625 153.395 73.975 153.645 ;
        RECT 74.610 153.295 74.960 153.945 ;
        RECT 73.270 152.575 73.770 153.185 ;
        RECT 75.130 153.125 75.360 154.115 ;
        RECT 74.695 152.955 75.360 153.125 ;
        RECT 74.695 152.665 74.865 152.955 ;
        RECT 75.035 152.405 75.365 152.785 ;
        RECT 75.535 152.665 75.720 154.785 ;
        RECT 75.960 154.495 76.225 154.955 ;
        RECT 76.395 154.360 76.645 154.785 ;
        RECT 76.855 154.510 77.960 154.680 ;
        RECT 76.340 154.230 76.645 154.360 ;
        RECT 75.890 153.035 76.170 153.985 ;
        RECT 76.340 153.125 76.510 154.230 ;
        RECT 76.680 153.445 76.920 154.040 ;
        RECT 77.090 153.975 77.620 154.340 ;
        RECT 77.090 153.275 77.260 153.975 ;
        RECT 77.790 153.895 77.960 154.510 ;
        RECT 78.130 154.155 78.300 154.955 ;
        RECT 78.470 154.455 78.720 154.785 ;
        RECT 78.945 154.485 79.830 154.655 ;
        RECT 77.790 153.805 78.300 153.895 ;
        RECT 76.340 152.995 76.565 153.125 ;
        RECT 76.735 153.055 77.260 153.275 ;
        RECT 77.430 153.635 78.300 153.805 ;
        RECT 75.975 152.405 76.225 152.865 ;
        RECT 76.395 152.855 76.565 152.995 ;
        RECT 77.430 152.855 77.600 153.635 ;
        RECT 78.130 153.565 78.300 153.635 ;
        RECT 77.810 153.385 78.010 153.415 ;
        RECT 78.470 153.385 78.640 154.455 ;
        RECT 78.810 153.565 79.000 154.285 ;
        RECT 77.810 153.085 78.640 153.385 ;
        RECT 79.170 153.355 79.490 154.315 ;
        RECT 76.395 152.685 76.730 152.855 ;
        RECT 76.925 152.685 77.600 152.855 ;
        RECT 77.920 152.405 78.290 152.905 ;
        RECT 78.470 152.855 78.640 153.085 ;
        RECT 79.025 153.025 79.490 153.355 ;
        RECT 79.660 153.645 79.830 154.485 ;
        RECT 80.010 154.455 80.325 154.955 ;
        RECT 80.555 154.225 80.895 154.785 ;
        RECT 80.000 153.850 80.895 154.225 ;
        RECT 81.065 153.945 81.235 154.955 ;
        RECT 80.705 153.645 80.895 153.850 ;
        RECT 81.405 153.895 81.735 154.740 ;
        RECT 81.405 153.815 81.795 153.895 ;
        RECT 81.580 153.765 81.795 153.815 ;
        RECT 79.660 153.315 80.535 153.645 ;
        RECT 80.705 153.315 81.455 153.645 ;
        RECT 79.660 152.855 79.830 153.315 ;
        RECT 80.705 153.145 80.905 153.315 ;
        RECT 81.625 153.185 81.795 153.765 ;
        RECT 81.965 153.865 83.175 154.955 ;
        RECT 81.965 153.325 82.485 153.865 ;
        RECT 81.570 153.145 81.795 153.185 ;
        RECT 82.655 153.155 83.175 153.695 ;
        RECT 78.470 152.685 78.875 152.855 ;
        RECT 79.045 152.685 79.830 152.855 ;
        RECT 80.105 152.405 80.315 152.935 ;
        RECT 80.575 152.620 80.905 153.145 ;
        RECT 81.415 153.060 81.795 153.145 ;
        RECT 81.075 152.405 81.245 153.015 ;
        RECT 81.415 152.625 81.745 153.060 ;
        RECT 81.965 152.405 83.175 153.155 ;
        RECT 5.520 152.235 83.260 152.405 ;
        RECT 5.605 151.485 6.815 152.235 ;
        RECT 6.985 151.690 12.330 152.235 ;
        RECT 12.505 151.690 17.850 152.235 ;
        RECT 18.025 151.690 23.370 152.235 ;
        RECT 5.605 150.945 6.125 151.485 ;
        RECT 6.295 150.775 6.815 151.315 ;
        RECT 8.570 150.860 8.910 151.690 ;
        RECT 5.605 149.685 6.815 150.775 ;
        RECT 10.390 150.120 10.740 151.370 ;
        RECT 14.090 150.860 14.430 151.690 ;
        RECT 15.910 150.120 16.260 151.370 ;
        RECT 19.610 150.860 19.950 151.690 ;
        RECT 23.545 151.465 27.055 152.235 ;
        RECT 21.430 150.120 21.780 151.370 ;
        RECT 23.545 150.945 25.195 151.465 ;
        RECT 27.225 151.435 27.535 152.235 ;
        RECT 27.740 151.435 28.435 152.065 ;
        RECT 25.365 150.775 27.055 151.295 ;
        RECT 27.235 150.995 27.570 151.265 ;
        RECT 27.740 150.835 27.910 151.435 ;
        RECT 28.080 150.995 28.415 151.245 ;
        RECT 6.985 149.685 12.330 150.120 ;
        RECT 12.505 149.685 17.850 150.120 ;
        RECT 18.025 149.685 23.370 150.120 ;
        RECT 23.545 149.685 27.055 150.775 ;
        RECT 27.225 149.685 27.505 150.825 ;
        RECT 27.675 149.855 28.005 150.835 ;
        RECT 28.175 149.685 28.435 150.825 ;
        RECT 28.615 149.865 28.875 152.055 ;
        RECT 29.135 151.865 29.805 152.235 ;
        RECT 29.985 151.685 30.295 152.055 ;
        RECT 29.065 151.485 30.295 151.685 ;
        RECT 29.065 150.815 29.355 151.485 ;
        RECT 30.475 151.305 30.705 151.945 ;
        RECT 30.885 151.505 31.175 152.235 ;
        RECT 31.365 151.510 31.655 152.235 ;
        RECT 31.915 151.685 32.085 151.975 ;
        RECT 32.255 151.855 32.585 152.235 ;
        RECT 31.915 151.515 32.580 151.685 ;
        RECT 29.535 150.995 30.000 151.305 ;
        RECT 30.180 150.995 30.705 151.305 ;
        RECT 30.885 150.995 31.185 151.325 ;
        RECT 29.065 150.595 29.835 150.815 ;
        RECT 29.045 149.685 29.385 150.415 ;
        RECT 29.565 149.865 29.835 150.595 ;
        RECT 30.015 150.575 31.175 150.815 ;
        RECT 30.015 149.865 30.245 150.575 ;
        RECT 30.415 149.685 30.745 150.395 ;
        RECT 30.915 149.865 31.175 150.575 ;
        RECT 31.365 149.685 31.655 150.850 ;
        RECT 31.830 150.695 32.180 151.345 ;
        RECT 32.350 150.525 32.580 151.515 ;
        RECT 31.915 150.355 32.580 150.525 ;
        RECT 31.915 149.855 32.085 150.355 ;
        RECT 32.255 149.685 32.585 150.185 ;
        RECT 32.755 149.855 32.940 151.975 ;
        RECT 33.195 151.775 33.445 152.235 ;
        RECT 33.615 151.785 33.950 151.955 ;
        RECT 34.145 151.785 34.820 151.955 ;
        RECT 33.615 151.645 33.785 151.785 ;
        RECT 33.110 150.655 33.390 151.605 ;
        RECT 33.560 151.515 33.785 151.645 ;
        RECT 33.560 150.410 33.730 151.515 ;
        RECT 33.955 151.365 34.480 151.585 ;
        RECT 33.900 150.600 34.140 151.195 ;
        RECT 34.310 150.665 34.480 151.365 ;
        RECT 34.650 151.005 34.820 151.785 ;
        RECT 35.140 151.735 35.510 152.235 ;
        RECT 35.690 151.785 36.095 151.955 ;
        RECT 36.265 151.785 37.050 151.955 ;
        RECT 35.690 151.555 35.860 151.785 ;
        RECT 35.030 151.255 35.860 151.555 ;
        RECT 36.245 151.285 36.710 151.615 ;
        RECT 35.030 151.225 35.230 151.255 ;
        RECT 35.350 151.005 35.520 151.075 ;
        RECT 34.650 150.835 35.520 151.005 ;
        RECT 35.010 150.745 35.520 150.835 ;
        RECT 33.560 150.280 33.865 150.410 ;
        RECT 34.310 150.300 34.840 150.665 ;
        RECT 33.180 149.685 33.445 150.145 ;
        RECT 33.615 149.855 33.865 150.280 ;
        RECT 35.010 150.130 35.180 150.745 ;
        RECT 34.075 149.960 35.180 150.130 ;
        RECT 35.350 149.685 35.520 150.485 ;
        RECT 35.690 150.185 35.860 151.255 ;
        RECT 36.030 150.355 36.220 151.075 ;
        RECT 36.390 150.325 36.710 151.285 ;
        RECT 36.880 151.325 37.050 151.785 ;
        RECT 37.325 151.705 37.535 152.235 ;
        RECT 37.795 151.495 38.125 152.020 ;
        RECT 38.295 151.625 38.465 152.235 ;
        RECT 38.635 151.580 38.965 152.015 ;
        RECT 39.735 151.685 39.905 151.975 ;
        RECT 40.075 151.855 40.405 152.235 ;
        RECT 38.635 151.495 39.015 151.580 ;
        RECT 39.735 151.515 40.400 151.685 ;
        RECT 37.925 151.325 38.125 151.495 ;
        RECT 38.790 151.455 39.015 151.495 ;
        RECT 36.880 150.995 37.755 151.325 ;
        RECT 37.925 150.995 38.675 151.325 ;
        RECT 35.690 149.855 35.940 150.185 ;
        RECT 36.880 150.155 37.050 150.995 ;
        RECT 37.925 150.790 38.115 150.995 ;
        RECT 38.845 150.875 39.015 151.455 ;
        RECT 38.800 150.825 39.015 150.875 ;
        RECT 37.220 150.415 38.115 150.790 ;
        RECT 38.625 150.745 39.015 150.825 ;
        RECT 36.165 149.985 37.050 150.155 ;
        RECT 37.230 149.685 37.545 150.185 ;
        RECT 37.775 149.855 38.115 150.415 ;
        RECT 38.285 149.685 38.455 150.695 ;
        RECT 38.625 149.900 38.955 150.745 ;
        RECT 39.650 150.695 40.000 151.345 ;
        RECT 40.170 150.525 40.400 151.515 ;
        RECT 39.735 150.355 40.400 150.525 ;
        RECT 39.735 149.855 39.905 150.355 ;
        RECT 40.075 149.685 40.405 150.185 ;
        RECT 40.575 149.855 40.760 151.975 ;
        RECT 41.015 151.775 41.265 152.235 ;
        RECT 41.435 151.785 41.770 151.955 ;
        RECT 41.965 151.785 42.640 151.955 ;
        RECT 41.435 151.645 41.605 151.785 ;
        RECT 40.930 150.655 41.210 151.605 ;
        RECT 41.380 151.515 41.605 151.645 ;
        RECT 41.380 150.410 41.550 151.515 ;
        RECT 41.775 151.365 42.300 151.585 ;
        RECT 41.720 150.600 41.960 151.195 ;
        RECT 42.130 150.665 42.300 151.365 ;
        RECT 42.470 151.005 42.640 151.785 ;
        RECT 42.960 151.735 43.330 152.235 ;
        RECT 43.510 151.785 43.915 151.955 ;
        RECT 44.085 151.785 44.870 151.955 ;
        RECT 43.510 151.555 43.680 151.785 ;
        RECT 42.850 151.255 43.680 151.555 ;
        RECT 44.065 151.285 44.530 151.615 ;
        RECT 42.850 151.225 43.050 151.255 ;
        RECT 43.170 151.005 43.340 151.075 ;
        RECT 42.470 150.835 43.340 151.005 ;
        RECT 42.830 150.745 43.340 150.835 ;
        RECT 41.380 150.280 41.685 150.410 ;
        RECT 42.130 150.300 42.660 150.665 ;
        RECT 41.000 149.685 41.265 150.145 ;
        RECT 41.435 149.855 41.685 150.280 ;
        RECT 42.830 150.130 43.000 150.745 ;
        RECT 41.895 149.960 43.000 150.130 ;
        RECT 43.170 149.685 43.340 150.485 ;
        RECT 43.510 150.185 43.680 151.255 ;
        RECT 43.850 150.355 44.040 151.075 ;
        RECT 44.210 150.325 44.530 151.285 ;
        RECT 44.700 151.325 44.870 151.785 ;
        RECT 45.145 151.705 45.355 152.235 ;
        RECT 45.615 151.495 45.945 152.020 ;
        RECT 46.115 151.625 46.285 152.235 ;
        RECT 46.455 151.580 46.785 152.015 ;
        RECT 47.005 151.735 47.345 152.235 ;
        RECT 46.455 151.495 46.835 151.580 ;
        RECT 45.745 151.325 45.945 151.495 ;
        RECT 46.610 151.455 46.835 151.495 ;
        RECT 44.700 150.995 45.575 151.325 ;
        RECT 45.745 150.995 46.495 151.325 ;
        RECT 43.510 149.855 43.760 150.185 ;
        RECT 44.700 150.155 44.870 150.995 ;
        RECT 45.745 150.790 45.935 150.995 ;
        RECT 46.665 150.875 46.835 151.455 ;
        RECT 47.005 150.995 47.345 151.565 ;
        RECT 47.515 151.325 47.760 152.015 ;
        RECT 47.955 151.735 48.285 152.235 ;
        RECT 48.485 151.665 48.655 152.015 ;
        RECT 48.830 151.835 49.160 152.235 ;
        RECT 49.330 151.665 49.500 152.015 ;
        RECT 49.670 151.835 50.050 152.235 ;
        RECT 48.485 151.495 50.070 151.665 ;
        RECT 50.240 151.560 50.515 151.905 ;
        RECT 49.900 151.325 50.070 151.495 ;
        RECT 47.515 150.995 48.170 151.325 ;
        RECT 46.620 150.825 46.835 150.875 ;
        RECT 45.040 150.415 45.935 150.790 ;
        RECT 46.445 150.745 46.835 150.825 ;
        RECT 43.985 149.985 44.870 150.155 ;
        RECT 45.050 149.685 45.365 150.185 ;
        RECT 45.595 149.855 45.935 150.415 ;
        RECT 46.105 149.685 46.275 150.695 ;
        RECT 46.445 149.900 46.775 150.745 ;
        RECT 47.005 149.685 47.345 150.760 ;
        RECT 47.515 150.400 47.755 150.995 ;
        RECT 47.950 150.535 48.270 150.825 ;
        RECT 48.440 150.705 49.180 151.325 ;
        RECT 49.350 150.995 49.730 151.325 ;
        RECT 49.900 150.995 50.175 151.325 ;
        RECT 49.900 150.825 50.070 150.995 ;
        RECT 50.345 150.825 50.515 151.560 ;
        RECT 49.410 150.655 50.070 150.825 ;
        RECT 49.410 150.535 49.580 150.655 ;
        RECT 47.950 150.365 49.580 150.535 ;
        RECT 47.530 149.905 49.580 150.195 ;
        RECT 49.750 149.685 50.030 150.485 ;
        RECT 50.240 149.855 50.515 150.825 ;
        RECT 50.685 151.585 50.945 152.065 ;
        RECT 51.115 151.775 51.445 152.235 ;
        RECT 51.635 151.595 51.835 152.015 ;
        RECT 50.685 150.555 50.855 151.585 ;
        RECT 51.025 150.895 51.255 151.325 ;
        RECT 51.425 151.075 51.835 151.595 ;
        RECT 52.005 151.750 52.795 152.015 ;
        RECT 52.005 150.895 52.260 151.750 ;
        RECT 52.975 151.415 53.305 151.835 ;
        RECT 53.475 151.415 53.735 152.235 ;
        RECT 53.925 151.545 54.165 152.065 ;
        RECT 54.335 151.740 54.730 152.235 ;
        RECT 55.295 151.905 55.465 152.050 ;
        RECT 55.090 151.710 55.465 151.905 ;
        RECT 52.975 151.325 53.225 151.415 ;
        RECT 52.430 151.075 53.225 151.325 ;
        RECT 51.025 150.725 52.815 150.895 ;
        RECT 50.685 149.855 50.960 150.555 ;
        RECT 51.130 150.430 51.845 150.725 ;
        RECT 52.065 150.365 52.395 150.555 ;
        RECT 51.170 149.685 51.385 150.230 ;
        RECT 51.555 149.855 52.030 150.195 ;
        RECT 52.200 150.190 52.395 150.365 ;
        RECT 52.565 150.360 52.815 150.725 ;
        RECT 52.200 149.685 52.815 150.190 ;
        RECT 53.055 149.855 53.225 151.075 ;
        RECT 53.395 150.365 53.735 151.245 ;
        RECT 53.925 150.875 54.100 151.545 ;
        RECT 55.090 151.375 55.260 151.710 ;
        RECT 55.745 151.665 55.985 152.040 ;
        RECT 56.155 151.730 56.490 152.235 ;
        RECT 55.745 151.515 55.965 151.665 ;
        RECT 54.275 151.015 55.260 151.375 ;
        RECT 55.430 151.185 55.965 151.515 ;
        RECT 54.275 150.995 55.560 151.015 ;
        RECT 53.925 150.740 54.135 150.875 ;
        RECT 54.700 150.845 55.560 150.995 ;
        RECT 53.475 149.685 53.735 150.195 ;
        RECT 53.925 149.955 54.230 150.740 ;
        RECT 54.405 150.365 55.100 150.675 ;
        RECT 54.410 149.685 55.095 150.155 ;
        RECT 55.275 149.900 55.560 150.845 ;
        RECT 55.730 150.535 55.965 151.185 ;
        RECT 56.135 150.705 56.435 151.555 ;
        RECT 57.125 151.510 57.415 152.235 ;
        RECT 57.590 151.495 57.845 152.065 ;
        RECT 58.015 151.835 58.345 152.235 ;
        RECT 58.770 151.700 59.300 152.065 ;
        RECT 59.490 151.895 59.765 152.065 ;
        RECT 59.485 151.725 59.765 151.895 ;
        RECT 58.770 151.665 58.945 151.700 ;
        RECT 58.015 151.495 58.945 151.665 ;
        RECT 55.730 150.305 56.405 150.535 ;
        RECT 55.735 149.685 56.065 150.135 ;
        RECT 56.235 149.875 56.405 150.305 ;
        RECT 57.125 149.685 57.415 150.850 ;
        RECT 57.590 150.825 57.760 151.495 ;
        RECT 58.015 151.325 58.185 151.495 ;
        RECT 57.930 150.995 58.185 151.325 ;
        RECT 58.410 150.995 58.605 151.325 ;
        RECT 57.590 149.855 57.925 150.825 ;
        RECT 58.095 149.685 58.265 150.825 ;
        RECT 58.435 150.025 58.605 150.995 ;
        RECT 58.775 150.365 58.945 151.495 ;
        RECT 59.115 150.705 59.285 151.505 ;
        RECT 59.490 150.905 59.765 151.725 ;
        RECT 59.935 150.705 60.125 152.065 ;
        RECT 60.305 151.700 60.815 152.235 ;
        RECT 61.035 151.425 61.280 152.030 ;
        RECT 61.730 151.495 61.985 152.065 ;
        RECT 62.155 151.835 62.485 152.235 ;
        RECT 62.910 151.700 63.440 152.065 ;
        RECT 63.630 151.895 63.905 152.065 ;
        RECT 63.625 151.725 63.905 151.895 ;
        RECT 62.910 151.665 63.085 151.700 ;
        RECT 62.155 151.495 63.085 151.665 ;
        RECT 60.325 151.255 61.555 151.425 ;
        RECT 59.115 150.535 60.125 150.705 ;
        RECT 60.295 150.690 61.045 150.880 ;
        RECT 58.775 150.195 59.900 150.365 ;
        RECT 60.295 150.025 60.465 150.690 ;
        RECT 61.215 150.445 61.555 151.255 ;
        RECT 58.435 149.855 60.465 150.025 ;
        RECT 60.635 149.685 60.805 150.445 ;
        RECT 61.040 150.035 61.555 150.445 ;
        RECT 61.730 150.825 61.900 151.495 ;
        RECT 62.155 151.325 62.325 151.495 ;
        RECT 62.070 150.995 62.325 151.325 ;
        RECT 62.550 150.995 62.745 151.325 ;
        RECT 61.730 149.855 62.065 150.825 ;
        RECT 62.235 149.685 62.405 150.825 ;
        RECT 62.575 150.025 62.745 150.995 ;
        RECT 62.915 150.365 63.085 151.495 ;
        RECT 63.255 150.705 63.425 151.505 ;
        RECT 63.630 150.905 63.905 151.725 ;
        RECT 64.075 150.705 64.265 152.065 ;
        RECT 64.445 151.700 64.955 152.235 ;
        RECT 65.175 151.425 65.420 152.030 ;
        RECT 65.865 151.495 66.250 152.065 ;
        RECT 66.420 151.775 66.745 152.235 ;
        RECT 67.265 151.605 67.545 152.065 ;
        RECT 64.465 151.255 65.695 151.425 ;
        RECT 63.255 150.535 64.265 150.705 ;
        RECT 64.435 150.690 65.185 150.880 ;
        RECT 62.915 150.195 64.040 150.365 ;
        RECT 64.435 150.025 64.605 150.690 ;
        RECT 65.355 150.445 65.695 151.255 ;
        RECT 62.575 149.855 64.605 150.025 ;
        RECT 64.775 149.685 64.945 150.445 ;
        RECT 65.180 150.035 65.695 150.445 ;
        RECT 65.865 150.825 66.145 151.495 ;
        RECT 66.420 151.435 67.545 151.605 ;
        RECT 66.420 151.325 66.870 151.435 ;
        RECT 66.315 150.995 66.870 151.325 ;
        RECT 67.735 151.265 68.135 152.065 ;
        RECT 68.535 151.775 68.805 152.235 ;
        RECT 68.975 151.605 69.260 152.065 ;
        RECT 65.865 149.855 66.250 150.825 ;
        RECT 66.420 150.535 66.870 150.995 ;
        RECT 67.040 150.705 68.135 151.265 ;
        RECT 66.420 150.315 67.545 150.535 ;
        RECT 66.420 149.685 66.745 150.145 ;
        RECT 67.265 149.855 67.545 150.315 ;
        RECT 67.735 149.855 68.135 150.705 ;
        RECT 68.305 151.435 69.260 151.605 ;
        RECT 69.545 151.435 69.885 152.065 ;
        RECT 70.055 151.435 70.305 152.235 ;
        RECT 70.495 151.585 70.825 152.065 ;
        RECT 70.995 151.775 71.220 152.235 ;
        RECT 71.390 151.585 71.720 152.065 ;
        RECT 68.305 150.535 68.515 151.435 ;
        RECT 69.545 151.385 69.775 151.435 ;
        RECT 70.495 151.415 71.720 151.585 ;
        RECT 72.350 151.455 72.850 152.065 ;
        RECT 73.225 151.560 73.485 152.065 ;
        RECT 73.665 151.855 73.995 152.235 ;
        RECT 74.175 151.685 74.345 152.065 ;
        RECT 68.685 150.705 69.375 151.265 ;
        RECT 69.545 150.825 69.720 151.385 ;
        RECT 69.890 151.075 70.585 151.245 ;
        RECT 70.415 150.825 70.585 151.075 ;
        RECT 70.760 151.045 71.180 151.245 ;
        RECT 71.350 151.045 71.680 151.245 ;
        RECT 71.850 151.045 72.180 151.245 ;
        RECT 72.350 150.825 72.520 151.455 ;
        RECT 72.705 150.995 73.055 151.245 ;
        RECT 68.305 150.315 69.260 150.535 ;
        RECT 68.535 149.685 68.805 150.145 ;
        RECT 68.975 149.855 69.260 150.315 ;
        RECT 69.545 149.855 69.885 150.825 ;
        RECT 70.055 149.685 70.225 150.825 ;
        RECT 70.415 150.655 72.850 150.825 ;
        RECT 70.495 149.685 70.745 150.485 ;
        RECT 71.390 149.855 71.720 150.655 ;
        RECT 72.020 149.685 72.350 150.485 ;
        RECT 72.520 149.855 72.850 150.655 ;
        RECT 73.225 150.760 73.395 151.560 ;
        RECT 73.680 151.515 74.345 151.685 ;
        RECT 74.695 151.685 74.865 151.975 ;
        RECT 75.035 151.855 75.365 152.235 ;
        RECT 74.695 151.515 75.360 151.685 ;
        RECT 73.680 151.260 73.850 151.515 ;
        RECT 73.565 150.930 73.850 151.260 ;
        RECT 74.085 150.965 74.415 151.335 ;
        RECT 73.680 150.785 73.850 150.930 ;
        RECT 73.225 149.855 73.495 150.760 ;
        RECT 73.680 150.615 74.345 150.785 ;
        RECT 74.610 150.695 74.960 151.345 ;
        RECT 73.665 149.685 73.995 150.445 ;
        RECT 74.175 149.855 74.345 150.615 ;
        RECT 75.130 150.525 75.360 151.515 ;
        RECT 74.695 150.355 75.360 150.525 ;
        RECT 74.695 149.855 74.865 150.355 ;
        RECT 75.035 149.685 75.365 150.185 ;
        RECT 75.535 149.855 75.720 151.975 ;
        RECT 75.975 151.775 76.225 152.235 ;
        RECT 76.395 151.785 76.730 151.955 ;
        RECT 76.925 151.785 77.600 151.955 ;
        RECT 76.395 151.645 76.565 151.785 ;
        RECT 75.890 150.655 76.170 151.605 ;
        RECT 76.340 151.515 76.565 151.645 ;
        RECT 76.340 150.410 76.510 151.515 ;
        RECT 76.735 151.365 77.260 151.585 ;
        RECT 76.680 150.600 76.920 151.195 ;
        RECT 77.090 150.665 77.260 151.365 ;
        RECT 77.430 151.005 77.600 151.785 ;
        RECT 77.920 151.735 78.290 152.235 ;
        RECT 78.470 151.785 78.875 151.955 ;
        RECT 79.045 151.785 79.830 151.955 ;
        RECT 78.470 151.555 78.640 151.785 ;
        RECT 77.810 151.255 78.640 151.555 ;
        RECT 79.025 151.285 79.490 151.615 ;
        RECT 77.810 151.225 78.010 151.255 ;
        RECT 78.130 151.005 78.300 151.075 ;
        RECT 77.430 150.835 78.300 151.005 ;
        RECT 77.790 150.745 78.300 150.835 ;
        RECT 76.340 150.280 76.645 150.410 ;
        RECT 77.090 150.300 77.620 150.665 ;
        RECT 75.960 149.685 76.225 150.145 ;
        RECT 76.395 149.855 76.645 150.280 ;
        RECT 77.790 150.130 77.960 150.745 ;
        RECT 76.855 149.960 77.960 150.130 ;
        RECT 78.130 149.685 78.300 150.485 ;
        RECT 78.470 150.185 78.640 151.255 ;
        RECT 78.810 150.355 79.000 151.075 ;
        RECT 79.170 150.325 79.490 151.285 ;
        RECT 79.660 151.325 79.830 151.785 ;
        RECT 80.105 151.705 80.315 152.235 ;
        RECT 80.575 151.495 80.905 152.020 ;
        RECT 81.075 151.625 81.245 152.235 ;
        RECT 81.415 151.580 81.745 152.015 ;
        RECT 81.415 151.495 81.795 151.580 ;
        RECT 80.705 151.325 80.905 151.495 ;
        RECT 81.570 151.455 81.795 151.495 ;
        RECT 81.965 151.485 83.175 152.235 ;
        RECT 79.660 150.995 80.535 151.325 ;
        RECT 80.705 150.995 81.455 151.325 ;
        RECT 78.470 149.855 78.720 150.185 ;
        RECT 79.660 150.155 79.830 150.995 ;
        RECT 80.705 150.790 80.895 150.995 ;
        RECT 81.625 150.875 81.795 151.455 ;
        RECT 81.580 150.825 81.795 150.875 ;
        RECT 80.000 150.415 80.895 150.790 ;
        RECT 81.405 150.745 81.795 150.825 ;
        RECT 81.965 150.775 82.485 151.315 ;
        RECT 82.655 150.945 83.175 151.485 ;
        RECT 78.945 149.985 79.830 150.155 ;
        RECT 80.010 149.685 80.325 150.185 ;
        RECT 80.555 149.855 80.895 150.415 ;
        RECT 81.065 149.685 81.235 150.695 ;
        RECT 81.405 149.900 81.735 150.745 ;
        RECT 81.965 149.685 83.175 150.775 ;
        RECT 5.520 149.515 83.260 149.685 ;
        RECT 5.605 148.425 6.815 149.515 ;
        RECT 6.985 149.080 12.330 149.515 ;
        RECT 12.505 149.080 17.850 149.515 ;
        RECT 5.605 147.715 6.125 148.255 ;
        RECT 6.295 147.885 6.815 148.425 ;
        RECT 5.605 146.965 6.815 147.715 ;
        RECT 8.570 147.510 8.910 148.340 ;
        RECT 10.390 147.830 10.740 149.080 ;
        RECT 14.090 147.510 14.430 148.340 ;
        RECT 15.910 147.830 16.260 149.080 ;
        RECT 18.485 148.350 18.775 149.515 ;
        RECT 18.945 149.080 24.290 149.515 ;
        RECT 6.985 146.965 12.330 147.510 ;
        RECT 12.505 146.965 17.850 147.510 ;
        RECT 18.485 146.965 18.775 147.690 ;
        RECT 20.530 147.510 20.870 148.340 ;
        RECT 22.350 147.830 22.700 149.080 ;
        RECT 24.465 148.425 27.975 149.515 ;
        RECT 24.465 147.735 26.115 148.255 ;
        RECT 26.285 147.905 27.975 148.425 ;
        RECT 28.610 148.375 28.885 149.345 ;
        RECT 29.095 148.715 29.375 149.515 ;
        RECT 29.545 149.005 30.735 149.295 ;
        RECT 29.545 148.665 30.715 148.835 ;
        RECT 29.545 148.545 29.715 148.665 ;
        RECT 29.055 148.375 29.715 148.545 ;
        RECT 18.945 146.965 24.290 147.510 ;
        RECT 24.465 146.965 27.975 147.735 ;
        RECT 28.610 147.640 28.780 148.375 ;
        RECT 29.055 148.205 29.225 148.375 ;
        RECT 30.025 148.205 30.220 148.495 ;
        RECT 30.390 148.375 30.715 148.665 ;
        RECT 31.090 148.545 31.480 148.720 ;
        RECT 31.965 148.715 32.295 149.515 ;
        RECT 32.465 148.725 33.000 149.345 ;
        RECT 31.090 148.375 32.515 148.545 ;
        RECT 28.950 147.875 29.225 148.205 ;
        RECT 29.395 147.875 30.220 148.205 ;
        RECT 30.390 147.875 30.735 148.205 ;
        RECT 29.055 147.705 29.225 147.875 ;
        RECT 28.610 147.295 28.885 147.640 ;
        RECT 29.055 147.535 30.720 147.705 ;
        RECT 30.965 147.645 31.320 148.205 ;
        RECT 29.075 146.965 29.455 147.365 ;
        RECT 29.625 147.185 29.795 147.535 ;
        RECT 29.965 146.965 30.295 147.365 ;
        RECT 30.465 147.185 30.720 147.535 ;
        RECT 31.490 147.475 31.660 148.375 ;
        RECT 31.830 147.645 32.095 148.205 ;
        RECT 32.345 147.875 32.515 148.375 ;
        RECT 32.685 147.705 33.000 148.725 ;
        RECT 31.070 146.965 31.310 147.475 ;
        RECT 31.490 147.145 31.770 147.475 ;
        RECT 32.000 146.965 32.215 147.475 ;
        RECT 32.385 147.135 33.000 147.705 ;
        RECT 33.205 148.375 33.480 149.345 ;
        RECT 33.690 148.715 33.970 149.515 ;
        RECT 34.140 149.005 35.755 149.335 ;
        RECT 34.140 148.665 35.315 148.835 ;
        RECT 34.140 148.545 34.310 148.665 ;
        RECT 33.650 148.375 34.310 148.545 ;
        RECT 33.205 147.640 33.375 148.375 ;
        RECT 33.650 148.205 33.820 148.375 ;
        RECT 34.570 148.205 34.815 148.495 ;
        RECT 34.985 148.375 35.315 148.665 ;
        RECT 35.575 148.205 35.745 148.765 ;
        RECT 35.995 148.375 36.255 149.515 ;
        RECT 36.425 148.375 36.810 149.345 ;
        RECT 36.980 149.055 37.305 149.515 ;
        RECT 37.825 148.885 38.105 149.345 ;
        RECT 36.980 148.665 38.105 148.885 ;
        RECT 33.545 147.875 33.820 148.205 ;
        RECT 33.990 147.875 34.815 148.205 ;
        RECT 35.030 147.875 35.745 148.205 ;
        RECT 35.915 147.955 36.250 148.205 ;
        RECT 33.650 147.705 33.820 147.875 ;
        RECT 35.495 147.785 35.745 147.875 ;
        RECT 33.205 147.295 33.480 147.640 ;
        RECT 33.650 147.535 35.315 147.705 ;
        RECT 33.670 146.965 34.045 147.365 ;
        RECT 34.215 147.185 34.385 147.535 ;
        RECT 34.555 146.965 34.885 147.365 ;
        RECT 35.055 147.135 35.315 147.535 ;
        RECT 35.495 147.365 35.825 147.785 ;
        RECT 35.995 146.965 36.255 147.785 ;
        RECT 36.425 147.705 36.705 148.375 ;
        RECT 36.980 148.205 37.430 148.665 ;
        RECT 38.295 148.495 38.695 149.345 ;
        RECT 39.095 149.055 39.365 149.515 ;
        RECT 39.535 148.885 39.820 149.345 ;
        RECT 36.875 147.875 37.430 148.205 ;
        RECT 37.600 147.935 38.695 148.495 ;
        RECT 36.980 147.765 37.430 147.875 ;
        RECT 36.425 147.135 36.810 147.705 ;
        RECT 36.980 147.595 38.105 147.765 ;
        RECT 36.980 146.965 37.305 147.425 ;
        RECT 37.825 147.135 38.105 147.595 ;
        RECT 38.295 147.135 38.695 147.935 ;
        RECT 38.865 148.665 39.820 148.885 ;
        RECT 40.220 148.885 40.505 149.345 ;
        RECT 40.675 149.055 40.945 149.515 ;
        RECT 40.220 148.665 41.175 148.885 ;
        RECT 38.865 147.765 39.075 148.665 ;
        RECT 39.245 147.935 39.935 148.495 ;
        RECT 40.105 147.935 40.795 148.495 ;
        RECT 40.965 147.765 41.175 148.665 ;
        RECT 38.865 147.595 39.820 147.765 ;
        RECT 39.095 146.965 39.365 147.425 ;
        RECT 39.535 147.135 39.820 147.595 ;
        RECT 40.220 147.595 41.175 147.765 ;
        RECT 41.345 148.495 41.745 149.345 ;
        RECT 41.935 148.885 42.215 149.345 ;
        RECT 42.735 149.055 43.060 149.515 ;
        RECT 41.935 148.665 43.060 148.885 ;
        RECT 41.345 147.935 42.440 148.495 ;
        RECT 42.610 148.205 43.060 148.665 ;
        RECT 43.230 148.375 43.615 149.345 ;
        RECT 40.220 147.135 40.505 147.595 ;
        RECT 40.675 146.965 40.945 147.425 ;
        RECT 41.345 147.135 41.745 147.935 ;
        RECT 42.610 147.875 43.165 148.205 ;
        RECT 42.610 147.765 43.060 147.875 ;
        RECT 41.935 147.595 43.060 147.765 ;
        RECT 43.335 147.705 43.615 148.375 ;
        RECT 44.245 148.350 44.535 149.515 ;
        RECT 44.705 148.375 44.965 149.515 ;
        RECT 45.135 148.365 45.465 149.345 ;
        RECT 45.635 148.375 45.915 149.515 ;
        RECT 46.085 148.375 46.425 149.345 ;
        RECT 46.595 148.375 46.765 149.515 ;
        RECT 47.035 148.715 47.285 149.515 ;
        RECT 47.930 148.545 48.260 149.345 ;
        RECT 48.560 148.715 48.890 149.515 ;
        RECT 49.060 148.545 49.390 149.345 ;
        RECT 46.955 148.375 49.390 148.545 ;
        RECT 49.765 148.645 50.040 149.345 ;
        RECT 50.250 148.970 50.465 149.515 ;
        RECT 50.635 149.005 51.110 149.345 ;
        RECT 51.280 149.010 51.895 149.515 ;
        RECT 51.280 148.835 51.475 149.010 ;
        RECT 44.725 147.955 45.060 148.205 ;
        RECT 45.230 147.765 45.400 148.365 ;
        RECT 45.570 147.935 45.905 148.205 ;
        RECT 46.085 147.765 46.260 148.375 ;
        RECT 46.955 148.125 47.125 148.375 ;
        RECT 46.430 147.955 47.125 148.125 ;
        RECT 47.300 147.955 47.720 148.155 ;
        RECT 47.890 147.955 48.220 148.155 ;
        RECT 48.390 147.955 48.720 148.155 ;
        RECT 41.935 147.135 42.215 147.595 ;
        RECT 42.735 146.965 43.060 147.425 ;
        RECT 43.230 147.135 43.615 147.705 ;
        RECT 44.245 146.965 44.535 147.690 ;
        RECT 44.705 147.135 45.400 147.765 ;
        RECT 45.605 146.965 45.915 147.765 ;
        RECT 46.085 147.135 46.425 147.765 ;
        RECT 46.595 146.965 46.845 147.765 ;
        RECT 47.035 147.615 48.260 147.785 ;
        RECT 47.035 147.135 47.365 147.615 ;
        RECT 47.535 146.965 47.760 147.425 ;
        RECT 47.930 147.135 48.260 147.615 ;
        RECT 48.890 147.745 49.060 148.375 ;
        RECT 49.245 147.955 49.595 148.205 ;
        RECT 48.890 147.135 49.390 147.745 ;
        RECT 49.765 147.615 49.935 148.645 ;
        RECT 50.210 148.475 50.925 148.770 ;
        RECT 51.145 148.645 51.475 148.835 ;
        RECT 51.645 148.475 51.895 148.840 ;
        RECT 50.105 148.305 51.895 148.475 ;
        RECT 50.105 147.875 50.335 148.305 ;
        RECT 49.765 147.135 50.025 147.615 ;
        RECT 50.505 147.605 50.915 148.125 ;
        RECT 50.195 146.965 50.525 147.425 ;
        RECT 50.715 147.185 50.915 147.605 ;
        RECT 51.085 147.450 51.340 148.305 ;
        RECT 52.135 148.125 52.305 149.345 ;
        RECT 52.555 149.005 52.815 149.515 ;
        RECT 51.510 147.875 52.305 148.125 ;
        RECT 52.475 147.955 52.815 148.835 ;
        RECT 53.005 148.460 53.310 149.245 ;
        RECT 53.490 149.045 54.175 149.515 ;
        RECT 53.485 148.525 54.180 148.835 ;
        RECT 52.055 147.785 52.305 147.875 ;
        RECT 51.085 147.185 51.875 147.450 ;
        RECT 52.055 147.365 52.385 147.785 ;
        RECT 52.555 146.965 52.815 147.785 ;
        RECT 53.005 147.655 53.180 148.460 ;
        RECT 54.355 148.355 54.640 149.300 ;
        RECT 54.815 149.065 55.145 149.515 ;
        RECT 55.315 148.895 55.485 149.325 ;
        RECT 53.780 148.205 54.640 148.355 ;
        RECT 53.355 148.185 54.640 148.205 ;
        RECT 54.810 148.665 55.485 148.895 ;
        RECT 53.355 147.825 54.340 148.185 ;
        RECT 54.810 148.015 55.045 148.665 ;
        RECT 55.750 148.565 56.015 149.335 ;
        RECT 56.185 148.795 56.515 149.515 ;
        RECT 56.705 148.975 56.965 149.335 ;
        RECT 57.135 149.145 57.465 149.515 ;
        RECT 57.635 148.975 57.895 149.335 ;
        RECT 56.705 148.745 57.895 148.975 ;
        RECT 58.465 148.565 58.755 149.335 ;
        RECT 53.005 147.135 53.245 147.655 ;
        RECT 54.170 147.490 54.340 147.825 ;
        RECT 54.510 147.685 55.045 148.015 ;
        RECT 54.825 147.535 55.045 147.685 ;
        RECT 55.215 147.645 55.515 148.495 ;
        RECT 53.415 146.965 53.810 147.460 ;
        RECT 54.170 147.295 54.545 147.490 ;
        RECT 54.375 147.150 54.545 147.295 ;
        RECT 54.825 147.160 55.065 147.535 ;
        RECT 55.235 146.965 55.570 147.470 ;
        RECT 55.750 147.145 56.085 148.565 ;
        RECT 56.260 148.385 58.755 148.565 ;
        RECT 56.260 147.695 56.485 148.385 ;
        RECT 58.970 148.375 59.305 149.345 ;
        RECT 59.475 148.375 59.645 149.515 ;
        RECT 59.815 149.175 61.845 149.345 ;
        RECT 56.685 147.875 56.965 148.205 ;
        RECT 57.145 147.875 57.720 148.205 ;
        RECT 57.900 147.875 58.335 148.205 ;
        RECT 58.515 147.875 58.785 148.205 ;
        RECT 58.970 147.705 59.140 148.375 ;
        RECT 59.815 148.205 59.985 149.175 ;
        RECT 59.310 147.875 59.565 148.205 ;
        RECT 59.790 147.875 59.985 148.205 ;
        RECT 60.155 148.835 61.280 149.005 ;
        RECT 59.395 147.705 59.565 147.875 ;
        RECT 60.155 147.705 60.325 148.835 ;
        RECT 56.260 147.505 58.745 147.695 ;
        RECT 56.265 146.965 57.010 147.335 ;
        RECT 57.575 147.145 57.830 147.505 ;
        RECT 58.010 146.965 58.340 147.335 ;
        RECT 58.520 147.145 58.745 147.505 ;
        RECT 58.970 147.135 59.225 147.705 ;
        RECT 59.395 147.535 60.325 147.705 ;
        RECT 60.495 148.495 61.505 148.665 ;
        RECT 60.495 147.695 60.665 148.495 ;
        RECT 60.870 148.155 61.145 148.295 ;
        RECT 60.865 147.985 61.145 148.155 ;
        RECT 60.150 147.500 60.325 147.535 ;
        RECT 59.395 146.965 59.725 147.365 ;
        RECT 60.150 147.135 60.680 147.500 ;
        RECT 60.870 147.135 61.145 147.985 ;
        RECT 61.315 147.135 61.505 148.495 ;
        RECT 61.675 148.510 61.845 149.175 ;
        RECT 62.015 148.755 62.185 149.515 ;
        RECT 62.420 148.755 62.935 149.165 ;
        RECT 61.675 148.320 62.425 148.510 ;
        RECT 62.595 147.945 62.935 148.755 ;
        RECT 61.705 147.775 62.935 147.945 ;
        RECT 63.110 148.375 63.445 149.345 ;
        RECT 63.615 148.375 63.785 149.515 ;
        RECT 63.955 149.175 65.985 149.345 ;
        RECT 61.685 146.965 62.195 147.500 ;
        RECT 62.415 147.170 62.660 147.775 ;
        RECT 63.110 147.705 63.280 148.375 ;
        RECT 63.955 148.205 64.125 149.175 ;
        RECT 63.450 147.875 63.705 148.205 ;
        RECT 63.930 147.875 64.125 148.205 ;
        RECT 64.295 148.835 65.420 149.005 ;
        RECT 63.535 147.705 63.705 147.875 ;
        RECT 64.295 147.705 64.465 148.835 ;
        RECT 63.110 147.135 63.365 147.705 ;
        RECT 63.535 147.535 64.465 147.705 ;
        RECT 64.635 148.495 65.645 148.665 ;
        RECT 64.635 147.695 64.805 148.495 ;
        RECT 65.010 148.155 65.285 148.295 ;
        RECT 65.005 147.985 65.285 148.155 ;
        RECT 64.290 147.500 64.465 147.535 ;
        RECT 63.535 146.965 63.865 147.365 ;
        RECT 64.290 147.135 64.820 147.500 ;
        RECT 65.010 147.135 65.285 147.985 ;
        RECT 65.455 147.135 65.645 148.495 ;
        RECT 65.815 148.510 65.985 149.175 ;
        RECT 66.155 148.755 66.325 149.515 ;
        RECT 66.560 148.755 67.075 149.165 ;
        RECT 65.815 148.320 66.565 148.510 ;
        RECT 66.735 147.945 67.075 148.755 ;
        RECT 67.890 148.545 68.280 148.720 ;
        RECT 68.765 148.715 69.095 149.515 ;
        RECT 69.265 148.725 69.800 149.345 ;
        RECT 67.890 148.375 69.315 148.545 ;
        RECT 65.845 147.775 67.075 147.945 ;
        RECT 65.825 146.965 66.335 147.500 ;
        RECT 66.555 147.170 66.800 147.775 ;
        RECT 67.765 147.645 68.120 148.205 ;
        RECT 68.290 147.475 68.460 148.375 ;
        RECT 68.630 147.645 68.895 148.205 ;
        RECT 69.145 147.875 69.315 148.375 ;
        RECT 69.485 147.705 69.800 148.725 ;
        RECT 70.005 148.350 70.295 149.515 ;
        RECT 70.465 148.375 70.850 149.345 ;
        RECT 71.020 149.055 71.345 149.515 ;
        RECT 71.865 148.885 72.145 149.345 ;
        RECT 71.020 148.665 72.145 148.885 ;
        RECT 67.870 146.965 68.110 147.475 ;
        RECT 68.290 147.145 68.570 147.475 ;
        RECT 68.800 146.965 69.015 147.475 ;
        RECT 69.185 147.135 69.800 147.705 ;
        RECT 70.465 147.705 70.745 148.375 ;
        RECT 71.020 148.205 71.470 148.665 ;
        RECT 72.335 148.495 72.735 149.345 ;
        RECT 73.135 149.055 73.405 149.515 ;
        RECT 73.575 148.885 73.860 149.345 ;
        RECT 70.915 147.875 71.470 148.205 ;
        RECT 71.640 147.935 72.735 148.495 ;
        RECT 71.020 147.765 71.470 147.875 ;
        RECT 70.005 146.965 70.295 147.690 ;
        RECT 70.465 147.135 70.850 147.705 ;
        RECT 71.020 147.595 72.145 147.765 ;
        RECT 71.020 146.965 71.345 147.425 ;
        RECT 71.865 147.135 72.145 147.595 ;
        RECT 72.335 147.135 72.735 147.935 ;
        RECT 72.905 148.665 73.860 148.885 ;
        RECT 72.905 147.765 73.115 148.665 ;
        RECT 73.285 147.935 73.975 148.495 ;
        RECT 74.145 148.375 74.485 149.345 ;
        RECT 74.655 148.375 74.825 149.515 ;
        RECT 75.095 148.715 75.345 149.515 ;
        RECT 75.990 148.545 76.320 149.345 ;
        RECT 76.620 148.715 76.950 149.515 ;
        RECT 77.120 148.545 77.450 149.345 ;
        RECT 75.015 148.375 77.450 148.545 ;
        RECT 77.825 148.375 78.165 149.345 ;
        RECT 78.335 148.375 78.505 149.515 ;
        RECT 78.775 148.715 79.025 149.515 ;
        RECT 79.670 148.545 80.000 149.345 ;
        RECT 80.300 148.715 80.630 149.515 ;
        RECT 80.800 148.545 81.130 149.345 ;
        RECT 78.695 148.375 81.130 148.545 ;
        RECT 81.965 148.425 83.175 149.515 ;
        RECT 74.145 147.765 74.320 148.375 ;
        RECT 75.015 148.125 75.185 148.375 ;
        RECT 74.490 147.955 75.185 148.125 ;
        RECT 75.360 147.955 75.780 148.155 ;
        RECT 75.950 147.955 76.280 148.155 ;
        RECT 76.450 147.955 76.780 148.155 ;
        RECT 72.905 147.595 73.860 147.765 ;
        RECT 73.135 146.965 73.405 147.425 ;
        RECT 73.575 147.135 73.860 147.595 ;
        RECT 74.145 147.135 74.485 147.765 ;
        RECT 74.655 146.965 74.905 147.765 ;
        RECT 75.095 147.615 76.320 147.785 ;
        RECT 75.095 147.135 75.425 147.615 ;
        RECT 75.595 146.965 75.820 147.425 ;
        RECT 75.990 147.135 76.320 147.615 ;
        RECT 76.950 147.745 77.120 148.375 ;
        RECT 77.305 147.955 77.655 148.205 ;
        RECT 77.825 147.765 78.000 148.375 ;
        RECT 78.695 148.125 78.865 148.375 ;
        RECT 78.170 147.955 78.865 148.125 ;
        RECT 79.040 147.955 79.460 148.155 ;
        RECT 79.630 147.955 79.960 148.155 ;
        RECT 80.130 147.955 80.460 148.155 ;
        RECT 76.950 147.135 77.450 147.745 ;
        RECT 77.825 147.135 78.165 147.765 ;
        RECT 78.335 146.965 78.585 147.765 ;
        RECT 78.775 147.615 80.000 147.785 ;
        RECT 78.775 147.135 79.105 147.615 ;
        RECT 79.275 146.965 79.500 147.425 ;
        RECT 79.670 147.135 80.000 147.615 ;
        RECT 80.630 147.745 80.800 148.375 ;
        RECT 80.985 147.955 81.335 148.205 ;
        RECT 81.965 147.885 82.485 148.425 ;
        RECT 80.630 147.135 81.130 147.745 ;
        RECT 82.655 147.715 83.175 148.255 ;
        RECT 81.965 146.965 83.175 147.715 ;
        RECT 5.520 146.795 83.260 146.965 ;
        RECT 5.605 146.045 6.815 146.795 ;
        RECT 6.985 146.250 12.330 146.795 ;
        RECT 12.505 146.250 17.850 146.795 ;
        RECT 18.025 146.250 23.370 146.795 ;
        RECT 23.545 146.250 28.890 146.795 ;
        RECT 5.605 145.505 6.125 146.045 ;
        RECT 6.295 145.335 6.815 145.875 ;
        RECT 8.570 145.420 8.910 146.250 ;
        RECT 5.605 144.245 6.815 145.335 ;
        RECT 10.390 144.680 10.740 145.930 ;
        RECT 14.090 145.420 14.430 146.250 ;
        RECT 15.910 144.680 16.260 145.930 ;
        RECT 19.610 145.420 19.950 146.250 ;
        RECT 21.430 144.680 21.780 145.930 ;
        RECT 25.130 145.420 25.470 146.250 ;
        RECT 29.065 146.025 30.735 146.795 ;
        RECT 31.365 146.070 31.655 146.795 ;
        RECT 32.755 146.070 33.085 146.580 ;
        RECT 33.255 146.395 33.585 146.795 ;
        RECT 34.635 146.225 34.965 146.565 ;
        RECT 35.135 146.395 35.465 146.795 ;
        RECT 26.950 144.680 27.300 145.930 ;
        RECT 29.065 145.505 29.815 146.025 ;
        RECT 29.985 145.335 30.735 145.855 ;
        RECT 6.985 144.245 12.330 144.680 ;
        RECT 12.505 144.245 17.850 144.680 ;
        RECT 18.025 144.245 23.370 144.680 ;
        RECT 23.545 144.245 28.890 144.680 ;
        RECT 29.065 144.245 30.735 145.335 ;
        RECT 31.365 144.245 31.655 145.410 ;
        RECT 32.755 145.305 32.945 146.070 ;
        RECT 33.255 146.055 35.620 146.225 ;
        RECT 36.475 146.140 36.805 146.575 ;
        RECT 36.975 146.185 37.145 146.795 ;
        RECT 33.255 145.885 33.425 146.055 ;
        RECT 33.115 145.555 33.425 145.885 ;
        RECT 33.595 145.555 33.900 145.885 ;
        RECT 32.755 144.455 33.085 145.305 ;
        RECT 33.255 144.245 33.505 145.385 ;
        RECT 33.685 145.225 33.900 145.555 ;
        RECT 34.075 145.225 34.360 145.885 ;
        RECT 34.555 145.225 34.820 145.885 ;
        RECT 35.035 145.225 35.280 145.885 ;
        RECT 35.450 145.055 35.620 146.055 ;
        RECT 36.425 146.055 36.805 146.140 ;
        RECT 37.315 146.055 37.645 146.580 ;
        RECT 37.905 146.265 38.115 146.795 ;
        RECT 38.390 146.345 39.175 146.515 ;
        RECT 39.345 146.345 39.750 146.515 ;
        RECT 36.425 146.015 36.650 146.055 ;
        RECT 36.425 145.435 36.595 146.015 ;
        RECT 37.315 145.885 37.515 146.055 ;
        RECT 38.390 145.885 38.560 146.345 ;
        RECT 36.765 145.555 37.515 145.885 ;
        RECT 37.685 145.555 38.560 145.885 ;
        RECT 36.425 145.385 36.640 145.435 ;
        RECT 36.425 145.305 36.815 145.385 ;
        RECT 33.695 144.885 34.985 145.055 ;
        RECT 33.695 144.465 33.945 144.885 ;
        RECT 34.175 144.245 34.505 144.715 ;
        RECT 34.735 144.465 34.985 144.885 ;
        RECT 35.165 144.885 35.620 145.055 ;
        RECT 35.165 144.455 35.495 144.885 ;
        RECT 36.485 144.460 36.815 145.305 ;
        RECT 37.325 145.350 37.515 145.555 ;
        RECT 36.985 144.245 37.155 145.255 ;
        RECT 37.325 144.975 38.220 145.350 ;
        RECT 37.325 144.415 37.665 144.975 ;
        RECT 37.895 144.245 38.210 144.745 ;
        RECT 38.390 144.715 38.560 145.555 ;
        RECT 38.730 145.845 39.195 146.175 ;
        RECT 39.580 146.115 39.750 146.345 ;
        RECT 39.930 146.295 40.300 146.795 ;
        RECT 40.620 146.345 41.295 146.515 ;
        RECT 41.490 146.345 41.825 146.515 ;
        RECT 38.730 144.885 39.050 145.845 ;
        RECT 39.580 145.815 40.410 146.115 ;
        RECT 39.220 144.915 39.410 145.635 ;
        RECT 39.580 144.745 39.750 145.815 ;
        RECT 40.210 145.785 40.410 145.815 ;
        RECT 39.920 145.565 40.090 145.635 ;
        RECT 40.620 145.565 40.790 146.345 ;
        RECT 41.655 146.205 41.825 146.345 ;
        RECT 41.995 146.335 42.245 146.795 ;
        RECT 39.920 145.395 40.790 145.565 ;
        RECT 40.960 145.925 41.485 146.145 ;
        RECT 41.655 146.075 41.880 146.205 ;
        RECT 39.920 145.305 40.430 145.395 ;
        RECT 38.390 144.545 39.275 144.715 ;
        RECT 39.500 144.415 39.750 144.745 ;
        RECT 39.920 144.245 40.090 145.045 ;
        RECT 40.260 144.690 40.430 145.305 ;
        RECT 40.960 145.225 41.130 145.925 ;
        RECT 40.600 144.860 41.130 145.225 ;
        RECT 41.300 145.160 41.540 145.755 ;
        RECT 41.710 144.970 41.880 146.075 ;
        RECT 42.050 145.215 42.330 146.165 ;
        RECT 41.575 144.840 41.880 144.970 ;
        RECT 40.260 144.520 41.365 144.690 ;
        RECT 41.575 144.415 41.825 144.840 ;
        RECT 41.995 144.245 42.260 144.705 ;
        RECT 42.500 144.415 42.685 146.535 ;
        RECT 42.855 146.415 43.185 146.795 ;
        RECT 43.355 146.245 43.525 146.535 ;
        RECT 42.860 146.075 43.525 146.245 ;
        RECT 42.860 145.085 43.090 146.075 ;
        RECT 43.260 145.255 43.610 145.905 ;
        RECT 42.860 144.915 43.525 145.085 ;
        RECT 42.855 144.245 43.185 144.745 ;
        RECT 43.355 144.415 43.525 144.915 ;
        RECT 43.795 144.425 44.055 146.615 ;
        RECT 44.315 146.425 44.985 146.795 ;
        RECT 45.165 146.245 45.475 146.615 ;
        RECT 44.245 146.045 45.475 146.245 ;
        RECT 44.245 145.375 44.535 146.045 ;
        RECT 45.655 145.865 45.885 146.505 ;
        RECT 46.065 146.065 46.355 146.795 ;
        RECT 47.555 146.245 47.725 146.535 ;
        RECT 47.895 146.415 48.225 146.795 ;
        RECT 47.555 146.075 48.220 146.245 ;
        RECT 44.715 145.555 45.180 145.865 ;
        RECT 45.360 145.555 45.885 145.865 ;
        RECT 46.065 145.555 46.365 145.885 ;
        RECT 44.245 145.155 45.015 145.375 ;
        RECT 44.225 144.245 44.565 144.975 ;
        RECT 44.745 144.425 45.015 145.155 ;
        RECT 45.195 145.135 46.355 145.375 ;
        RECT 47.470 145.255 47.820 145.905 ;
        RECT 45.195 144.425 45.425 145.135 ;
        RECT 45.595 144.245 45.925 144.955 ;
        RECT 46.095 144.425 46.355 145.135 ;
        RECT 47.990 145.085 48.220 146.075 ;
        RECT 47.555 144.915 48.220 145.085 ;
        RECT 47.555 144.415 47.725 144.915 ;
        RECT 47.895 144.245 48.225 144.745 ;
        RECT 48.395 144.415 48.580 146.535 ;
        RECT 48.835 146.335 49.085 146.795 ;
        RECT 49.255 146.345 49.590 146.515 ;
        RECT 49.785 146.345 50.460 146.515 ;
        RECT 49.255 146.205 49.425 146.345 ;
        RECT 48.750 145.215 49.030 146.165 ;
        RECT 49.200 146.075 49.425 146.205 ;
        RECT 49.200 144.970 49.370 146.075 ;
        RECT 49.595 145.925 50.120 146.145 ;
        RECT 49.540 145.160 49.780 145.755 ;
        RECT 49.950 145.225 50.120 145.925 ;
        RECT 50.290 145.565 50.460 146.345 ;
        RECT 50.780 146.295 51.150 146.795 ;
        RECT 51.330 146.345 51.735 146.515 ;
        RECT 51.905 146.345 52.690 146.515 ;
        RECT 51.330 146.115 51.500 146.345 ;
        RECT 50.670 145.815 51.500 146.115 ;
        RECT 51.885 145.845 52.350 146.175 ;
        RECT 50.670 145.785 50.870 145.815 ;
        RECT 50.990 145.565 51.160 145.635 ;
        RECT 50.290 145.395 51.160 145.565 ;
        RECT 50.650 145.305 51.160 145.395 ;
        RECT 49.200 144.840 49.505 144.970 ;
        RECT 49.950 144.860 50.480 145.225 ;
        RECT 48.820 144.245 49.085 144.705 ;
        RECT 49.255 144.415 49.505 144.840 ;
        RECT 50.650 144.690 50.820 145.305 ;
        RECT 49.715 144.520 50.820 144.690 ;
        RECT 50.990 144.245 51.160 145.045 ;
        RECT 51.330 144.745 51.500 145.815 ;
        RECT 51.670 144.915 51.860 145.635 ;
        RECT 52.030 144.885 52.350 145.845 ;
        RECT 52.520 145.885 52.690 146.345 ;
        RECT 52.965 146.265 53.175 146.795 ;
        RECT 53.435 146.055 53.765 146.580 ;
        RECT 53.935 146.185 54.105 146.795 ;
        RECT 54.275 146.140 54.605 146.575 ;
        RECT 54.825 146.145 55.085 146.625 ;
        RECT 55.255 146.255 55.505 146.795 ;
        RECT 54.275 146.055 54.655 146.140 ;
        RECT 53.565 145.885 53.765 146.055 ;
        RECT 54.430 146.015 54.655 146.055 ;
        RECT 52.520 145.555 53.395 145.885 ;
        RECT 53.565 145.555 54.315 145.885 ;
        RECT 51.330 144.415 51.580 144.745 ;
        RECT 52.520 144.715 52.690 145.555 ;
        RECT 53.565 145.350 53.755 145.555 ;
        RECT 54.485 145.435 54.655 146.015 ;
        RECT 54.440 145.385 54.655 145.435 ;
        RECT 52.860 144.975 53.755 145.350 ;
        RECT 54.265 145.305 54.655 145.385 ;
        RECT 51.805 144.545 52.690 144.715 ;
        RECT 52.870 144.245 53.185 144.745 ;
        RECT 53.415 144.415 53.755 144.975 ;
        RECT 53.925 144.245 54.095 145.255 ;
        RECT 54.265 144.460 54.595 145.305 ;
        RECT 54.825 145.115 54.995 146.145 ;
        RECT 55.675 146.090 55.895 146.575 ;
        RECT 55.165 145.495 55.395 145.890 ;
        RECT 55.565 145.665 55.895 146.090 ;
        RECT 56.065 146.415 56.955 146.585 ;
        RECT 56.065 145.690 56.235 146.415 ;
        RECT 56.405 145.860 56.955 146.245 ;
        RECT 57.125 146.070 57.415 146.795 ;
        RECT 57.585 146.055 57.970 146.625 ;
        RECT 58.140 146.335 58.465 146.795 ;
        RECT 58.985 146.165 59.265 146.625 ;
        RECT 56.065 145.620 56.955 145.690 ;
        RECT 56.060 145.595 56.955 145.620 ;
        RECT 56.050 145.580 56.955 145.595 ;
        RECT 56.045 145.565 56.955 145.580 ;
        RECT 56.035 145.560 56.955 145.565 ;
        RECT 56.030 145.550 56.955 145.560 ;
        RECT 56.025 145.540 56.955 145.550 ;
        RECT 56.015 145.535 56.955 145.540 ;
        RECT 56.005 145.525 56.955 145.535 ;
        RECT 55.995 145.520 56.955 145.525 ;
        RECT 55.995 145.515 56.330 145.520 ;
        RECT 55.980 145.510 56.330 145.515 ;
        RECT 55.965 145.500 56.330 145.510 ;
        RECT 55.940 145.495 56.330 145.500 ;
        RECT 55.165 145.490 56.330 145.495 ;
        RECT 55.165 145.455 56.300 145.490 ;
        RECT 55.165 145.430 56.265 145.455 ;
        RECT 55.165 145.400 56.235 145.430 ;
        RECT 55.165 145.370 56.215 145.400 ;
        RECT 55.165 145.340 56.195 145.370 ;
        RECT 55.165 145.330 56.125 145.340 ;
        RECT 55.165 145.320 56.100 145.330 ;
        RECT 55.165 145.305 56.080 145.320 ;
        RECT 55.165 145.290 56.060 145.305 ;
        RECT 55.270 145.280 56.055 145.290 ;
        RECT 55.270 145.245 56.040 145.280 ;
        RECT 54.825 144.415 55.100 145.115 ;
        RECT 55.270 144.995 56.025 145.245 ;
        RECT 56.195 144.925 56.525 145.170 ;
        RECT 56.695 145.070 56.955 145.520 ;
        RECT 56.340 144.900 56.525 144.925 ;
        RECT 56.340 144.800 56.955 144.900 ;
        RECT 55.270 144.245 55.525 144.790 ;
        RECT 55.695 144.415 56.175 144.755 ;
        RECT 56.350 144.245 56.955 144.800 ;
        RECT 57.125 144.245 57.415 145.410 ;
        RECT 57.585 145.385 57.865 146.055 ;
        RECT 58.140 145.995 59.265 146.165 ;
        RECT 58.140 145.885 58.590 145.995 ;
        RECT 58.035 145.555 58.590 145.885 ;
        RECT 59.455 145.825 59.855 146.625 ;
        RECT 60.255 146.335 60.525 146.795 ;
        RECT 60.695 146.165 60.980 146.625 ;
        RECT 57.585 144.415 57.970 145.385 ;
        RECT 58.140 145.095 58.590 145.555 ;
        RECT 58.760 145.265 59.855 145.825 ;
        RECT 58.140 144.875 59.265 145.095 ;
        RECT 58.140 144.245 58.465 144.705 ;
        RECT 58.985 144.415 59.265 144.875 ;
        RECT 59.455 144.415 59.855 145.265 ;
        RECT 60.025 145.995 60.980 146.165 ;
        RECT 61.355 146.245 61.525 146.535 ;
        RECT 61.695 146.415 62.025 146.795 ;
        RECT 61.355 146.075 62.020 146.245 ;
        RECT 60.025 145.095 60.235 145.995 ;
        RECT 60.405 145.265 61.095 145.825 ;
        RECT 61.270 145.255 61.620 145.905 ;
        RECT 60.025 144.875 60.980 145.095 ;
        RECT 61.790 145.085 62.020 146.075 ;
        RECT 60.255 144.245 60.525 144.705 ;
        RECT 60.695 144.415 60.980 144.875 ;
        RECT 61.355 144.915 62.020 145.085 ;
        RECT 61.355 144.415 61.525 144.915 ;
        RECT 61.695 144.245 62.025 144.745 ;
        RECT 62.195 144.415 62.380 146.535 ;
        RECT 62.635 146.335 62.885 146.795 ;
        RECT 63.055 146.345 63.390 146.515 ;
        RECT 63.585 146.345 64.260 146.515 ;
        RECT 63.055 146.205 63.225 146.345 ;
        RECT 62.550 145.215 62.830 146.165 ;
        RECT 63.000 146.075 63.225 146.205 ;
        RECT 63.000 144.970 63.170 146.075 ;
        RECT 63.395 145.925 63.920 146.145 ;
        RECT 63.340 145.160 63.580 145.755 ;
        RECT 63.750 145.225 63.920 145.925 ;
        RECT 64.090 145.565 64.260 146.345 ;
        RECT 64.580 146.295 64.950 146.795 ;
        RECT 65.130 146.345 65.535 146.515 ;
        RECT 65.705 146.345 66.490 146.515 ;
        RECT 65.130 146.115 65.300 146.345 ;
        RECT 64.470 145.815 65.300 146.115 ;
        RECT 65.685 145.845 66.150 146.175 ;
        RECT 64.470 145.785 64.670 145.815 ;
        RECT 64.790 145.565 64.960 145.635 ;
        RECT 64.090 145.395 64.960 145.565 ;
        RECT 64.450 145.305 64.960 145.395 ;
        RECT 63.000 144.840 63.305 144.970 ;
        RECT 63.750 144.860 64.280 145.225 ;
        RECT 62.620 144.245 62.885 144.705 ;
        RECT 63.055 144.415 63.305 144.840 ;
        RECT 64.450 144.690 64.620 145.305 ;
        RECT 63.515 144.520 64.620 144.690 ;
        RECT 64.790 144.245 64.960 145.045 ;
        RECT 65.130 144.745 65.300 145.815 ;
        RECT 65.470 144.915 65.660 145.635 ;
        RECT 65.830 144.885 66.150 145.845 ;
        RECT 66.320 145.885 66.490 146.345 ;
        RECT 66.765 146.265 66.975 146.795 ;
        RECT 67.235 146.055 67.565 146.580 ;
        RECT 67.735 146.185 67.905 146.795 ;
        RECT 68.075 146.140 68.405 146.575 ;
        RECT 68.075 146.055 68.455 146.140 ;
        RECT 67.365 145.885 67.565 146.055 ;
        RECT 68.230 146.015 68.455 146.055 ;
        RECT 66.320 145.555 67.195 145.885 ;
        RECT 67.365 145.555 68.115 145.885 ;
        RECT 65.130 144.415 65.380 144.745 ;
        RECT 66.320 144.715 66.490 145.555 ;
        RECT 67.365 145.350 67.555 145.555 ;
        RECT 68.285 145.435 68.455 146.015 ;
        RECT 68.240 145.385 68.455 145.435 ;
        RECT 66.660 144.975 67.555 145.350 ;
        RECT 68.065 145.305 68.455 145.385 ;
        RECT 68.625 146.055 69.010 146.625 ;
        RECT 69.180 146.335 69.505 146.795 ;
        RECT 70.025 146.165 70.305 146.625 ;
        RECT 68.625 145.385 68.905 146.055 ;
        RECT 69.180 145.995 70.305 146.165 ;
        RECT 69.180 145.885 69.630 145.995 ;
        RECT 69.075 145.555 69.630 145.885 ;
        RECT 70.495 145.825 70.895 146.625 ;
        RECT 71.295 146.335 71.565 146.795 ;
        RECT 71.735 146.165 72.020 146.625 ;
        RECT 65.605 144.545 66.490 144.715 ;
        RECT 66.670 144.245 66.985 144.745 ;
        RECT 67.215 144.415 67.555 144.975 ;
        RECT 67.725 144.245 67.895 145.255 ;
        RECT 68.065 144.460 68.395 145.305 ;
        RECT 68.625 144.415 69.010 145.385 ;
        RECT 69.180 145.095 69.630 145.555 ;
        RECT 69.800 145.265 70.895 145.825 ;
        RECT 69.180 144.875 70.305 145.095 ;
        RECT 69.180 144.245 69.505 144.705 ;
        RECT 70.025 144.415 70.305 144.875 ;
        RECT 70.495 144.415 70.895 145.265 ;
        RECT 71.065 145.995 72.020 146.165 ;
        RECT 71.065 145.095 71.275 145.995 ;
        RECT 71.445 145.265 72.135 145.825 ;
        RECT 72.310 145.195 72.645 146.615 ;
        RECT 72.825 146.425 73.570 146.795 ;
        RECT 74.135 146.255 74.390 146.615 ;
        RECT 74.570 146.425 74.900 146.795 ;
        RECT 75.080 146.255 75.305 146.615 ;
        RECT 72.820 146.065 75.305 146.255 ;
        RECT 75.615 146.245 75.785 146.625 ;
        RECT 76.000 146.415 76.330 146.795 ;
        RECT 75.615 146.075 76.330 146.245 ;
        RECT 72.820 145.375 73.045 146.065 ;
        RECT 73.245 145.555 73.525 145.885 ;
        RECT 73.705 145.555 74.280 145.885 ;
        RECT 74.460 145.555 74.895 145.885 ;
        RECT 75.075 145.555 75.345 145.885 ;
        RECT 75.525 145.525 75.880 145.895 ;
        RECT 76.160 145.885 76.330 146.075 ;
        RECT 76.500 146.050 76.755 146.625 ;
        RECT 76.160 145.555 76.415 145.885 ;
        RECT 72.820 145.195 75.315 145.375 ;
        RECT 76.160 145.345 76.330 145.555 ;
        RECT 71.065 144.875 72.020 145.095 ;
        RECT 71.295 144.245 71.565 144.705 ;
        RECT 71.735 144.415 72.020 144.875 ;
        RECT 72.310 144.425 72.575 145.195 ;
        RECT 72.745 144.245 73.075 144.965 ;
        RECT 73.265 144.785 74.455 145.015 ;
        RECT 73.265 144.425 73.525 144.785 ;
        RECT 73.695 144.245 74.025 144.615 ;
        RECT 74.195 144.425 74.455 144.785 ;
        RECT 75.025 144.425 75.315 145.195 ;
        RECT 75.615 145.175 76.330 145.345 ;
        RECT 76.585 145.320 76.755 146.050 ;
        RECT 76.930 145.955 77.190 146.795 ;
        RECT 75.615 144.415 75.785 145.175 ;
        RECT 76.000 144.245 76.330 145.005 ;
        RECT 76.500 144.415 76.755 145.320 ;
        RECT 76.930 144.245 77.190 145.395 ;
        RECT 77.370 145.195 77.705 146.615 ;
        RECT 77.885 146.425 78.630 146.795 ;
        RECT 79.195 146.255 79.450 146.615 ;
        RECT 79.630 146.425 79.960 146.795 ;
        RECT 80.140 146.255 80.365 146.615 ;
        RECT 77.880 146.065 80.365 146.255 ;
        RECT 80.585 146.120 80.845 146.625 ;
        RECT 81.025 146.415 81.355 146.795 ;
        RECT 81.535 146.245 81.705 146.625 ;
        RECT 77.880 145.375 78.105 146.065 ;
        RECT 78.305 145.555 78.585 145.885 ;
        RECT 78.765 145.555 79.340 145.885 ;
        RECT 79.520 145.555 79.955 145.885 ;
        RECT 80.135 145.555 80.405 145.885 ;
        RECT 77.880 145.195 80.375 145.375 ;
        RECT 77.370 144.425 77.635 145.195 ;
        RECT 77.805 144.245 78.135 144.965 ;
        RECT 78.325 144.785 79.515 145.015 ;
        RECT 78.325 144.425 78.585 144.785 ;
        RECT 78.755 144.245 79.085 144.615 ;
        RECT 79.255 144.425 79.515 144.785 ;
        RECT 80.085 144.425 80.375 145.195 ;
        RECT 80.585 145.320 80.765 146.120 ;
        RECT 81.040 146.075 81.705 146.245 ;
        RECT 81.040 145.820 81.210 146.075 ;
        RECT 81.965 146.045 83.175 146.795 ;
        RECT 80.935 145.490 81.210 145.820 ;
        RECT 81.435 145.525 81.775 145.895 ;
        RECT 81.040 145.345 81.210 145.490 ;
        RECT 80.585 144.415 80.855 145.320 ;
        RECT 81.040 145.175 81.715 145.345 ;
        RECT 81.025 144.245 81.355 145.005 ;
        RECT 81.535 144.415 81.715 145.175 ;
        RECT 81.965 145.335 82.485 145.875 ;
        RECT 82.655 145.505 83.175 146.045 ;
        RECT 81.965 144.245 83.175 145.335 ;
        RECT 5.520 144.075 83.260 144.245 ;
        RECT 5.605 142.985 6.815 144.075 ;
        RECT 6.985 143.640 12.330 144.075 ;
        RECT 5.605 142.275 6.125 142.815 ;
        RECT 6.295 142.445 6.815 142.985 ;
        RECT 5.605 141.525 6.815 142.275 ;
        RECT 8.570 142.070 8.910 142.900 ;
        RECT 10.390 142.390 10.740 143.640 ;
        RECT 12.505 142.985 16.015 144.075 ;
        RECT 16.650 143.650 16.985 144.075 ;
        RECT 17.155 143.470 17.340 143.875 ;
        RECT 12.505 142.295 14.155 142.815 ;
        RECT 14.325 142.465 16.015 142.985 ;
        RECT 16.675 143.295 17.340 143.470 ;
        RECT 17.545 143.295 17.875 144.075 ;
        RECT 6.985 141.525 12.330 142.070 ;
        RECT 12.505 141.525 16.015 142.295 ;
        RECT 16.675 142.265 17.015 143.295 ;
        RECT 18.045 143.105 18.315 143.875 ;
        RECT 17.185 142.935 18.315 143.105 ;
        RECT 17.185 142.435 17.435 142.935 ;
        RECT 16.675 142.095 17.360 142.265 ;
        RECT 17.615 142.185 17.975 142.765 ;
        RECT 16.650 141.525 16.985 141.925 ;
        RECT 17.155 141.695 17.360 142.095 ;
        RECT 18.145 142.025 18.315 142.935 ;
        RECT 18.485 142.910 18.775 144.075 ;
        RECT 18.945 143.640 24.290 144.075 ;
        RECT 24.465 143.640 29.810 144.075 ;
        RECT 17.570 141.525 17.845 142.005 ;
        RECT 18.055 141.695 18.315 142.025 ;
        RECT 18.485 141.525 18.775 142.250 ;
        RECT 20.530 142.070 20.870 142.900 ;
        RECT 22.350 142.390 22.700 143.640 ;
        RECT 26.050 142.070 26.390 142.900 ;
        RECT 27.870 142.390 28.220 143.640 ;
        RECT 29.985 142.985 33.495 144.075 ;
        RECT 29.985 142.295 31.635 142.815 ;
        RECT 31.805 142.465 33.495 142.985 ;
        RECT 33.705 142.935 33.935 144.075 ;
        RECT 34.105 142.925 34.435 143.905 ;
        RECT 34.605 142.935 34.815 144.075 ;
        RECT 35.045 142.935 35.305 144.075 ;
        RECT 35.475 142.925 35.805 143.905 ;
        RECT 35.975 142.935 36.255 144.075 ;
        RECT 36.425 142.985 37.635 144.075 ;
        RECT 33.685 142.515 34.015 142.765 ;
        RECT 18.945 141.525 24.290 142.070 ;
        RECT 24.465 141.525 29.810 142.070 ;
        RECT 29.985 141.525 33.495 142.295 ;
        RECT 33.705 141.525 33.935 142.345 ;
        RECT 34.185 142.325 34.435 142.925 ;
        RECT 35.065 142.515 35.400 142.765 ;
        RECT 34.105 141.695 34.435 142.325 ;
        RECT 34.605 141.525 34.815 142.345 ;
        RECT 35.570 142.325 35.740 142.925 ;
        RECT 35.910 142.495 36.245 142.765 ;
        RECT 35.045 141.695 35.740 142.325 ;
        RECT 35.945 141.525 36.255 142.325 ;
        RECT 36.425 142.275 36.945 142.815 ;
        RECT 37.115 142.445 37.635 142.985 ;
        RECT 37.805 142.935 38.190 143.905 ;
        RECT 38.360 143.615 38.685 144.075 ;
        RECT 39.205 143.445 39.485 143.905 ;
        RECT 38.360 143.225 39.485 143.445 ;
        RECT 36.425 141.525 37.635 142.275 ;
        RECT 37.805 142.265 38.085 142.935 ;
        RECT 38.360 142.765 38.810 143.225 ;
        RECT 39.675 143.055 40.075 143.905 ;
        RECT 40.475 143.615 40.745 144.075 ;
        RECT 40.915 143.445 41.200 143.905 ;
        RECT 38.255 142.435 38.810 142.765 ;
        RECT 38.980 142.495 40.075 143.055 ;
        RECT 38.360 142.325 38.810 142.435 ;
        RECT 37.805 141.695 38.190 142.265 ;
        RECT 38.360 142.155 39.485 142.325 ;
        RECT 38.360 141.525 38.685 141.985 ;
        RECT 39.205 141.695 39.485 142.155 ;
        RECT 39.675 141.695 40.075 142.495 ;
        RECT 40.245 143.225 41.200 143.445 ;
        RECT 40.245 142.325 40.455 143.225 ;
        RECT 40.625 142.495 41.315 143.055 ;
        RECT 41.485 142.985 42.695 144.075 ;
        RECT 40.245 142.155 41.200 142.325 ;
        RECT 40.475 141.525 40.745 141.985 ;
        RECT 40.915 141.695 41.200 142.155 ;
        RECT 41.485 142.275 42.005 142.815 ;
        RECT 42.175 142.445 42.695 142.985 ;
        RECT 42.875 142.935 43.205 144.075 ;
        RECT 43.735 143.105 44.065 143.890 ;
        RECT 43.385 142.935 44.065 143.105 ;
        RECT 42.865 142.515 43.215 142.765 ;
        RECT 43.385 142.335 43.555 142.935 ;
        RECT 44.245 142.910 44.535 144.075 ;
        RECT 44.705 143.520 45.310 144.075 ;
        RECT 45.485 143.565 45.965 143.905 ;
        RECT 46.135 143.530 46.390 144.075 ;
        RECT 44.705 143.420 45.320 143.520 ;
        RECT 45.135 143.395 45.320 143.420 ;
        RECT 44.705 142.800 44.965 143.250 ;
        RECT 45.135 143.150 45.465 143.395 ;
        RECT 45.635 143.075 46.390 143.325 ;
        RECT 46.560 143.205 46.835 143.905 ;
        RECT 45.620 143.040 46.390 143.075 ;
        RECT 45.605 143.030 46.390 143.040 ;
        RECT 45.600 143.015 46.495 143.030 ;
        RECT 45.580 143.000 46.495 143.015 ;
        RECT 45.560 142.990 46.495 143.000 ;
        RECT 45.535 142.980 46.495 142.990 ;
        RECT 45.465 142.950 46.495 142.980 ;
        RECT 45.445 142.920 46.495 142.950 ;
        RECT 45.425 142.890 46.495 142.920 ;
        RECT 45.395 142.865 46.495 142.890 ;
        RECT 45.360 142.830 46.495 142.865 ;
        RECT 45.330 142.825 46.495 142.830 ;
        RECT 45.330 142.820 45.720 142.825 ;
        RECT 45.330 142.810 45.695 142.820 ;
        RECT 45.330 142.805 45.680 142.810 ;
        RECT 45.330 142.800 45.665 142.805 ;
        RECT 44.705 142.795 45.665 142.800 ;
        RECT 44.705 142.785 45.655 142.795 ;
        RECT 44.705 142.780 45.645 142.785 ;
        RECT 44.705 142.770 45.635 142.780 ;
        RECT 43.725 142.515 44.075 142.765 ;
        RECT 44.705 142.760 45.630 142.770 ;
        RECT 44.705 142.755 45.625 142.760 ;
        RECT 44.705 142.740 45.615 142.755 ;
        RECT 44.705 142.725 45.610 142.740 ;
        RECT 44.705 142.700 45.600 142.725 ;
        RECT 44.705 142.630 45.595 142.700 ;
        RECT 41.485 141.525 42.695 142.275 ;
        RECT 42.875 141.525 43.145 142.335 ;
        RECT 43.315 141.695 43.645 142.335 ;
        RECT 43.815 141.525 44.055 142.335 ;
        RECT 44.245 141.525 44.535 142.250 ;
        RECT 44.705 142.075 45.255 142.460 ;
        RECT 45.425 141.905 45.595 142.630 ;
        RECT 44.705 141.735 45.595 141.905 ;
        RECT 45.765 142.230 46.095 142.655 ;
        RECT 46.265 142.430 46.495 142.825 ;
        RECT 45.765 141.745 45.985 142.230 ;
        RECT 46.665 142.175 46.835 143.205 ;
        RECT 47.005 142.985 48.675 144.075 ;
        RECT 46.155 141.525 46.405 142.065 ;
        RECT 46.575 141.695 46.835 142.175 ;
        RECT 47.005 142.295 47.755 142.815 ;
        RECT 47.925 142.465 48.675 142.985 ;
        RECT 48.850 142.925 49.110 144.075 ;
        RECT 49.285 143.000 49.540 143.905 ;
        RECT 49.710 143.315 50.040 144.075 ;
        RECT 50.255 143.145 50.425 143.905 ;
        RECT 47.005 141.525 48.675 142.295 ;
        RECT 48.850 141.525 49.110 142.365 ;
        RECT 49.285 142.270 49.455 143.000 ;
        RECT 49.710 142.975 50.425 143.145 ;
        RECT 49.710 142.765 49.880 142.975 ;
        RECT 50.690 142.935 51.025 143.905 ;
        RECT 51.195 142.935 51.365 144.075 ;
        RECT 51.535 143.735 53.565 143.905 ;
        RECT 49.625 142.435 49.880 142.765 ;
        RECT 49.285 141.695 49.540 142.270 ;
        RECT 49.710 142.245 49.880 142.435 ;
        RECT 50.160 142.425 50.515 142.795 ;
        RECT 50.690 142.265 50.860 142.935 ;
        RECT 51.535 142.765 51.705 143.735 ;
        RECT 51.030 142.435 51.285 142.765 ;
        RECT 51.510 142.435 51.705 142.765 ;
        RECT 51.875 143.395 53.000 143.565 ;
        RECT 51.115 142.265 51.285 142.435 ;
        RECT 51.875 142.265 52.045 143.395 ;
        RECT 49.710 142.075 50.425 142.245 ;
        RECT 49.710 141.525 50.040 141.905 ;
        RECT 50.255 141.695 50.425 142.075 ;
        RECT 50.690 141.695 50.945 142.265 ;
        RECT 51.115 142.095 52.045 142.265 ;
        RECT 52.215 143.055 53.225 143.225 ;
        RECT 52.215 142.255 52.385 143.055 ;
        RECT 51.870 142.060 52.045 142.095 ;
        RECT 51.115 141.525 51.445 141.925 ;
        RECT 51.870 141.695 52.400 142.060 ;
        RECT 52.590 142.035 52.865 142.855 ;
        RECT 52.585 141.865 52.865 142.035 ;
        RECT 52.590 141.695 52.865 141.865 ;
        RECT 53.035 141.695 53.225 143.055 ;
        RECT 53.395 143.070 53.565 143.735 ;
        RECT 53.735 143.315 53.905 144.075 ;
        RECT 54.140 143.315 54.655 143.725 ;
        RECT 53.395 142.880 54.145 143.070 ;
        RECT 54.315 142.505 54.655 143.315 ;
        RECT 54.835 142.935 55.165 144.075 ;
        RECT 53.425 142.335 54.655 142.505 ;
        RECT 53.405 141.525 53.915 142.060 ;
        RECT 54.135 141.730 54.380 142.335 ;
        RECT 54.825 142.185 55.165 142.765 ;
        RECT 55.335 142.735 55.695 143.905 ;
        RECT 55.895 142.905 56.225 144.075 ;
        RECT 56.425 142.735 56.755 143.905 ;
        RECT 56.955 142.905 57.285 144.075 ;
        RECT 58.160 143.445 58.445 143.905 ;
        RECT 58.615 143.615 58.885 144.075 ;
        RECT 58.160 143.225 59.115 143.445 ;
        RECT 55.335 142.455 56.755 142.735 ;
        RECT 58.045 142.495 58.735 143.055 ;
        RECT 55.335 142.120 55.695 142.455 ;
        RECT 58.905 142.325 59.115 143.225 ;
        RECT 54.835 141.525 55.165 142.015 ;
        RECT 55.335 141.695 55.955 142.120 ;
        RECT 56.415 141.525 56.745 142.215 ;
        RECT 58.160 142.155 59.115 142.325 ;
        RECT 59.285 143.055 59.685 143.905 ;
        RECT 59.875 143.445 60.155 143.905 ;
        RECT 60.675 143.615 61.000 144.075 ;
        RECT 59.875 143.225 61.000 143.445 ;
        RECT 59.285 142.495 60.380 143.055 ;
        RECT 60.550 142.765 61.000 143.225 ;
        RECT 61.170 142.935 61.555 143.905 ;
        RECT 61.815 143.405 61.985 143.905 ;
        RECT 62.155 143.575 62.485 144.075 ;
        RECT 61.815 143.235 62.480 143.405 ;
        RECT 58.160 141.695 58.445 142.155 ;
        RECT 58.615 141.525 58.885 141.985 ;
        RECT 59.285 141.695 59.685 142.495 ;
        RECT 60.550 142.435 61.105 142.765 ;
        RECT 60.550 142.325 61.000 142.435 ;
        RECT 59.875 142.155 61.000 142.325 ;
        RECT 61.275 142.265 61.555 142.935 ;
        RECT 61.730 142.415 62.080 143.065 ;
        RECT 59.875 141.695 60.155 142.155 ;
        RECT 60.675 141.525 61.000 141.985 ;
        RECT 61.170 141.695 61.555 142.265 ;
        RECT 62.250 142.245 62.480 143.235 ;
        RECT 61.815 142.075 62.480 142.245 ;
        RECT 61.815 141.785 61.985 142.075 ;
        RECT 62.155 141.525 62.485 141.905 ;
        RECT 62.655 141.785 62.840 143.905 ;
        RECT 63.080 143.615 63.345 144.075 ;
        RECT 63.515 143.480 63.765 143.905 ;
        RECT 63.975 143.630 65.080 143.800 ;
        RECT 63.460 143.350 63.765 143.480 ;
        RECT 63.010 142.155 63.290 143.105 ;
        RECT 63.460 142.245 63.630 143.350 ;
        RECT 63.800 142.565 64.040 143.160 ;
        RECT 64.210 143.095 64.740 143.460 ;
        RECT 64.210 142.395 64.380 143.095 ;
        RECT 64.910 143.015 65.080 143.630 ;
        RECT 65.250 143.275 65.420 144.075 ;
        RECT 65.590 143.575 65.840 143.905 ;
        RECT 66.065 143.605 66.950 143.775 ;
        RECT 64.910 142.925 65.420 143.015 ;
        RECT 63.460 142.115 63.685 142.245 ;
        RECT 63.855 142.175 64.380 142.395 ;
        RECT 64.550 142.755 65.420 142.925 ;
        RECT 63.095 141.525 63.345 141.985 ;
        RECT 63.515 141.975 63.685 142.115 ;
        RECT 64.550 141.975 64.720 142.755 ;
        RECT 65.250 142.685 65.420 142.755 ;
        RECT 64.930 142.505 65.130 142.535 ;
        RECT 65.590 142.505 65.760 143.575 ;
        RECT 65.930 142.685 66.120 143.405 ;
        RECT 64.930 142.205 65.760 142.505 ;
        RECT 66.290 142.475 66.610 143.435 ;
        RECT 63.515 141.805 63.850 141.975 ;
        RECT 64.045 141.805 64.720 141.975 ;
        RECT 65.040 141.525 65.410 142.025 ;
        RECT 65.590 141.975 65.760 142.205 ;
        RECT 66.145 142.145 66.610 142.475 ;
        RECT 66.780 142.765 66.950 143.605 ;
        RECT 67.130 143.575 67.445 144.075 ;
        RECT 67.675 143.345 68.015 143.905 ;
        RECT 67.120 142.970 68.015 143.345 ;
        RECT 68.185 143.065 68.355 144.075 ;
        RECT 67.825 142.765 68.015 142.970 ;
        RECT 68.525 143.015 68.855 143.860 ;
        RECT 68.525 142.935 68.915 143.015 ;
        RECT 68.700 142.885 68.915 142.935 ;
        RECT 70.005 142.910 70.295 144.075 ;
        RECT 70.670 143.105 71.000 143.905 ;
        RECT 71.170 143.275 71.500 144.075 ;
        RECT 71.800 143.105 72.130 143.905 ;
        RECT 72.775 143.275 73.025 144.075 ;
        RECT 70.670 142.935 73.105 143.105 ;
        RECT 73.295 142.935 73.465 144.075 ;
        RECT 73.635 142.935 73.975 143.905 ;
        RECT 74.695 143.405 74.865 143.905 ;
        RECT 75.035 143.575 75.365 144.075 ;
        RECT 74.695 143.235 75.360 143.405 ;
        RECT 66.780 142.435 67.655 142.765 ;
        RECT 67.825 142.435 68.575 142.765 ;
        RECT 66.780 141.975 66.950 142.435 ;
        RECT 67.825 142.265 68.025 142.435 ;
        RECT 68.745 142.305 68.915 142.885 ;
        RECT 70.465 142.515 70.815 142.765 ;
        RECT 71.000 142.305 71.170 142.935 ;
        RECT 71.340 142.515 71.670 142.715 ;
        RECT 71.840 142.515 72.170 142.715 ;
        RECT 72.340 142.515 72.760 142.715 ;
        RECT 72.935 142.685 73.105 142.935 ;
        RECT 72.935 142.515 73.630 142.685 ;
        RECT 68.690 142.265 68.915 142.305 ;
        RECT 65.590 141.805 65.995 141.975 ;
        RECT 66.165 141.805 66.950 141.975 ;
        RECT 67.225 141.525 67.435 142.055 ;
        RECT 67.695 141.740 68.025 142.265 ;
        RECT 68.535 142.180 68.915 142.265 ;
        RECT 68.195 141.525 68.365 142.135 ;
        RECT 68.535 141.745 68.865 142.180 ;
        RECT 70.005 141.525 70.295 142.250 ;
        RECT 70.670 141.695 71.170 142.305 ;
        RECT 71.800 142.175 73.025 142.345 ;
        RECT 73.800 142.325 73.975 142.935 ;
        RECT 74.610 142.415 74.960 143.065 ;
        RECT 71.800 141.695 72.130 142.175 ;
        RECT 72.300 141.525 72.525 141.985 ;
        RECT 72.695 141.695 73.025 142.175 ;
        RECT 73.215 141.525 73.465 142.325 ;
        RECT 73.635 141.695 73.975 142.325 ;
        RECT 75.130 142.245 75.360 143.235 ;
        RECT 74.695 142.075 75.360 142.245 ;
        RECT 74.695 141.785 74.865 142.075 ;
        RECT 75.035 141.525 75.365 141.905 ;
        RECT 75.535 141.785 75.720 143.905 ;
        RECT 75.960 143.615 76.225 144.075 ;
        RECT 76.395 143.480 76.645 143.905 ;
        RECT 76.855 143.630 77.960 143.800 ;
        RECT 76.340 143.350 76.645 143.480 ;
        RECT 75.890 142.155 76.170 143.105 ;
        RECT 76.340 142.245 76.510 143.350 ;
        RECT 76.680 142.565 76.920 143.160 ;
        RECT 77.090 143.095 77.620 143.460 ;
        RECT 77.090 142.395 77.260 143.095 ;
        RECT 77.790 143.015 77.960 143.630 ;
        RECT 78.130 143.275 78.300 144.075 ;
        RECT 78.470 143.575 78.720 143.905 ;
        RECT 78.945 143.605 79.830 143.775 ;
        RECT 77.790 142.925 78.300 143.015 ;
        RECT 76.340 142.115 76.565 142.245 ;
        RECT 76.735 142.175 77.260 142.395 ;
        RECT 77.430 142.755 78.300 142.925 ;
        RECT 75.975 141.525 76.225 141.985 ;
        RECT 76.395 141.975 76.565 142.115 ;
        RECT 77.430 141.975 77.600 142.755 ;
        RECT 78.130 142.685 78.300 142.755 ;
        RECT 77.810 142.505 78.010 142.535 ;
        RECT 78.470 142.505 78.640 143.575 ;
        RECT 78.810 142.685 79.000 143.405 ;
        RECT 77.810 142.205 78.640 142.505 ;
        RECT 79.170 142.475 79.490 143.435 ;
        RECT 76.395 141.805 76.730 141.975 ;
        RECT 76.925 141.805 77.600 141.975 ;
        RECT 77.920 141.525 78.290 142.025 ;
        RECT 78.470 141.975 78.640 142.205 ;
        RECT 79.025 142.145 79.490 142.475 ;
        RECT 79.660 142.765 79.830 143.605 ;
        RECT 80.010 143.575 80.325 144.075 ;
        RECT 80.555 143.345 80.895 143.905 ;
        RECT 80.000 142.970 80.895 143.345 ;
        RECT 81.065 143.065 81.235 144.075 ;
        RECT 80.705 142.765 80.895 142.970 ;
        RECT 81.405 143.015 81.735 143.860 ;
        RECT 81.405 142.935 81.795 143.015 ;
        RECT 81.580 142.885 81.795 142.935 ;
        RECT 79.660 142.435 80.535 142.765 ;
        RECT 80.705 142.435 81.455 142.765 ;
        RECT 79.660 141.975 79.830 142.435 ;
        RECT 80.705 142.265 80.905 142.435 ;
        RECT 81.625 142.305 81.795 142.885 ;
        RECT 81.965 142.985 83.175 144.075 ;
        RECT 81.965 142.445 82.485 142.985 ;
        RECT 81.570 142.265 81.795 142.305 ;
        RECT 82.655 142.275 83.175 142.815 ;
        RECT 78.470 141.805 78.875 141.975 ;
        RECT 79.045 141.805 79.830 141.975 ;
        RECT 80.105 141.525 80.315 142.055 ;
        RECT 80.575 141.740 80.905 142.265 ;
        RECT 81.415 142.180 81.795 142.265 ;
        RECT 81.075 141.525 81.245 142.135 ;
        RECT 81.415 141.745 81.745 142.180 ;
        RECT 81.965 141.525 83.175 142.275 ;
        RECT 5.520 141.355 83.260 141.525 ;
        RECT 5.605 140.605 6.815 141.355 ;
        RECT 6.985 140.810 12.330 141.355 ;
        RECT 5.605 140.065 6.125 140.605 ;
        RECT 6.295 139.895 6.815 140.435 ;
        RECT 8.570 139.980 8.910 140.810 ;
        RECT 12.505 140.605 13.715 141.355 ;
        RECT 13.975 140.805 14.145 141.095 ;
        RECT 14.315 140.975 14.645 141.355 ;
        RECT 13.975 140.635 14.640 140.805 ;
        RECT 5.605 138.805 6.815 139.895 ;
        RECT 10.390 139.240 10.740 140.490 ;
        RECT 12.505 140.065 13.025 140.605 ;
        RECT 13.195 139.895 13.715 140.435 ;
        RECT 6.985 138.805 12.330 139.240 ;
        RECT 12.505 138.805 13.715 139.895 ;
        RECT 13.890 139.815 14.240 140.465 ;
        RECT 14.410 139.645 14.640 140.635 ;
        RECT 13.975 139.475 14.640 139.645 ;
        RECT 13.975 138.975 14.145 139.475 ;
        RECT 14.315 138.805 14.645 139.305 ;
        RECT 14.815 138.975 15.000 141.095 ;
        RECT 15.255 140.895 15.505 141.355 ;
        RECT 15.675 140.905 16.010 141.075 ;
        RECT 16.205 140.905 16.880 141.075 ;
        RECT 15.675 140.765 15.845 140.905 ;
        RECT 15.170 139.775 15.450 140.725 ;
        RECT 15.620 140.635 15.845 140.765 ;
        RECT 15.620 139.530 15.790 140.635 ;
        RECT 16.015 140.485 16.540 140.705 ;
        RECT 15.960 139.720 16.200 140.315 ;
        RECT 16.370 139.785 16.540 140.485 ;
        RECT 16.710 140.125 16.880 140.905 ;
        RECT 17.200 140.855 17.570 141.355 ;
        RECT 17.750 140.905 18.155 141.075 ;
        RECT 18.325 140.905 19.110 141.075 ;
        RECT 17.750 140.675 17.920 140.905 ;
        RECT 17.090 140.375 17.920 140.675 ;
        RECT 18.305 140.405 18.770 140.735 ;
        RECT 17.090 140.345 17.290 140.375 ;
        RECT 17.410 140.125 17.580 140.195 ;
        RECT 16.710 139.955 17.580 140.125 ;
        RECT 17.070 139.865 17.580 139.955 ;
        RECT 15.620 139.400 15.925 139.530 ;
        RECT 16.370 139.420 16.900 139.785 ;
        RECT 15.240 138.805 15.505 139.265 ;
        RECT 15.675 138.975 15.925 139.400 ;
        RECT 17.070 139.250 17.240 139.865 ;
        RECT 16.135 139.080 17.240 139.250 ;
        RECT 17.410 138.805 17.580 139.605 ;
        RECT 17.750 139.305 17.920 140.375 ;
        RECT 18.090 139.475 18.280 140.195 ;
        RECT 18.450 139.445 18.770 140.405 ;
        RECT 18.940 140.445 19.110 140.905 ;
        RECT 19.385 140.825 19.595 141.355 ;
        RECT 19.855 140.615 20.185 141.140 ;
        RECT 20.355 140.745 20.525 141.355 ;
        RECT 20.695 140.700 21.025 141.135 ;
        RECT 20.695 140.615 21.075 140.700 ;
        RECT 19.985 140.445 20.185 140.615 ;
        RECT 20.850 140.575 21.075 140.615 ;
        RECT 18.940 140.115 19.815 140.445 ;
        RECT 19.985 140.115 20.735 140.445 ;
        RECT 17.750 138.975 18.000 139.305 ;
        RECT 18.940 139.275 19.110 140.115 ;
        RECT 19.985 139.910 20.175 140.115 ;
        RECT 20.905 139.995 21.075 140.575 ;
        RECT 21.265 140.545 21.505 141.355 ;
        RECT 21.675 140.545 22.005 141.185 ;
        RECT 22.175 140.545 22.445 141.355 ;
        RECT 22.625 140.810 27.970 141.355 ;
        RECT 21.245 140.115 21.595 140.365 ;
        RECT 20.860 139.945 21.075 139.995 ;
        RECT 21.765 139.945 21.935 140.545 ;
        RECT 22.105 140.115 22.455 140.365 ;
        RECT 24.210 139.980 24.550 140.810 ;
        RECT 28.145 140.585 30.735 141.355 ;
        RECT 31.365 140.630 31.655 141.355 ;
        RECT 31.825 140.585 33.495 141.355 ;
        RECT 19.280 139.535 20.175 139.910 ;
        RECT 20.685 139.865 21.075 139.945 ;
        RECT 18.225 139.105 19.110 139.275 ;
        RECT 19.290 138.805 19.605 139.305 ;
        RECT 19.835 138.975 20.175 139.535 ;
        RECT 20.345 138.805 20.515 139.815 ;
        RECT 20.685 139.020 21.015 139.865 ;
        RECT 21.255 139.775 21.935 139.945 ;
        RECT 21.255 138.990 21.585 139.775 ;
        RECT 22.115 138.805 22.445 139.945 ;
        RECT 26.030 139.240 26.380 140.490 ;
        RECT 28.145 140.065 29.355 140.585 ;
        RECT 29.525 139.895 30.735 140.415 ;
        RECT 31.825 140.065 32.575 140.585 ;
        RECT 33.665 140.555 33.975 141.355 ;
        RECT 34.180 140.555 34.875 141.185 ;
        RECT 35.045 140.630 35.305 141.185 ;
        RECT 35.475 140.910 35.905 141.355 ;
        RECT 36.140 140.785 36.310 141.185 ;
        RECT 36.480 140.955 37.200 141.355 ;
        RECT 34.180 140.505 34.355 140.555 ;
        RECT 22.625 138.805 27.970 139.240 ;
        RECT 28.145 138.805 30.735 139.895 ;
        RECT 31.365 138.805 31.655 139.970 ;
        RECT 32.745 139.895 33.495 140.415 ;
        RECT 33.675 140.115 34.010 140.385 ;
        RECT 34.180 139.955 34.350 140.505 ;
        RECT 34.520 140.115 34.855 140.365 ;
        RECT 31.825 138.805 33.495 139.895 ;
        RECT 33.665 138.805 33.945 139.945 ;
        RECT 34.115 138.975 34.445 139.955 ;
        RECT 34.615 138.805 34.875 139.945 ;
        RECT 35.045 139.915 35.220 140.630 ;
        RECT 36.140 140.615 37.020 140.785 ;
        RECT 37.370 140.740 37.540 141.185 ;
        RECT 38.115 140.845 38.515 141.355 ;
        RECT 35.390 140.115 35.645 140.445 ;
        RECT 35.045 138.975 35.305 139.915 ;
        RECT 35.475 139.635 35.645 140.115 ;
        RECT 35.870 139.825 36.200 140.445 ;
        RECT 36.370 140.065 36.660 140.445 ;
        RECT 36.850 139.895 37.020 140.615 ;
        RECT 36.500 139.725 37.020 139.895 ;
        RECT 37.190 140.570 37.540 140.740 ;
        RECT 35.475 139.465 36.235 139.635 ;
        RECT 36.500 139.535 36.670 139.725 ;
        RECT 37.190 139.545 37.360 140.570 ;
        RECT 37.780 140.085 38.040 140.675 ;
        RECT 37.560 139.785 38.040 140.085 ;
        RECT 38.240 139.785 38.500 140.675 ;
        RECT 38.760 140.615 39.375 141.185 ;
        RECT 39.545 140.845 39.760 141.355 ;
        RECT 39.990 140.845 40.270 141.175 ;
        RECT 40.450 140.845 40.690 141.355 ;
        RECT 36.065 139.240 36.235 139.465 ;
        RECT 36.950 139.375 37.360 139.545 ;
        RECT 37.535 139.435 38.475 139.605 ;
        RECT 36.950 139.240 37.205 139.375 ;
        RECT 35.475 138.805 35.805 139.205 ;
        RECT 36.065 139.070 37.205 139.240 ;
        RECT 37.535 139.185 37.705 139.435 ;
        RECT 36.950 138.975 37.205 139.070 ;
        RECT 37.375 139.015 37.705 139.185 ;
        RECT 37.875 138.805 38.125 139.265 ;
        RECT 38.295 138.975 38.475 139.435 ;
        RECT 38.760 139.595 39.075 140.615 ;
        RECT 39.245 139.945 39.415 140.445 ;
        RECT 39.665 140.115 39.930 140.675 ;
        RECT 40.100 139.945 40.270 140.845 ;
        RECT 41.025 140.680 41.285 141.185 ;
        RECT 41.465 140.975 41.795 141.355 ;
        RECT 41.975 140.805 42.145 141.185 ;
        RECT 40.440 140.115 40.795 140.675 ;
        RECT 39.245 139.775 40.670 139.945 ;
        RECT 38.760 138.975 39.295 139.595 ;
        RECT 39.465 138.805 39.795 139.605 ;
        RECT 40.280 139.600 40.670 139.775 ;
        RECT 41.025 139.880 41.205 140.680 ;
        RECT 41.480 140.635 42.145 140.805 ;
        RECT 41.480 140.380 41.650 140.635 ;
        RECT 42.405 140.605 43.615 141.355 ;
        RECT 43.790 140.615 44.045 141.185 ;
        RECT 44.215 140.955 44.545 141.355 ;
        RECT 44.970 140.820 45.500 141.185 ;
        RECT 44.970 140.785 45.145 140.820 ;
        RECT 44.215 140.615 45.145 140.785 ;
        RECT 41.375 140.050 41.650 140.380 ;
        RECT 41.875 140.085 42.215 140.455 ;
        RECT 42.405 140.065 42.925 140.605 ;
        RECT 41.480 139.905 41.650 140.050 ;
        RECT 41.025 138.975 41.295 139.880 ;
        RECT 41.480 139.735 42.155 139.905 ;
        RECT 43.095 139.895 43.615 140.435 ;
        RECT 41.465 138.805 41.795 139.565 ;
        RECT 41.975 138.975 42.155 139.735 ;
        RECT 42.405 138.805 43.615 139.895 ;
        RECT 43.790 139.945 43.960 140.615 ;
        RECT 44.215 140.445 44.385 140.615 ;
        RECT 44.130 140.115 44.385 140.445 ;
        RECT 44.610 140.115 44.805 140.445 ;
        RECT 43.790 138.975 44.125 139.945 ;
        RECT 44.295 138.805 44.465 139.945 ;
        RECT 44.635 139.145 44.805 140.115 ;
        RECT 44.975 139.485 45.145 140.615 ;
        RECT 45.315 139.825 45.485 140.625 ;
        RECT 45.690 140.335 45.965 141.185 ;
        RECT 45.685 140.165 45.965 140.335 ;
        RECT 45.690 140.025 45.965 140.165 ;
        RECT 46.135 139.825 46.325 141.185 ;
        RECT 46.505 140.820 47.015 141.355 ;
        RECT 47.235 140.545 47.480 141.150 ;
        RECT 47.925 140.585 51.435 141.355 ;
        RECT 51.605 140.605 52.815 141.355 ;
        RECT 52.990 140.615 53.245 141.185 ;
        RECT 53.415 140.955 53.745 141.355 ;
        RECT 54.170 140.820 54.700 141.185 ;
        RECT 54.890 141.015 55.165 141.185 ;
        RECT 54.885 140.845 55.165 141.015 ;
        RECT 54.170 140.785 54.345 140.820 ;
        RECT 53.415 140.615 54.345 140.785 ;
        RECT 46.525 140.375 47.755 140.545 ;
        RECT 45.315 139.655 46.325 139.825 ;
        RECT 46.495 139.810 47.245 140.000 ;
        RECT 44.975 139.315 46.100 139.485 ;
        RECT 46.495 139.145 46.665 139.810 ;
        RECT 47.415 139.565 47.755 140.375 ;
        RECT 47.925 140.065 49.575 140.585 ;
        RECT 49.745 139.895 51.435 140.415 ;
        RECT 51.605 140.065 52.125 140.605 ;
        RECT 52.295 139.895 52.815 140.435 ;
        RECT 44.635 138.975 46.665 139.145 ;
        RECT 46.835 138.805 47.005 139.565 ;
        RECT 47.240 139.155 47.755 139.565 ;
        RECT 47.925 138.805 51.435 139.895 ;
        RECT 51.605 138.805 52.815 139.895 ;
        RECT 52.990 139.945 53.160 140.615 ;
        RECT 53.415 140.445 53.585 140.615 ;
        RECT 53.330 140.115 53.585 140.445 ;
        RECT 53.810 140.115 54.005 140.445 ;
        RECT 52.990 138.975 53.325 139.945 ;
        RECT 53.495 138.805 53.665 139.945 ;
        RECT 53.835 139.145 54.005 140.115 ;
        RECT 54.175 139.485 54.345 140.615 ;
        RECT 54.515 139.825 54.685 140.625 ;
        RECT 54.890 140.025 55.165 140.845 ;
        RECT 55.335 139.825 55.525 141.185 ;
        RECT 55.705 140.820 56.215 141.355 ;
        RECT 56.435 140.545 56.680 141.150 ;
        RECT 57.125 140.630 57.415 141.355 ;
        RECT 57.635 140.700 57.965 141.135 ;
        RECT 58.135 140.745 58.305 141.355 ;
        RECT 57.585 140.615 57.965 140.700 ;
        RECT 58.475 140.615 58.805 141.140 ;
        RECT 59.065 140.825 59.275 141.355 ;
        RECT 59.550 140.905 60.335 141.075 ;
        RECT 60.505 140.905 60.910 141.075 ;
        RECT 57.585 140.575 57.810 140.615 ;
        RECT 55.725 140.375 56.955 140.545 ;
        RECT 54.515 139.655 55.525 139.825 ;
        RECT 55.695 139.810 56.445 140.000 ;
        RECT 54.175 139.315 55.300 139.485 ;
        RECT 55.695 139.145 55.865 139.810 ;
        RECT 56.615 139.565 56.955 140.375 ;
        RECT 57.585 139.995 57.755 140.575 ;
        RECT 58.475 140.445 58.675 140.615 ;
        RECT 59.550 140.445 59.720 140.905 ;
        RECT 57.925 140.115 58.675 140.445 ;
        RECT 58.845 140.115 59.720 140.445 ;
        RECT 53.835 138.975 55.865 139.145 ;
        RECT 56.035 138.805 56.205 139.565 ;
        RECT 56.440 139.155 56.955 139.565 ;
        RECT 57.125 138.805 57.415 139.970 ;
        RECT 57.585 139.945 57.800 139.995 ;
        RECT 57.585 139.865 57.975 139.945 ;
        RECT 57.645 139.020 57.975 139.865 ;
        RECT 58.485 139.910 58.675 140.115 ;
        RECT 58.145 138.805 58.315 139.815 ;
        RECT 58.485 139.535 59.380 139.910 ;
        RECT 58.485 138.975 58.825 139.535 ;
        RECT 59.055 138.805 59.370 139.305 ;
        RECT 59.550 139.275 59.720 140.115 ;
        RECT 59.890 140.405 60.355 140.735 ;
        RECT 60.740 140.675 60.910 140.905 ;
        RECT 61.090 140.855 61.460 141.355 ;
        RECT 61.780 140.905 62.455 141.075 ;
        RECT 62.650 140.905 62.985 141.075 ;
        RECT 59.890 139.445 60.210 140.405 ;
        RECT 60.740 140.375 61.570 140.675 ;
        RECT 60.380 139.475 60.570 140.195 ;
        RECT 60.740 139.305 60.910 140.375 ;
        RECT 61.370 140.345 61.570 140.375 ;
        RECT 61.080 140.125 61.250 140.195 ;
        RECT 61.780 140.125 61.950 140.905 ;
        RECT 62.815 140.765 62.985 140.905 ;
        RECT 63.155 140.895 63.405 141.355 ;
        RECT 61.080 139.955 61.950 140.125 ;
        RECT 62.120 140.485 62.645 140.705 ;
        RECT 62.815 140.635 63.040 140.765 ;
        RECT 61.080 139.865 61.590 139.955 ;
        RECT 59.550 139.105 60.435 139.275 ;
        RECT 60.660 138.975 60.910 139.305 ;
        RECT 61.080 138.805 61.250 139.605 ;
        RECT 61.420 139.250 61.590 139.865 ;
        RECT 62.120 139.785 62.290 140.485 ;
        RECT 61.760 139.420 62.290 139.785 ;
        RECT 62.460 139.720 62.700 140.315 ;
        RECT 62.870 139.530 63.040 140.635 ;
        RECT 63.210 139.775 63.490 140.725 ;
        RECT 62.735 139.400 63.040 139.530 ;
        RECT 61.420 139.080 62.525 139.250 ;
        RECT 62.735 138.975 62.985 139.400 ;
        RECT 63.155 138.805 63.420 139.265 ;
        RECT 63.660 138.975 63.845 141.095 ;
        RECT 64.015 140.975 64.345 141.355 ;
        RECT 64.515 140.805 64.685 141.095 ;
        RECT 64.020 140.635 64.685 140.805 ;
        RECT 64.020 139.645 64.250 140.635 ;
        RECT 64.950 140.615 65.205 141.185 ;
        RECT 65.375 140.955 65.705 141.355 ;
        RECT 66.130 140.820 66.660 141.185 ;
        RECT 66.850 141.015 67.125 141.185 ;
        RECT 66.845 140.845 67.125 141.015 ;
        RECT 66.130 140.785 66.305 140.820 ;
        RECT 65.375 140.615 66.305 140.785 ;
        RECT 64.420 139.815 64.770 140.465 ;
        RECT 64.950 139.945 65.120 140.615 ;
        RECT 65.375 140.445 65.545 140.615 ;
        RECT 65.290 140.115 65.545 140.445 ;
        RECT 65.770 140.115 65.965 140.445 ;
        RECT 64.020 139.475 64.685 139.645 ;
        RECT 64.015 138.805 64.345 139.305 ;
        RECT 64.515 138.975 64.685 139.475 ;
        RECT 64.950 138.975 65.285 139.945 ;
        RECT 65.455 138.805 65.625 139.945 ;
        RECT 65.795 139.145 65.965 140.115 ;
        RECT 66.135 139.485 66.305 140.615 ;
        RECT 66.475 139.825 66.645 140.625 ;
        RECT 66.850 140.025 67.125 140.845 ;
        RECT 67.295 139.825 67.485 141.185 ;
        RECT 67.665 140.820 68.175 141.355 ;
        RECT 68.395 140.545 68.640 141.150 ;
        RECT 69.085 140.615 69.470 141.185 ;
        RECT 69.640 140.895 69.965 141.355 ;
        RECT 70.485 140.725 70.765 141.185 ;
        RECT 67.685 140.375 68.915 140.545 ;
        RECT 66.475 139.655 67.485 139.825 ;
        RECT 67.655 139.810 68.405 140.000 ;
        RECT 66.135 139.315 67.260 139.485 ;
        RECT 67.655 139.145 67.825 139.810 ;
        RECT 68.575 139.565 68.915 140.375 ;
        RECT 65.795 138.975 67.825 139.145 ;
        RECT 67.995 138.805 68.165 139.565 ;
        RECT 68.400 139.155 68.915 139.565 ;
        RECT 69.085 139.945 69.365 140.615 ;
        RECT 69.640 140.555 70.765 140.725 ;
        RECT 69.640 140.445 70.090 140.555 ;
        RECT 69.535 140.115 70.090 140.445 ;
        RECT 70.955 140.385 71.355 141.185 ;
        RECT 71.755 140.895 72.025 141.355 ;
        RECT 72.195 140.725 72.480 141.185 ;
        RECT 69.085 138.975 69.470 139.945 ;
        RECT 69.640 139.655 70.090 140.115 ;
        RECT 70.260 139.825 71.355 140.385 ;
        RECT 69.640 139.435 70.765 139.655 ;
        RECT 69.640 138.805 69.965 139.265 ;
        RECT 70.485 138.975 70.765 139.435 ;
        RECT 70.955 138.975 71.355 139.825 ;
        RECT 71.525 140.555 72.480 140.725 ;
        RECT 72.765 140.615 73.150 141.185 ;
        RECT 73.320 140.895 73.645 141.355 ;
        RECT 74.165 140.725 74.445 141.185 ;
        RECT 71.525 139.655 71.735 140.555 ;
        RECT 71.905 139.825 72.595 140.385 ;
        RECT 72.765 139.945 73.045 140.615 ;
        RECT 73.320 140.555 74.445 140.725 ;
        RECT 73.320 140.445 73.770 140.555 ;
        RECT 73.215 140.115 73.770 140.445 ;
        RECT 74.635 140.385 75.035 141.185 ;
        RECT 75.435 140.895 75.705 141.355 ;
        RECT 75.875 140.725 76.160 141.185 ;
        RECT 71.525 139.435 72.480 139.655 ;
        RECT 71.755 138.805 72.025 139.265 ;
        RECT 72.195 138.975 72.480 139.435 ;
        RECT 72.765 138.975 73.150 139.945 ;
        RECT 73.320 139.655 73.770 140.115 ;
        RECT 73.940 139.825 75.035 140.385 ;
        RECT 73.320 139.435 74.445 139.655 ;
        RECT 73.320 138.805 73.645 139.265 ;
        RECT 74.165 138.975 74.445 139.435 ;
        RECT 74.635 138.975 75.035 139.825 ;
        RECT 75.205 140.555 76.160 140.725 ;
        RECT 76.445 140.555 76.785 141.185 ;
        RECT 76.955 140.555 77.205 141.355 ;
        RECT 77.395 140.705 77.725 141.185 ;
        RECT 77.895 140.895 78.120 141.355 ;
        RECT 78.290 140.705 78.620 141.185 ;
        RECT 75.205 139.655 75.415 140.555 ;
        RECT 75.585 139.825 76.275 140.385 ;
        RECT 76.445 139.945 76.620 140.555 ;
        RECT 77.395 140.535 78.620 140.705 ;
        RECT 79.250 140.575 79.750 141.185 ;
        RECT 80.215 140.805 80.385 141.185 ;
        RECT 80.600 140.975 80.930 141.355 ;
        RECT 80.215 140.635 80.930 140.805 ;
        RECT 76.790 140.195 77.485 140.365 ;
        RECT 77.315 139.945 77.485 140.195 ;
        RECT 77.660 140.165 78.080 140.365 ;
        RECT 78.250 140.165 78.580 140.365 ;
        RECT 78.750 140.165 79.080 140.365 ;
        RECT 79.250 139.945 79.420 140.575 ;
        RECT 79.605 140.115 79.955 140.365 ;
        RECT 80.125 140.085 80.480 140.455 ;
        RECT 80.760 140.445 80.930 140.635 ;
        RECT 81.100 140.610 81.355 141.185 ;
        RECT 80.760 140.115 81.015 140.445 ;
        RECT 75.205 139.435 76.160 139.655 ;
        RECT 75.435 138.805 75.705 139.265 ;
        RECT 75.875 138.975 76.160 139.435 ;
        RECT 76.445 138.975 76.785 139.945 ;
        RECT 76.955 138.805 77.125 139.945 ;
        RECT 77.315 139.775 79.750 139.945 ;
        RECT 80.760 139.905 80.930 140.115 ;
        RECT 77.395 138.805 77.645 139.605 ;
        RECT 78.290 138.975 78.620 139.775 ;
        RECT 78.920 138.805 79.250 139.605 ;
        RECT 79.420 138.975 79.750 139.775 ;
        RECT 80.215 139.735 80.930 139.905 ;
        RECT 81.185 139.880 81.355 140.610 ;
        RECT 81.530 140.515 81.790 141.355 ;
        RECT 81.965 140.605 83.175 141.355 ;
        RECT 80.215 138.975 80.385 139.735 ;
        RECT 80.600 138.805 80.930 139.565 ;
        RECT 81.100 138.975 81.355 139.880 ;
        RECT 81.530 138.805 81.790 139.955 ;
        RECT 81.965 139.895 82.485 140.435 ;
        RECT 82.655 140.065 83.175 140.605 ;
        RECT 81.965 138.805 83.175 139.895 ;
        RECT 5.520 138.635 83.260 138.805 ;
        RECT 5.605 137.545 6.815 138.635 ;
        RECT 6.985 137.545 9.575 138.635 ;
        RECT 10.295 137.965 10.465 138.465 ;
        RECT 10.635 138.135 10.965 138.635 ;
        RECT 10.295 137.795 10.960 137.965 ;
        RECT 5.605 136.835 6.125 137.375 ;
        RECT 6.295 137.005 6.815 137.545 ;
        RECT 6.985 136.855 8.195 137.375 ;
        RECT 8.365 137.025 9.575 137.545 ;
        RECT 10.210 136.975 10.560 137.625 ;
        RECT 5.605 136.085 6.815 136.835 ;
        RECT 6.985 136.085 9.575 136.855 ;
        RECT 10.730 136.805 10.960 137.795 ;
        RECT 10.295 136.635 10.960 136.805 ;
        RECT 10.295 136.345 10.465 136.635 ;
        RECT 10.635 136.085 10.965 136.465 ;
        RECT 11.135 136.345 11.320 138.465 ;
        RECT 11.560 138.175 11.825 138.635 ;
        RECT 11.995 138.040 12.245 138.465 ;
        RECT 12.455 138.190 13.560 138.360 ;
        RECT 11.940 137.910 12.245 138.040 ;
        RECT 11.490 136.715 11.770 137.665 ;
        RECT 11.940 136.805 12.110 137.910 ;
        RECT 12.280 137.125 12.520 137.720 ;
        RECT 12.690 137.655 13.220 138.020 ;
        RECT 12.690 136.955 12.860 137.655 ;
        RECT 13.390 137.575 13.560 138.190 ;
        RECT 13.730 137.835 13.900 138.635 ;
        RECT 14.070 138.135 14.320 138.465 ;
        RECT 14.545 138.165 15.430 138.335 ;
        RECT 13.390 137.485 13.900 137.575 ;
        RECT 11.940 136.675 12.165 136.805 ;
        RECT 12.335 136.735 12.860 136.955 ;
        RECT 13.030 137.315 13.900 137.485 ;
        RECT 11.575 136.085 11.825 136.545 ;
        RECT 11.995 136.535 12.165 136.675 ;
        RECT 13.030 136.535 13.200 137.315 ;
        RECT 13.730 137.245 13.900 137.315 ;
        RECT 13.410 137.065 13.610 137.095 ;
        RECT 14.070 137.065 14.240 138.135 ;
        RECT 14.410 137.245 14.600 137.965 ;
        RECT 13.410 136.765 14.240 137.065 ;
        RECT 14.770 137.035 15.090 137.995 ;
        RECT 11.995 136.365 12.330 136.535 ;
        RECT 12.525 136.365 13.200 136.535 ;
        RECT 13.520 136.085 13.890 136.585 ;
        RECT 14.070 136.535 14.240 136.765 ;
        RECT 14.625 136.705 15.090 137.035 ;
        RECT 15.260 137.325 15.430 138.165 ;
        RECT 15.610 138.135 15.925 138.635 ;
        RECT 16.155 137.905 16.495 138.465 ;
        RECT 15.600 137.530 16.495 137.905 ;
        RECT 16.665 137.625 16.835 138.635 ;
        RECT 16.305 137.325 16.495 137.530 ;
        RECT 17.005 137.575 17.335 138.420 ;
        RECT 17.005 137.495 17.395 137.575 ;
        RECT 17.180 137.445 17.395 137.495 ;
        RECT 18.485 137.470 18.775 138.635 ;
        RECT 18.955 137.665 19.285 138.450 ;
        RECT 18.955 137.495 19.635 137.665 ;
        RECT 19.815 137.495 20.145 138.635 ;
        RECT 20.415 137.965 20.585 138.465 ;
        RECT 20.755 138.135 21.085 138.635 ;
        RECT 20.415 137.795 21.080 137.965 ;
        RECT 15.260 136.995 16.135 137.325 ;
        RECT 16.305 136.995 17.055 137.325 ;
        RECT 15.260 136.535 15.430 136.995 ;
        RECT 16.305 136.825 16.505 136.995 ;
        RECT 17.225 136.865 17.395 137.445 ;
        RECT 18.945 137.075 19.295 137.325 ;
        RECT 19.465 136.895 19.635 137.495 ;
        RECT 19.805 137.075 20.155 137.325 ;
        RECT 20.330 136.975 20.680 137.625 ;
        RECT 17.170 136.825 17.395 136.865 ;
        RECT 14.070 136.365 14.475 136.535 ;
        RECT 14.645 136.365 15.430 136.535 ;
        RECT 15.705 136.085 15.915 136.615 ;
        RECT 16.175 136.300 16.505 136.825 ;
        RECT 17.015 136.740 17.395 136.825 ;
        RECT 16.675 136.085 16.845 136.695 ;
        RECT 17.015 136.305 17.345 136.740 ;
        RECT 18.485 136.085 18.775 136.810 ;
        RECT 18.965 136.085 19.205 136.895 ;
        RECT 19.375 136.255 19.705 136.895 ;
        RECT 19.875 136.085 20.145 136.895 ;
        RECT 20.850 136.805 21.080 137.795 ;
        RECT 20.415 136.635 21.080 136.805 ;
        RECT 20.415 136.345 20.585 136.635 ;
        RECT 20.755 136.085 21.085 136.465 ;
        RECT 21.255 136.345 21.440 138.465 ;
        RECT 21.680 138.175 21.945 138.635 ;
        RECT 22.115 138.040 22.365 138.465 ;
        RECT 22.575 138.190 23.680 138.360 ;
        RECT 22.060 137.910 22.365 138.040 ;
        RECT 21.610 136.715 21.890 137.665 ;
        RECT 22.060 136.805 22.230 137.910 ;
        RECT 22.400 137.125 22.640 137.720 ;
        RECT 22.810 137.655 23.340 138.020 ;
        RECT 22.810 136.955 22.980 137.655 ;
        RECT 23.510 137.575 23.680 138.190 ;
        RECT 23.850 137.835 24.020 138.635 ;
        RECT 24.190 138.135 24.440 138.465 ;
        RECT 24.665 138.165 25.550 138.335 ;
        RECT 23.510 137.485 24.020 137.575 ;
        RECT 22.060 136.675 22.285 136.805 ;
        RECT 22.455 136.735 22.980 136.955 ;
        RECT 23.150 137.315 24.020 137.485 ;
        RECT 21.695 136.085 21.945 136.545 ;
        RECT 22.115 136.535 22.285 136.675 ;
        RECT 23.150 136.535 23.320 137.315 ;
        RECT 23.850 137.245 24.020 137.315 ;
        RECT 23.530 137.065 23.730 137.095 ;
        RECT 24.190 137.065 24.360 138.135 ;
        RECT 24.530 137.245 24.720 137.965 ;
        RECT 23.530 136.765 24.360 137.065 ;
        RECT 24.890 137.035 25.210 137.995 ;
        RECT 22.115 136.365 22.450 136.535 ;
        RECT 22.645 136.365 23.320 136.535 ;
        RECT 23.640 136.085 24.010 136.585 ;
        RECT 24.190 136.535 24.360 136.765 ;
        RECT 24.745 136.705 25.210 137.035 ;
        RECT 25.380 137.325 25.550 138.165 ;
        RECT 25.730 138.135 26.045 138.635 ;
        RECT 26.275 137.905 26.615 138.465 ;
        RECT 25.720 137.530 26.615 137.905 ;
        RECT 26.785 137.625 26.955 138.635 ;
        RECT 26.425 137.325 26.615 137.530 ;
        RECT 27.125 137.575 27.455 138.420 ;
        RECT 27.775 137.965 27.945 138.465 ;
        RECT 28.115 138.135 28.445 138.635 ;
        RECT 27.775 137.795 28.440 137.965 ;
        RECT 27.125 137.495 27.515 137.575 ;
        RECT 27.300 137.445 27.515 137.495 ;
        RECT 25.380 136.995 26.255 137.325 ;
        RECT 26.425 136.995 27.175 137.325 ;
        RECT 25.380 136.535 25.550 136.995 ;
        RECT 26.425 136.825 26.625 136.995 ;
        RECT 27.345 136.865 27.515 137.445 ;
        RECT 27.690 136.975 28.040 137.625 ;
        RECT 27.290 136.825 27.515 136.865 ;
        RECT 24.190 136.365 24.595 136.535 ;
        RECT 24.765 136.365 25.550 136.535 ;
        RECT 25.825 136.085 26.035 136.615 ;
        RECT 26.295 136.300 26.625 136.825 ;
        RECT 27.135 136.740 27.515 136.825 ;
        RECT 28.210 136.805 28.440 137.795 ;
        RECT 26.795 136.085 26.965 136.695 ;
        RECT 27.135 136.305 27.465 136.740 ;
        RECT 27.775 136.635 28.440 136.805 ;
        RECT 27.775 136.345 27.945 136.635 ;
        RECT 28.115 136.085 28.445 136.465 ;
        RECT 28.615 136.345 28.800 138.465 ;
        RECT 29.040 138.175 29.305 138.635 ;
        RECT 29.475 138.040 29.725 138.465 ;
        RECT 29.935 138.190 31.040 138.360 ;
        RECT 29.420 137.910 29.725 138.040 ;
        RECT 28.970 136.715 29.250 137.665 ;
        RECT 29.420 136.805 29.590 137.910 ;
        RECT 29.760 137.125 30.000 137.720 ;
        RECT 30.170 137.655 30.700 138.020 ;
        RECT 30.170 136.955 30.340 137.655 ;
        RECT 30.870 137.575 31.040 138.190 ;
        RECT 31.210 137.835 31.380 138.635 ;
        RECT 31.550 138.135 31.800 138.465 ;
        RECT 32.025 138.165 32.910 138.335 ;
        RECT 30.870 137.485 31.380 137.575 ;
        RECT 29.420 136.675 29.645 136.805 ;
        RECT 29.815 136.735 30.340 136.955 ;
        RECT 30.510 137.315 31.380 137.485 ;
        RECT 29.055 136.085 29.305 136.545 ;
        RECT 29.475 136.535 29.645 136.675 ;
        RECT 30.510 136.535 30.680 137.315 ;
        RECT 31.210 137.245 31.380 137.315 ;
        RECT 30.890 137.065 31.090 137.095 ;
        RECT 31.550 137.065 31.720 138.135 ;
        RECT 31.890 137.245 32.080 137.965 ;
        RECT 30.890 136.765 31.720 137.065 ;
        RECT 32.250 137.035 32.570 137.995 ;
        RECT 29.475 136.365 29.810 136.535 ;
        RECT 30.005 136.365 30.680 136.535 ;
        RECT 31.000 136.085 31.370 136.585 ;
        RECT 31.550 136.535 31.720 136.765 ;
        RECT 32.105 136.705 32.570 137.035 ;
        RECT 32.740 137.325 32.910 138.165 ;
        RECT 33.090 138.135 33.405 138.635 ;
        RECT 33.635 137.905 33.975 138.465 ;
        RECT 33.080 137.530 33.975 137.905 ;
        RECT 34.145 137.625 34.315 138.635 ;
        RECT 33.785 137.325 33.975 137.530 ;
        RECT 34.485 137.575 34.815 138.420 ;
        RECT 34.485 137.495 34.875 137.575 ;
        RECT 34.660 137.445 34.875 137.495 ;
        RECT 32.740 136.995 33.615 137.325 ;
        RECT 33.785 136.995 34.535 137.325 ;
        RECT 32.740 136.535 32.910 136.995 ;
        RECT 33.785 136.825 33.985 136.995 ;
        RECT 34.705 136.865 34.875 137.445 ;
        RECT 34.650 136.825 34.875 136.865 ;
        RECT 31.550 136.365 31.955 136.535 ;
        RECT 32.125 136.365 32.910 136.535 ;
        RECT 33.185 136.085 33.395 136.615 ;
        RECT 33.655 136.300 33.985 136.825 ;
        RECT 34.495 136.740 34.875 136.825 ;
        RECT 35.045 137.495 35.430 138.465 ;
        RECT 35.600 138.175 35.925 138.635 ;
        RECT 36.445 138.005 36.725 138.465 ;
        RECT 35.600 137.785 36.725 138.005 ;
        RECT 35.045 136.825 35.325 137.495 ;
        RECT 35.600 137.325 36.050 137.785 ;
        RECT 36.915 137.615 37.315 138.465 ;
        RECT 37.715 138.175 37.985 138.635 ;
        RECT 38.155 138.005 38.440 138.465 ;
        RECT 35.495 136.995 36.050 137.325 ;
        RECT 36.220 137.055 37.315 137.615 ;
        RECT 35.600 136.885 36.050 136.995 ;
        RECT 34.155 136.085 34.325 136.695 ;
        RECT 34.495 136.305 34.825 136.740 ;
        RECT 35.045 136.255 35.430 136.825 ;
        RECT 35.600 136.715 36.725 136.885 ;
        RECT 35.600 136.085 35.925 136.545 ;
        RECT 36.445 136.255 36.725 136.715 ;
        RECT 36.915 136.255 37.315 137.055 ;
        RECT 37.485 137.785 38.440 138.005 ;
        RECT 37.485 136.885 37.695 137.785 ;
        RECT 37.865 137.055 38.555 137.615 ;
        RECT 38.725 137.545 40.395 138.635 ;
        RECT 37.485 136.715 38.440 136.885 ;
        RECT 37.715 136.085 37.985 136.545 ;
        RECT 38.155 136.255 38.440 136.715 ;
        RECT 38.725 136.855 39.475 137.375 ;
        RECT 39.645 137.025 40.395 137.545 ;
        RECT 40.565 137.495 40.950 138.465 ;
        RECT 41.120 138.175 41.445 138.635 ;
        RECT 41.965 138.005 42.245 138.465 ;
        RECT 41.120 137.785 42.245 138.005 ;
        RECT 38.725 136.085 40.395 136.855 ;
        RECT 40.565 136.825 40.845 137.495 ;
        RECT 41.120 137.325 41.570 137.785 ;
        RECT 42.435 137.615 42.835 138.465 ;
        RECT 43.235 138.175 43.505 138.635 ;
        RECT 43.675 138.005 43.960 138.465 ;
        RECT 41.015 136.995 41.570 137.325 ;
        RECT 41.740 137.055 42.835 137.615 ;
        RECT 41.120 136.885 41.570 136.995 ;
        RECT 40.565 136.255 40.950 136.825 ;
        RECT 41.120 136.715 42.245 136.885 ;
        RECT 41.120 136.085 41.445 136.545 ;
        RECT 41.965 136.255 42.245 136.715 ;
        RECT 42.435 136.255 42.835 137.055 ;
        RECT 43.005 137.785 43.960 138.005 ;
        RECT 43.005 136.885 43.215 137.785 ;
        RECT 43.385 137.055 44.075 137.615 ;
        RECT 44.245 137.470 44.535 138.635 ;
        RECT 44.715 137.665 45.045 138.450 ;
        RECT 44.715 137.495 45.395 137.665 ;
        RECT 45.575 137.495 45.905 138.635 ;
        RECT 46.085 137.545 47.755 138.635 ;
        RECT 48.015 137.965 48.185 138.465 ;
        RECT 48.355 138.135 48.685 138.635 ;
        RECT 48.015 137.795 48.680 137.965 ;
        RECT 44.705 137.075 45.055 137.325 ;
        RECT 45.225 136.895 45.395 137.495 ;
        RECT 45.565 137.075 45.915 137.325 ;
        RECT 43.005 136.715 43.960 136.885 ;
        RECT 43.235 136.085 43.505 136.545 ;
        RECT 43.675 136.255 43.960 136.715 ;
        RECT 44.245 136.085 44.535 136.810 ;
        RECT 44.725 136.085 44.965 136.895 ;
        RECT 45.135 136.255 45.465 136.895 ;
        RECT 45.635 136.085 45.905 136.895 ;
        RECT 46.085 136.855 46.835 137.375 ;
        RECT 47.005 137.025 47.755 137.545 ;
        RECT 47.930 136.975 48.280 137.625 ;
        RECT 46.085 136.085 47.755 136.855 ;
        RECT 48.450 136.805 48.680 137.795 ;
        RECT 48.015 136.635 48.680 136.805 ;
        RECT 48.015 136.345 48.185 136.635 ;
        RECT 48.355 136.085 48.685 136.465 ;
        RECT 48.855 136.345 49.040 138.465 ;
        RECT 49.280 138.175 49.545 138.635 ;
        RECT 49.715 138.040 49.965 138.465 ;
        RECT 50.175 138.190 51.280 138.360 ;
        RECT 49.660 137.910 49.965 138.040 ;
        RECT 49.210 136.715 49.490 137.665 ;
        RECT 49.660 136.805 49.830 137.910 ;
        RECT 50.000 137.125 50.240 137.720 ;
        RECT 50.410 137.655 50.940 138.020 ;
        RECT 50.410 136.955 50.580 137.655 ;
        RECT 51.110 137.575 51.280 138.190 ;
        RECT 51.450 137.835 51.620 138.635 ;
        RECT 51.790 138.135 52.040 138.465 ;
        RECT 52.265 138.165 53.150 138.335 ;
        RECT 51.110 137.485 51.620 137.575 ;
        RECT 49.660 136.675 49.885 136.805 ;
        RECT 50.055 136.735 50.580 136.955 ;
        RECT 50.750 137.315 51.620 137.485 ;
        RECT 49.295 136.085 49.545 136.545 ;
        RECT 49.715 136.535 49.885 136.675 ;
        RECT 50.750 136.535 50.920 137.315 ;
        RECT 51.450 137.245 51.620 137.315 ;
        RECT 51.130 137.065 51.330 137.095 ;
        RECT 51.790 137.065 51.960 138.135 ;
        RECT 52.130 137.245 52.320 137.965 ;
        RECT 51.130 136.765 51.960 137.065 ;
        RECT 52.490 137.035 52.810 137.995 ;
        RECT 49.715 136.365 50.050 136.535 ;
        RECT 50.245 136.365 50.920 136.535 ;
        RECT 51.240 136.085 51.610 136.585 ;
        RECT 51.790 136.535 51.960 136.765 ;
        RECT 52.345 136.705 52.810 137.035 ;
        RECT 52.980 137.325 53.150 138.165 ;
        RECT 53.330 138.135 53.645 138.635 ;
        RECT 53.875 137.905 54.215 138.465 ;
        RECT 53.320 137.530 54.215 137.905 ;
        RECT 54.385 137.625 54.555 138.635 ;
        RECT 54.025 137.325 54.215 137.530 ;
        RECT 54.725 137.575 55.055 138.420 ;
        RECT 54.725 137.495 55.115 137.575 ;
        RECT 54.900 137.445 55.115 137.495 ;
        RECT 55.750 137.485 56.010 138.635 ;
        RECT 56.185 137.560 56.440 138.465 ;
        RECT 56.610 137.875 56.940 138.635 ;
        RECT 57.155 137.705 57.325 138.465 ;
        RECT 52.980 136.995 53.855 137.325 ;
        RECT 54.025 136.995 54.775 137.325 ;
        RECT 52.980 136.535 53.150 136.995 ;
        RECT 54.025 136.825 54.225 136.995 ;
        RECT 54.945 136.865 55.115 137.445 ;
        RECT 54.890 136.825 55.115 136.865 ;
        RECT 51.790 136.365 52.195 136.535 ;
        RECT 52.365 136.365 53.150 136.535 ;
        RECT 53.425 136.085 53.635 136.615 ;
        RECT 53.895 136.300 54.225 136.825 ;
        RECT 54.735 136.740 55.115 136.825 ;
        RECT 54.395 136.085 54.565 136.695 ;
        RECT 54.735 136.305 55.065 136.740 ;
        RECT 55.750 136.085 56.010 136.925 ;
        RECT 56.185 136.830 56.355 137.560 ;
        RECT 56.610 137.535 57.325 137.705 ;
        RECT 57.585 137.875 58.100 138.285 ;
        RECT 58.335 137.875 58.505 138.635 ;
        RECT 58.675 138.295 60.705 138.465 ;
        RECT 56.610 137.325 56.780 137.535 ;
        RECT 56.525 136.995 56.780 137.325 ;
        RECT 56.185 136.255 56.440 136.830 ;
        RECT 56.610 136.805 56.780 136.995 ;
        RECT 57.060 136.985 57.415 137.355 ;
        RECT 57.585 137.065 57.925 137.875 ;
        RECT 58.675 137.630 58.845 138.295 ;
        RECT 59.240 137.955 60.365 138.125 ;
        RECT 58.095 137.440 58.845 137.630 ;
        RECT 59.015 137.615 60.025 137.785 ;
        RECT 57.585 136.895 58.815 137.065 ;
        RECT 56.610 136.635 57.325 136.805 ;
        RECT 56.610 136.085 56.940 136.465 ;
        RECT 57.155 136.255 57.325 136.635 ;
        RECT 57.860 136.290 58.105 136.895 ;
        RECT 58.325 136.085 58.835 136.620 ;
        RECT 59.015 136.255 59.205 137.615 ;
        RECT 59.375 136.595 59.650 137.415 ;
        RECT 59.855 136.815 60.025 137.615 ;
        RECT 60.195 136.825 60.365 137.955 ;
        RECT 60.535 137.325 60.705 138.295 ;
        RECT 60.875 137.495 61.045 138.635 ;
        RECT 61.215 137.495 61.550 138.465 ;
        RECT 60.535 136.995 60.730 137.325 ;
        RECT 60.955 136.995 61.210 137.325 ;
        RECT 60.955 136.825 61.125 136.995 ;
        RECT 61.380 136.825 61.550 137.495 ;
        RECT 60.195 136.655 61.125 136.825 ;
        RECT 60.195 136.620 60.370 136.655 ;
        RECT 59.375 136.425 59.655 136.595 ;
        RECT 59.375 136.255 59.650 136.425 ;
        RECT 59.840 136.255 60.370 136.620 ;
        RECT 60.795 136.085 61.125 136.485 ;
        RECT 61.295 136.255 61.550 136.825 ;
        RECT 61.730 137.495 62.065 138.465 ;
        RECT 62.235 137.495 62.405 138.635 ;
        RECT 62.575 138.295 64.605 138.465 ;
        RECT 61.730 136.825 61.900 137.495 ;
        RECT 62.575 137.325 62.745 138.295 ;
        RECT 62.070 136.995 62.325 137.325 ;
        RECT 62.550 136.995 62.745 137.325 ;
        RECT 62.915 137.955 64.040 138.125 ;
        RECT 62.155 136.825 62.325 136.995 ;
        RECT 62.915 136.825 63.085 137.955 ;
        RECT 61.730 136.255 61.985 136.825 ;
        RECT 62.155 136.655 63.085 136.825 ;
        RECT 63.255 137.615 64.265 137.785 ;
        RECT 63.255 136.815 63.425 137.615 ;
        RECT 63.630 136.935 63.905 137.415 ;
        RECT 63.625 136.765 63.905 136.935 ;
        RECT 62.910 136.620 63.085 136.655 ;
        RECT 62.155 136.085 62.485 136.485 ;
        RECT 62.910 136.255 63.440 136.620 ;
        RECT 63.630 136.255 63.905 136.765 ;
        RECT 64.075 136.255 64.265 137.615 ;
        RECT 64.435 137.630 64.605 138.295 ;
        RECT 64.775 137.875 64.945 138.635 ;
        RECT 65.180 137.875 65.695 138.285 ;
        RECT 64.435 137.440 65.185 137.630 ;
        RECT 65.355 137.065 65.695 137.875 ;
        RECT 64.465 136.895 65.695 137.065 ;
        RECT 65.870 137.495 66.205 138.465 ;
        RECT 66.375 137.495 66.545 138.635 ;
        RECT 66.715 138.295 68.745 138.465 ;
        RECT 64.445 136.085 64.955 136.620 ;
        RECT 65.175 136.290 65.420 136.895 ;
        RECT 65.870 136.825 66.040 137.495 ;
        RECT 66.715 137.325 66.885 138.295 ;
        RECT 66.210 136.995 66.465 137.325 ;
        RECT 66.690 136.995 66.885 137.325 ;
        RECT 67.055 137.955 68.180 138.125 ;
        RECT 66.295 136.825 66.465 136.995 ;
        RECT 67.055 136.825 67.225 137.955 ;
        RECT 65.870 136.255 66.125 136.825 ;
        RECT 66.295 136.655 67.225 136.825 ;
        RECT 67.395 137.615 68.405 137.785 ;
        RECT 67.395 136.815 67.565 137.615 ;
        RECT 67.770 137.275 68.045 137.415 ;
        RECT 67.765 137.105 68.045 137.275 ;
        RECT 67.050 136.620 67.225 136.655 ;
        RECT 66.295 136.085 66.625 136.485 ;
        RECT 67.050 136.255 67.580 136.620 ;
        RECT 67.770 136.255 68.045 137.105 ;
        RECT 68.215 136.255 68.405 137.615 ;
        RECT 68.575 137.630 68.745 138.295 ;
        RECT 68.915 137.875 69.085 138.635 ;
        RECT 69.320 137.875 69.835 138.285 ;
        RECT 68.575 137.440 69.325 137.630 ;
        RECT 69.495 137.065 69.835 137.875 ;
        RECT 70.005 137.470 70.295 138.635 ;
        RECT 70.555 137.965 70.725 138.465 ;
        RECT 70.895 138.135 71.225 138.635 ;
        RECT 70.555 137.795 71.220 137.965 ;
        RECT 68.605 136.895 69.835 137.065 ;
        RECT 70.470 136.975 70.820 137.625 ;
        RECT 68.585 136.085 69.095 136.620 ;
        RECT 69.315 136.290 69.560 136.895 ;
        RECT 70.005 136.085 70.295 136.810 ;
        RECT 70.990 136.805 71.220 137.795 ;
        RECT 70.555 136.635 71.220 136.805 ;
        RECT 70.555 136.345 70.725 136.635 ;
        RECT 70.895 136.085 71.225 136.465 ;
        RECT 71.395 136.345 71.580 138.465 ;
        RECT 71.820 138.175 72.085 138.635 ;
        RECT 72.255 138.040 72.505 138.465 ;
        RECT 72.715 138.190 73.820 138.360 ;
        RECT 72.200 137.910 72.505 138.040 ;
        RECT 71.750 136.715 72.030 137.665 ;
        RECT 72.200 136.805 72.370 137.910 ;
        RECT 72.540 137.125 72.780 137.720 ;
        RECT 72.950 137.655 73.480 138.020 ;
        RECT 72.950 136.955 73.120 137.655 ;
        RECT 73.650 137.575 73.820 138.190 ;
        RECT 73.990 137.835 74.160 138.635 ;
        RECT 74.330 138.135 74.580 138.465 ;
        RECT 74.805 138.165 75.690 138.335 ;
        RECT 73.650 137.485 74.160 137.575 ;
        RECT 72.200 136.675 72.425 136.805 ;
        RECT 72.595 136.735 73.120 136.955 ;
        RECT 73.290 137.315 74.160 137.485 ;
        RECT 71.835 136.085 72.085 136.545 ;
        RECT 72.255 136.535 72.425 136.675 ;
        RECT 73.290 136.535 73.460 137.315 ;
        RECT 73.990 137.245 74.160 137.315 ;
        RECT 73.670 137.065 73.870 137.095 ;
        RECT 74.330 137.065 74.500 138.135 ;
        RECT 74.670 137.245 74.860 137.965 ;
        RECT 73.670 136.765 74.500 137.065 ;
        RECT 75.030 137.035 75.350 137.995 ;
        RECT 72.255 136.365 72.590 136.535 ;
        RECT 72.785 136.365 73.460 136.535 ;
        RECT 73.780 136.085 74.150 136.585 ;
        RECT 74.330 136.535 74.500 136.765 ;
        RECT 74.885 136.705 75.350 137.035 ;
        RECT 75.520 137.325 75.690 138.165 ;
        RECT 75.870 138.135 76.185 138.635 ;
        RECT 76.415 137.905 76.755 138.465 ;
        RECT 75.860 137.530 76.755 137.905 ;
        RECT 76.925 137.625 77.095 138.635 ;
        RECT 76.565 137.325 76.755 137.530 ;
        RECT 77.265 137.575 77.595 138.420 ;
        RECT 77.265 137.495 77.655 137.575 ;
        RECT 77.440 137.445 77.655 137.495 ;
        RECT 75.520 136.995 76.395 137.325 ;
        RECT 76.565 136.995 77.315 137.325 ;
        RECT 75.520 136.535 75.690 136.995 ;
        RECT 76.565 136.825 76.765 136.995 ;
        RECT 77.485 136.865 77.655 137.445 ;
        RECT 77.430 136.825 77.655 136.865 ;
        RECT 74.330 136.365 74.735 136.535 ;
        RECT 74.905 136.365 75.690 136.535 ;
        RECT 75.965 136.085 76.175 136.615 ;
        RECT 76.435 136.300 76.765 136.825 ;
        RECT 77.275 136.740 77.655 136.825 ;
        RECT 77.825 137.495 78.165 138.465 ;
        RECT 78.335 137.495 78.505 138.635 ;
        RECT 78.775 137.835 79.025 138.635 ;
        RECT 79.670 137.665 80.000 138.465 ;
        RECT 80.300 137.835 80.630 138.635 ;
        RECT 80.800 137.665 81.130 138.465 ;
        RECT 78.695 137.495 81.130 137.665 ;
        RECT 81.965 137.545 83.175 138.635 ;
        RECT 77.825 136.885 78.000 137.495 ;
        RECT 78.695 137.245 78.865 137.495 ;
        RECT 78.170 137.075 78.865 137.245 ;
        RECT 79.040 137.075 79.460 137.275 ;
        RECT 79.630 137.075 79.960 137.275 ;
        RECT 80.130 137.075 80.460 137.275 ;
        RECT 76.935 136.085 77.105 136.695 ;
        RECT 77.275 136.305 77.605 136.740 ;
        RECT 77.825 136.255 78.165 136.885 ;
        RECT 78.335 136.085 78.585 136.885 ;
        RECT 78.775 136.735 80.000 136.905 ;
        RECT 78.775 136.255 79.105 136.735 ;
        RECT 79.275 136.085 79.500 136.545 ;
        RECT 79.670 136.255 80.000 136.735 ;
        RECT 80.630 136.865 80.800 137.495 ;
        RECT 80.985 137.075 81.335 137.325 ;
        RECT 81.965 137.005 82.485 137.545 ;
        RECT 80.630 136.255 81.130 136.865 ;
        RECT 82.655 136.835 83.175 137.375 ;
        RECT 81.965 136.085 83.175 136.835 ;
        RECT 5.520 135.915 83.260 136.085 ;
        RECT 5.605 135.165 6.815 135.915 ;
        RECT 5.605 134.625 6.125 135.165 ;
        RECT 7.455 135.105 7.725 135.915 ;
        RECT 7.895 135.105 8.225 135.745 ;
        RECT 8.395 135.105 8.635 135.915 ;
        RECT 8.910 135.345 9.085 135.745 ;
        RECT 9.255 135.535 9.585 135.915 ;
        RECT 9.830 135.415 10.060 135.745 ;
        RECT 8.910 135.175 9.540 135.345 ;
        RECT 6.295 134.455 6.815 134.995 ;
        RECT 7.445 134.675 7.795 134.925 ;
        RECT 7.965 134.505 8.135 135.105 ;
        RECT 9.370 135.005 9.540 135.175 ;
        RECT 8.305 134.675 8.655 134.925 ;
        RECT 5.605 133.365 6.815 134.455 ;
        RECT 7.455 133.365 7.785 134.505 ;
        RECT 7.965 134.335 8.645 134.505 ;
        RECT 8.315 133.550 8.645 134.335 ;
        RECT 8.825 134.325 9.190 135.005 ;
        RECT 9.370 134.675 9.720 135.005 ;
        RECT 9.370 134.155 9.540 134.675 ;
        RECT 8.910 133.985 9.540 134.155 ;
        RECT 9.890 134.125 10.060 135.415 ;
        RECT 10.260 134.305 10.540 135.580 ;
        RECT 10.765 135.575 11.035 135.580 ;
        RECT 10.725 135.405 11.035 135.575 ;
        RECT 11.495 135.535 11.825 135.915 ;
        RECT 11.995 135.660 12.330 135.705 ;
        RECT 10.765 134.305 11.035 135.405 ;
        RECT 11.225 134.305 11.565 135.335 ;
        RECT 11.995 135.195 12.335 135.660 ;
        RECT 11.735 134.675 11.995 135.005 ;
        RECT 11.735 134.125 11.905 134.675 ;
        RECT 12.165 134.505 12.335 135.195 ;
        RECT 12.590 135.345 12.765 135.745 ;
        RECT 12.935 135.535 13.265 135.915 ;
        RECT 13.510 135.415 13.740 135.745 ;
        RECT 12.590 135.175 13.220 135.345 ;
        RECT 13.050 135.005 13.220 135.175 ;
        RECT 8.910 133.535 9.085 133.985 ;
        RECT 9.890 133.955 11.905 134.125 ;
        RECT 9.255 133.365 9.585 133.805 ;
        RECT 9.890 133.535 10.060 133.955 ;
        RECT 10.295 133.365 10.965 133.775 ;
        RECT 11.180 133.535 11.350 133.955 ;
        RECT 11.550 133.365 11.880 133.775 ;
        RECT 12.075 133.535 12.335 134.505 ;
        RECT 12.505 134.325 12.870 135.005 ;
        RECT 13.050 134.675 13.400 135.005 ;
        RECT 13.050 134.155 13.220 134.675 ;
        RECT 12.590 133.985 13.220 134.155 ;
        RECT 13.570 134.125 13.740 135.415 ;
        RECT 13.940 134.305 14.220 135.580 ;
        RECT 14.445 135.575 14.715 135.580 ;
        RECT 14.405 135.405 14.715 135.575 ;
        RECT 15.175 135.535 15.505 135.915 ;
        RECT 15.675 135.660 16.010 135.705 ;
        RECT 14.445 134.305 14.715 135.405 ;
        RECT 14.905 134.305 15.245 135.335 ;
        RECT 15.675 135.195 16.015 135.660 ;
        RECT 16.275 135.365 16.445 135.655 ;
        RECT 16.615 135.535 16.945 135.915 ;
        RECT 16.275 135.195 16.940 135.365 ;
        RECT 15.415 134.675 15.675 135.005 ;
        RECT 15.415 134.125 15.585 134.675 ;
        RECT 15.845 134.505 16.015 135.195 ;
        RECT 12.590 133.535 12.765 133.985 ;
        RECT 13.570 133.955 15.585 134.125 ;
        RECT 12.935 133.365 13.265 133.805 ;
        RECT 13.570 133.535 13.740 133.955 ;
        RECT 13.975 133.365 14.645 133.775 ;
        RECT 14.860 133.535 15.030 133.955 ;
        RECT 15.230 133.365 15.560 133.775 ;
        RECT 15.755 133.535 16.015 134.505 ;
        RECT 16.190 134.375 16.540 135.025 ;
        RECT 16.710 134.205 16.940 135.195 ;
        RECT 16.275 134.035 16.940 134.205 ;
        RECT 16.275 133.535 16.445 134.035 ;
        RECT 16.615 133.365 16.945 133.865 ;
        RECT 17.115 133.535 17.300 135.655 ;
        RECT 17.555 135.455 17.805 135.915 ;
        RECT 17.975 135.465 18.310 135.635 ;
        RECT 18.505 135.465 19.180 135.635 ;
        RECT 17.975 135.325 18.145 135.465 ;
        RECT 17.470 134.335 17.750 135.285 ;
        RECT 17.920 135.195 18.145 135.325 ;
        RECT 17.920 134.090 18.090 135.195 ;
        RECT 18.315 135.045 18.840 135.265 ;
        RECT 18.260 134.280 18.500 134.875 ;
        RECT 18.670 134.345 18.840 135.045 ;
        RECT 19.010 134.685 19.180 135.465 ;
        RECT 19.500 135.415 19.870 135.915 ;
        RECT 20.050 135.465 20.455 135.635 ;
        RECT 20.625 135.465 21.410 135.635 ;
        RECT 20.050 135.235 20.220 135.465 ;
        RECT 19.390 134.935 20.220 135.235 ;
        RECT 20.605 134.965 21.070 135.295 ;
        RECT 19.390 134.905 19.590 134.935 ;
        RECT 19.710 134.685 19.880 134.755 ;
        RECT 19.010 134.515 19.880 134.685 ;
        RECT 19.370 134.425 19.880 134.515 ;
        RECT 17.920 133.960 18.225 134.090 ;
        RECT 18.670 133.980 19.200 134.345 ;
        RECT 17.540 133.365 17.805 133.825 ;
        RECT 17.975 133.535 18.225 133.960 ;
        RECT 19.370 133.810 19.540 134.425 ;
        RECT 18.435 133.640 19.540 133.810 ;
        RECT 19.710 133.365 19.880 134.165 ;
        RECT 20.050 133.865 20.220 134.935 ;
        RECT 20.390 134.035 20.580 134.755 ;
        RECT 20.750 134.005 21.070 134.965 ;
        RECT 21.240 135.005 21.410 135.465 ;
        RECT 21.685 135.385 21.895 135.915 ;
        RECT 22.155 135.175 22.485 135.700 ;
        RECT 22.655 135.305 22.825 135.915 ;
        RECT 22.995 135.260 23.325 135.695 ;
        RECT 23.635 135.365 23.805 135.655 ;
        RECT 23.975 135.535 24.305 135.915 ;
        RECT 22.995 135.175 23.375 135.260 ;
        RECT 23.635 135.195 24.300 135.365 ;
        RECT 22.285 135.005 22.485 135.175 ;
        RECT 23.150 135.135 23.375 135.175 ;
        RECT 21.240 134.675 22.115 135.005 ;
        RECT 22.285 134.675 23.035 135.005 ;
        RECT 20.050 133.535 20.300 133.865 ;
        RECT 21.240 133.835 21.410 134.675 ;
        RECT 22.285 134.470 22.475 134.675 ;
        RECT 23.205 134.555 23.375 135.135 ;
        RECT 23.160 134.505 23.375 134.555 ;
        RECT 21.580 134.095 22.475 134.470 ;
        RECT 22.985 134.425 23.375 134.505 ;
        RECT 20.525 133.665 21.410 133.835 ;
        RECT 21.590 133.365 21.905 133.865 ;
        RECT 22.135 133.535 22.475 134.095 ;
        RECT 22.645 133.365 22.815 134.375 ;
        RECT 22.985 133.580 23.315 134.425 ;
        RECT 23.550 134.375 23.900 135.025 ;
        RECT 24.070 134.205 24.300 135.195 ;
        RECT 23.635 134.035 24.300 134.205 ;
        RECT 23.635 133.535 23.805 134.035 ;
        RECT 23.975 133.365 24.305 133.865 ;
        RECT 24.475 133.535 24.660 135.655 ;
        RECT 24.915 135.455 25.165 135.915 ;
        RECT 25.335 135.465 25.670 135.635 ;
        RECT 25.865 135.465 26.540 135.635 ;
        RECT 25.335 135.325 25.505 135.465 ;
        RECT 24.830 134.335 25.110 135.285 ;
        RECT 25.280 135.195 25.505 135.325 ;
        RECT 25.280 134.090 25.450 135.195 ;
        RECT 25.675 135.045 26.200 135.265 ;
        RECT 25.620 134.280 25.860 134.875 ;
        RECT 26.030 134.345 26.200 135.045 ;
        RECT 26.370 134.685 26.540 135.465 ;
        RECT 26.860 135.415 27.230 135.915 ;
        RECT 27.410 135.465 27.815 135.635 ;
        RECT 27.985 135.465 28.770 135.635 ;
        RECT 27.410 135.235 27.580 135.465 ;
        RECT 26.750 134.935 27.580 135.235 ;
        RECT 27.965 134.965 28.430 135.295 ;
        RECT 26.750 134.905 26.950 134.935 ;
        RECT 27.070 134.685 27.240 134.755 ;
        RECT 26.370 134.515 27.240 134.685 ;
        RECT 26.730 134.425 27.240 134.515 ;
        RECT 25.280 133.960 25.585 134.090 ;
        RECT 26.030 133.980 26.560 134.345 ;
        RECT 24.900 133.365 25.165 133.825 ;
        RECT 25.335 133.535 25.585 133.960 ;
        RECT 26.730 133.810 26.900 134.425 ;
        RECT 25.795 133.640 26.900 133.810 ;
        RECT 27.070 133.365 27.240 134.165 ;
        RECT 27.410 133.865 27.580 134.935 ;
        RECT 27.750 134.035 27.940 134.755 ;
        RECT 28.110 134.005 28.430 134.965 ;
        RECT 28.600 135.005 28.770 135.465 ;
        RECT 29.045 135.385 29.255 135.915 ;
        RECT 29.515 135.175 29.845 135.700 ;
        RECT 30.015 135.305 30.185 135.915 ;
        RECT 30.355 135.260 30.685 135.695 ;
        RECT 30.855 135.400 31.025 135.915 ;
        RECT 30.355 135.175 30.735 135.260 ;
        RECT 31.365 135.190 31.655 135.915 ;
        RECT 31.915 135.365 32.085 135.655 ;
        RECT 32.255 135.535 32.585 135.915 ;
        RECT 31.915 135.195 32.580 135.365 ;
        RECT 29.645 135.005 29.845 135.175 ;
        RECT 30.510 135.135 30.735 135.175 ;
        RECT 28.600 134.675 29.475 135.005 ;
        RECT 29.645 134.675 30.395 135.005 ;
        RECT 27.410 133.535 27.660 133.865 ;
        RECT 28.600 133.835 28.770 134.675 ;
        RECT 29.645 134.470 29.835 134.675 ;
        RECT 30.565 134.555 30.735 135.135 ;
        RECT 30.520 134.505 30.735 134.555 ;
        RECT 28.940 134.095 29.835 134.470 ;
        RECT 30.345 134.425 30.735 134.505 ;
        RECT 27.885 133.665 28.770 133.835 ;
        RECT 28.950 133.365 29.265 133.865 ;
        RECT 29.495 133.535 29.835 134.095 ;
        RECT 30.005 133.365 30.175 134.375 ;
        RECT 30.345 133.580 30.675 134.425 ;
        RECT 30.845 133.365 31.015 134.280 ;
        RECT 31.365 133.365 31.655 134.530 ;
        RECT 31.830 134.375 32.180 135.025 ;
        RECT 32.350 134.205 32.580 135.195 ;
        RECT 31.915 134.035 32.580 134.205 ;
        RECT 31.915 133.535 32.085 134.035 ;
        RECT 32.255 133.365 32.585 133.865 ;
        RECT 32.755 133.535 32.940 135.655 ;
        RECT 33.195 135.455 33.445 135.915 ;
        RECT 33.615 135.465 33.950 135.635 ;
        RECT 34.145 135.465 34.820 135.635 ;
        RECT 33.615 135.325 33.785 135.465 ;
        RECT 33.110 134.335 33.390 135.285 ;
        RECT 33.560 135.195 33.785 135.325 ;
        RECT 33.560 134.090 33.730 135.195 ;
        RECT 33.955 135.045 34.480 135.265 ;
        RECT 33.900 134.280 34.140 134.875 ;
        RECT 34.310 134.345 34.480 135.045 ;
        RECT 34.650 134.685 34.820 135.465 ;
        RECT 35.140 135.415 35.510 135.915 ;
        RECT 35.690 135.465 36.095 135.635 ;
        RECT 36.265 135.465 37.050 135.635 ;
        RECT 35.690 135.235 35.860 135.465 ;
        RECT 35.030 134.935 35.860 135.235 ;
        RECT 36.245 134.965 36.710 135.295 ;
        RECT 35.030 134.905 35.230 134.935 ;
        RECT 35.350 134.685 35.520 134.755 ;
        RECT 34.650 134.515 35.520 134.685 ;
        RECT 35.010 134.425 35.520 134.515 ;
        RECT 33.560 133.960 33.865 134.090 ;
        RECT 34.310 133.980 34.840 134.345 ;
        RECT 33.180 133.365 33.445 133.825 ;
        RECT 33.615 133.535 33.865 133.960 ;
        RECT 35.010 133.810 35.180 134.425 ;
        RECT 34.075 133.640 35.180 133.810 ;
        RECT 35.350 133.365 35.520 134.165 ;
        RECT 35.690 133.865 35.860 134.935 ;
        RECT 36.030 134.035 36.220 134.755 ;
        RECT 36.390 134.005 36.710 134.965 ;
        RECT 36.880 135.005 37.050 135.465 ;
        RECT 37.325 135.385 37.535 135.915 ;
        RECT 37.795 135.175 38.125 135.700 ;
        RECT 38.295 135.305 38.465 135.915 ;
        RECT 38.635 135.260 38.965 135.695 ;
        RECT 40.195 135.365 40.365 135.655 ;
        RECT 40.535 135.535 40.865 135.915 ;
        RECT 38.635 135.175 39.015 135.260 ;
        RECT 40.195 135.195 40.860 135.365 ;
        RECT 37.925 135.005 38.125 135.175 ;
        RECT 38.790 135.135 39.015 135.175 ;
        RECT 36.880 134.675 37.755 135.005 ;
        RECT 37.925 134.675 38.675 135.005 ;
        RECT 35.690 133.535 35.940 133.865 ;
        RECT 36.880 133.835 37.050 134.675 ;
        RECT 37.925 134.470 38.115 134.675 ;
        RECT 38.845 134.555 39.015 135.135 ;
        RECT 38.800 134.505 39.015 134.555 ;
        RECT 37.220 134.095 38.115 134.470 ;
        RECT 38.625 134.425 39.015 134.505 ;
        RECT 36.165 133.665 37.050 133.835 ;
        RECT 37.230 133.365 37.545 133.865 ;
        RECT 37.775 133.535 38.115 134.095 ;
        RECT 38.285 133.365 38.455 134.375 ;
        RECT 38.625 133.580 38.955 134.425 ;
        RECT 40.110 134.375 40.460 135.025 ;
        RECT 40.630 134.205 40.860 135.195 ;
        RECT 40.195 134.035 40.860 134.205 ;
        RECT 40.195 133.535 40.365 134.035 ;
        RECT 40.535 133.365 40.865 133.865 ;
        RECT 41.035 133.535 41.220 135.655 ;
        RECT 41.475 135.455 41.725 135.915 ;
        RECT 41.895 135.465 42.230 135.635 ;
        RECT 42.425 135.465 43.100 135.635 ;
        RECT 41.895 135.325 42.065 135.465 ;
        RECT 41.390 134.335 41.670 135.285 ;
        RECT 41.840 135.195 42.065 135.325 ;
        RECT 41.840 134.090 42.010 135.195 ;
        RECT 42.235 135.045 42.760 135.265 ;
        RECT 42.180 134.280 42.420 134.875 ;
        RECT 42.590 134.345 42.760 135.045 ;
        RECT 42.930 134.685 43.100 135.465 ;
        RECT 43.420 135.415 43.790 135.915 ;
        RECT 43.970 135.465 44.375 135.635 ;
        RECT 44.545 135.465 45.330 135.635 ;
        RECT 43.970 135.235 44.140 135.465 ;
        RECT 43.310 134.935 44.140 135.235 ;
        RECT 44.525 134.965 44.990 135.295 ;
        RECT 43.310 134.905 43.510 134.935 ;
        RECT 43.630 134.685 43.800 134.755 ;
        RECT 42.930 134.515 43.800 134.685 ;
        RECT 43.290 134.425 43.800 134.515 ;
        RECT 41.840 133.960 42.145 134.090 ;
        RECT 42.590 133.980 43.120 134.345 ;
        RECT 41.460 133.365 41.725 133.825 ;
        RECT 41.895 133.535 42.145 133.960 ;
        RECT 43.290 133.810 43.460 134.425 ;
        RECT 42.355 133.640 43.460 133.810 ;
        RECT 43.630 133.365 43.800 134.165 ;
        RECT 43.970 133.865 44.140 134.935 ;
        RECT 44.310 134.035 44.500 134.755 ;
        RECT 44.670 134.005 44.990 134.965 ;
        RECT 45.160 135.005 45.330 135.465 ;
        RECT 45.605 135.385 45.815 135.915 ;
        RECT 46.075 135.175 46.405 135.700 ;
        RECT 46.575 135.305 46.745 135.915 ;
        RECT 46.915 135.260 47.245 135.695 ;
        RECT 46.915 135.175 47.295 135.260 ;
        RECT 46.205 135.005 46.405 135.175 ;
        RECT 47.070 135.135 47.295 135.175 ;
        RECT 45.160 134.675 46.035 135.005 ;
        RECT 46.205 134.675 46.955 135.005 ;
        RECT 43.970 133.535 44.220 133.865 ;
        RECT 45.160 133.835 45.330 134.675 ;
        RECT 46.205 134.470 46.395 134.675 ;
        RECT 47.125 134.555 47.295 135.135 ;
        RECT 47.080 134.505 47.295 134.555 ;
        RECT 45.500 134.095 46.395 134.470 ;
        RECT 46.905 134.425 47.295 134.505 ;
        RECT 47.930 135.175 48.185 135.745 ;
        RECT 48.355 135.515 48.685 135.915 ;
        RECT 49.110 135.380 49.640 135.745 ;
        RECT 49.110 135.345 49.285 135.380 ;
        RECT 48.355 135.175 49.285 135.345 ;
        RECT 47.930 134.505 48.100 135.175 ;
        RECT 48.355 135.005 48.525 135.175 ;
        RECT 48.270 134.675 48.525 135.005 ;
        RECT 48.750 134.675 48.945 135.005 ;
        RECT 44.445 133.665 45.330 133.835 ;
        RECT 45.510 133.365 45.825 133.865 ;
        RECT 46.055 133.535 46.395 134.095 ;
        RECT 46.565 133.365 46.735 134.375 ;
        RECT 46.905 133.580 47.235 134.425 ;
        RECT 47.930 133.535 48.265 134.505 ;
        RECT 48.435 133.365 48.605 134.505 ;
        RECT 48.775 133.705 48.945 134.675 ;
        RECT 49.115 134.045 49.285 135.175 ;
        RECT 49.455 134.385 49.625 135.185 ;
        RECT 49.830 134.895 50.105 135.745 ;
        RECT 49.825 134.725 50.105 134.895 ;
        RECT 49.830 134.585 50.105 134.725 ;
        RECT 50.275 134.385 50.465 135.745 ;
        RECT 50.645 135.380 51.155 135.915 ;
        RECT 51.375 135.105 51.620 135.710 ;
        RECT 52.065 135.175 52.450 135.745 ;
        RECT 52.620 135.455 52.945 135.915 ;
        RECT 53.465 135.285 53.745 135.745 ;
        RECT 50.665 134.935 51.895 135.105 ;
        RECT 49.455 134.215 50.465 134.385 ;
        RECT 50.635 134.370 51.385 134.560 ;
        RECT 49.115 133.875 50.240 134.045 ;
        RECT 50.635 133.705 50.805 134.370 ;
        RECT 51.555 134.125 51.895 134.935 ;
        RECT 48.775 133.535 50.805 133.705 ;
        RECT 50.975 133.365 51.145 134.125 ;
        RECT 51.380 133.715 51.895 134.125 ;
        RECT 52.065 134.505 52.345 135.175 ;
        RECT 52.620 135.115 53.745 135.285 ;
        RECT 52.620 135.005 53.070 135.115 ;
        RECT 52.515 134.675 53.070 135.005 ;
        RECT 53.935 134.945 54.335 135.745 ;
        RECT 54.735 135.455 55.005 135.915 ;
        RECT 55.175 135.285 55.460 135.745 ;
        RECT 52.065 133.535 52.450 134.505 ;
        RECT 52.620 134.215 53.070 134.675 ;
        RECT 53.240 134.385 54.335 134.945 ;
        RECT 52.620 133.995 53.745 134.215 ;
        RECT 52.620 133.365 52.945 133.825 ;
        RECT 53.465 133.535 53.745 133.995 ;
        RECT 53.935 133.535 54.335 134.385 ;
        RECT 54.505 135.115 55.460 135.285 ;
        RECT 55.745 135.165 56.955 135.915 ;
        RECT 57.125 135.190 57.415 135.915 ;
        RECT 57.830 135.435 58.130 135.915 ;
        RECT 58.300 135.265 58.560 135.720 ;
        RECT 58.730 135.435 58.990 135.915 ;
        RECT 59.160 135.265 59.420 135.720 ;
        RECT 59.590 135.435 59.850 135.915 ;
        RECT 60.020 135.265 60.280 135.720 ;
        RECT 60.450 135.435 60.710 135.915 ;
        RECT 60.880 135.265 61.140 135.720 ;
        RECT 61.310 135.390 61.570 135.915 ;
        RECT 54.505 134.215 54.715 135.115 ;
        RECT 54.885 134.385 55.575 134.945 ;
        RECT 55.745 134.625 56.265 135.165 ;
        RECT 57.830 135.095 61.140 135.265 ;
        RECT 56.435 134.455 56.955 134.995 ;
        RECT 54.505 133.995 55.460 134.215 ;
        RECT 54.735 133.365 55.005 133.825 ;
        RECT 55.175 133.535 55.460 133.995 ;
        RECT 55.745 133.365 56.955 134.455 ;
        RECT 57.125 133.365 57.415 134.530 ;
        RECT 57.830 134.505 58.800 135.095 ;
        RECT 61.740 134.925 61.990 135.735 ;
        RECT 62.170 135.455 62.415 135.915 ;
        RECT 58.970 134.675 61.990 134.925 ;
        RECT 62.160 134.675 62.475 135.285 ;
        RECT 62.650 135.175 62.905 135.745 ;
        RECT 63.075 135.515 63.405 135.915 ;
        RECT 63.830 135.380 64.360 135.745 ;
        RECT 64.550 135.575 64.825 135.745 ;
        RECT 64.545 135.405 64.825 135.575 ;
        RECT 63.830 135.345 64.005 135.380 ;
        RECT 63.075 135.175 64.005 135.345 ;
        RECT 57.830 134.265 61.140 134.505 ;
        RECT 57.835 133.365 58.130 134.095 ;
        RECT 58.300 133.540 58.560 134.265 ;
        RECT 58.730 133.365 58.990 134.095 ;
        RECT 59.160 133.540 59.420 134.265 ;
        RECT 59.590 133.365 59.850 134.095 ;
        RECT 60.020 133.540 60.280 134.265 ;
        RECT 60.450 133.365 60.710 134.095 ;
        RECT 60.880 133.540 61.140 134.265 ;
        RECT 61.310 133.365 61.570 134.475 ;
        RECT 61.740 133.540 61.990 134.675 ;
        RECT 62.650 134.505 62.820 135.175 ;
        RECT 63.075 135.005 63.245 135.175 ;
        RECT 62.990 134.675 63.245 135.005 ;
        RECT 63.470 134.675 63.665 135.005 ;
        RECT 62.170 133.365 62.465 134.475 ;
        RECT 62.650 133.535 62.985 134.505 ;
        RECT 63.155 133.365 63.325 134.505 ;
        RECT 63.495 133.705 63.665 134.675 ;
        RECT 63.835 134.045 64.005 135.175 ;
        RECT 64.175 134.385 64.345 135.185 ;
        RECT 64.550 134.585 64.825 135.405 ;
        RECT 64.995 134.385 65.185 135.745 ;
        RECT 65.365 135.380 65.875 135.915 ;
        RECT 66.095 135.105 66.340 135.710 ;
        RECT 67.295 135.260 67.625 135.695 ;
        RECT 67.795 135.305 67.965 135.915 ;
        RECT 67.245 135.175 67.625 135.260 ;
        RECT 68.135 135.175 68.465 135.700 ;
        RECT 68.725 135.385 68.935 135.915 ;
        RECT 69.210 135.465 69.995 135.635 ;
        RECT 70.165 135.465 70.570 135.635 ;
        RECT 67.245 135.135 67.470 135.175 ;
        RECT 65.385 134.935 66.615 135.105 ;
        RECT 64.175 134.215 65.185 134.385 ;
        RECT 65.355 134.370 66.105 134.560 ;
        RECT 63.835 133.875 64.960 134.045 ;
        RECT 65.355 133.705 65.525 134.370 ;
        RECT 66.275 134.125 66.615 134.935 ;
        RECT 67.245 134.555 67.415 135.135 ;
        RECT 68.135 135.005 68.335 135.175 ;
        RECT 69.210 135.005 69.380 135.465 ;
        RECT 67.585 134.675 68.335 135.005 ;
        RECT 68.505 134.675 69.380 135.005 ;
        RECT 67.245 134.505 67.460 134.555 ;
        RECT 67.245 134.425 67.635 134.505 ;
        RECT 63.495 133.535 65.525 133.705 ;
        RECT 65.695 133.365 65.865 134.125 ;
        RECT 66.100 133.715 66.615 134.125 ;
        RECT 67.305 133.580 67.635 134.425 ;
        RECT 68.145 134.470 68.335 134.675 ;
        RECT 67.805 133.365 67.975 134.375 ;
        RECT 68.145 134.095 69.040 134.470 ;
        RECT 68.145 133.535 68.485 134.095 ;
        RECT 68.715 133.365 69.030 133.865 ;
        RECT 69.210 133.835 69.380 134.675 ;
        RECT 69.550 134.965 70.015 135.295 ;
        RECT 70.400 135.235 70.570 135.465 ;
        RECT 70.750 135.415 71.120 135.915 ;
        RECT 71.440 135.465 72.115 135.635 ;
        RECT 72.310 135.465 72.645 135.635 ;
        RECT 69.550 134.005 69.870 134.965 ;
        RECT 70.400 134.935 71.230 135.235 ;
        RECT 70.040 134.035 70.230 134.755 ;
        RECT 70.400 133.865 70.570 134.935 ;
        RECT 71.030 134.905 71.230 134.935 ;
        RECT 70.740 134.685 70.910 134.755 ;
        RECT 71.440 134.685 71.610 135.465 ;
        RECT 72.475 135.325 72.645 135.465 ;
        RECT 72.815 135.455 73.065 135.915 ;
        RECT 70.740 134.515 71.610 134.685 ;
        RECT 71.780 135.045 72.305 135.265 ;
        RECT 72.475 135.195 72.700 135.325 ;
        RECT 70.740 134.425 71.250 134.515 ;
        RECT 69.210 133.665 70.095 133.835 ;
        RECT 70.320 133.535 70.570 133.865 ;
        RECT 70.740 133.365 70.910 134.165 ;
        RECT 71.080 133.810 71.250 134.425 ;
        RECT 71.780 134.345 71.950 135.045 ;
        RECT 71.420 133.980 71.950 134.345 ;
        RECT 72.120 134.280 72.360 134.875 ;
        RECT 72.530 134.090 72.700 135.195 ;
        RECT 72.870 134.335 73.150 135.285 ;
        RECT 72.395 133.960 72.700 134.090 ;
        RECT 71.080 133.640 72.185 133.810 ;
        RECT 72.395 133.535 72.645 133.960 ;
        RECT 72.815 133.365 73.080 133.825 ;
        RECT 73.320 133.535 73.505 135.655 ;
        RECT 73.675 135.535 74.005 135.915 ;
        RECT 74.175 135.365 74.345 135.655 ;
        RECT 73.680 135.195 74.345 135.365 ;
        RECT 74.695 135.365 74.865 135.655 ;
        RECT 75.035 135.535 75.365 135.915 ;
        RECT 74.695 135.195 75.360 135.365 ;
        RECT 73.680 134.205 73.910 135.195 ;
        RECT 74.080 134.375 74.430 135.025 ;
        RECT 74.610 134.375 74.960 135.025 ;
        RECT 75.130 134.205 75.360 135.195 ;
        RECT 73.680 134.035 74.345 134.205 ;
        RECT 73.675 133.365 74.005 133.865 ;
        RECT 74.175 133.535 74.345 134.035 ;
        RECT 74.695 134.035 75.360 134.205 ;
        RECT 74.695 133.535 74.865 134.035 ;
        RECT 75.035 133.365 75.365 133.865 ;
        RECT 75.535 133.535 75.720 135.655 ;
        RECT 75.975 135.455 76.225 135.915 ;
        RECT 76.395 135.465 76.730 135.635 ;
        RECT 76.925 135.465 77.600 135.635 ;
        RECT 76.395 135.325 76.565 135.465 ;
        RECT 75.890 134.335 76.170 135.285 ;
        RECT 76.340 135.195 76.565 135.325 ;
        RECT 76.340 134.090 76.510 135.195 ;
        RECT 76.735 135.045 77.260 135.265 ;
        RECT 76.680 134.280 76.920 134.875 ;
        RECT 77.090 134.345 77.260 135.045 ;
        RECT 77.430 134.685 77.600 135.465 ;
        RECT 77.920 135.415 78.290 135.915 ;
        RECT 78.470 135.465 78.875 135.635 ;
        RECT 79.045 135.465 79.830 135.635 ;
        RECT 78.470 135.235 78.640 135.465 ;
        RECT 77.810 134.935 78.640 135.235 ;
        RECT 79.025 134.965 79.490 135.295 ;
        RECT 77.810 134.905 78.010 134.935 ;
        RECT 78.130 134.685 78.300 134.755 ;
        RECT 77.430 134.515 78.300 134.685 ;
        RECT 77.790 134.425 78.300 134.515 ;
        RECT 76.340 133.960 76.645 134.090 ;
        RECT 77.090 133.980 77.620 134.345 ;
        RECT 75.960 133.365 76.225 133.825 ;
        RECT 76.395 133.535 76.645 133.960 ;
        RECT 77.790 133.810 77.960 134.425 ;
        RECT 76.855 133.640 77.960 133.810 ;
        RECT 78.130 133.365 78.300 134.165 ;
        RECT 78.470 133.865 78.640 134.935 ;
        RECT 78.810 134.035 79.000 134.755 ;
        RECT 79.170 134.005 79.490 134.965 ;
        RECT 79.660 135.005 79.830 135.465 ;
        RECT 80.105 135.385 80.315 135.915 ;
        RECT 80.575 135.175 80.905 135.700 ;
        RECT 81.075 135.305 81.245 135.915 ;
        RECT 81.415 135.260 81.745 135.695 ;
        RECT 81.415 135.175 81.795 135.260 ;
        RECT 80.705 135.005 80.905 135.175 ;
        RECT 81.570 135.135 81.795 135.175 ;
        RECT 81.965 135.165 83.175 135.915 ;
        RECT 79.660 134.675 80.535 135.005 ;
        RECT 80.705 134.675 81.455 135.005 ;
        RECT 78.470 133.535 78.720 133.865 ;
        RECT 79.660 133.835 79.830 134.675 ;
        RECT 80.705 134.470 80.895 134.675 ;
        RECT 81.625 134.555 81.795 135.135 ;
        RECT 81.580 134.505 81.795 134.555 ;
        RECT 80.000 134.095 80.895 134.470 ;
        RECT 81.405 134.425 81.795 134.505 ;
        RECT 81.965 134.455 82.485 134.995 ;
        RECT 82.655 134.625 83.175 135.165 ;
        RECT 78.945 133.665 79.830 133.835 ;
        RECT 80.010 133.365 80.325 133.865 ;
        RECT 80.555 133.535 80.895 134.095 ;
        RECT 81.065 133.365 81.235 134.375 ;
        RECT 81.405 133.580 81.735 134.425 ;
        RECT 81.965 133.365 83.175 134.455 ;
        RECT 5.520 133.195 83.260 133.365 ;
        RECT 5.605 132.105 6.815 133.195 ;
        RECT 6.985 132.105 9.575 133.195 ;
        RECT 5.605 131.395 6.125 131.935 ;
        RECT 6.295 131.565 6.815 132.105 ;
        RECT 6.985 131.415 8.195 131.935 ;
        RECT 8.365 131.585 9.575 132.105 ;
        RECT 9.745 132.095 10.065 133.025 ;
        RECT 10.245 132.515 10.645 133.025 ;
        RECT 10.815 132.685 10.985 133.195 ;
        RECT 11.155 132.515 11.485 133.025 ;
        RECT 10.245 132.345 11.485 132.515 ;
        RECT 11.655 132.345 11.825 133.195 ;
        RECT 12.415 132.345 12.795 133.025 ;
        RECT 9.745 131.925 10.375 132.095 ;
        RECT 5.605 130.645 6.815 131.395 ;
        RECT 6.985 130.645 9.575 131.415 ;
        RECT 9.745 130.645 10.035 131.480 ;
        RECT 10.205 131.045 10.375 131.925 ;
        RECT 11.150 132.005 12.455 132.175 ;
        RECT 10.545 131.385 10.775 131.885 ;
        RECT 11.150 131.805 11.320 132.005 ;
        RECT 10.945 131.635 11.320 131.805 ;
        RECT 11.490 131.635 12.040 131.835 ;
        RECT 12.210 131.555 12.455 132.005 ;
        RECT 12.625 131.385 12.795 132.345 ;
        RECT 10.545 131.215 12.795 131.385 ;
        RECT 12.965 132.055 13.225 133.025 ;
        RECT 13.420 132.785 13.750 133.195 ;
        RECT 13.950 132.605 14.120 133.025 ;
        RECT 14.335 132.785 15.005 133.195 ;
        RECT 15.240 132.605 15.410 133.025 ;
        RECT 15.715 132.755 16.045 133.195 ;
        RECT 13.395 132.435 15.410 132.605 ;
        RECT 16.215 132.575 16.390 133.025 ;
        RECT 12.965 131.365 13.135 132.055 ;
        RECT 13.395 131.885 13.565 132.435 ;
        RECT 13.305 131.555 13.565 131.885 ;
        RECT 10.205 130.875 11.160 131.045 ;
        RECT 11.575 130.645 11.905 131.035 ;
        RECT 12.075 130.895 12.245 131.215 ;
        RECT 12.415 130.645 12.745 131.035 ;
        RECT 12.965 130.900 13.305 131.365 ;
        RECT 13.735 131.225 14.075 132.255 ;
        RECT 14.265 131.155 14.535 132.255 ;
        RECT 12.970 130.855 13.305 130.900 ;
        RECT 13.475 130.645 13.805 131.025 ;
        RECT 14.265 130.985 14.575 131.155 ;
        RECT 14.265 130.980 14.535 130.985 ;
        RECT 14.760 130.980 15.040 132.255 ;
        RECT 15.240 131.145 15.410 132.435 ;
        RECT 15.760 132.405 16.390 132.575 ;
        RECT 16.655 132.585 16.985 133.015 ;
        RECT 17.165 132.755 17.360 133.195 ;
        RECT 17.530 132.585 17.860 133.015 ;
        RECT 16.655 132.415 17.860 132.585 ;
        RECT 15.760 131.885 15.930 132.405 ;
        RECT 15.580 131.555 15.930 131.885 ;
        RECT 16.110 131.555 16.475 132.235 ;
        RECT 16.655 132.085 17.550 132.415 ;
        RECT 18.030 132.245 18.305 133.015 ;
        RECT 17.720 132.055 18.305 132.245 ;
        RECT 16.660 131.555 16.955 131.885 ;
        RECT 17.135 131.555 17.550 131.885 ;
        RECT 15.760 131.385 15.930 131.555 ;
        RECT 15.760 131.215 16.390 131.385 ;
        RECT 15.240 130.815 15.470 131.145 ;
        RECT 15.715 130.645 16.045 131.025 ;
        RECT 16.215 130.815 16.390 131.215 ;
        RECT 16.655 130.645 16.955 131.375 ;
        RECT 17.135 130.935 17.365 131.555 ;
        RECT 17.720 131.385 17.895 132.055 ;
        RECT 18.485 132.030 18.775 133.195 ;
        RECT 19.950 132.575 20.125 133.025 ;
        RECT 20.295 132.755 20.625 133.195 ;
        RECT 20.930 132.605 21.100 133.025 ;
        RECT 21.335 132.785 22.005 133.195 ;
        RECT 22.220 132.605 22.390 133.025 ;
        RECT 22.590 132.785 22.920 133.195 ;
        RECT 19.950 132.405 20.580 132.575 ;
        RECT 17.565 131.205 17.895 131.385 ;
        RECT 18.065 131.235 18.305 131.885 ;
        RECT 19.865 131.555 20.230 132.235 ;
        RECT 20.410 131.885 20.580 132.405 ;
        RECT 20.930 132.435 22.945 132.605 ;
        RECT 20.410 131.555 20.760 131.885 ;
        RECT 20.410 131.385 20.580 131.555 ;
        RECT 17.565 130.825 17.790 131.205 ;
        RECT 17.960 130.645 18.290 131.035 ;
        RECT 18.485 130.645 18.775 131.370 ;
        RECT 19.950 131.215 20.580 131.385 ;
        RECT 19.950 130.815 20.125 131.215 ;
        RECT 20.930 131.145 21.100 132.435 ;
        RECT 20.295 130.645 20.625 131.025 ;
        RECT 20.870 130.815 21.100 131.145 ;
        RECT 21.300 130.980 21.580 132.255 ;
        RECT 21.805 131.495 22.075 132.255 ;
        RECT 21.765 131.325 22.075 131.495 ;
        RECT 21.805 130.980 22.075 131.325 ;
        RECT 22.265 131.225 22.605 132.255 ;
        RECT 22.775 131.885 22.945 132.435 ;
        RECT 23.115 132.055 23.375 133.025 ;
        RECT 23.630 132.575 23.805 133.025 ;
        RECT 23.975 132.755 24.305 133.195 ;
        RECT 24.610 132.605 24.780 133.025 ;
        RECT 25.015 132.785 25.685 133.195 ;
        RECT 25.900 132.605 26.070 133.025 ;
        RECT 26.270 132.785 26.600 133.195 ;
        RECT 23.630 132.405 24.260 132.575 ;
        RECT 22.775 131.555 23.035 131.885 ;
        RECT 23.205 131.365 23.375 132.055 ;
        RECT 23.545 131.555 23.910 132.235 ;
        RECT 24.090 131.885 24.260 132.405 ;
        RECT 24.610 132.435 26.625 132.605 ;
        RECT 24.090 131.555 24.440 131.885 ;
        RECT 24.090 131.385 24.260 131.555 ;
        RECT 22.535 130.645 22.865 131.025 ;
        RECT 23.035 130.900 23.375 131.365 ;
        RECT 23.630 131.215 24.260 131.385 ;
        RECT 23.035 130.855 23.370 130.900 ;
        RECT 23.630 130.815 23.805 131.215 ;
        RECT 24.610 131.145 24.780 132.435 ;
        RECT 23.975 130.645 24.305 131.025 ;
        RECT 24.550 130.815 24.780 131.145 ;
        RECT 24.980 130.980 25.260 132.255 ;
        RECT 25.485 132.175 25.755 132.255 ;
        RECT 25.445 132.005 25.755 132.175 ;
        RECT 25.485 130.980 25.755 132.005 ;
        RECT 25.945 131.225 26.285 132.255 ;
        RECT 26.455 131.885 26.625 132.435 ;
        RECT 26.795 132.055 27.055 133.025 ;
        RECT 27.235 132.585 27.565 133.015 ;
        RECT 27.745 132.755 27.940 133.195 ;
        RECT 28.110 132.585 28.440 133.015 ;
        RECT 27.235 132.415 28.440 132.585 ;
        RECT 27.235 132.085 28.130 132.415 ;
        RECT 28.610 132.245 28.885 133.015 ;
        RECT 26.455 131.555 26.715 131.885 ;
        RECT 26.885 131.365 27.055 132.055 ;
        RECT 28.300 132.055 28.885 132.245 ;
        RECT 29.075 132.245 29.350 133.015 ;
        RECT 29.520 132.585 29.850 133.015 ;
        RECT 30.020 132.755 30.215 133.195 ;
        RECT 30.395 132.585 30.725 133.015 ;
        RECT 29.520 132.415 30.725 132.585 ;
        RECT 29.075 132.055 29.660 132.245 ;
        RECT 29.830 132.085 30.725 132.415 ;
        RECT 31.365 132.055 31.645 133.195 ;
        RECT 27.240 131.555 27.535 131.885 ;
        RECT 27.715 131.555 28.130 131.885 ;
        RECT 26.215 130.645 26.545 131.025 ;
        RECT 26.715 130.900 27.055 131.365 ;
        RECT 26.715 130.855 27.050 130.900 ;
        RECT 27.235 130.645 27.535 131.375 ;
        RECT 27.715 130.935 27.945 131.555 ;
        RECT 28.300 131.385 28.475 132.055 ;
        RECT 28.145 131.205 28.475 131.385 ;
        RECT 28.645 131.235 28.885 131.885 ;
        RECT 29.075 131.235 29.315 131.885 ;
        RECT 29.485 131.385 29.660 132.055 ;
        RECT 31.815 132.045 32.145 133.025 ;
        RECT 32.315 132.055 32.575 133.195 ;
        RECT 32.835 132.525 33.005 133.025 ;
        RECT 33.175 132.695 33.505 133.195 ;
        RECT 32.835 132.355 33.500 132.525 ;
        RECT 29.830 131.555 30.245 131.885 ;
        RECT 30.425 131.555 30.720 131.885 ;
        RECT 31.375 131.615 31.710 131.885 ;
        RECT 29.485 131.205 29.815 131.385 ;
        RECT 28.145 130.825 28.370 131.205 ;
        RECT 28.540 130.645 28.870 131.035 ;
        RECT 29.090 130.645 29.420 131.035 ;
        RECT 29.590 130.825 29.815 131.205 ;
        RECT 30.015 130.935 30.245 131.555 ;
        RECT 31.880 131.445 32.050 132.045 ;
        RECT 32.220 131.635 32.555 131.885 ;
        RECT 32.750 131.535 33.100 132.185 ;
        RECT 30.425 130.645 30.725 131.375 ;
        RECT 31.365 130.645 31.675 131.445 ;
        RECT 31.880 130.815 32.575 131.445 ;
        RECT 33.270 131.365 33.500 132.355 ;
        RECT 32.835 131.195 33.500 131.365 ;
        RECT 32.835 130.905 33.005 131.195 ;
        RECT 33.175 130.645 33.505 131.025 ;
        RECT 33.675 130.905 33.860 133.025 ;
        RECT 34.100 132.735 34.365 133.195 ;
        RECT 34.535 132.600 34.785 133.025 ;
        RECT 34.995 132.750 36.100 132.920 ;
        RECT 34.480 132.470 34.785 132.600 ;
        RECT 34.030 131.275 34.310 132.225 ;
        RECT 34.480 131.365 34.650 132.470 ;
        RECT 34.820 131.685 35.060 132.280 ;
        RECT 35.230 132.215 35.760 132.580 ;
        RECT 35.230 131.515 35.400 132.215 ;
        RECT 35.930 132.135 36.100 132.750 ;
        RECT 36.270 132.395 36.440 133.195 ;
        RECT 36.610 132.695 36.860 133.025 ;
        RECT 37.085 132.725 37.970 132.895 ;
        RECT 35.930 132.045 36.440 132.135 ;
        RECT 34.480 131.235 34.705 131.365 ;
        RECT 34.875 131.295 35.400 131.515 ;
        RECT 35.570 131.875 36.440 132.045 ;
        RECT 34.115 130.645 34.365 131.105 ;
        RECT 34.535 131.095 34.705 131.235 ;
        RECT 35.570 131.095 35.740 131.875 ;
        RECT 36.270 131.805 36.440 131.875 ;
        RECT 35.950 131.625 36.150 131.655 ;
        RECT 36.610 131.625 36.780 132.695 ;
        RECT 36.950 131.805 37.140 132.525 ;
        RECT 35.950 131.325 36.780 131.625 ;
        RECT 37.310 131.595 37.630 132.555 ;
        RECT 34.535 130.925 34.870 131.095 ;
        RECT 35.065 130.925 35.740 131.095 ;
        RECT 36.060 130.645 36.430 131.145 ;
        RECT 36.610 131.095 36.780 131.325 ;
        RECT 37.165 131.265 37.630 131.595 ;
        RECT 37.800 131.885 37.970 132.725 ;
        RECT 38.150 132.695 38.465 133.195 ;
        RECT 38.695 132.465 39.035 133.025 ;
        RECT 38.140 132.090 39.035 132.465 ;
        RECT 39.205 132.185 39.375 133.195 ;
        RECT 38.845 131.885 39.035 132.090 ;
        RECT 39.545 132.135 39.875 132.980 ;
        RECT 39.545 132.055 39.935 132.135 ;
        RECT 39.720 132.005 39.935 132.055 ;
        RECT 37.800 131.555 38.675 131.885 ;
        RECT 38.845 131.555 39.595 131.885 ;
        RECT 37.800 131.095 37.970 131.555 ;
        RECT 38.845 131.385 39.045 131.555 ;
        RECT 39.765 131.425 39.935 132.005 ;
        RECT 39.710 131.385 39.935 131.425 ;
        RECT 36.610 130.925 37.015 131.095 ;
        RECT 37.185 130.925 37.970 131.095 ;
        RECT 38.245 130.645 38.455 131.175 ;
        RECT 38.715 130.860 39.045 131.385 ;
        RECT 39.555 131.300 39.935 131.385 ;
        RECT 40.110 132.055 40.445 133.025 ;
        RECT 40.615 132.055 40.785 133.195 ;
        RECT 40.955 132.855 42.985 133.025 ;
        RECT 40.110 131.385 40.280 132.055 ;
        RECT 40.955 131.885 41.125 132.855 ;
        RECT 40.450 131.555 40.705 131.885 ;
        RECT 40.930 131.555 41.125 131.885 ;
        RECT 41.295 132.515 42.420 132.685 ;
        RECT 40.535 131.385 40.705 131.555 ;
        RECT 41.295 131.385 41.465 132.515 ;
        RECT 39.215 130.645 39.385 131.255 ;
        RECT 39.555 130.865 39.885 131.300 ;
        RECT 40.110 130.815 40.365 131.385 ;
        RECT 40.535 131.215 41.465 131.385 ;
        RECT 41.635 132.175 42.645 132.345 ;
        RECT 41.635 131.375 41.805 132.175 ;
        RECT 42.010 131.495 42.285 131.975 ;
        RECT 42.005 131.325 42.285 131.495 ;
        RECT 41.290 131.180 41.465 131.215 ;
        RECT 40.535 130.645 40.865 131.045 ;
        RECT 41.290 130.815 41.820 131.180 ;
        RECT 42.010 130.815 42.285 131.325 ;
        RECT 42.455 130.815 42.645 132.175 ;
        RECT 42.815 132.190 42.985 132.855 ;
        RECT 43.155 132.435 43.325 133.195 ;
        RECT 43.560 132.435 44.075 132.845 ;
        RECT 42.815 132.000 43.565 132.190 ;
        RECT 43.735 131.625 44.075 132.435 ;
        RECT 44.245 132.030 44.535 133.195 ;
        RECT 44.795 132.525 44.965 133.025 ;
        RECT 45.135 132.695 45.465 133.195 ;
        RECT 44.795 132.355 45.460 132.525 ;
        RECT 42.845 131.455 44.075 131.625 ;
        RECT 44.710 131.535 45.060 132.185 ;
        RECT 42.825 130.645 43.335 131.180 ;
        RECT 43.555 130.850 43.800 131.455 ;
        RECT 44.245 130.645 44.535 131.370 ;
        RECT 45.230 131.365 45.460 132.355 ;
        RECT 44.795 131.195 45.460 131.365 ;
        RECT 44.795 130.905 44.965 131.195 ;
        RECT 45.135 130.645 45.465 131.025 ;
        RECT 45.635 130.905 45.820 133.025 ;
        RECT 46.060 132.735 46.325 133.195 ;
        RECT 46.495 132.600 46.745 133.025 ;
        RECT 46.955 132.750 48.060 132.920 ;
        RECT 46.440 132.470 46.745 132.600 ;
        RECT 45.990 131.275 46.270 132.225 ;
        RECT 46.440 131.365 46.610 132.470 ;
        RECT 46.780 131.685 47.020 132.280 ;
        RECT 47.190 132.215 47.720 132.580 ;
        RECT 47.190 131.515 47.360 132.215 ;
        RECT 47.890 132.135 48.060 132.750 ;
        RECT 48.230 132.395 48.400 133.195 ;
        RECT 48.570 132.695 48.820 133.025 ;
        RECT 49.045 132.725 49.930 132.895 ;
        RECT 47.890 132.045 48.400 132.135 ;
        RECT 46.440 131.235 46.665 131.365 ;
        RECT 46.835 131.295 47.360 131.515 ;
        RECT 47.530 131.875 48.400 132.045 ;
        RECT 46.075 130.645 46.325 131.105 ;
        RECT 46.495 131.095 46.665 131.235 ;
        RECT 47.530 131.095 47.700 131.875 ;
        RECT 48.230 131.805 48.400 131.875 ;
        RECT 47.910 131.625 48.110 131.655 ;
        RECT 48.570 131.625 48.740 132.695 ;
        RECT 48.910 131.805 49.100 132.525 ;
        RECT 47.910 131.325 48.740 131.625 ;
        RECT 49.270 131.595 49.590 132.555 ;
        RECT 46.495 130.925 46.830 131.095 ;
        RECT 47.025 130.925 47.700 131.095 ;
        RECT 48.020 130.645 48.390 131.145 ;
        RECT 48.570 131.095 48.740 131.325 ;
        RECT 49.125 131.265 49.590 131.595 ;
        RECT 49.760 131.885 49.930 132.725 ;
        RECT 50.110 132.695 50.425 133.195 ;
        RECT 50.655 132.465 50.995 133.025 ;
        RECT 50.100 132.090 50.995 132.465 ;
        RECT 51.165 132.185 51.335 133.195 ;
        RECT 50.805 131.885 50.995 132.090 ;
        RECT 51.505 132.135 51.835 132.980 ;
        RECT 52.155 132.525 52.325 133.025 ;
        RECT 52.495 132.695 52.825 133.195 ;
        RECT 52.155 132.355 52.820 132.525 ;
        RECT 51.505 132.055 51.895 132.135 ;
        RECT 51.680 132.005 51.895 132.055 ;
        RECT 49.760 131.555 50.635 131.885 ;
        RECT 50.805 131.555 51.555 131.885 ;
        RECT 49.760 131.095 49.930 131.555 ;
        RECT 50.805 131.385 51.005 131.555 ;
        RECT 51.725 131.425 51.895 132.005 ;
        RECT 52.070 131.535 52.420 132.185 ;
        RECT 51.670 131.385 51.895 131.425 ;
        RECT 48.570 130.925 48.975 131.095 ;
        RECT 49.145 130.925 49.930 131.095 ;
        RECT 50.205 130.645 50.415 131.175 ;
        RECT 50.675 130.860 51.005 131.385 ;
        RECT 51.515 131.300 51.895 131.385 ;
        RECT 52.590 131.365 52.820 132.355 ;
        RECT 51.175 130.645 51.345 131.255 ;
        RECT 51.515 130.865 51.845 131.300 ;
        RECT 52.155 131.195 52.820 131.365 ;
        RECT 52.155 130.905 52.325 131.195 ;
        RECT 52.495 130.645 52.825 131.025 ;
        RECT 52.995 130.905 53.180 133.025 ;
        RECT 53.420 132.735 53.685 133.195 ;
        RECT 53.855 132.600 54.105 133.025 ;
        RECT 54.315 132.750 55.420 132.920 ;
        RECT 53.800 132.470 54.105 132.600 ;
        RECT 53.350 131.275 53.630 132.225 ;
        RECT 53.800 131.365 53.970 132.470 ;
        RECT 54.140 131.685 54.380 132.280 ;
        RECT 54.550 132.215 55.080 132.580 ;
        RECT 54.550 131.515 54.720 132.215 ;
        RECT 55.250 132.135 55.420 132.750 ;
        RECT 55.590 132.395 55.760 133.195 ;
        RECT 55.930 132.695 56.180 133.025 ;
        RECT 56.405 132.725 57.290 132.895 ;
        RECT 55.250 132.045 55.760 132.135 ;
        RECT 53.800 131.235 54.025 131.365 ;
        RECT 54.195 131.295 54.720 131.515 ;
        RECT 54.890 131.875 55.760 132.045 ;
        RECT 53.435 130.645 53.685 131.105 ;
        RECT 53.855 131.095 54.025 131.235 ;
        RECT 54.890 131.095 55.060 131.875 ;
        RECT 55.590 131.805 55.760 131.875 ;
        RECT 55.270 131.625 55.470 131.655 ;
        RECT 55.930 131.625 56.100 132.695 ;
        RECT 56.270 131.805 56.460 132.525 ;
        RECT 55.270 131.325 56.100 131.625 ;
        RECT 56.630 131.595 56.950 132.555 ;
        RECT 53.855 130.925 54.190 131.095 ;
        RECT 54.385 130.925 55.060 131.095 ;
        RECT 55.380 130.645 55.750 131.145 ;
        RECT 55.930 131.095 56.100 131.325 ;
        RECT 56.485 131.265 56.950 131.595 ;
        RECT 57.120 131.885 57.290 132.725 ;
        RECT 57.470 132.695 57.785 133.195 ;
        RECT 58.015 132.465 58.355 133.025 ;
        RECT 57.460 132.090 58.355 132.465 ;
        RECT 58.525 132.185 58.695 133.195 ;
        RECT 58.165 131.885 58.355 132.090 ;
        RECT 58.865 132.135 59.195 132.980 ;
        RECT 59.485 132.135 59.815 132.980 ;
        RECT 59.985 132.185 60.155 133.195 ;
        RECT 60.325 132.465 60.665 133.025 ;
        RECT 60.895 132.695 61.210 133.195 ;
        RECT 61.390 132.725 62.275 132.895 ;
        RECT 58.865 132.055 59.255 132.135 ;
        RECT 59.040 132.005 59.255 132.055 ;
        RECT 57.120 131.555 57.995 131.885 ;
        RECT 58.165 131.555 58.915 131.885 ;
        RECT 57.120 131.095 57.290 131.555 ;
        RECT 58.165 131.385 58.365 131.555 ;
        RECT 59.085 131.425 59.255 132.005 ;
        RECT 59.030 131.385 59.255 131.425 ;
        RECT 55.930 130.925 56.335 131.095 ;
        RECT 56.505 130.925 57.290 131.095 ;
        RECT 57.565 130.645 57.775 131.175 ;
        RECT 58.035 130.860 58.365 131.385 ;
        RECT 58.875 131.300 59.255 131.385 ;
        RECT 59.425 132.055 59.815 132.135 ;
        RECT 60.325 132.090 61.220 132.465 ;
        RECT 59.425 132.005 59.640 132.055 ;
        RECT 59.425 131.425 59.595 132.005 ;
        RECT 60.325 131.885 60.515 132.090 ;
        RECT 61.390 131.885 61.560 132.725 ;
        RECT 62.500 132.695 62.750 133.025 ;
        RECT 59.765 131.555 60.515 131.885 ;
        RECT 60.685 131.555 61.560 131.885 ;
        RECT 59.425 131.385 59.650 131.425 ;
        RECT 60.315 131.385 60.515 131.555 ;
        RECT 59.425 131.300 59.805 131.385 ;
        RECT 58.535 130.645 58.705 131.255 ;
        RECT 58.875 130.865 59.205 131.300 ;
        RECT 59.475 130.865 59.805 131.300 ;
        RECT 59.975 130.645 60.145 131.255 ;
        RECT 60.315 130.860 60.645 131.385 ;
        RECT 60.905 130.645 61.115 131.175 ;
        RECT 61.390 131.095 61.560 131.555 ;
        RECT 61.730 131.595 62.050 132.555 ;
        RECT 62.220 131.805 62.410 132.525 ;
        RECT 62.580 131.625 62.750 132.695 ;
        RECT 62.920 132.395 63.090 133.195 ;
        RECT 63.260 132.750 64.365 132.920 ;
        RECT 63.260 132.135 63.430 132.750 ;
        RECT 64.575 132.600 64.825 133.025 ;
        RECT 64.995 132.735 65.260 133.195 ;
        RECT 63.600 132.215 64.130 132.580 ;
        RECT 64.575 132.470 64.880 132.600 ;
        RECT 62.920 132.045 63.430 132.135 ;
        RECT 62.920 131.875 63.790 132.045 ;
        RECT 62.920 131.805 63.090 131.875 ;
        RECT 63.210 131.625 63.410 131.655 ;
        RECT 61.730 131.265 62.195 131.595 ;
        RECT 62.580 131.325 63.410 131.625 ;
        RECT 62.580 131.095 62.750 131.325 ;
        RECT 61.390 130.925 62.175 131.095 ;
        RECT 62.345 130.925 62.750 131.095 ;
        RECT 62.930 130.645 63.300 131.145 ;
        RECT 63.620 131.095 63.790 131.875 ;
        RECT 63.960 131.515 64.130 132.215 ;
        RECT 64.300 131.685 64.540 132.280 ;
        RECT 63.960 131.295 64.485 131.515 ;
        RECT 64.710 131.365 64.880 132.470 ;
        RECT 64.655 131.235 64.880 131.365 ;
        RECT 65.050 131.275 65.330 132.225 ;
        RECT 64.655 131.095 64.825 131.235 ;
        RECT 63.620 130.925 64.295 131.095 ;
        RECT 64.490 130.925 64.825 131.095 ;
        RECT 64.995 130.645 65.245 131.105 ;
        RECT 65.500 130.905 65.685 133.025 ;
        RECT 65.855 132.695 66.185 133.195 ;
        RECT 66.355 132.525 66.525 133.025 ;
        RECT 65.860 132.355 66.525 132.525 ;
        RECT 65.860 131.365 66.090 132.355 ;
        RECT 67.890 132.225 68.280 132.400 ;
        RECT 68.765 132.395 69.095 133.195 ;
        RECT 69.265 132.405 69.800 133.025 ;
        RECT 66.260 131.535 66.610 132.185 ;
        RECT 67.890 132.055 69.315 132.225 ;
        RECT 65.860 131.195 66.525 131.365 ;
        RECT 67.765 131.325 68.120 131.885 ;
        RECT 65.855 130.645 66.185 131.025 ;
        RECT 66.355 130.905 66.525 131.195 ;
        RECT 68.290 131.155 68.460 132.055 ;
        RECT 68.630 131.325 68.895 131.885 ;
        RECT 69.145 131.555 69.315 132.055 ;
        RECT 69.485 131.385 69.800 132.405 ;
        RECT 70.005 132.030 70.295 133.195 ;
        RECT 70.465 132.055 70.850 133.025 ;
        RECT 71.020 132.735 71.345 133.195 ;
        RECT 71.865 132.565 72.145 133.025 ;
        RECT 71.020 132.345 72.145 132.565 ;
        RECT 67.870 130.645 68.110 131.155 ;
        RECT 68.290 130.825 68.570 131.155 ;
        RECT 68.800 130.645 69.015 131.155 ;
        RECT 69.185 130.815 69.800 131.385 ;
        RECT 70.465 131.385 70.745 132.055 ;
        RECT 71.020 131.885 71.470 132.345 ;
        RECT 72.335 132.175 72.735 133.025 ;
        RECT 73.135 132.735 73.405 133.195 ;
        RECT 73.575 132.565 73.860 133.025 ;
        RECT 70.915 131.555 71.470 131.885 ;
        RECT 71.640 131.615 72.735 132.175 ;
        RECT 71.020 131.445 71.470 131.555 ;
        RECT 70.005 130.645 70.295 131.370 ;
        RECT 70.465 130.815 70.850 131.385 ;
        RECT 71.020 131.275 72.145 131.445 ;
        RECT 71.020 130.645 71.345 131.105 ;
        RECT 71.865 130.815 72.145 131.275 ;
        RECT 72.335 130.815 72.735 131.615 ;
        RECT 72.905 132.345 73.860 132.565 ;
        RECT 72.905 131.445 73.115 132.345 ;
        RECT 73.285 131.615 73.975 132.175 ;
        RECT 74.145 132.055 74.530 133.025 ;
        RECT 74.700 132.735 75.025 133.195 ;
        RECT 75.545 132.565 75.825 133.025 ;
        RECT 74.700 132.345 75.825 132.565 ;
        RECT 72.905 131.275 73.860 131.445 ;
        RECT 73.135 130.645 73.405 131.105 ;
        RECT 73.575 130.815 73.860 131.275 ;
        RECT 74.145 131.385 74.425 132.055 ;
        RECT 74.700 131.885 75.150 132.345 ;
        RECT 76.015 132.175 76.415 133.025 ;
        RECT 76.815 132.735 77.085 133.195 ;
        RECT 77.255 132.565 77.540 133.025 ;
        RECT 74.595 131.555 75.150 131.885 ;
        RECT 75.320 131.615 76.415 132.175 ;
        RECT 74.700 131.445 75.150 131.555 ;
        RECT 74.145 130.815 74.530 131.385 ;
        RECT 74.700 131.275 75.825 131.445 ;
        RECT 74.700 130.645 75.025 131.105 ;
        RECT 75.545 130.815 75.825 131.275 ;
        RECT 76.015 130.815 76.415 131.615 ;
        RECT 76.585 132.345 77.540 132.565 ;
        RECT 76.585 131.445 76.795 132.345 ;
        RECT 76.965 131.615 77.655 132.175 ;
        RECT 77.825 132.055 78.165 133.025 ;
        RECT 78.335 132.055 78.505 133.195 ;
        RECT 78.775 132.395 79.025 133.195 ;
        RECT 79.670 132.225 80.000 133.025 ;
        RECT 80.300 132.395 80.630 133.195 ;
        RECT 80.800 132.225 81.130 133.025 ;
        RECT 78.695 132.055 81.130 132.225 ;
        RECT 81.965 132.105 83.175 133.195 ;
        RECT 77.825 131.445 78.000 132.055 ;
        RECT 78.695 131.805 78.865 132.055 ;
        RECT 78.170 131.635 78.865 131.805 ;
        RECT 79.040 131.635 79.460 131.835 ;
        RECT 79.630 131.635 79.960 131.835 ;
        RECT 80.130 131.635 80.460 131.835 ;
        RECT 76.585 131.275 77.540 131.445 ;
        RECT 76.815 130.645 77.085 131.105 ;
        RECT 77.255 130.815 77.540 131.275 ;
        RECT 77.825 130.815 78.165 131.445 ;
        RECT 78.335 130.645 78.585 131.445 ;
        RECT 78.775 131.295 80.000 131.465 ;
        RECT 78.775 130.815 79.105 131.295 ;
        RECT 79.275 130.645 79.500 131.105 ;
        RECT 79.670 130.815 80.000 131.295 ;
        RECT 80.630 131.425 80.800 132.055 ;
        RECT 80.985 131.635 81.335 131.885 ;
        RECT 81.965 131.565 82.485 132.105 ;
        RECT 80.630 130.815 81.130 131.425 ;
        RECT 82.655 131.395 83.175 131.935 ;
        RECT 81.965 130.645 83.175 131.395 ;
        RECT 5.520 130.475 83.260 130.645 ;
        RECT 5.605 129.725 6.815 130.475 ;
        RECT 6.985 129.930 12.330 130.475 ;
        RECT 5.605 129.185 6.125 129.725 ;
        RECT 6.295 129.015 6.815 129.555 ;
        RECT 8.570 129.100 8.910 129.930 ;
        RECT 12.505 129.705 15.095 130.475 ;
        RECT 15.725 129.825 15.985 130.305 ;
        RECT 16.155 129.935 16.405 130.475 ;
        RECT 5.605 127.925 6.815 129.015 ;
        RECT 10.390 128.360 10.740 129.610 ;
        RECT 12.505 129.185 13.715 129.705 ;
        RECT 13.885 129.015 15.095 129.535 ;
        RECT 6.985 127.925 12.330 128.360 ;
        RECT 12.505 127.925 15.095 129.015 ;
        RECT 15.725 128.795 15.895 129.825 ;
        RECT 16.575 129.795 16.795 130.255 ;
        RECT 16.545 129.770 16.795 129.795 ;
        RECT 16.065 129.175 16.295 129.570 ;
        RECT 16.465 129.345 16.795 129.770 ;
        RECT 16.965 130.095 17.855 130.265 ;
        RECT 16.965 129.370 17.135 130.095 ;
        RECT 17.305 129.540 17.855 129.925 ;
        RECT 18.025 129.755 18.365 130.265 ;
        RECT 16.965 129.300 17.855 129.370 ;
        RECT 16.960 129.275 17.855 129.300 ;
        RECT 16.950 129.260 17.855 129.275 ;
        RECT 16.945 129.245 17.855 129.260 ;
        RECT 16.935 129.240 17.855 129.245 ;
        RECT 16.930 129.230 17.855 129.240 ;
        RECT 16.925 129.220 17.855 129.230 ;
        RECT 16.915 129.215 17.855 129.220 ;
        RECT 16.905 129.205 17.855 129.215 ;
        RECT 16.895 129.200 17.855 129.205 ;
        RECT 16.895 129.195 17.230 129.200 ;
        RECT 16.880 129.190 17.230 129.195 ;
        RECT 16.865 129.180 17.230 129.190 ;
        RECT 16.840 129.175 17.230 129.180 ;
        RECT 16.065 129.170 17.230 129.175 ;
        RECT 16.065 129.135 17.200 129.170 ;
        RECT 16.065 129.110 17.165 129.135 ;
        RECT 16.065 129.080 17.135 129.110 ;
        RECT 16.065 129.050 17.115 129.080 ;
        RECT 16.065 129.020 17.095 129.050 ;
        RECT 16.065 129.010 17.025 129.020 ;
        RECT 16.065 129.000 17.000 129.010 ;
        RECT 16.065 128.985 16.980 129.000 ;
        RECT 16.065 128.970 16.960 128.985 ;
        RECT 16.170 128.960 16.955 128.970 ;
        RECT 16.170 128.925 16.940 128.960 ;
        RECT 15.725 128.095 16.000 128.795 ;
        RECT 16.170 128.675 16.925 128.925 ;
        RECT 17.095 128.605 17.425 128.850 ;
        RECT 17.595 128.750 17.855 129.200 ;
        RECT 17.240 128.580 17.425 128.605 ;
        RECT 17.240 128.480 17.855 128.580 ;
        RECT 16.170 127.925 16.425 128.470 ;
        RECT 16.595 128.095 17.075 128.435 ;
        RECT 17.250 127.925 17.855 128.480 ;
        RECT 18.025 128.355 18.285 129.755 ;
        RECT 18.535 129.675 18.805 130.475 ;
        RECT 18.460 129.235 18.790 129.485 ;
        RECT 18.985 129.235 19.265 130.205 ;
        RECT 19.445 129.235 19.745 130.205 ;
        RECT 19.925 129.235 20.275 130.200 ;
        RECT 20.495 129.975 20.990 130.305 ;
        RECT 18.475 129.065 18.790 129.235 ;
        RECT 20.495 129.065 20.665 129.975 ;
        RECT 18.475 128.895 20.665 129.065 ;
        RECT 18.025 128.095 18.365 128.355 ;
        RECT 18.535 127.925 18.865 128.725 ;
        RECT 19.330 128.095 19.580 128.895 ;
        RECT 19.765 127.925 20.095 128.645 ;
        RECT 20.315 128.095 20.565 128.895 ;
        RECT 20.835 128.485 21.075 129.795 ;
        RECT 21.245 129.640 21.535 130.475 ;
        RECT 21.705 130.075 22.660 130.245 ;
        RECT 23.075 130.085 23.405 130.475 ;
        RECT 21.705 129.195 21.875 130.075 ;
        RECT 23.575 129.905 23.745 130.225 ;
        RECT 23.915 130.085 24.245 130.475 ;
        RECT 22.045 129.735 24.295 129.905 ;
        RECT 22.045 129.235 22.275 129.735 ;
        RECT 22.445 129.315 22.820 129.485 ;
        RECT 21.245 129.025 21.875 129.195 ;
        RECT 22.650 129.115 22.820 129.315 ;
        RECT 22.990 129.285 23.540 129.485 ;
        RECT 23.710 129.115 23.955 129.565 ;
        RECT 20.735 127.925 21.070 128.305 ;
        RECT 21.245 128.095 21.565 129.025 ;
        RECT 22.650 128.945 23.955 129.115 ;
        RECT 24.125 128.775 24.295 129.735 ;
        RECT 24.465 129.725 25.675 130.475 ;
        RECT 25.845 130.095 26.735 130.265 ;
        RECT 24.465 129.185 24.985 129.725 ;
        RECT 25.155 129.015 25.675 129.555 ;
        RECT 25.845 129.540 26.395 129.925 ;
        RECT 26.565 129.370 26.735 130.095 ;
        RECT 21.745 128.605 22.985 128.775 ;
        RECT 21.745 128.095 22.145 128.605 ;
        RECT 22.315 127.925 22.485 128.435 ;
        RECT 22.655 128.095 22.985 128.605 ;
        RECT 23.155 127.925 23.325 128.775 ;
        RECT 23.915 128.095 24.295 128.775 ;
        RECT 24.465 127.925 25.675 129.015 ;
        RECT 25.845 129.300 26.735 129.370 ;
        RECT 26.905 129.770 27.125 130.255 ;
        RECT 27.295 129.935 27.545 130.475 ;
        RECT 27.715 129.825 27.975 130.305 ;
        RECT 26.905 129.345 27.235 129.770 ;
        RECT 25.845 129.275 26.740 129.300 ;
        RECT 25.845 129.260 26.750 129.275 ;
        RECT 25.845 129.245 26.755 129.260 ;
        RECT 25.845 129.240 26.765 129.245 ;
        RECT 25.845 129.230 26.770 129.240 ;
        RECT 25.845 129.220 26.775 129.230 ;
        RECT 25.845 129.215 26.785 129.220 ;
        RECT 25.845 129.205 26.795 129.215 ;
        RECT 25.845 129.200 26.805 129.205 ;
        RECT 25.845 128.750 26.105 129.200 ;
        RECT 26.470 129.195 26.805 129.200 ;
        RECT 26.470 129.190 26.820 129.195 ;
        RECT 26.470 129.180 26.835 129.190 ;
        RECT 26.470 129.175 26.860 129.180 ;
        RECT 27.405 129.175 27.635 129.570 ;
        RECT 26.470 129.170 27.635 129.175 ;
        RECT 26.500 129.135 27.635 129.170 ;
        RECT 26.535 129.110 27.635 129.135 ;
        RECT 26.565 129.080 27.635 129.110 ;
        RECT 26.585 129.050 27.635 129.080 ;
        RECT 26.605 129.020 27.635 129.050 ;
        RECT 26.675 129.010 27.635 129.020 ;
        RECT 26.700 129.000 27.635 129.010 ;
        RECT 26.720 128.985 27.635 129.000 ;
        RECT 26.740 128.970 27.635 128.985 ;
        RECT 26.745 128.960 27.530 128.970 ;
        RECT 26.760 128.925 27.530 128.960 ;
        RECT 26.275 128.605 26.605 128.850 ;
        RECT 26.775 128.675 27.530 128.925 ;
        RECT 27.805 128.795 27.975 129.825 ;
        RECT 28.165 129.665 28.405 130.475 ;
        RECT 28.575 129.665 28.905 130.305 ;
        RECT 29.075 129.665 29.345 130.475 ;
        RECT 28.145 129.235 28.495 129.485 ;
        RECT 28.665 129.065 28.835 129.665 ;
        RECT 30.045 129.655 30.255 130.475 ;
        RECT 30.425 129.675 30.755 130.305 ;
        RECT 29.005 129.235 29.355 129.485 ;
        RECT 30.425 129.075 30.675 129.675 ;
        RECT 30.925 129.655 31.155 130.475 ;
        RECT 31.365 129.750 31.655 130.475 ;
        RECT 32.400 129.845 32.685 130.305 ;
        RECT 32.855 130.015 33.125 130.475 ;
        RECT 32.400 129.675 33.355 129.845 ;
        RECT 30.845 129.235 31.175 129.485 ;
        RECT 26.275 128.580 26.460 128.605 ;
        RECT 25.845 128.480 26.460 128.580 ;
        RECT 25.845 127.925 26.450 128.480 ;
        RECT 26.625 128.095 27.105 128.435 ;
        RECT 27.275 127.925 27.530 128.470 ;
        RECT 27.700 128.095 27.975 128.795 ;
        RECT 28.155 128.895 28.835 129.065 ;
        RECT 28.155 128.110 28.485 128.895 ;
        RECT 29.015 127.925 29.345 129.065 ;
        RECT 30.045 127.925 30.255 129.065 ;
        RECT 30.425 128.095 30.755 129.075 ;
        RECT 30.925 127.925 31.155 129.065 ;
        RECT 31.365 127.925 31.655 129.090 ;
        RECT 32.285 128.945 32.975 129.505 ;
        RECT 33.145 128.775 33.355 129.675 ;
        RECT 32.400 128.555 33.355 128.775 ;
        RECT 33.525 129.505 33.925 130.305 ;
        RECT 34.115 129.845 34.395 130.305 ;
        RECT 34.915 130.015 35.240 130.475 ;
        RECT 34.115 129.675 35.240 129.845 ;
        RECT 35.410 129.735 35.795 130.305 ;
        RECT 36.025 130.015 36.270 130.475 ;
        RECT 34.790 129.565 35.240 129.675 ;
        RECT 33.525 128.945 34.620 129.505 ;
        RECT 34.790 129.235 35.345 129.565 ;
        RECT 32.400 128.095 32.685 128.555 ;
        RECT 32.855 127.925 33.125 128.385 ;
        RECT 33.525 128.095 33.925 128.945 ;
        RECT 34.790 128.775 35.240 129.235 ;
        RECT 35.515 129.065 35.795 129.735 ;
        RECT 35.965 129.235 36.280 129.845 ;
        RECT 36.450 129.485 36.700 130.295 ;
        RECT 36.870 129.950 37.130 130.475 ;
        RECT 37.300 129.825 37.560 130.280 ;
        RECT 37.730 129.995 37.990 130.475 ;
        RECT 38.160 129.825 38.420 130.280 ;
        RECT 38.590 129.995 38.850 130.475 ;
        RECT 39.020 129.825 39.280 130.280 ;
        RECT 39.450 129.995 39.710 130.475 ;
        RECT 39.880 129.825 40.140 130.280 ;
        RECT 40.310 129.995 40.610 130.475 ;
        RECT 41.115 129.925 41.285 130.215 ;
        RECT 41.455 130.095 41.785 130.475 ;
        RECT 37.300 129.655 40.610 129.825 ;
        RECT 41.115 129.755 41.780 129.925 ;
        RECT 36.450 129.235 39.470 129.485 ;
        RECT 34.115 128.555 35.240 128.775 ;
        RECT 34.115 128.095 34.395 128.555 ;
        RECT 34.915 127.925 35.240 128.385 ;
        RECT 35.410 128.095 35.795 129.065 ;
        RECT 35.975 127.925 36.270 129.035 ;
        RECT 36.450 128.100 36.700 129.235 ;
        RECT 39.640 129.065 40.610 129.655 ;
        RECT 36.870 127.925 37.130 129.035 ;
        RECT 37.300 128.825 40.610 129.065 ;
        RECT 41.030 128.935 41.380 129.585 ;
        RECT 37.300 128.100 37.560 128.825 ;
        RECT 37.730 127.925 37.990 128.655 ;
        RECT 38.160 128.100 38.420 128.825 ;
        RECT 38.590 127.925 38.850 128.655 ;
        RECT 39.020 128.100 39.280 128.825 ;
        RECT 39.450 127.925 39.710 128.655 ;
        RECT 39.880 128.100 40.140 128.825 ;
        RECT 41.550 128.765 41.780 129.755 ;
        RECT 40.310 127.925 40.605 128.655 ;
        RECT 41.115 128.595 41.780 128.765 ;
        RECT 41.115 128.095 41.285 128.595 ;
        RECT 41.455 127.925 41.785 128.425 ;
        RECT 41.955 128.095 42.140 130.215 ;
        RECT 42.395 130.015 42.645 130.475 ;
        RECT 42.815 130.025 43.150 130.195 ;
        RECT 43.345 130.025 44.020 130.195 ;
        RECT 42.815 129.885 42.985 130.025 ;
        RECT 42.310 128.895 42.590 129.845 ;
        RECT 42.760 129.755 42.985 129.885 ;
        RECT 42.760 128.650 42.930 129.755 ;
        RECT 43.155 129.605 43.680 129.825 ;
        RECT 43.100 128.840 43.340 129.435 ;
        RECT 43.510 128.905 43.680 129.605 ;
        RECT 43.850 129.245 44.020 130.025 ;
        RECT 44.340 129.975 44.710 130.475 ;
        RECT 44.890 130.025 45.295 130.195 ;
        RECT 45.465 130.025 46.250 130.195 ;
        RECT 44.890 129.795 45.060 130.025 ;
        RECT 44.230 129.495 45.060 129.795 ;
        RECT 45.445 129.525 45.910 129.855 ;
        RECT 44.230 129.465 44.430 129.495 ;
        RECT 44.550 129.245 44.720 129.315 ;
        RECT 43.850 129.075 44.720 129.245 ;
        RECT 44.210 128.985 44.720 129.075 ;
        RECT 42.760 128.520 43.065 128.650 ;
        RECT 43.510 128.540 44.040 128.905 ;
        RECT 42.380 127.925 42.645 128.385 ;
        RECT 42.815 128.095 43.065 128.520 ;
        RECT 44.210 128.370 44.380 128.985 ;
        RECT 43.275 128.200 44.380 128.370 ;
        RECT 44.550 127.925 44.720 128.725 ;
        RECT 44.890 128.425 45.060 129.495 ;
        RECT 45.230 128.595 45.420 129.315 ;
        RECT 45.590 128.565 45.910 129.525 ;
        RECT 46.080 129.565 46.250 130.025 ;
        RECT 46.525 129.945 46.735 130.475 ;
        RECT 46.995 129.735 47.325 130.260 ;
        RECT 47.495 129.865 47.665 130.475 ;
        RECT 47.835 129.820 48.165 130.255 ;
        RECT 47.835 129.735 48.215 129.820 ;
        RECT 47.125 129.565 47.325 129.735 ;
        RECT 47.990 129.695 48.215 129.735 ;
        RECT 46.080 129.235 46.955 129.565 ;
        RECT 47.125 129.235 47.875 129.565 ;
        RECT 44.890 128.095 45.140 128.425 ;
        RECT 46.080 128.395 46.250 129.235 ;
        RECT 47.125 129.030 47.315 129.235 ;
        RECT 48.045 129.115 48.215 129.695 ;
        RECT 48.000 129.065 48.215 129.115 ;
        RECT 46.420 128.655 47.315 129.030 ;
        RECT 47.825 128.985 48.215 129.065 ;
        RECT 48.390 129.735 48.645 130.305 ;
        RECT 48.815 130.075 49.145 130.475 ;
        RECT 49.570 129.940 50.100 130.305 ;
        RECT 49.570 129.905 49.745 129.940 ;
        RECT 48.815 129.735 49.745 129.905 ;
        RECT 50.290 129.795 50.565 130.305 ;
        RECT 48.390 129.065 48.560 129.735 ;
        RECT 48.815 129.565 48.985 129.735 ;
        RECT 48.730 129.235 48.985 129.565 ;
        RECT 49.210 129.235 49.405 129.565 ;
        RECT 45.365 128.225 46.250 128.395 ;
        RECT 46.430 127.925 46.745 128.425 ;
        RECT 46.975 128.095 47.315 128.655 ;
        RECT 47.485 127.925 47.655 128.935 ;
        RECT 47.825 128.140 48.155 128.985 ;
        RECT 48.390 128.095 48.725 129.065 ;
        RECT 48.895 127.925 49.065 129.065 ;
        RECT 49.235 128.265 49.405 129.235 ;
        RECT 49.575 128.605 49.745 129.735 ;
        RECT 49.915 128.945 50.085 129.745 ;
        RECT 50.285 129.625 50.565 129.795 ;
        RECT 50.290 129.145 50.565 129.625 ;
        RECT 50.735 128.945 50.925 130.305 ;
        RECT 51.105 129.940 51.615 130.475 ;
        RECT 51.835 129.665 52.080 130.270 ;
        RECT 52.990 129.735 53.245 130.305 ;
        RECT 53.415 130.075 53.745 130.475 ;
        RECT 54.170 129.940 54.700 130.305 ;
        RECT 54.890 130.135 55.165 130.305 ;
        RECT 54.885 129.965 55.165 130.135 ;
        RECT 54.170 129.905 54.345 129.940 ;
        RECT 53.415 129.735 54.345 129.905 ;
        RECT 51.125 129.495 52.355 129.665 ;
        RECT 49.915 128.775 50.925 128.945 ;
        RECT 51.095 128.930 51.845 129.120 ;
        RECT 49.575 128.435 50.700 128.605 ;
        RECT 51.095 128.265 51.265 128.930 ;
        RECT 52.015 128.685 52.355 129.495 ;
        RECT 49.235 128.095 51.265 128.265 ;
        RECT 51.435 127.925 51.605 128.685 ;
        RECT 51.840 128.275 52.355 128.685 ;
        RECT 52.990 129.065 53.160 129.735 ;
        RECT 53.415 129.565 53.585 129.735 ;
        RECT 53.330 129.235 53.585 129.565 ;
        RECT 53.810 129.235 54.005 129.565 ;
        RECT 52.990 128.095 53.325 129.065 ;
        RECT 53.495 127.925 53.665 129.065 ;
        RECT 53.835 128.265 54.005 129.235 ;
        RECT 54.175 128.605 54.345 129.735 ;
        RECT 54.515 128.945 54.685 129.745 ;
        RECT 54.890 129.145 55.165 129.965 ;
        RECT 55.335 128.945 55.525 130.305 ;
        RECT 55.705 129.940 56.215 130.475 ;
        RECT 56.435 129.665 56.680 130.270 ;
        RECT 57.125 129.750 57.415 130.475 ;
        RECT 57.585 129.725 58.795 130.475 ;
        RECT 59.015 129.820 59.345 130.255 ;
        RECT 59.515 129.865 59.685 130.475 ;
        RECT 58.965 129.735 59.345 129.820 ;
        RECT 59.855 129.735 60.185 130.260 ;
        RECT 60.445 129.945 60.655 130.475 ;
        RECT 60.930 130.025 61.715 130.195 ;
        RECT 61.885 130.025 62.290 130.195 ;
        RECT 55.725 129.495 56.955 129.665 ;
        RECT 54.515 128.775 55.525 128.945 ;
        RECT 55.695 128.930 56.445 129.120 ;
        RECT 54.175 128.435 55.300 128.605 ;
        RECT 55.695 128.265 55.865 128.930 ;
        RECT 56.615 128.685 56.955 129.495 ;
        RECT 57.585 129.185 58.105 129.725 ;
        RECT 58.965 129.695 59.190 129.735 ;
        RECT 53.835 128.095 55.865 128.265 ;
        RECT 56.035 127.925 56.205 128.685 ;
        RECT 56.440 128.275 56.955 128.685 ;
        RECT 57.125 127.925 57.415 129.090 ;
        RECT 58.275 129.015 58.795 129.555 ;
        RECT 57.585 127.925 58.795 129.015 ;
        RECT 58.965 129.115 59.135 129.695 ;
        RECT 59.855 129.565 60.055 129.735 ;
        RECT 60.930 129.565 61.100 130.025 ;
        RECT 59.305 129.235 60.055 129.565 ;
        RECT 60.225 129.235 61.100 129.565 ;
        RECT 58.965 129.065 59.180 129.115 ;
        RECT 58.965 128.985 59.355 129.065 ;
        RECT 59.025 128.140 59.355 128.985 ;
        RECT 59.865 129.030 60.055 129.235 ;
        RECT 59.525 127.925 59.695 128.935 ;
        RECT 59.865 128.655 60.760 129.030 ;
        RECT 59.865 128.095 60.205 128.655 ;
        RECT 60.435 127.925 60.750 128.425 ;
        RECT 60.930 128.395 61.100 129.235 ;
        RECT 61.270 129.525 61.735 129.855 ;
        RECT 62.120 129.795 62.290 130.025 ;
        RECT 62.470 129.975 62.840 130.475 ;
        RECT 63.160 130.025 63.835 130.195 ;
        RECT 64.030 130.025 64.365 130.195 ;
        RECT 61.270 128.565 61.590 129.525 ;
        RECT 62.120 129.495 62.950 129.795 ;
        RECT 61.760 128.595 61.950 129.315 ;
        RECT 62.120 128.425 62.290 129.495 ;
        RECT 62.750 129.465 62.950 129.495 ;
        RECT 62.460 129.245 62.630 129.315 ;
        RECT 63.160 129.245 63.330 130.025 ;
        RECT 64.195 129.885 64.365 130.025 ;
        RECT 64.535 130.015 64.785 130.475 ;
        RECT 62.460 129.075 63.330 129.245 ;
        RECT 63.500 129.605 64.025 129.825 ;
        RECT 64.195 129.755 64.420 129.885 ;
        RECT 62.460 128.985 62.970 129.075 ;
        RECT 60.930 128.225 61.815 128.395 ;
        RECT 62.040 128.095 62.290 128.425 ;
        RECT 62.460 127.925 62.630 128.725 ;
        RECT 62.800 128.370 62.970 128.985 ;
        RECT 63.500 128.905 63.670 129.605 ;
        RECT 63.140 128.540 63.670 128.905 ;
        RECT 63.840 128.840 64.080 129.435 ;
        RECT 64.250 128.650 64.420 129.755 ;
        RECT 64.590 128.895 64.870 129.845 ;
        RECT 64.115 128.520 64.420 128.650 ;
        RECT 62.800 128.200 63.905 128.370 ;
        RECT 64.115 128.095 64.365 128.520 ;
        RECT 64.535 127.925 64.800 128.385 ;
        RECT 65.040 128.095 65.225 130.215 ;
        RECT 65.395 130.095 65.725 130.475 ;
        RECT 65.895 129.925 66.065 130.215 ;
        RECT 66.385 130.015 66.630 130.475 ;
        RECT 65.400 129.755 66.065 129.925 ;
        RECT 65.400 128.765 65.630 129.755 ;
        RECT 65.800 128.935 66.150 129.585 ;
        RECT 66.325 129.235 66.640 129.845 ;
        RECT 66.810 129.485 67.060 130.295 ;
        RECT 67.230 129.950 67.490 130.475 ;
        RECT 67.660 129.825 67.920 130.280 ;
        RECT 68.090 129.995 68.350 130.475 ;
        RECT 68.520 129.825 68.780 130.280 ;
        RECT 68.950 129.995 69.210 130.475 ;
        RECT 69.380 129.825 69.640 130.280 ;
        RECT 69.810 129.995 70.070 130.475 ;
        RECT 70.240 129.825 70.500 130.280 ;
        RECT 70.670 129.995 70.970 130.475 ;
        RECT 67.660 129.655 70.970 129.825 ;
        RECT 66.810 129.235 69.830 129.485 ;
        RECT 65.400 128.595 66.065 128.765 ;
        RECT 65.395 127.925 65.725 128.425 ;
        RECT 65.895 128.095 66.065 128.595 ;
        RECT 66.335 127.925 66.630 129.035 ;
        RECT 66.810 128.100 67.060 129.235 ;
        RECT 70.000 129.065 70.970 129.655 ;
        RECT 67.230 127.925 67.490 129.035 ;
        RECT 67.660 128.825 70.970 129.065 ;
        RECT 71.390 129.735 71.645 130.305 ;
        RECT 71.815 130.075 72.145 130.475 ;
        RECT 72.570 129.940 73.100 130.305 ;
        RECT 73.290 130.135 73.565 130.305 ;
        RECT 73.285 129.965 73.565 130.135 ;
        RECT 72.570 129.905 72.745 129.940 ;
        RECT 71.815 129.735 72.745 129.905 ;
        RECT 71.390 129.065 71.560 129.735 ;
        RECT 71.815 129.565 71.985 129.735 ;
        RECT 71.730 129.235 71.985 129.565 ;
        RECT 72.210 129.235 72.405 129.565 ;
        RECT 67.660 128.100 67.920 128.825 ;
        RECT 68.090 127.925 68.350 128.655 ;
        RECT 68.520 128.100 68.780 128.825 ;
        RECT 68.950 127.925 69.210 128.655 ;
        RECT 69.380 128.100 69.640 128.825 ;
        RECT 69.810 127.925 70.070 128.655 ;
        RECT 70.240 128.100 70.500 128.825 ;
        RECT 70.670 127.925 70.965 128.655 ;
        RECT 71.390 128.095 71.725 129.065 ;
        RECT 71.895 127.925 72.065 129.065 ;
        RECT 72.235 128.265 72.405 129.235 ;
        RECT 72.575 128.605 72.745 129.735 ;
        RECT 72.915 128.945 73.085 129.745 ;
        RECT 73.290 129.145 73.565 129.965 ;
        RECT 73.735 128.945 73.925 130.305 ;
        RECT 74.105 129.940 74.615 130.475 ;
        RECT 74.835 129.665 75.080 130.270 ;
        RECT 74.125 129.495 75.355 129.665 ;
        RECT 72.915 128.775 73.925 128.945 ;
        RECT 74.095 128.930 74.845 129.120 ;
        RECT 72.575 128.435 73.700 128.605 ;
        RECT 74.095 128.265 74.265 128.930 ;
        RECT 75.015 128.685 75.355 129.495 ;
        RECT 72.235 128.095 74.265 128.265 ;
        RECT 74.435 127.925 74.605 128.685 ;
        RECT 74.840 128.275 75.355 128.685 ;
        RECT 75.530 128.875 75.865 130.295 ;
        RECT 76.045 130.105 76.790 130.475 ;
        RECT 77.355 129.935 77.610 130.295 ;
        RECT 77.790 130.105 78.120 130.475 ;
        RECT 78.300 129.935 78.525 130.295 ;
        RECT 76.040 129.745 78.525 129.935 ;
        RECT 76.040 129.055 76.265 129.745 ;
        RECT 78.780 129.735 79.395 130.305 ;
        RECT 79.565 129.965 79.780 130.475 ;
        RECT 80.010 129.965 80.290 130.295 ;
        RECT 80.470 129.965 80.710 130.475 ;
        RECT 76.465 129.235 76.745 129.565 ;
        RECT 76.925 129.235 77.500 129.565 ;
        RECT 77.680 129.235 78.115 129.565 ;
        RECT 78.295 129.235 78.565 129.565 ;
        RECT 76.040 128.875 78.535 129.055 ;
        RECT 75.530 128.105 75.795 128.875 ;
        RECT 75.965 127.925 76.295 128.645 ;
        RECT 76.485 128.465 77.675 128.695 ;
        RECT 76.485 128.105 76.745 128.465 ;
        RECT 76.915 127.925 77.245 128.295 ;
        RECT 77.415 128.105 77.675 128.465 ;
        RECT 78.245 128.105 78.535 128.875 ;
        RECT 78.780 128.715 79.095 129.735 ;
        RECT 79.265 129.065 79.435 129.565 ;
        RECT 79.685 129.235 79.950 129.795 ;
        RECT 80.120 129.065 80.290 129.965 ;
        RECT 80.460 129.235 80.815 129.795 ;
        RECT 81.965 129.725 83.175 130.475 ;
        RECT 79.265 128.895 80.690 129.065 ;
        RECT 78.780 128.095 79.315 128.715 ;
        RECT 79.485 127.925 79.815 128.725 ;
        RECT 80.300 128.720 80.690 128.895 ;
        RECT 81.965 129.015 82.485 129.555 ;
        RECT 82.655 129.185 83.175 129.725 ;
        RECT 81.965 127.925 83.175 129.015 ;
        RECT 5.520 127.755 83.260 127.925 ;
        RECT 5.605 126.665 6.815 127.755 ;
        RECT 5.605 125.955 6.125 126.495 ;
        RECT 6.295 126.125 6.815 126.665 ;
        RECT 7.075 126.825 7.245 127.585 ;
        RECT 7.425 126.995 7.755 127.755 ;
        RECT 7.075 126.655 7.740 126.825 ;
        RECT 7.925 126.680 8.195 127.585 ;
        RECT 8.365 127.320 13.710 127.755 ;
        RECT 7.570 126.510 7.740 126.655 ;
        RECT 7.005 126.105 7.335 126.475 ;
        RECT 7.570 126.180 7.855 126.510 ;
        RECT 5.605 125.205 6.815 125.955 ;
        RECT 7.570 125.925 7.740 126.180 ;
        RECT 7.075 125.755 7.740 125.925 ;
        RECT 8.025 125.880 8.195 126.680 ;
        RECT 7.075 125.375 7.245 125.755 ;
        RECT 7.425 125.205 7.755 125.585 ;
        RECT 7.935 125.375 8.195 125.880 ;
        RECT 9.950 125.750 10.290 126.580 ;
        RECT 11.770 126.070 12.120 127.320 ;
        RECT 13.885 126.665 17.395 127.755 ;
        RECT 13.885 125.975 15.535 126.495 ;
        RECT 15.705 126.145 17.395 126.665 ;
        RECT 18.485 126.590 18.775 127.755 ;
        RECT 18.945 127.320 24.290 127.755 ;
        RECT 8.365 125.205 13.710 125.750 ;
        RECT 13.885 125.205 17.395 125.975 ;
        RECT 18.485 125.205 18.775 125.930 ;
        RECT 20.530 125.750 20.870 126.580 ;
        RECT 22.350 126.070 22.700 127.320 ;
        RECT 24.465 126.665 27.055 127.755 ;
        RECT 27.935 127.025 28.230 127.755 ;
        RECT 28.400 126.855 28.660 127.580 ;
        RECT 28.830 127.025 29.090 127.755 ;
        RECT 29.260 126.855 29.520 127.580 ;
        RECT 29.690 127.025 29.950 127.755 ;
        RECT 30.120 126.855 30.380 127.580 ;
        RECT 30.550 127.025 30.810 127.755 ;
        RECT 30.980 126.855 31.240 127.580 ;
        RECT 24.465 125.975 25.675 126.495 ;
        RECT 25.845 126.145 27.055 126.665 ;
        RECT 27.930 126.615 31.240 126.855 ;
        RECT 31.410 126.645 31.670 127.755 ;
        RECT 27.930 126.025 28.900 126.615 ;
        RECT 31.840 126.445 32.090 127.580 ;
        RECT 32.270 126.645 32.565 127.755 ;
        RECT 33.205 127.165 33.905 127.585 ;
        RECT 34.105 127.395 34.435 127.755 ;
        RECT 34.605 127.165 34.935 127.565 ;
        RECT 33.205 126.935 34.935 127.165 ;
        RECT 29.070 126.195 32.090 126.445 ;
        RECT 18.945 125.205 24.290 125.750 ;
        RECT 24.465 125.205 27.055 125.975 ;
        RECT 27.930 125.855 31.240 126.025 ;
        RECT 27.930 125.205 28.230 125.685 ;
        RECT 28.400 125.400 28.660 125.855 ;
        RECT 28.830 125.205 29.090 125.685 ;
        RECT 29.260 125.400 29.520 125.855 ;
        RECT 29.690 125.205 29.950 125.685 ;
        RECT 30.120 125.400 30.380 125.855 ;
        RECT 30.550 125.205 30.810 125.685 ;
        RECT 30.980 125.400 31.240 125.855 ;
        RECT 31.410 125.205 31.670 125.730 ;
        RECT 31.840 125.385 32.090 126.195 ;
        RECT 32.260 125.835 32.575 126.445 ;
        RECT 33.205 125.965 33.410 126.935 ;
        RECT 33.580 126.195 33.910 126.735 ;
        RECT 34.085 126.445 34.410 126.735 ;
        RECT 34.605 126.715 34.935 126.935 ;
        RECT 35.105 126.445 35.275 127.415 ;
        RECT 35.455 126.695 35.785 127.755 ;
        RECT 36.495 126.750 36.750 127.555 ;
        RECT 36.920 126.920 37.180 127.755 ;
        RECT 37.350 126.750 37.610 127.555 ;
        RECT 37.780 126.920 38.035 127.755 ;
        RECT 36.495 126.580 38.095 126.750 ;
        RECT 34.085 126.115 34.580 126.445 ;
        RECT 34.900 126.115 35.275 126.445 ;
        RECT 35.485 126.115 35.795 126.445 ;
        RECT 36.425 126.185 37.645 126.410 ;
        RECT 37.815 126.015 38.095 126.580 ;
        RECT 32.270 125.205 32.515 125.665 ;
        RECT 33.205 125.375 33.915 125.965 ;
        RECT 34.425 125.735 35.785 125.945 ;
        RECT 34.425 125.375 34.755 125.735 ;
        RECT 34.955 125.205 35.285 125.565 ;
        RECT 35.455 125.375 35.785 125.735 ;
        RECT 37.365 125.845 38.095 126.015 ;
        RECT 38.270 126.615 38.545 127.585 ;
        RECT 38.755 126.955 39.035 127.755 ;
        RECT 39.205 127.245 40.395 127.535 ;
        RECT 39.205 126.905 40.375 127.075 ;
        RECT 39.205 126.785 39.375 126.905 ;
        RECT 38.715 126.615 39.375 126.785 ;
        RECT 38.270 125.880 38.440 126.615 ;
        RECT 38.715 126.445 38.885 126.615 ;
        RECT 39.685 126.445 39.880 126.735 ;
        RECT 40.050 126.615 40.375 126.905 ;
        RECT 40.565 126.615 40.950 127.585 ;
        RECT 41.120 127.295 41.445 127.755 ;
        RECT 41.965 127.125 42.245 127.585 ;
        RECT 41.120 126.905 42.245 127.125 ;
        RECT 38.610 126.115 38.885 126.445 ;
        RECT 39.055 126.115 39.880 126.445 ;
        RECT 40.050 126.115 40.395 126.445 ;
        RECT 38.715 125.945 38.885 126.115 ;
        RECT 40.565 125.945 40.845 126.615 ;
        RECT 41.120 126.445 41.570 126.905 ;
        RECT 42.435 126.735 42.835 127.585 ;
        RECT 43.235 127.295 43.505 127.755 ;
        RECT 43.675 127.125 43.960 127.585 ;
        RECT 41.015 126.115 41.570 126.445 ;
        RECT 41.740 126.175 42.835 126.735 ;
        RECT 41.120 126.005 41.570 126.115 ;
        RECT 36.900 125.205 37.195 125.730 ;
        RECT 37.365 125.400 37.590 125.845 ;
        RECT 37.760 125.205 38.090 125.675 ;
        RECT 38.270 125.535 38.545 125.880 ;
        RECT 38.715 125.775 40.380 125.945 ;
        RECT 38.735 125.205 39.115 125.605 ;
        RECT 39.285 125.425 39.455 125.775 ;
        RECT 39.625 125.205 39.955 125.605 ;
        RECT 40.125 125.425 40.380 125.775 ;
        RECT 40.565 125.375 40.950 125.945 ;
        RECT 41.120 125.835 42.245 126.005 ;
        RECT 41.120 125.205 41.445 125.665 ;
        RECT 41.965 125.375 42.245 125.835 ;
        RECT 42.435 125.375 42.835 126.175 ;
        RECT 43.005 126.905 43.960 127.125 ;
        RECT 43.005 126.005 43.215 126.905 ;
        RECT 43.385 126.175 44.075 126.735 ;
        RECT 44.245 126.590 44.535 127.755 ;
        RECT 45.170 126.615 45.505 127.585 ;
        RECT 45.675 126.615 45.845 127.755 ;
        RECT 46.015 127.415 48.045 127.585 ;
        RECT 43.005 125.835 43.960 126.005 ;
        RECT 45.170 125.945 45.340 126.615 ;
        RECT 46.015 126.445 46.185 127.415 ;
        RECT 45.510 126.115 45.765 126.445 ;
        RECT 45.990 126.115 46.185 126.445 ;
        RECT 46.355 127.075 47.480 127.245 ;
        RECT 45.595 125.945 45.765 126.115 ;
        RECT 46.355 125.945 46.525 127.075 ;
        RECT 43.235 125.205 43.505 125.665 ;
        RECT 43.675 125.375 43.960 125.835 ;
        RECT 44.245 125.205 44.535 125.930 ;
        RECT 45.170 125.375 45.425 125.945 ;
        RECT 45.595 125.775 46.525 125.945 ;
        RECT 46.695 126.735 47.705 126.905 ;
        RECT 46.695 125.935 46.865 126.735 ;
        RECT 47.070 126.055 47.345 126.535 ;
        RECT 47.065 125.885 47.345 126.055 ;
        RECT 46.350 125.740 46.525 125.775 ;
        RECT 45.595 125.205 45.925 125.605 ;
        RECT 46.350 125.375 46.880 125.740 ;
        RECT 47.070 125.375 47.345 125.885 ;
        RECT 47.515 125.375 47.705 126.735 ;
        RECT 47.875 126.750 48.045 127.415 ;
        RECT 48.215 126.995 48.385 127.755 ;
        RECT 48.620 126.995 49.135 127.405 ;
        RECT 47.875 126.560 48.625 126.750 ;
        RECT 48.795 126.185 49.135 126.995 ;
        RECT 47.905 126.015 49.135 126.185 ;
        RECT 49.305 126.615 49.690 127.585 ;
        RECT 49.860 127.295 50.185 127.755 ;
        RECT 50.705 127.125 50.985 127.585 ;
        RECT 49.860 126.905 50.985 127.125 ;
        RECT 47.885 125.205 48.395 125.740 ;
        RECT 48.615 125.410 48.860 126.015 ;
        RECT 49.305 125.945 49.585 126.615 ;
        RECT 49.860 126.445 50.310 126.905 ;
        RECT 51.175 126.735 51.575 127.585 ;
        RECT 51.975 127.295 52.245 127.755 ;
        RECT 52.415 127.125 52.700 127.585 ;
        RECT 49.755 126.115 50.310 126.445 ;
        RECT 50.480 126.175 51.575 126.735 ;
        RECT 49.860 126.005 50.310 126.115 ;
        RECT 49.305 125.375 49.690 125.945 ;
        RECT 49.860 125.835 50.985 126.005 ;
        RECT 49.860 125.205 50.185 125.665 ;
        RECT 50.705 125.375 50.985 125.835 ;
        RECT 51.175 125.375 51.575 126.175 ;
        RECT 51.745 126.905 52.700 127.125 ;
        RECT 51.745 126.005 51.955 126.905 ;
        RECT 52.125 126.175 52.815 126.735 ;
        RECT 52.985 126.665 54.655 127.755 ;
        RECT 51.745 125.835 52.700 126.005 ;
        RECT 51.975 125.205 52.245 125.665 ;
        RECT 52.415 125.375 52.700 125.835 ;
        RECT 52.985 125.975 53.735 126.495 ;
        RECT 53.905 126.145 54.655 126.665 ;
        RECT 54.830 126.605 55.090 127.755 ;
        RECT 55.265 126.680 55.520 127.585 ;
        RECT 55.690 126.995 56.020 127.755 ;
        RECT 56.235 126.825 56.405 127.585 ;
        RECT 56.780 127.125 57.065 127.585 ;
        RECT 57.235 127.295 57.505 127.755 ;
        RECT 56.780 126.905 57.735 127.125 ;
        RECT 52.985 125.205 54.655 125.975 ;
        RECT 54.830 125.205 55.090 126.045 ;
        RECT 55.265 125.950 55.435 126.680 ;
        RECT 55.690 126.655 56.405 126.825 ;
        RECT 55.690 126.445 55.860 126.655 ;
        RECT 55.605 126.115 55.860 126.445 ;
        RECT 55.265 125.375 55.520 125.950 ;
        RECT 55.690 125.925 55.860 126.115 ;
        RECT 56.140 126.105 56.495 126.475 ;
        RECT 56.665 126.175 57.355 126.735 ;
        RECT 57.525 126.005 57.735 126.905 ;
        RECT 55.690 125.755 56.405 125.925 ;
        RECT 55.690 125.205 56.020 125.585 ;
        RECT 56.235 125.375 56.405 125.755 ;
        RECT 56.780 125.835 57.735 126.005 ;
        RECT 57.905 126.735 58.305 127.585 ;
        RECT 58.495 127.125 58.775 127.585 ;
        RECT 59.295 127.295 59.620 127.755 ;
        RECT 58.495 126.905 59.620 127.125 ;
        RECT 57.905 126.175 59.000 126.735 ;
        RECT 59.170 126.445 59.620 126.905 ;
        RECT 59.790 126.615 60.175 127.585 ;
        RECT 56.780 125.375 57.065 125.835 ;
        RECT 57.235 125.205 57.505 125.665 ;
        RECT 57.905 125.375 58.305 126.175 ;
        RECT 59.170 126.115 59.725 126.445 ;
        RECT 59.170 126.005 59.620 126.115 ;
        RECT 58.495 125.835 59.620 126.005 ;
        RECT 59.895 125.945 60.175 126.615 ;
        RECT 60.350 126.605 60.610 127.755 ;
        RECT 60.785 126.680 61.040 127.585 ;
        RECT 61.210 126.995 61.540 127.755 ;
        RECT 61.755 126.825 61.925 127.585 ;
        RECT 58.495 125.375 58.775 125.835 ;
        RECT 59.295 125.205 59.620 125.665 ;
        RECT 59.790 125.375 60.175 125.945 ;
        RECT 60.350 125.205 60.610 126.045 ;
        RECT 60.785 125.950 60.955 126.680 ;
        RECT 61.210 126.655 61.925 126.825 ;
        RECT 61.210 126.445 61.380 126.655 ;
        RECT 62.185 126.615 62.570 127.585 ;
        RECT 62.740 127.295 63.065 127.755 ;
        RECT 63.585 127.125 63.865 127.585 ;
        RECT 62.740 126.905 63.865 127.125 ;
        RECT 61.125 126.115 61.380 126.445 ;
        RECT 60.785 125.375 61.040 125.950 ;
        RECT 61.210 125.925 61.380 126.115 ;
        RECT 61.660 126.105 62.015 126.475 ;
        RECT 62.185 125.945 62.465 126.615 ;
        RECT 62.740 126.445 63.190 126.905 ;
        RECT 64.055 126.735 64.455 127.585 ;
        RECT 64.855 127.295 65.125 127.755 ;
        RECT 65.295 127.125 65.580 127.585 ;
        RECT 62.635 126.115 63.190 126.445 ;
        RECT 63.360 126.175 64.455 126.735 ;
        RECT 62.740 126.005 63.190 126.115 ;
        RECT 61.210 125.755 61.925 125.925 ;
        RECT 61.210 125.205 61.540 125.585 ;
        RECT 61.755 125.375 61.925 125.755 ;
        RECT 62.185 125.375 62.570 125.945 ;
        RECT 62.740 125.835 63.865 126.005 ;
        RECT 62.740 125.205 63.065 125.665 ;
        RECT 63.585 125.375 63.865 125.835 ;
        RECT 64.055 125.375 64.455 126.175 ;
        RECT 64.625 126.905 65.580 127.125 ;
        RECT 65.980 127.125 66.265 127.585 ;
        RECT 66.435 127.295 66.705 127.755 ;
        RECT 65.980 126.905 66.935 127.125 ;
        RECT 64.625 126.005 64.835 126.905 ;
        RECT 65.005 126.175 65.695 126.735 ;
        RECT 65.865 126.175 66.555 126.735 ;
        RECT 66.725 126.005 66.935 126.905 ;
        RECT 64.625 125.835 65.580 126.005 ;
        RECT 64.855 125.205 65.125 125.665 ;
        RECT 65.295 125.375 65.580 125.835 ;
        RECT 65.980 125.835 66.935 126.005 ;
        RECT 67.105 126.735 67.505 127.585 ;
        RECT 67.695 127.125 67.975 127.585 ;
        RECT 68.495 127.295 68.820 127.755 ;
        RECT 67.695 126.905 68.820 127.125 ;
        RECT 67.105 126.175 68.200 126.735 ;
        RECT 68.370 126.445 68.820 126.905 ;
        RECT 68.990 126.615 69.375 127.585 ;
        RECT 65.980 125.375 66.265 125.835 ;
        RECT 66.435 125.205 66.705 125.665 ;
        RECT 67.105 125.375 67.505 126.175 ;
        RECT 68.370 126.115 68.925 126.445 ;
        RECT 68.370 126.005 68.820 126.115 ;
        RECT 67.695 125.835 68.820 126.005 ;
        RECT 69.095 125.945 69.375 126.615 ;
        RECT 70.005 126.590 70.295 127.755 ;
        RECT 70.470 126.805 70.735 127.575 ;
        RECT 70.905 127.035 71.235 127.755 ;
        RECT 71.425 127.215 71.685 127.575 ;
        RECT 71.855 127.385 72.185 127.755 ;
        RECT 72.355 127.215 72.615 127.575 ;
        RECT 71.425 126.985 72.615 127.215 ;
        RECT 73.185 126.805 73.475 127.575 ;
        RECT 74.695 127.085 74.865 127.585 ;
        RECT 75.035 127.255 75.365 127.755 ;
        RECT 74.695 126.915 75.360 127.085 ;
        RECT 67.695 125.375 67.975 125.835 ;
        RECT 68.495 125.205 68.820 125.665 ;
        RECT 68.990 125.375 69.375 125.945 ;
        RECT 70.005 125.205 70.295 125.930 ;
        RECT 70.470 125.385 70.805 126.805 ;
        RECT 70.980 126.625 73.475 126.805 ;
        RECT 70.980 125.935 71.205 126.625 ;
        RECT 71.405 126.115 71.685 126.445 ;
        RECT 71.865 126.115 72.440 126.445 ;
        RECT 72.620 126.115 73.055 126.445 ;
        RECT 73.235 126.115 73.505 126.445 ;
        RECT 74.610 126.095 74.960 126.745 ;
        RECT 70.980 125.745 73.465 125.935 ;
        RECT 75.130 125.925 75.360 126.915 ;
        RECT 70.985 125.205 71.730 125.575 ;
        RECT 72.295 125.385 72.550 125.745 ;
        RECT 72.730 125.205 73.060 125.575 ;
        RECT 73.240 125.385 73.465 125.745 ;
        RECT 74.695 125.755 75.360 125.925 ;
        RECT 74.695 125.465 74.865 125.755 ;
        RECT 75.035 125.205 75.365 125.585 ;
        RECT 75.535 125.465 75.720 127.585 ;
        RECT 75.960 127.295 76.225 127.755 ;
        RECT 76.395 127.160 76.645 127.585 ;
        RECT 76.855 127.310 77.960 127.480 ;
        RECT 76.340 127.030 76.645 127.160 ;
        RECT 75.890 125.835 76.170 126.785 ;
        RECT 76.340 125.925 76.510 127.030 ;
        RECT 76.680 126.245 76.920 126.840 ;
        RECT 77.090 126.775 77.620 127.140 ;
        RECT 77.090 126.075 77.260 126.775 ;
        RECT 77.790 126.695 77.960 127.310 ;
        RECT 78.130 126.955 78.300 127.755 ;
        RECT 78.470 127.255 78.720 127.585 ;
        RECT 78.945 127.285 79.830 127.455 ;
        RECT 77.790 126.605 78.300 126.695 ;
        RECT 76.340 125.795 76.565 125.925 ;
        RECT 76.735 125.855 77.260 126.075 ;
        RECT 77.430 126.435 78.300 126.605 ;
        RECT 75.975 125.205 76.225 125.665 ;
        RECT 76.395 125.655 76.565 125.795 ;
        RECT 77.430 125.655 77.600 126.435 ;
        RECT 78.130 126.365 78.300 126.435 ;
        RECT 77.810 126.185 78.010 126.215 ;
        RECT 78.470 126.185 78.640 127.255 ;
        RECT 78.810 126.365 79.000 127.085 ;
        RECT 77.810 125.885 78.640 126.185 ;
        RECT 79.170 126.155 79.490 127.115 ;
        RECT 76.395 125.485 76.730 125.655 ;
        RECT 76.925 125.485 77.600 125.655 ;
        RECT 77.920 125.205 78.290 125.705 ;
        RECT 78.470 125.655 78.640 125.885 ;
        RECT 79.025 125.825 79.490 126.155 ;
        RECT 79.660 126.445 79.830 127.285 ;
        RECT 80.010 127.255 80.325 127.755 ;
        RECT 80.555 127.025 80.895 127.585 ;
        RECT 80.000 126.650 80.895 127.025 ;
        RECT 81.065 126.745 81.235 127.755 ;
        RECT 80.705 126.445 80.895 126.650 ;
        RECT 81.405 126.695 81.735 127.540 ;
        RECT 81.405 126.615 81.795 126.695 ;
        RECT 81.580 126.565 81.795 126.615 ;
        RECT 79.660 126.115 80.535 126.445 ;
        RECT 80.705 126.115 81.455 126.445 ;
        RECT 79.660 125.655 79.830 126.115 ;
        RECT 80.705 125.945 80.905 126.115 ;
        RECT 81.625 125.985 81.795 126.565 ;
        RECT 81.965 126.665 83.175 127.755 ;
        RECT 81.965 126.125 82.485 126.665 ;
        RECT 81.570 125.945 81.795 125.985 ;
        RECT 82.655 125.955 83.175 126.495 ;
        RECT 78.470 125.485 78.875 125.655 ;
        RECT 79.045 125.485 79.830 125.655 ;
        RECT 80.105 125.205 80.315 125.735 ;
        RECT 80.575 125.420 80.905 125.945 ;
        RECT 81.415 125.860 81.795 125.945 ;
        RECT 81.075 125.205 81.245 125.815 ;
        RECT 81.415 125.425 81.745 125.860 ;
        RECT 81.965 125.205 83.175 125.955 ;
        RECT 5.520 125.035 83.260 125.205 ;
        RECT 5.605 124.285 6.815 125.035 ;
        RECT 6.985 124.285 8.195 125.035 ;
        RECT 8.370 124.780 8.705 124.825 ;
        RECT 8.365 124.315 8.705 124.780 ;
        RECT 8.875 124.655 9.205 125.035 ;
        RECT 5.605 123.745 6.125 124.285 ;
        RECT 6.295 123.575 6.815 124.115 ;
        RECT 6.985 123.745 7.505 124.285 ;
        RECT 7.675 123.575 8.195 124.115 ;
        RECT 5.605 122.485 6.815 123.575 ;
        RECT 6.985 122.485 8.195 123.575 ;
        RECT 8.365 123.625 8.535 124.315 ;
        RECT 8.705 123.795 8.965 124.125 ;
        RECT 8.365 122.655 8.625 123.625 ;
        RECT 8.795 123.245 8.965 123.795 ;
        RECT 9.135 123.425 9.475 124.455 ;
        RECT 9.665 124.015 9.935 124.700 ;
        RECT 9.665 123.845 9.975 124.015 ;
        RECT 9.665 123.425 9.935 123.845 ;
        RECT 10.160 123.425 10.440 124.700 ;
        RECT 10.640 124.535 10.870 124.865 ;
        RECT 11.115 124.655 11.445 125.035 ;
        RECT 10.640 123.245 10.810 124.535 ;
        RECT 11.615 124.465 11.790 124.865 ;
        RECT 12.045 124.490 17.390 125.035 ;
        RECT 11.160 124.295 11.790 124.465 ;
        RECT 11.160 124.125 11.330 124.295 ;
        RECT 10.980 123.795 11.330 124.125 ;
        RECT 8.795 123.075 10.810 123.245 ;
        RECT 11.160 123.275 11.330 123.795 ;
        RECT 11.510 123.445 11.875 124.125 ;
        RECT 13.630 123.660 13.970 124.490 ;
        RECT 17.655 124.485 17.825 124.865 ;
        RECT 18.040 124.655 18.370 125.035 ;
        RECT 17.655 124.315 18.370 124.485 ;
        RECT 11.160 123.105 11.790 123.275 ;
        RECT 8.820 122.485 9.150 122.895 ;
        RECT 9.350 122.655 9.520 123.075 ;
        RECT 9.735 122.485 10.405 122.895 ;
        RECT 10.640 122.655 10.810 123.075 ;
        RECT 11.115 122.485 11.445 122.925 ;
        RECT 11.615 122.655 11.790 123.105 ;
        RECT 15.450 122.920 15.800 124.170 ;
        RECT 17.565 123.765 17.920 124.135 ;
        RECT 18.200 124.125 18.370 124.315 ;
        RECT 18.540 124.290 18.795 124.865 ;
        RECT 18.200 123.795 18.455 124.125 ;
        RECT 18.200 123.585 18.370 123.795 ;
        RECT 17.655 123.415 18.370 123.585 ;
        RECT 18.625 123.560 18.795 124.290 ;
        RECT 18.970 124.195 19.230 125.035 ;
        RECT 19.405 124.405 19.745 124.865 ;
        RECT 19.915 124.575 20.085 125.035 ;
        RECT 20.715 124.600 21.075 124.865 ;
        RECT 20.720 124.595 21.075 124.600 ;
        RECT 20.725 124.585 21.075 124.595 ;
        RECT 20.730 124.580 21.075 124.585 ;
        RECT 20.735 124.570 21.075 124.580 ;
        RECT 21.315 124.575 21.485 125.035 ;
        RECT 20.740 124.565 21.075 124.570 ;
        RECT 20.750 124.555 21.075 124.565 ;
        RECT 20.760 124.545 21.075 124.555 ;
        RECT 20.255 124.405 20.585 124.485 ;
        RECT 19.405 124.215 20.585 124.405 ;
        RECT 20.775 124.405 21.075 124.545 ;
        RECT 20.775 124.215 21.485 124.405 ;
        RECT 19.405 123.845 19.735 124.045 ;
        RECT 20.045 124.025 20.375 124.045 ;
        RECT 19.925 123.845 20.375 124.025 ;
        RECT 12.045 122.485 17.390 122.920 ;
        RECT 17.655 122.655 17.825 123.415 ;
        RECT 18.040 122.485 18.370 123.245 ;
        RECT 18.540 122.655 18.795 123.560 ;
        RECT 18.970 122.485 19.230 123.635 ;
        RECT 19.405 123.505 19.635 123.845 ;
        RECT 19.415 122.485 19.745 123.205 ;
        RECT 19.925 122.730 20.140 123.845 ;
        RECT 20.545 123.815 21.015 124.045 ;
        RECT 21.200 123.645 21.485 124.215 ;
        RECT 21.655 124.090 21.995 124.865 ;
        RECT 20.335 123.430 21.485 123.645 ;
        RECT 20.335 122.655 20.665 123.430 ;
        RECT 20.835 122.485 21.545 123.260 ;
        RECT 21.715 122.655 21.995 124.090 ;
        RECT 22.165 124.575 22.725 124.865 ;
        RECT 22.895 124.575 23.145 125.035 ;
        RECT 22.165 123.205 22.415 124.575 ;
        RECT 23.765 124.405 24.095 124.765 ;
        RECT 22.705 124.215 24.095 124.405 ;
        RECT 24.465 124.265 26.135 125.035 ;
        RECT 22.705 124.125 22.875 124.215 ;
        RECT 22.585 123.795 22.875 124.125 ;
        RECT 23.045 123.795 23.385 124.045 ;
        RECT 23.605 123.795 24.280 124.045 ;
        RECT 22.705 123.545 22.875 123.795 ;
        RECT 22.705 123.375 23.645 123.545 ;
        RECT 24.015 123.435 24.280 123.795 ;
        RECT 24.465 123.745 25.215 124.265 ;
        RECT 26.315 124.225 26.585 125.035 ;
        RECT 26.755 124.225 27.085 124.865 ;
        RECT 27.255 124.225 27.495 125.035 ;
        RECT 28.165 124.565 28.460 125.035 ;
        RECT 28.630 124.395 28.890 124.840 ;
        RECT 29.060 124.565 29.320 125.035 ;
        RECT 29.490 124.395 29.745 124.840 ;
        RECT 29.915 124.565 30.215 125.035 ;
        RECT 27.705 124.225 30.735 124.395 ;
        RECT 31.365 124.310 31.655 125.035 ;
        RECT 31.845 124.225 32.085 125.035 ;
        RECT 32.255 124.225 32.585 124.865 ;
        RECT 32.755 124.225 33.025 125.035 ;
        RECT 34.215 124.485 34.385 124.775 ;
        RECT 34.555 124.655 34.885 125.035 ;
        RECT 34.215 124.315 34.880 124.485 ;
        RECT 25.385 123.575 26.135 124.095 ;
        RECT 26.305 123.795 26.655 124.045 ;
        RECT 26.825 123.625 26.995 124.225 ;
        RECT 27.165 123.795 27.515 124.045 ;
        RECT 27.705 123.660 27.875 124.225 ;
        RECT 28.045 123.830 30.260 124.055 ;
        RECT 30.435 123.660 30.735 124.225 ;
        RECT 31.825 123.795 32.175 124.045 ;
        RECT 22.165 122.655 22.625 123.205 ;
        RECT 22.815 122.485 23.145 123.205 ;
        RECT 23.345 122.825 23.645 123.375 ;
        RECT 23.815 122.485 24.095 123.155 ;
        RECT 24.465 122.485 26.135 123.575 ;
        RECT 26.315 122.485 26.645 123.625 ;
        RECT 26.825 123.455 27.505 123.625 ;
        RECT 27.705 123.490 30.735 123.660 ;
        RECT 27.175 122.670 27.505 123.455 ;
        RECT 27.685 122.485 28.030 123.320 ;
        RECT 28.205 122.685 28.460 123.490 ;
        RECT 28.630 122.485 28.890 123.320 ;
        RECT 29.065 122.685 29.320 123.490 ;
        RECT 29.490 122.485 29.750 123.320 ;
        RECT 29.920 122.685 30.180 123.490 ;
        RECT 30.350 122.485 30.735 123.320 ;
        RECT 31.365 122.485 31.655 123.650 ;
        RECT 32.345 123.625 32.515 124.225 ;
        RECT 32.685 123.795 33.035 124.045 ;
        RECT 31.835 123.455 32.515 123.625 ;
        RECT 31.835 122.670 32.165 123.455 ;
        RECT 32.695 122.485 33.025 123.625 ;
        RECT 34.130 123.495 34.480 124.145 ;
        RECT 34.650 123.325 34.880 124.315 ;
        RECT 34.215 123.155 34.880 123.325 ;
        RECT 34.215 122.655 34.385 123.155 ;
        RECT 34.555 122.485 34.885 122.985 ;
        RECT 35.055 122.655 35.240 124.775 ;
        RECT 35.495 124.575 35.745 125.035 ;
        RECT 35.915 124.585 36.250 124.755 ;
        RECT 36.445 124.585 37.120 124.755 ;
        RECT 35.915 124.445 36.085 124.585 ;
        RECT 35.410 123.455 35.690 124.405 ;
        RECT 35.860 124.315 36.085 124.445 ;
        RECT 35.860 123.210 36.030 124.315 ;
        RECT 36.255 124.165 36.780 124.385 ;
        RECT 36.200 123.400 36.440 123.995 ;
        RECT 36.610 123.465 36.780 124.165 ;
        RECT 36.950 123.805 37.120 124.585 ;
        RECT 37.440 124.535 37.810 125.035 ;
        RECT 37.990 124.585 38.395 124.755 ;
        RECT 38.565 124.585 39.350 124.755 ;
        RECT 37.990 124.355 38.160 124.585 ;
        RECT 37.330 124.055 38.160 124.355 ;
        RECT 38.545 124.085 39.010 124.415 ;
        RECT 37.330 124.025 37.530 124.055 ;
        RECT 37.650 123.805 37.820 123.875 ;
        RECT 36.950 123.635 37.820 123.805 ;
        RECT 37.310 123.545 37.820 123.635 ;
        RECT 35.860 123.080 36.165 123.210 ;
        RECT 36.610 123.100 37.140 123.465 ;
        RECT 35.480 122.485 35.745 122.945 ;
        RECT 35.915 122.655 36.165 123.080 ;
        RECT 37.310 122.930 37.480 123.545 ;
        RECT 36.375 122.760 37.480 122.930 ;
        RECT 37.650 122.485 37.820 123.285 ;
        RECT 37.990 122.985 38.160 124.055 ;
        RECT 38.330 123.155 38.520 123.875 ;
        RECT 38.690 123.125 39.010 124.085 ;
        RECT 39.180 124.125 39.350 124.585 ;
        RECT 39.625 124.505 39.835 125.035 ;
        RECT 40.095 124.295 40.425 124.820 ;
        RECT 40.595 124.425 40.765 125.035 ;
        RECT 40.935 124.380 41.265 124.815 ;
        RECT 40.935 124.295 41.315 124.380 ;
        RECT 40.225 124.125 40.425 124.295 ;
        RECT 41.090 124.255 41.315 124.295 ;
        RECT 39.180 123.795 40.055 124.125 ;
        RECT 40.225 123.795 40.975 124.125 ;
        RECT 37.990 122.655 38.240 122.985 ;
        RECT 39.180 122.955 39.350 123.795 ;
        RECT 40.225 123.590 40.415 123.795 ;
        RECT 41.145 123.675 41.315 124.255 ;
        RECT 41.100 123.625 41.315 123.675 ;
        RECT 39.520 123.215 40.415 123.590 ;
        RECT 40.925 123.545 41.315 123.625 ;
        RECT 41.490 124.295 41.745 124.865 ;
        RECT 41.915 124.635 42.245 125.035 ;
        RECT 42.670 124.500 43.200 124.865 ;
        RECT 42.670 124.465 42.845 124.500 ;
        RECT 41.915 124.295 42.845 124.465 ;
        RECT 43.390 124.355 43.665 124.865 ;
        RECT 41.490 123.625 41.660 124.295 ;
        RECT 41.915 124.125 42.085 124.295 ;
        RECT 41.830 123.795 42.085 124.125 ;
        RECT 42.310 123.795 42.505 124.125 ;
        RECT 38.465 122.785 39.350 122.955 ;
        RECT 39.530 122.485 39.845 122.985 ;
        RECT 40.075 122.655 40.415 123.215 ;
        RECT 40.585 122.485 40.755 123.495 ;
        RECT 40.925 122.700 41.255 123.545 ;
        RECT 41.490 122.655 41.825 123.625 ;
        RECT 41.995 122.485 42.165 123.625 ;
        RECT 42.335 122.825 42.505 123.795 ;
        RECT 42.675 123.165 42.845 124.295 ;
        RECT 43.015 123.505 43.185 124.305 ;
        RECT 43.385 124.185 43.665 124.355 ;
        RECT 43.390 123.705 43.665 124.185 ;
        RECT 43.835 123.505 44.025 124.865 ;
        RECT 44.205 124.500 44.715 125.035 ;
        RECT 44.935 124.225 45.180 124.830 ;
        RECT 45.625 124.535 45.925 124.865 ;
        RECT 46.095 124.555 46.370 125.035 ;
        RECT 44.225 124.055 45.455 124.225 ;
        RECT 43.015 123.335 44.025 123.505 ;
        RECT 44.195 123.490 44.945 123.680 ;
        RECT 42.675 122.995 43.800 123.165 ;
        RECT 44.195 122.825 44.365 123.490 ;
        RECT 45.115 123.245 45.455 124.055 ;
        RECT 42.335 122.655 44.365 122.825 ;
        RECT 44.535 122.485 44.705 123.245 ;
        RECT 44.940 122.835 45.455 123.245 ;
        RECT 45.625 123.625 45.795 124.535 ;
        RECT 46.550 124.385 46.845 124.775 ;
        RECT 47.015 124.555 47.270 125.035 ;
        RECT 47.445 124.385 47.705 124.775 ;
        RECT 47.875 124.555 48.155 125.035 ;
        RECT 45.965 123.795 46.315 124.365 ;
        RECT 46.550 124.215 48.200 124.385 ;
        RECT 46.485 123.875 47.625 124.045 ;
        RECT 46.485 123.625 46.655 123.875 ;
        RECT 47.795 123.705 48.200 124.215 ;
        RECT 48.385 124.285 49.595 125.035 ;
        RECT 49.855 124.485 50.025 124.775 ;
        RECT 50.195 124.655 50.525 125.035 ;
        RECT 49.855 124.315 50.520 124.485 ;
        RECT 48.385 123.745 48.905 124.285 ;
        RECT 45.625 123.455 46.655 123.625 ;
        RECT 47.445 123.535 48.200 123.705 ;
        RECT 49.075 123.575 49.595 124.115 ;
        RECT 45.625 122.655 45.935 123.455 ;
        RECT 47.445 123.285 47.705 123.535 ;
        RECT 46.105 122.485 46.415 123.285 ;
        RECT 46.585 123.115 47.705 123.285 ;
        RECT 46.585 122.655 46.845 123.115 ;
        RECT 47.015 122.485 47.270 122.945 ;
        RECT 47.445 122.655 47.705 123.115 ;
        RECT 47.875 122.485 48.160 123.355 ;
        RECT 48.385 122.485 49.595 123.575 ;
        RECT 49.770 123.495 50.120 124.145 ;
        RECT 50.290 123.325 50.520 124.315 ;
        RECT 49.855 123.155 50.520 123.325 ;
        RECT 49.855 122.655 50.025 123.155 ;
        RECT 50.195 122.485 50.525 122.985 ;
        RECT 50.695 122.655 50.880 124.775 ;
        RECT 51.135 124.575 51.385 125.035 ;
        RECT 51.555 124.585 51.890 124.755 ;
        RECT 52.085 124.585 52.760 124.755 ;
        RECT 51.555 124.445 51.725 124.585 ;
        RECT 51.050 123.455 51.330 124.405 ;
        RECT 51.500 124.315 51.725 124.445 ;
        RECT 51.500 123.210 51.670 124.315 ;
        RECT 51.895 124.165 52.420 124.385 ;
        RECT 51.840 123.400 52.080 123.995 ;
        RECT 52.250 123.465 52.420 124.165 ;
        RECT 52.590 123.805 52.760 124.585 ;
        RECT 53.080 124.535 53.450 125.035 ;
        RECT 53.630 124.585 54.035 124.755 ;
        RECT 54.205 124.585 54.990 124.755 ;
        RECT 53.630 124.355 53.800 124.585 ;
        RECT 52.970 124.055 53.800 124.355 ;
        RECT 54.185 124.085 54.650 124.415 ;
        RECT 52.970 124.025 53.170 124.055 ;
        RECT 53.290 123.805 53.460 123.875 ;
        RECT 52.590 123.635 53.460 123.805 ;
        RECT 52.950 123.545 53.460 123.635 ;
        RECT 51.500 123.080 51.805 123.210 ;
        RECT 52.250 123.100 52.780 123.465 ;
        RECT 51.120 122.485 51.385 122.945 ;
        RECT 51.555 122.655 51.805 123.080 ;
        RECT 52.950 122.930 53.120 123.545 ;
        RECT 52.015 122.760 53.120 122.930 ;
        RECT 53.290 122.485 53.460 123.285 ;
        RECT 53.630 122.985 53.800 124.055 ;
        RECT 53.970 123.155 54.160 123.875 ;
        RECT 54.330 123.125 54.650 124.085 ;
        RECT 54.820 124.125 54.990 124.585 ;
        RECT 55.265 124.505 55.475 125.035 ;
        RECT 55.735 124.295 56.065 124.820 ;
        RECT 56.235 124.425 56.405 125.035 ;
        RECT 56.575 124.380 56.905 124.815 ;
        RECT 56.575 124.295 56.955 124.380 ;
        RECT 57.125 124.310 57.415 125.035 ;
        RECT 57.675 124.485 57.845 124.775 ;
        RECT 58.015 124.655 58.345 125.035 ;
        RECT 57.675 124.315 58.340 124.485 ;
        RECT 55.865 124.125 56.065 124.295 ;
        RECT 56.730 124.255 56.955 124.295 ;
        RECT 54.820 123.795 55.695 124.125 ;
        RECT 55.865 123.795 56.615 124.125 ;
        RECT 53.630 122.655 53.880 122.985 ;
        RECT 54.820 122.955 54.990 123.795 ;
        RECT 55.865 123.590 56.055 123.795 ;
        RECT 56.785 123.675 56.955 124.255 ;
        RECT 56.740 123.625 56.955 123.675 ;
        RECT 55.160 123.215 56.055 123.590 ;
        RECT 56.565 123.545 56.955 123.625 ;
        RECT 54.105 122.785 54.990 122.955 ;
        RECT 55.170 122.485 55.485 122.985 ;
        RECT 55.715 122.655 56.055 123.215 ;
        RECT 56.225 122.485 56.395 123.495 ;
        RECT 56.565 122.700 56.895 123.545 ;
        RECT 57.125 122.485 57.415 123.650 ;
        RECT 57.590 123.495 57.940 124.145 ;
        RECT 58.110 123.325 58.340 124.315 ;
        RECT 57.675 123.155 58.340 123.325 ;
        RECT 57.675 122.655 57.845 123.155 ;
        RECT 58.015 122.485 58.345 122.985 ;
        RECT 58.515 122.655 58.700 124.775 ;
        RECT 58.955 124.575 59.205 125.035 ;
        RECT 59.375 124.585 59.710 124.755 ;
        RECT 59.905 124.585 60.580 124.755 ;
        RECT 59.375 124.445 59.545 124.585 ;
        RECT 58.870 123.455 59.150 124.405 ;
        RECT 59.320 124.315 59.545 124.445 ;
        RECT 59.320 123.210 59.490 124.315 ;
        RECT 59.715 124.165 60.240 124.385 ;
        RECT 59.660 123.400 59.900 123.995 ;
        RECT 60.070 123.465 60.240 124.165 ;
        RECT 60.410 123.805 60.580 124.585 ;
        RECT 60.900 124.535 61.270 125.035 ;
        RECT 61.450 124.585 61.855 124.755 ;
        RECT 62.025 124.585 62.810 124.755 ;
        RECT 61.450 124.355 61.620 124.585 ;
        RECT 60.790 124.055 61.620 124.355 ;
        RECT 62.005 124.085 62.470 124.415 ;
        RECT 60.790 124.025 60.990 124.055 ;
        RECT 61.110 123.805 61.280 123.875 ;
        RECT 60.410 123.635 61.280 123.805 ;
        RECT 60.770 123.545 61.280 123.635 ;
        RECT 59.320 123.080 59.625 123.210 ;
        RECT 60.070 123.100 60.600 123.465 ;
        RECT 58.940 122.485 59.205 122.945 ;
        RECT 59.375 122.655 59.625 123.080 ;
        RECT 60.770 122.930 60.940 123.545 ;
        RECT 59.835 122.760 60.940 122.930 ;
        RECT 61.110 122.485 61.280 123.285 ;
        RECT 61.450 122.985 61.620 124.055 ;
        RECT 61.790 123.155 61.980 123.875 ;
        RECT 62.150 123.125 62.470 124.085 ;
        RECT 62.640 124.125 62.810 124.585 ;
        RECT 63.085 124.505 63.295 125.035 ;
        RECT 63.555 124.295 63.885 124.820 ;
        RECT 64.055 124.425 64.225 125.035 ;
        RECT 64.395 124.380 64.725 124.815 ;
        RECT 64.395 124.295 64.775 124.380 ;
        RECT 63.685 124.125 63.885 124.295 ;
        RECT 64.550 124.255 64.775 124.295 ;
        RECT 62.640 123.795 63.515 124.125 ;
        RECT 63.685 123.795 64.435 124.125 ;
        RECT 61.450 122.655 61.700 122.985 ;
        RECT 62.640 122.955 62.810 123.795 ;
        RECT 63.685 123.590 63.875 123.795 ;
        RECT 64.605 123.675 64.775 124.255 ;
        RECT 64.560 123.625 64.775 123.675 ;
        RECT 62.980 123.215 63.875 123.590 ;
        RECT 64.385 123.545 64.775 123.625 ;
        RECT 64.950 124.295 65.205 124.865 ;
        RECT 65.375 124.635 65.705 125.035 ;
        RECT 66.130 124.500 66.660 124.865 ;
        RECT 66.850 124.695 67.125 124.865 ;
        RECT 66.845 124.525 67.125 124.695 ;
        RECT 66.130 124.465 66.305 124.500 ;
        RECT 65.375 124.295 66.305 124.465 ;
        RECT 64.950 123.625 65.120 124.295 ;
        RECT 65.375 124.125 65.545 124.295 ;
        RECT 65.290 123.795 65.545 124.125 ;
        RECT 65.770 123.795 65.965 124.125 ;
        RECT 61.925 122.785 62.810 122.955 ;
        RECT 62.990 122.485 63.305 122.985 ;
        RECT 63.535 122.655 63.875 123.215 ;
        RECT 64.045 122.485 64.215 123.495 ;
        RECT 64.385 122.700 64.715 123.545 ;
        RECT 64.950 122.655 65.285 123.625 ;
        RECT 65.455 122.485 65.625 123.625 ;
        RECT 65.795 122.825 65.965 123.795 ;
        RECT 66.135 123.165 66.305 124.295 ;
        RECT 66.475 123.505 66.645 124.305 ;
        RECT 66.850 123.705 67.125 124.525 ;
        RECT 67.295 123.505 67.485 124.865 ;
        RECT 67.665 124.500 68.175 125.035 ;
        RECT 68.395 124.225 68.640 124.830 ;
        RECT 67.685 124.055 68.915 124.225 ;
        RECT 69.090 124.195 69.350 125.035 ;
        RECT 69.525 124.290 69.780 124.865 ;
        RECT 69.950 124.655 70.280 125.035 ;
        RECT 70.495 124.485 70.665 124.865 ;
        RECT 69.950 124.315 70.665 124.485 ;
        RECT 66.475 123.335 67.485 123.505 ;
        RECT 67.655 123.490 68.405 123.680 ;
        RECT 66.135 122.995 67.260 123.165 ;
        RECT 67.655 122.825 67.825 123.490 ;
        RECT 68.575 123.245 68.915 124.055 ;
        RECT 65.795 122.655 67.825 122.825 ;
        RECT 67.995 122.485 68.165 123.245 ;
        RECT 68.400 122.835 68.915 123.245 ;
        RECT 69.090 122.485 69.350 123.635 ;
        RECT 69.525 123.560 69.695 124.290 ;
        RECT 69.950 124.125 70.120 124.315 ;
        RECT 71.130 124.255 71.630 124.865 ;
        RECT 69.865 123.795 70.120 124.125 ;
        RECT 69.950 123.585 70.120 123.795 ;
        RECT 70.400 123.765 70.755 124.135 ;
        RECT 70.925 123.795 71.275 124.045 ;
        RECT 71.460 123.625 71.630 124.255 ;
        RECT 72.260 124.385 72.590 124.865 ;
        RECT 72.760 124.575 72.985 125.035 ;
        RECT 73.155 124.385 73.485 124.865 ;
        RECT 72.260 124.215 73.485 124.385 ;
        RECT 73.675 124.235 73.925 125.035 ;
        RECT 74.095 124.235 74.435 124.865 ;
        RECT 74.695 124.485 74.865 124.775 ;
        RECT 75.035 124.655 75.365 125.035 ;
        RECT 74.695 124.315 75.360 124.485 ;
        RECT 71.800 123.845 72.130 124.045 ;
        RECT 72.300 123.845 72.630 124.045 ;
        RECT 72.800 123.845 73.220 124.045 ;
        RECT 73.395 123.875 74.090 124.045 ;
        RECT 73.395 123.625 73.565 123.875 ;
        RECT 74.260 123.625 74.435 124.235 ;
        RECT 69.525 122.655 69.780 123.560 ;
        RECT 69.950 123.415 70.665 123.585 ;
        RECT 69.950 122.485 70.280 123.245 ;
        RECT 70.495 122.655 70.665 123.415 ;
        RECT 71.130 123.455 73.565 123.625 ;
        RECT 71.130 122.655 71.460 123.455 ;
        RECT 71.630 122.485 71.960 123.285 ;
        RECT 72.260 122.655 72.590 123.455 ;
        RECT 73.235 122.485 73.485 123.285 ;
        RECT 73.755 122.485 73.925 123.625 ;
        RECT 74.095 122.655 74.435 123.625 ;
        RECT 74.610 123.495 74.960 124.145 ;
        RECT 75.130 123.325 75.360 124.315 ;
        RECT 74.695 123.155 75.360 123.325 ;
        RECT 74.695 122.655 74.865 123.155 ;
        RECT 75.035 122.485 75.365 122.985 ;
        RECT 75.535 122.655 75.720 124.775 ;
        RECT 75.975 124.575 76.225 125.035 ;
        RECT 76.395 124.585 76.730 124.755 ;
        RECT 76.925 124.585 77.600 124.755 ;
        RECT 76.395 124.445 76.565 124.585 ;
        RECT 75.890 123.455 76.170 124.405 ;
        RECT 76.340 124.315 76.565 124.445 ;
        RECT 76.340 123.210 76.510 124.315 ;
        RECT 76.735 124.165 77.260 124.385 ;
        RECT 76.680 123.400 76.920 123.995 ;
        RECT 77.090 123.465 77.260 124.165 ;
        RECT 77.430 123.805 77.600 124.585 ;
        RECT 77.920 124.535 78.290 125.035 ;
        RECT 78.470 124.585 78.875 124.755 ;
        RECT 79.045 124.585 79.830 124.755 ;
        RECT 78.470 124.355 78.640 124.585 ;
        RECT 77.810 124.055 78.640 124.355 ;
        RECT 79.025 124.085 79.490 124.415 ;
        RECT 77.810 124.025 78.010 124.055 ;
        RECT 78.130 123.805 78.300 123.875 ;
        RECT 77.430 123.635 78.300 123.805 ;
        RECT 77.790 123.545 78.300 123.635 ;
        RECT 76.340 123.080 76.645 123.210 ;
        RECT 77.090 123.100 77.620 123.465 ;
        RECT 75.960 122.485 76.225 122.945 ;
        RECT 76.395 122.655 76.645 123.080 ;
        RECT 77.790 122.930 77.960 123.545 ;
        RECT 76.855 122.760 77.960 122.930 ;
        RECT 78.130 122.485 78.300 123.285 ;
        RECT 78.470 122.985 78.640 124.055 ;
        RECT 78.810 123.155 79.000 123.875 ;
        RECT 79.170 123.125 79.490 124.085 ;
        RECT 79.660 124.125 79.830 124.585 ;
        RECT 80.105 124.505 80.315 125.035 ;
        RECT 80.575 124.295 80.905 124.820 ;
        RECT 81.075 124.425 81.245 125.035 ;
        RECT 81.415 124.380 81.745 124.815 ;
        RECT 81.415 124.295 81.795 124.380 ;
        RECT 80.705 124.125 80.905 124.295 ;
        RECT 81.570 124.255 81.795 124.295 ;
        RECT 81.965 124.285 83.175 125.035 ;
        RECT 79.660 123.795 80.535 124.125 ;
        RECT 80.705 123.795 81.455 124.125 ;
        RECT 78.470 122.655 78.720 122.985 ;
        RECT 79.660 122.955 79.830 123.795 ;
        RECT 80.705 123.590 80.895 123.795 ;
        RECT 81.625 123.675 81.795 124.255 ;
        RECT 81.580 123.625 81.795 123.675 ;
        RECT 80.000 123.215 80.895 123.590 ;
        RECT 81.405 123.545 81.795 123.625 ;
        RECT 81.965 123.575 82.485 124.115 ;
        RECT 82.655 123.745 83.175 124.285 ;
        RECT 78.945 122.785 79.830 122.955 ;
        RECT 80.010 122.485 80.325 122.985 ;
        RECT 80.555 122.655 80.895 123.215 ;
        RECT 81.065 122.485 81.235 123.495 ;
        RECT 81.405 122.700 81.735 123.545 ;
        RECT 81.965 122.485 83.175 123.575 ;
        RECT 5.520 122.315 83.260 122.485 ;
        RECT 5.605 121.225 6.815 122.315 ;
        RECT 7.535 121.645 7.705 122.145 ;
        RECT 7.875 121.815 8.205 122.315 ;
        RECT 7.535 121.475 8.200 121.645 ;
        RECT 5.605 120.515 6.125 121.055 ;
        RECT 6.295 120.685 6.815 121.225 ;
        RECT 7.450 120.655 7.800 121.305 ;
        RECT 5.605 119.765 6.815 120.515 ;
        RECT 7.970 120.485 8.200 121.475 ;
        RECT 7.535 120.315 8.200 120.485 ;
        RECT 7.535 120.025 7.705 120.315 ;
        RECT 7.875 119.765 8.205 120.145 ;
        RECT 8.375 120.025 8.560 122.145 ;
        RECT 8.800 121.855 9.065 122.315 ;
        RECT 9.235 121.720 9.485 122.145 ;
        RECT 9.695 121.870 10.800 122.040 ;
        RECT 9.180 121.590 9.485 121.720 ;
        RECT 8.730 120.395 9.010 121.345 ;
        RECT 9.180 120.485 9.350 121.590 ;
        RECT 9.520 120.805 9.760 121.400 ;
        RECT 9.930 121.335 10.460 121.700 ;
        RECT 9.930 120.635 10.100 121.335 ;
        RECT 10.630 121.255 10.800 121.870 ;
        RECT 10.970 121.515 11.140 122.315 ;
        RECT 11.310 121.815 11.560 122.145 ;
        RECT 11.785 121.845 12.670 122.015 ;
        RECT 10.630 121.165 11.140 121.255 ;
        RECT 9.180 120.355 9.405 120.485 ;
        RECT 9.575 120.415 10.100 120.635 ;
        RECT 10.270 120.995 11.140 121.165 ;
        RECT 8.815 119.765 9.065 120.225 ;
        RECT 9.235 120.215 9.405 120.355 ;
        RECT 10.270 120.215 10.440 120.995 ;
        RECT 10.970 120.925 11.140 120.995 ;
        RECT 10.650 120.745 10.850 120.775 ;
        RECT 11.310 120.745 11.480 121.815 ;
        RECT 11.650 120.925 11.840 121.645 ;
        RECT 10.650 120.445 11.480 120.745 ;
        RECT 12.010 120.715 12.330 121.675 ;
        RECT 9.235 120.045 9.570 120.215 ;
        RECT 9.765 120.045 10.440 120.215 ;
        RECT 10.760 119.765 11.130 120.265 ;
        RECT 11.310 120.215 11.480 120.445 ;
        RECT 11.865 120.385 12.330 120.715 ;
        RECT 12.500 121.005 12.670 121.845 ;
        RECT 12.850 121.815 13.165 122.315 ;
        RECT 13.395 121.585 13.735 122.145 ;
        RECT 12.840 121.210 13.735 121.585 ;
        RECT 13.905 121.305 14.075 122.315 ;
        RECT 13.545 121.005 13.735 121.210 ;
        RECT 14.245 121.255 14.575 122.100 ;
        RECT 14.815 121.345 15.145 122.130 ;
        RECT 14.245 121.175 14.635 121.255 ;
        RECT 14.815 121.175 15.495 121.345 ;
        RECT 15.675 121.175 16.005 122.315 ;
        RECT 16.685 121.855 16.900 122.315 ;
        RECT 17.070 121.685 17.400 122.145 ;
        RECT 16.230 121.515 17.400 121.685 ;
        RECT 17.570 121.515 17.820 122.315 ;
        RECT 14.420 121.125 14.635 121.175 ;
        RECT 12.500 120.675 13.375 121.005 ;
        RECT 13.545 120.675 14.295 121.005 ;
        RECT 12.500 120.215 12.670 120.675 ;
        RECT 13.545 120.505 13.745 120.675 ;
        RECT 14.465 120.545 14.635 121.125 ;
        RECT 14.805 120.755 15.155 121.005 ;
        RECT 15.325 120.575 15.495 121.175 ;
        RECT 15.665 120.755 16.015 121.005 ;
        RECT 14.410 120.505 14.635 120.545 ;
        RECT 11.310 120.045 11.715 120.215 ;
        RECT 11.885 120.045 12.670 120.215 ;
        RECT 12.945 119.765 13.155 120.295 ;
        RECT 13.415 119.980 13.745 120.505 ;
        RECT 14.255 120.420 14.635 120.505 ;
        RECT 13.915 119.765 14.085 120.375 ;
        RECT 14.255 119.985 14.585 120.420 ;
        RECT 14.825 119.765 15.065 120.575 ;
        RECT 15.235 119.935 15.565 120.575 ;
        RECT 15.735 119.765 16.005 120.575 ;
        RECT 16.230 120.225 16.600 121.515 ;
        RECT 18.030 121.345 18.310 121.505 ;
        RECT 16.975 121.175 18.310 121.345 ;
        RECT 16.975 121.005 17.145 121.175 ;
        RECT 18.485 121.150 18.775 122.315 ;
        RECT 18.945 121.175 19.225 122.315 ;
        RECT 19.395 121.165 19.725 122.145 ;
        RECT 19.895 121.175 20.155 122.315 ;
        RECT 20.325 121.345 20.635 122.145 ;
        RECT 20.805 121.515 21.115 122.315 ;
        RECT 21.285 121.685 21.545 122.145 ;
        RECT 21.715 121.855 21.970 122.315 ;
        RECT 22.145 121.685 22.405 122.145 ;
        RECT 21.285 121.515 22.405 121.685 ;
        RECT 20.325 121.175 21.355 121.345 ;
        RECT 16.770 120.755 17.145 121.005 ;
        RECT 17.315 120.755 17.790 120.995 ;
        RECT 17.960 120.755 18.310 120.995 ;
        RECT 16.975 120.585 17.145 120.755 ;
        RECT 18.955 120.735 19.290 121.005 ;
        RECT 16.975 120.415 18.310 120.585 ;
        RECT 19.460 120.565 19.630 121.165 ;
        RECT 19.800 120.755 20.135 121.005 ;
        RECT 16.230 119.935 16.980 120.225 ;
        RECT 17.490 119.765 17.820 120.225 ;
        RECT 18.040 120.205 18.310 120.415 ;
        RECT 18.485 119.765 18.775 120.490 ;
        RECT 18.945 119.765 19.255 120.565 ;
        RECT 19.460 119.935 20.155 120.565 ;
        RECT 20.325 120.265 20.495 121.175 ;
        RECT 20.665 120.435 21.015 121.005 ;
        RECT 21.185 120.925 21.355 121.175 ;
        RECT 22.145 121.265 22.405 121.515 ;
        RECT 22.575 121.445 22.860 122.315 ;
        RECT 23.170 121.695 23.345 122.145 ;
        RECT 23.515 121.875 23.845 122.315 ;
        RECT 24.150 121.725 24.320 122.145 ;
        RECT 24.555 121.905 25.225 122.315 ;
        RECT 25.440 121.725 25.610 122.145 ;
        RECT 25.810 121.905 26.140 122.315 ;
        RECT 23.170 121.525 23.800 121.695 ;
        RECT 22.145 121.095 22.900 121.265 ;
        RECT 21.185 120.755 22.325 120.925 ;
        RECT 22.495 120.585 22.900 121.095 ;
        RECT 23.085 120.675 23.450 121.355 ;
        RECT 23.630 121.005 23.800 121.525 ;
        RECT 24.150 121.555 26.165 121.725 ;
        RECT 23.630 120.675 23.980 121.005 ;
        RECT 21.250 120.415 22.900 120.585 ;
        RECT 23.630 120.505 23.800 120.675 ;
        RECT 20.325 119.935 20.625 120.265 ;
        RECT 20.795 119.765 21.070 120.245 ;
        RECT 21.250 120.025 21.545 120.415 ;
        RECT 21.715 119.765 21.970 120.245 ;
        RECT 22.145 120.025 22.405 120.415 ;
        RECT 23.170 120.335 23.800 120.505 ;
        RECT 22.575 119.765 22.855 120.245 ;
        RECT 23.170 119.935 23.345 120.335 ;
        RECT 24.150 120.265 24.320 121.555 ;
        RECT 23.515 119.765 23.845 120.145 ;
        RECT 24.090 119.935 24.320 120.265 ;
        RECT 24.520 120.100 24.800 121.375 ;
        RECT 25.025 121.295 25.295 121.375 ;
        RECT 24.985 121.125 25.295 121.295 ;
        RECT 25.025 120.100 25.295 121.125 ;
        RECT 25.485 120.345 25.825 121.375 ;
        RECT 25.995 121.005 26.165 121.555 ;
        RECT 26.335 121.175 26.595 122.145 ;
        RECT 26.850 121.695 27.025 122.145 ;
        RECT 27.195 121.875 27.525 122.315 ;
        RECT 27.830 121.725 28.000 122.145 ;
        RECT 28.235 121.905 28.905 122.315 ;
        RECT 29.120 121.725 29.290 122.145 ;
        RECT 29.490 121.905 29.820 122.315 ;
        RECT 26.850 121.525 27.480 121.695 ;
        RECT 25.995 120.675 26.255 121.005 ;
        RECT 26.425 120.485 26.595 121.175 ;
        RECT 26.765 120.675 27.130 121.355 ;
        RECT 27.310 121.005 27.480 121.525 ;
        RECT 27.830 121.555 29.845 121.725 ;
        RECT 27.310 120.675 27.660 121.005 ;
        RECT 27.310 120.505 27.480 120.675 ;
        RECT 25.755 119.765 26.085 120.145 ;
        RECT 26.255 120.020 26.595 120.485 ;
        RECT 26.850 120.335 27.480 120.505 ;
        RECT 26.255 119.975 26.590 120.020 ;
        RECT 26.850 119.935 27.025 120.335 ;
        RECT 27.830 120.265 28.000 121.555 ;
        RECT 27.195 119.765 27.525 120.145 ;
        RECT 27.770 119.935 28.000 120.265 ;
        RECT 28.200 120.100 28.480 121.375 ;
        RECT 28.705 120.275 28.975 121.375 ;
        RECT 29.165 120.345 29.505 121.375 ;
        RECT 29.675 121.005 29.845 121.555 ;
        RECT 30.015 121.175 30.275 122.145 ;
        RECT 30.450 121.935 30.785 122.315 ;
        RECT 29.675 120.675 29.935 121.005 ;
        RECT 30.105 120.485 30.275 121.175 ;
        RECT 28.665 120.105 28.975 120.275 ;
        RECT 28.705 120.100 28.975 120.105 ;
        RECT 29.435 119.765 29.765 120.145 ;
        RECT 29.935 120.020 30.275 120.485 ;
        RECT 30.445 120.445 30.685 121.755 ;
        RECT 30.955 121.345 31.205 122.145 ;
        RECT 31.425 121.595 31.755 122.315 ;
        RECT 31.940 121.345 32.190 122.145 ;
        RECT 32.655 121.515 32.985 122.315 ;
        RECT 33.155 121.885 33.495 122.145 ;
        RECT 30.855 121.175 33.045 121.345 ;
        RECT 30.855 120.265 31.025 121.175 ;
        RECT 32.730 121.005 33.045 121.175 ;
        RECT 29.935 119.975 30.270 120.020 ;
        RECT 30.530 119.935 31.025 120.265 ;
        RECT 31.245 120.040 31.595 121.005 ;
        RECT 31.775 120.035 32.075 121.005 ;
        RECT 32.255 120.035 32.535 121.005 ;
        RECT 32.730 120.755 33.060 121.005 ;
        RECT 32.715 119.765 32.985 120.565 ;
        RECT 33.235 120.485 33.495 121.885 ;
        RECT 33.665 121.805 33.965 122.315 ;
        RECT 34.135 121.635 34.465 122.145 ;
        RECT 34.635 121.805 35.265 122.315 ;
        RECT 35.845 121.805 36.225 121.975 ;
        RECT 36.395 121.805 36.695 122.315 ;
        RECT 36.055 121.635 36.225 121.805 ;
        RECT 33.155 119.975 33.495 120.485 ;
        RECT 33.665 121.465 35.885 121.635 ;
        RECT 33.665 120.505 33.835 121.465 ;
        RECT 34.005 121.125 35.545 121.295 ;
        RECT 34.005 120.675 34.250 121.125 ;
        RECT 34.510 120.755 35.205 120.955 ;
        RECT 35.375 120.925 35.545 121.125 ;
        RECT 35.715 121.265 35.885 121.465 ;
        RECT 36.055 121.435 36.715 121.635 ;
        RECT 35.715 121.095 36.375 121.265 ;
        RECT 35.375 120.755 35.975 120.925 ;
        RECT 36.205 120.675 36.375 121.095 ;
        RECT 33.665 119.960 34.130 120.505 ;
        RECT 34.635 119.765 34.805 120.585 ;
        RECT 34.975 120.505 35.885 120.585 ;
        RECT 36.545 120.505 36.715 121.435 ;
        RECT 36.945 121.255 37.275 122.100 ;
        RECT 37.445 121.305 37.615 122.315 ;
        RECT 37.785 121.585 38.125 122.145 ;
        RECT 38.355 121.815 38.670 122.315 ;
        RECT 38.850 121.845 39.735 122.015 ;
        RECT 34.975 120.415 36.225 120.505 ;
        RECT 34.975 119.935 35.305 120.415 ;
        RECT 35.715 120.335 36.225 120.415 ;
        RECT 35.475 119.765 35.825 120.155 ;
        RECT 35.995 119.935 36.225 120.335 ;
        RECT 36.395 120.025 36.715 120.505 ;
        RECT 36.885 121.175 37.275 121.255 ;
        RECT 37.785 121.210 38.680 121.585 ;
        RECT 36.885 121.125 37.100 121.175 ;
        RECT 36.885 120.545 37.055 121.125 ;
        RECT 37.785 121.005 37.975 121.210 ;
        RECT 38.850 121.005 39.020 121.845 ;
        RECT 39.960 121.815 40.210 122.145 ;
        RECT 37.225 120.675 37.975 121.005 ;
        RECT 38.145 120.675 39.020 121.005 ;
        RECT 36.885 120.505 37.110 120.545 ;
        RECT 37.775 120.505 37.975 120.675 ;
        RECT 36.885 120.420 37.265 120.505 ;
        RECT 36.935 119.985 37.265 120.420 ;
        RECT 37.435 119.765 37.605 120.375 ;
        RECT 37.775 119.980 38.105 120.505 ;
        RECT 38.365 119.765 38.575 120.295 ;
        RECT 38.850 120.215 39.020 120.675 ;
        RECT 39.190 120.715 39.510 121.675 ;
        RECT 39.680 120.925 39.870 121.645 ;
        RECT 40.040 120.745 40.210 121.815 ;
        RECT 40.380 121.515 40.550 122.315 ;
        RECT 40.720 121.870 41.825 122.040 ;
        RECT 40.720 121.255 40.890 121.870 ;
        RECT 42.035 121.720 42.285 122.145 ;
        RECT 42.455 121.855 42.720 122.315 ;
        RECT 41.060 121.335 41.590 121.700 ;
        RECT 42.035 121.590 42.340 121.720 ;
        RECT 40.380 121.165 40.890 121.255 ;
        RECT 40.380 120.995 41.250 121.165 ;
        RECT 40.380 120.925 40.550 120.995 ;
        RECT 40.670 120.745 40.870 120.775 ;
        RECT 39.190 120.385 39.655 120.715 ;
        RECT 40.040 120.445 40.870 120.745 ;
        RECT 40.040 120.215 40.210 120.445 ;
        RECT 38.850 120.045 39.635 120.215 ;
        RECT 39.805 120.045 40.210 120.215 ;
        RECT 40.390 119.765 40.760 120.265 ;
        RECT 41.080 120.215 41.250 120.995 ;
        RECT 41.420 120.635 41.590 121.335 ;
        RECT 41.760 120.805 42.000 121.400 ;
        RECT 41.420 120.415 41.945 120.635 ;
        RECT 42.170 120.485 42.340 121.590 ;
        RECT 42.115 120.355 42.340 120.485 ;
        RECT 42.510 120.395 42.790 121.345 ;
        RECT 42.115 120.215 42.285 120.355 ;
        RECT 41.080 120.045 41.755 120.215 ;
        RECT 41.950 120.045 42.285 120.215 ;
        RECT 42.455 119.765 42.705 120.225 ;
        RECT 42.960 120.025 43.145 122.145 ;
        RECT 43.315 121.815 43.645 122.315 ;
        RECT 43.815 121.645 43.985 122.145 ;
        RECT 43.320 121.475 43.985 121.645 ;
        RECT 43.320 120.485 43.550 121.475 ;
        RECT 43.720 120.655 44.070 121.305 ;
        RECT 44.245 121.150 44.535 122.315 ;
        RECT 44.705 121.225 47.295 122.315 ;
        RECT 44.705 120.535 45.915 121.055 ;
        RECT 46.085 120.705 47.295 121.225 ;
        RECT 47.985 121.175 48.195 122.315 ;
        RECT 48.365 121.165 48.695 122.145 ;
        RECT 48.865 121.175 49.095 122.315 ;
        RECT 49.305 121.175 49.585 122.315 ;
        RECT 49.755 121.165 50.085 122.145 ;
        RECT 50.255 121.175 50.515 122.315 ;
        RECT 50.690 121.175 51.025 122.145 ;
        RECT 51.195 121.175 51.365 122.315 ;
        RECT 51.535 121.975 53.565 122.145 ;
        RECT 43.320 120.315 43.985 120.485 ;
        RECT 43.315 119.765 43.645 120.145 ;
        RECT 43.815 120.025 43.985 120.315 ;
        RECT 44.245 119.765 44.535 120.490 ;
        RECT 44.705 119.765 47.295 120.535 ;
        RECT 47.985 119.765 48.195 120.585 ;
        RECT 48.365 120.565 48.615 121.165 ;
        RECT 48.785 120.755 49.115 121.005 ;
        RECT 49.315 120.735 49.650 121.005 ;
        RECT 49.820 120.615 49.990 121.165 ;
        RECT 50.160 120.755 50.495 121.005 ;
        RECT 48.365 119.935 48.695 120.565 ;
        RECT 48.865 119.765 49.095 120.585 ;
        RECT 49.820 120.565 49.995 120.615 ;
        RECT 49.305 119.765 49.615 120.565 ;
        RECT 49.820 119.935 50.515 120.565 ;
        RECT 50.690 120.505 50.860 121.175 ;
        RECT 51.535 121.005 51.705 121.975 ;
        RECT 51.030 120.675 51.285 121.005 ;
        RECT 51.510 120.675 51.705 121.005 ;
        RECT 51.875 121.635 53.000 121.805 ;
        RECT 51.115 120.505 51.285 120.675 ;
        RECT 51.875 120.505 52.045 121.635 ;
        RECT 50.690 119.935 50.945 120.505 ;
        RECT 51.115 120.335 52.045 120.505 ;
        RECT 52.215 121.295 53.225 121.465 ;
        RECT 52.215 120.495 52.385 121.295 ;
        RECT 51.870 120.300 52.045 120.335 ;
        RECT 51.115 119.765 51.445 120.165 ;
        RECT 51.870 119.935 52.400 120.300 ;
        RECT 52.590 120.275 52.865 121.095 ;
        RECT 52.585 120.105 52.865 120.275 ;
        RECT 52.590 119.935 52.865 120.105 ;
        RECT 53.035 119.935 53.225 121.295 ;
        RECT 53.395 121.310 53.565 121.975 ;
        RECT 53.735 121.555 53.905 122.315 ;
        RECT 54.140 121.555 54.655 121.965 ;
        RECT 53.395 121.120 54.145 121.310 ;
        RECT 54.315 120.745 54.655 121.555 ;
        RECT 54.830 121.165 55.090 122.315 ;
        RECT 55.265 121.240 55.520 122.145 ;
        RECT 55.690 121.555 56.020 122.315 ;
        RECT 56.235 121.385 56.405 122.145 ;
        RECT 53.425 120.575 54.655 120.745 ;
        RECT 53.405 119.765 53.915 120.300 ;
        RECT 54.135 119.970 54.380 120.575 ;
        RECT 54.830 119.765 55.090 120.605 ;
        RECT 55.265 120.510 55.435 121.240 ;
        RECT 55.690 121.215 56.405 121.385 ;
        RECT 55.690 121.005 55.860 121.215 ;
        RECT 56.665 121.175 56.925 122.315 ;
        RECT 57.095 121.165 57.425 122.145 ;
        RECT 57.595 121.175 57.875 122.315 ;
        RECT 58.045 121.175 58.305 122.315 ;
        RECT 58.475 121.165 58.805 122.145 ;
        RECT 58.975 121.175 59.255 122.315 ;
        RECT 59.945 121.255 60.275 122.100 ;
        RECT 60.445 121.305 60.615 122.315 ;
        RECT 60.785 121.585 61.125 122.145 ;
        RECT 61.355 121.815 61.670 122.315 ;
        RECT 61.850 121.845 62.735 122.015 ;
        RECT 59.885 121.175 60.275 121.255 ;
        RECT 60.785 121.210 61.680 121.585 ;
        RECT 55.605 120.675 55.860 121.005 ;
        RECT 55.265 119.935 55.520 120.510 ;
        RECT 55.690 120.485 55.860 120.675 ;
        RECT 56.140 120.665 56.495 121.035 ;
        RECT 56.685 120.755 57.020 121.005 ;
        RECT 57.190 120.565 57.360 121.165 ;
        RECT 57.530 120.735 57.865 121.005 ;
        RECT 58.065 120.755 58.400 121.005 ;
        RECT 58.570 120.565 58.740 121.165 ;
        RECT 59.885 121.125 60.100 121.175 ;
        RECT 58.910 120.735 59.245 121.005 ;
        RECT 55.690 120.315 56.405 120.485 ;
        RECT 55.690 119.765 56.020 120.145 ;
        RECT 56.235 119.935 56.405 120.315 ;
        RECT 56.665 119.935 57.360 120.565 ;
        RECT 57.565 119.765 57.875 120.565 ;
        RECT 58.045 119.935 58.740 120.565 ;
        RECT 58.945 119.765 59.255 120.565 ;
        RECT 59.885 120.545 60.055 121.125 ;
        RECT 60.785 121.005 60.975 121.210 ;
        RECT 61.850 121.005 62.020 121.845 ;
        RECT 62.960 121.815 63.210 122.145 ;
        RECT 60.225 120.675 60.975 121.005 ;
        RECT 61.145 120.675 62.020 121.005 ;
        RECT 59.885 120.505 60.110 120.545 ;
        RECT 60.775 120.505 60.975 120.675 ;
        RECT 59.885 120.420 60.265 120.505 ;
        RECT 59.935 119.985 60.265 120.420 ;
        RECT 60.435 119.765 60.605 120.375 ;
        RECT 60.775 119.980 61.105 120.505 ;
        RECT 61.365 119.765 61.575 120.295 ;
        RECT 61.850 120.215 62.020 120.675 ;
        RECT 62.190 120.715 62.510 121.675 ;
        RECT 62.680 120.925 62.870 121.645 ;
        RECT 63.040 120.745 63.210 121.815 ;
        RECT 63.380 121.515 63.550 122.315 ;
        RECT 63.720 121.870 64.825 122.040 ;
        RECT 63.720 121.255 63.890 121.870 ;
        RECT 65.035 121.720 65.285 122.145 ;
        RECT 65.455 121.855 65.720 122.315 ;
        RECT 64.060 121.335 64.590 121.700 ;
        RECT 65.035 121.590 65.340 121.720 ;
        RECT 63.380 121.165 63.890 121.255 ;
        RECT 63.380 120.995 64.250 121.165 ;
        RECT 63.380 120.925 63.550 120.995 ;
        RECT 63.670 120.745 63.870 120.775 ;
        RECT 62.190 120.385 62.655 120.715 ;
        RECT 63.040 120.445 63.870 120.745 ;
        RECT 63.040 120.215 63.210 120.445 ;
        RECT 61.850 120.045 62.635 120.215 ;
        RECT 62.805 120.045 63.210 120.215 ;
        RECT 63.390 119.765 63.760 120.265 ;
        RECT 64.080 120.215 64.250 120.995 ;
        RECT 64.420 120.635 64.590 121.335 ;
        RECT 64.760 120.805 65.000 121.400 ;
        RECT 64.420 120.415 64.945 120.635 ;
        RECT 65.170 120.485 65.340 121.590 ;
        RECT 65.115 120.355 65.340 120.485 ;
        RECT 65.510 120.395 65.790 121.345 ;
        RECT 65.115 120.215 65.285 120.355 ;
        RECT 64.080 120.045 64.755 120.215 ;
        RECT 64.950 120.045 65.285 120.215 ;
        RECT 65.455 119.765 65.705 120.225 ;
        RECT 65.960 120.025 66.145 122.145 ;
        RECT 66.315 121.815 66.645 122.315 ;
        RECT 66.815 121.645 66.985 122.145 ;
        RECT 66.320 121.475 66.985 121.645 ;
        RECT 66.320 120.485 66.550 121.475 ;
        RECT 67.890 121.345 68.280 121.520 ;
        RECT 68.765 121.515 69.095 122.315 ;
        RECT 69.265 121.525 69.800 122.145 ;
        RECT 66.720 120.655 67.070 121.305 ;
        RECT 67.890 121.175 69.315 121.345 ;
        RECT 66.320 120.315 66.985 120.485 ;
        RECT 67.765 120.445 68.120 121.005 ;
        RECT 66.315 119.765 66.645 120.145 ;
        RECT 66.815 120.025 66.985 120.315 ;
        RECT 68.290 120.275 68.460 121.175 ;
        RECT 68.630 120.445 68.895 121.005 ;
        RECT 69.145 120.675 69.315 121.175 ;
        RECT 69.485 120.505 69.800 121.525 ;
        RECT 70.005 121.150 70.295 122.315 ;
        RECT 70.465 121.175 70.805 122.145 ;
        RECT 70.975 121.175 71.145 122.315 ;
        RECT 71.415 121.515 71.665 122.315 ;
        RECT 72.310 121.345 72.640 122.145 ;
        RECT 72.940 121.515 73.270 122.315 ;
        RECT 73.440 121.345 73.770 122.145 ;
        RECT 71.335 121.175 73.770 121.345 ;
        RECT 74.350 121.345 74.680 122.145 ;
        RECT 74.850 121.515 75.180 122.315 ;
        RECT 75.480 121.345 75.810 122.145 ;
        RECT 76.455 121.515 76.705 122.315 ;
        RECT 74.350 121.175 76.785 121.345 ;
        RECT 76.975 121.175 77.145 122.315 ;
        RECT 77.315 121.175 77.655 122.145 ;
        RECT 67.870 119.765 68.110 120.275 ;
        RECT 68.290 119.945 68.570 120.275 ;
        RECT 68.800 119.765 69.015 120.275 ;
        RECT 69.185 119.935 69.800 120.505 ;
        RECT 70.465 120.565 70.640 121.175 ;
        RECT 71.335 120.925 71.505 121.175 ;
        RECT 70.810 120.755 71.505 120.925 ;
        RECT 71.680 120.755 72.100 120.955 ;
        RECT 72.270 120.755 72.600 120.955 ;
        RECT 72.770 120.755 73.100 120.955 ;
        RECT 70.005 119.765 70.295 120.490 ;
        RECT 70.465 119.935 70.805 120.565 ;
        RECT 70.975 119.765 71.225 120.565 ;
        RECT 71.415 120.415 72.640 120.585 ;
        RECT 71.415 119.935 71.745 120.415 ;
        RECT 71.915 119.765 72.140 120.225 ;
        RECT 72.310 119.935 72.640 120.415 ;
        RECT 73.270 120.545 73.440 121.175 ;
        RECT 73.625 120.755 73.975 121.005 ;
        RECT 74.145 120.755 74.495 121.005 ;
        RECT 74.680 120.545 74.850 121.175 ;
        RECT 75.020 120.755 75.350 120.955 ;
        RECT 75.520 120.755 75.850 120.955 ;
        RECT 76.020 120.755 76.440 120.955 ;
        RECT 76.615 120.925 76.785 121.175 ;
        RECT 76.615 120.755 77.310 120.925 ;
        RECT 73.270 119.935 73.770 120.545 ;
        RECT 74.350 119.935 74.850 120.545 ;
        RECT 75.480 120.415 76.705 120.585 ;
        RECT 77.480 120.565 77.655 121.175 ;
        RECT 75.480 119.935 75.810 120.415 ;
        RECT 75.980 119.765 76.205 120.225 ;
        RECT 76.375 119.935 76.705 120.415 ;
        RECT 76.895 119.765 77.145 120.565 ;
        RECT 77.315 119.935 77.655 120.565 ;
        RECT 77.825 121.465 78.085 122.145 ;
        RECT 78.255 121.535 78.505 122.315 ;
        RECT 78.755 121.765 79.005 122.145 ;
        RECT 79.175 121.935 79.530 122.315 ;
        RECT 80.535 121.925 80.870 122.145 ;
        RECT 80.135 121.765 80.365 121.805 ;
        RECT 78.755 121.565 80.365 121.765 ;
        RECT 78.755 121.555 79.590 121.565 ;
        RECT 80.180 121.475 80.365 121.565 ;
        RECT 77.825 120.265 77.995 121.465 ;
        RECT 79.695 121.365 80.025 121.395 ;
        RECT 78.225 121.305 80.025 121.365 ;
        RECT 80.615 121.305 80.870 121.925 ;
        RECT 78.165 121.195 80.870 121.305 ;
        RECT 78.165 121.160 78.365 121.195 ;
        RECT 78.165 120.585 78.335 121.160 ;
        RECT 79.695 121.135 80.870 121.195 ;
        RECT 81.965 121.225 83.175 122.315 ;
        RECT 78.565 120.720 78.975 121.025 ;
        RECT 79.145 120.755 79.475 120.965 ;
        RECT 78.165 120.465 78.435 120.585 ;
        RECT 78.165 120.420 79.010 120.465 ;
        RECT 78.255 120.295 79.010 120.420 ;
        RECT 79.265 120.355 79.475 120.755 ;
        RECT 79.720 120.755 80.195 120.965 ;
        RECT 80.385 120.755 80.875 120.955 ;
        RECT 79.720 120.355 79.940 120.755 ;
        RECT 81.965 120.685 82.485 121.225 ;
        RECT 77.825 119.935 78.085 120.265 ;
        RECT 78.840 120.145 79.010 120.295 ;
        RECT 78.255 119.765 78.585 120.125 ;
        RECT 78.840 119.935 80.140 120.145 ;
        RECT 80.415 119.765 80.870 120.530 ;
        RECT 82.655 120.515 83.175 121.055 ;
        RECT 81.965 119.765 83.175 120.515 ;
        RECT 5.520 119.595 83.260 119.765 ;
        RECT 5.605 118.845 6.815 119.595 ;
        RECT 7.075 119.045 7.245 119.335 ;
        RECT 7.415 119.215 7.745 119.595 ;
        RECT 7.075 118.875 7.740 119.045 ;
        RECT 5.605 118.305 6.125 118.845 ;
        RECT 6.295 118.135 6.815 118.675 ;
        RECT 5.605 117.045 6.815 118.135 ;
        RECT 6.990 118.055 7.340 118.705 ;
        RECT 7.510 117.885 7.740 118.875 ;
        RECT 7.075 117.715 7.740 117.885 ;
        RECT 7.075 117.215 7.245 117.715 ;
        RECT 7.415 117.045 7.745 117.545 ;
        RECT 7.915 117.215 8.100 119.335 ;
        RECT 8.355 119.135 8.605 119.595 ;
        RECT 8.775 119.145 9.110 119.315 ;
        RECT 9.305 119.145 9.980 119.315 ;
        RECT 8.775 119.005 8.945 119.145 ;
        RECT 8.270 118.015 8.550 118.965 ;
        RECT 8.720 118.875 8.945 119.005 ;
        RECT 8.720 117.770 8.890 118.875 ;
        RECT 9.115 118.725 9.640 118.945 ;
        RECT 9.060 117.960 9.300 118.555 ;
        RECT 9.470 118.025 9.640 118.725 ;
        RECT 9.810 118.365 9.980 119.145 ;
        RECT 10.300 119.095 10.670 119.595 ;
        RECT 10.850 119.145 11.255 119.315 ;
        RECT 11.425 119.145 12.210 119.315 ;
        RECT 10.850 118.915 11.020 119.145 ;
        RECT 10.190 118.615 11.020 118.915 ;
        RECT 11.405 118.645 11.870 118.975 ;
        RECT 10.190 118.585 10.390 118.615 ;
        RECT 10.510 118.365 10.680 118.435 ;
        RECT 9.810 118.195 10.680 118.365 ;
        RECT 10.170 118.105 10.680 118.195 ;
        RECT 8.720 117.640 9.025 117.770 ;
        RECT 9.470 117.660 10.000 118.025 ;
        RECT 8.340 117.045 8.605 117.505 ;
        RECT 8.775 117.215 9.025 117.640 ;
        RECT 10.170 117.490 10.340 118.105 ;
        RECT 9.235 117.320 10.340 117.490 ;
        RECT 10.510 117.045 10.680 117.845 ;
        RECT 10.850 117.545 11.020 118.615 ;
        RECT 11.190 117.715 11.380 118.435 ;
        RECT 11.550 117.685 11.870 118.645 ;
        RECT 12.040 118.685 12.210 119.145 ;
        RECT 12.485 119.065 12.695 119.595 ;
        RECT 12.955 118.855 13.285 119.380 ;
        RECT 13.455 118.985 13.625 119.595 ;
        RECT 13.795 118.940 14.125 119.375 ;
        RECT 13.795 118.855 14.175 118.940 ;
        RECT 13.085 118.685 13.285 118.855 ;
        RECT 13.950 118.815 14.175 118.855 ;
        RECT 12.040 118.355 12.915 118.685 ;
        RECT 13.085 118.355 13.835 118.685 ;
        RECT 10.850 117.215 11.100 117.545 ;
        RECT 12.040 117.515 12.210 118.355 ;
        RECT 13.085 118.150 13.275 118.355 ;
        RECT 14.005 118.235 14.175 118.815 ;
        RECT 14.365 118.785 14.605 119.595 ;
        RECT 14.775 118.785 15.105 119.425 ;
        RECT 15.275 118.785 15.545 119.595 ;
        RECT 15.930 118.815 16.430 119.425 ;
        RECT 14.345 118.355 14.695 118.605 ;
        RECT 13.960 118.185 14.175 118.235 ;
        RECT 14.865 118.185 15.035 118.785 ;
        RECT 15.205 118.355 15.555 118.605 ;
        RECT 15.725 118.355 16.075 118.605 ;
        RECT 16.260 118.185 16.430 118.815 ;
        RECT 17.060 118.945 17.390 119.425 ;
        RECT 17.560 119.135 17.785 119.595 ;
        RECT 17.955 118.945 18.285 119.425 ;
        RECT 17.060 118.775 18.285 118.945 ;
        RECT 18.475 118.795 18.725 119.595 ;
        RECT 18.895 118.795 19.235 119.425 ;
        RECT 16.600 118.405 16.930 118.605 ;
        RECT 17.100 118.405 17.430 118.605 ;
        RECT 17.600 118.405 18.020 118.605 ;
        RECT 18.195 118.435 18.890 118.605 ;
        RECT 18.195 118.185 18.365 118.435 ;
        RECT 19.060 118.185 19.235 118.795 ;
        RECT 12.380 117.775 13.275 118.150 ;
        RECT 13.785 118.105 14.175 118.185 ;
        RECT 11.325 117.345 12.210 117.515 ;
        RECT 12.390 117.045 12.705 117.545 ;
        RECT 12.935 117.215 13.275 117.775 ;
        RECT 13.445 117.045 13.615 118.055 ;
        RECT 13.785 117.260 14.115 118.105 ;
        RECT 14.355 118.015 15.035 118.185 ;
        RECT 14.355 117.230 14.685 118.015 ;
        RECT 15.215 117.045 15.545 118.185 ;
        RECT 15.930 118.015 18.365 118.185 ;
        RECT 15.930 117.215 16.260 118.015 ;
        RECT 16.430 117.045 16.760 117.845 ;
        RECT 17.060 117.215 17.390 118.015 ;
        RECT 18.035 117.045 18.285 117.845 ;
        RECT 18.555 117.045 18.725 118.185 ;
        RECT 18.895 117.215 19.235 118.185 ;
        RECT 19.865 117.215 20.145 119.315 ;
        RECT 20.375 119.135 20.545 119.595 ;
        RECT 20.815 119.205 22.065 119.385 ;
        RECT 21.200 118.965 21.565 119.035 ;
        RECT 20.315 118.785 21.565 118.965 ;
        RECT 21.735 118.985 22.065 119.205 ;
        RECT 22.235 119.155 22.405 119.595 ;
        RECT 22.575 118.985 22.915 119.400 ;
        RECT 21.735 118.815 22.915 118.985 ;
        RECT 24.095 119.045 24.265 119.335 ;
        RECT 24.435 119.215 24.765 119.595 ;
        RECT 24.095 118.875 24.760 119.045 ;
        RECT 20.315 118.185 20.590 118.785 ;
        RECT 20.760 118.355 21.115 118.605 ;
        RECT 21.310 118.575 21.775 118.605 ;
        RECT 21.305 118.405 21.775 118.575 ;
        RECT 21.310 118.355 21.775 118.405 ;
        RECT 21.945 118.355 22.275 118.605 ;
        RECT 22.450 118.405 22.915 118.605 ;
        RECT 22.095 118.235 22.275 118.355 ;
        RECT 20.315 117.975 21.925 118.185 ;
        RECT 22.095 118.065 22.425 118.235 ;
        RECT 21.515 117.875 21.925 117.975 ;
        RECT 20.335 117.045 21.120 117.805 ;
        RECT 21.515 117.215 21.900 117.875 ;
        RECT 22.225 117.275 22.425 118.065 ;
        RECT 22.595 117.045 22.915 118.225 ;
        RECT 24.010 118.055 24.360 118.705 ;
        RECT 24.530 117.885 24.760 118.875 ;
        RECT 24.095 117.715 24.760 117.885 ;
        RECT 24.095 117.215 24.265 117.715 ;
        RECT 24.435 117.045 24.765 117.545 ;
        RECT 24.935 117.215 25.120 119.335 ;
        RECT 25.375 119.135 25.625 119.595 ;
        RECT 25.795 119.145 26.130 119.315 ;
        RECT 26.325 119.145 27.000 119.315 ;
        RECT 25.795 119.005 25.965 119.145 ;
        RECT 25.290 118.015 25.570 118.965 ;
        RECT 25.740 118.875 25.965 119.005 ;
        RECT 25.740 117.770 25.910 118.875 ;
        RECT 26.135 118.725 26.660 118.945 ;
        RECT 26.080 117.960 26.320 118.555 ;
        RECT 26.490 118.025 26.660 118.725 ;
        RECT 26.830 118.365 27.000 119.145 ;
        RECT 27.320 119.095 27.690 119.595 ;
        RECT 27.870 119.145 28.275 119.315 ;
        RECT 28.445 119.145 29.230 119.315 ;
        RECT 27.870 118.915 28.040 119.145 ;
        RECT 27.210 118.615 28.040 118.915 ;
        RECT 28.425 118.645 28.890 118.975 ;
        RECT 27.210 118.585 27.410 118.615 ;
        RECT 27.530 118.365 27.700 118.435 ;
        RECT 26.830 118.195 27.700 118.365 ;
        RECT 27.190 118.105 27.700 118.195 ;
        RECT 25.740 117.640 26.045 117.770 ;
        RECT 26.490 117.660 27.020 118.025 ;
        RECT 25.360 117.045 25.625 117.505 ;
        RECT 25.795 117.215 26.045 117.640 ;
        RECT 27.190 117.490 27.360 118.105 ;
        RECT 26.255 117.320 27.360 117.490 ;
        RECT 27.530 117.045 27.700 117.845 ;
        RECT 27.870 117.545 28.040 118.615 ;
        RECT 28.210 117.715 28.400 118.435 ;
        RECT 28.570 117.685 28.890 118.645 ;
        RECT 29.060 118.685 29.230 119.145 ;
        RECT 29.505 119.065 29.715 119.595 ;
        RECT 29.975 118.855 30.305 119.380 ;
        RECT 30.475 118.985 30.645 119.595 ;
        RECT 30.815 118.940 31.145 119.375 ;
        RECT 30.815 118.855 31.195 118.940 ;
        RECT 31.365 118.870 31.655 119.595 ;
        RECT 31.825 119.050 37.170 119.595 ;
        RECT 37.345 119.050 42.690 119.595 ;
        RECT 30.105 118.685 30.305 118.855 ;
        RECT 30.970 118.815 31.195 118.855 ;
        RECT 29.060 118.355 29.935 118.685 ;
        RECT 30.105 118.355 30.855 118.685 ;
        RECT 27.870 117.215 28.120 117.545 ;
        RECT 29.060 117.515 29.230 118.355 ;
        RECT 30.105 118.150 30.295 118.355 ;
        RECT 31.025 118.235 31.195 118.815 ;
        RECT 30.980 118.185 31.195 118.235 ;
        RECT 33.410 118.220 33.750 119.050 ;
        RECT 29.400 117.775 30.295 118.150 ;
        RECT 30.805 118.105 31.195 118.185 ;
        RECT 28.345 117.345 29.230 117.515 ;
        RECT 29.410 117.045 29.725 117.545 ;
        RECT 29.955 117.215 30.295 117.775 ;
        RECT 30.465 117.045 30.635 118.055 ;
        RECT 30.805 117.260 31.135 118.105 ;
        RECT 31.365 117.045 31.655 118.210 ;
        RECT 35.230 117.480 35.580 118.730 ;
        RECT 38.930 118.220 39.270 119.050 ;
        RECT 42.865 118.825 45.455 119.595 ;
        RECT 46.175 119.045 46.345 119.335 ;
        RECT 46.515 119.215 46.845 119.595 ;
        RECT 46.175 118.875 46.840 119.045 ;
        RECT 40.750 117.480 41.100 118.730 ;
        RECT 42.865 118.305 44.075 118.825 ;
        RECT 44.245 118.135 45.455 118.655 ;
        RECT 31.825 117.045 37.170 117.480 ;
        RECT 37.345 117.045 42.690 117.480 ;
        RECT 42.865 117.045 45.455 118.135 ;
        RECT 46.090 118.055 46.440 118.705 ;
        RECT 46.610 117.885 46.840 118.875 ;
        RECT 46.175 117.715 46.840 117.885 ;
        RECT 46.175 117.215 46.345 117.715 ;
        RECT 46.515 117.045 46.845 117.545 ;
        RECT 47.015 117.215 47.200 119.335 ;
        RECT 47.455 119.135 47.705 119.595 ;
        RECT 47.875 119.145 48.210 119.315 ;
        RECT 48.405 119.145 49.080 119.315 ;
        RECT 47.875 119.005 48.045 119.145 ;
        RECT 47.370 118.015 47.650 118.965 ;
        RECT 47.820 118.875 48.045 119.005 ;
        RECT 47.820 117.770 47.990 118.875 ;
        RECT 48.215 118.725 48.740 118.945 ;
        RECT 48.160 117.960 48.400 118.555 ;
        RECT 48.570 118.025 48.740 118.725 ;
        RECT 48.910 118.365 49.080 119.145 ;
        RECT 49.400 119.095 49.770 119.595 ;
        RECT 49.950 119.145 50.355 119.315 ;
        RECT 50.525 119.145 51.310 119.315 ;
        RECT 49.950 118.915 50.120 119.145 ;
        RECT 49.290 118.615 50.120 118.915 ;
        RECT 50.505 118.645 50.970 118.975 ;
        RECT 49.290 118.585 49.490 118.615 ;
        RECT 49.610 118.365 49.780 118.435 ;
        RECT 48.910 118.195 49.780 118.365 ;
        RECT 49.270 118.105 49.780 118.195 ;
        RECT 47.820 117.640 48.125 117.770 ;
        RECT 48.570 117.660 49.100 118.025 ;
        RECT 47.440 117.045 47.705 117.505 ;
        RECT 47.875 117.215 48.125 117.640 ;
        RECT 49.270 117.490 49.440 118.105 ;
        RECT 48.335 117.320 49.440 117.490 ;
        RECT 49.610 117.045 49.780 117.845 ;
        RECT 49.950 117.545 50.120 118.615 ;
        RECT 50.290 117.715 50.480 118.435 ;
        RECT 50.650 117.685 50.970 118.645 ;
        RECT 51.140 118.685 51.310 119.145 ;
        RECT 51.585 119.065 51.795 119.595 ;
        RECT 52.055 118.855 52.385 119.380 ;
        RECT 52.555 118.985 52.725 119.595 ;
        RECT 52.895 118.940 53.225 119.375 ;
        RECT 53.560 118.965 53.845 119.425 ;
        RECT 54.015 119.135 54.285 119.595 ;
        RECT 52.895 118.855 53.275 118.940 ;
        RECT 52.185 118.685 52.385 118.855 ;
        RECT 53.050 118.815 53.275 118.855 ;
        RECT 51.140 118.355 52.015 118.685 ;
        RECT 52.185 118.355 52.935 118.685 ;
        RECT 49.950 117.215 50.200 117.545 ;
        RECT 51.140 117.515 51.310 118.355 ;
        RECT 52.185 118.150 52.375 118.355 ;
        RECT 53.105 118.235 53.275 118.815 ;
        RECT 53.560 118.795 54.515 118.965 ;
        RECT 53.060 118.185 53.275 118.235 ;
        RECT 51.480 117.775 52.375 118.150 ;
        RECT 52.885 118.105 53.275 118.185 ;
        RECT 50.425 117.345 51.310 117.515 ;
        RECT 51.490 117.045 51.805 117.545 ;
        RECT 52.035 117.215 52.375 117.775 ;
        RECT 52.545 117.045 52.715 118.055 ;
        RECT 52.885 117.260 53.215 118.105 ;
        RECT 53.445 118.065 54.135 118.625 ;
        RECT 54.305 117.895 54.515 118.795 ;
        RECT 53.560 117.675 54.515 117.895 ;
        RECT 54.685 118.625 55.085 119.425 ;
        RECT 55.275 118.965 55.555 119.425 ;
        RECT 56.075 119.135 56.400 119.595 ;
        RECT 55.275 118.795 56.400 118.965 ;
        RECT 56.570 118.855 56.955 119.425 ;
        RECT 57.125 118.870 57.415 119.595 ;
        RECT 57.585 119.095 57.845 119.425 ;
        RECT 58.015 119.235 58.345 119.595 ;
        RECT 58.600 119.215 59.900 119.425 ;
        RECT 55.950 118.685 56.400 118.795 ;
        RECT 54.685 118.065 55.780 118.625 ;
        RECT 55.950 118.355 56.505 118.685 ;
        RECT 53.560 117.215 53.845 117.675 ;
        RECT 54.015 117.045 54.285 117.505 ;
        RECT 54.685 117.215 55.085 118.065 ;
        RECT 55.950 117.895 56.400 118.355 ;
        RECT 56.675 118.185 56.955 118.855 ;
        RECT 55.275 117.675 56.400 117.895 ;
        RECT 55.275 117.215 55.555 117.675 ;
        RECT 56.075 117.045 56.400 117.505 ;
        RECT 56.570 117.215 56.955 118.185 ;
        RECT 57.125 117.045 57.415 118.210 ;
        RECT 57.585 117.895 57.755 119.095 ;
        RECT 58.600 119.065 58.770 119.215 ;
        RECT 58.015 118.940 58.770 119.065 ;
        RECT 57.925 118.895 58.770 118.940 ;
        RECT 57.925 118.775 58.195 118.895 ;
        RECT 57.925 118.200 58.095 118.775 ;
        RECT 58.325 118.335 58.735 118.640 ;
        RECT 59.025 118.605 59.235 119.005 ;
        RECT 58.905 118.395 59.235 118.605 ;
        RECT 59.480 118.605 59.700 119.005 ;
        RECT 60.175 118.830 60.630 119.595 ;
        RECT 60.810 118.755 61.070 119.595 ;
        RECT 61.245 118.850 61.500 119.425 ;
        RECT 61.670 119.215 62.000 119.595 ;
        RECT 62.215 119.045 62.385 119.425 ;
        RECT 61.670 118.875 62.385 119.045 ;
        RECT 59.480 118.395 59.955 118.605 ;
        RECT 60.145 118.405 60.635 118.605 ;
        RECT 57.925 118.165 58.125 118.200 ;
        RECT 59.455 118.165 60.630 118.225 ;
        RECT 57.925 118.055 60.630 118.165 ;
        RECT 57.985 117.995 59.785 118.055 ;
        RECT 59.455 117.965 59.785 117.995 ;
        RECT 57.585 117.215 57.845 117.895 ;
        RECT 58.015 117.045 58.265 117.825 ;
        RECT 58.515 117.795 59.350 117.805 ;
        RECT 59.940 117.795 60.125 117.885 ;
        RECT 58.515 117.595 60.125 117.795 ;
        RECT 58.515 117.215 58.765 117.595 ;
        RECT 59.895 117.555 60.125 117.595 ;
        RECT 60.375 117.435 60.630 118.055 ;
        RECT 58.935 117.045 59.290 117.425 ;
        RECT 60.295 117.215 60.630 117.435 ;
        RECT 60.810 117.045 61.070 118.195 ;
        RECT 61.245 118.120 61.415 118.850 ;
        RECT 61.670 118.685 61.840 118.875 ;
        RECT 62.650 118.830 63.105 119.595 ;
        RECT 63.380 119.215 64.680 119.425 ;
        RECT 64.935 119.235 65.265 119.595 ;
        RECT 64.510 119.065 64.680 119.215 ;
        RECT 65.435 119.095 65.695 119.425 ;
        RECT 65.465 119.085 65.695 119.095 ;
        RECT 61.585 118.355 61.840 118.685 ;
        RECT 61.670 118.145 61.840 118.355 ;
        RECT 62.120 118.325 62.475 118.695 ;
        RECT 63.580 118.605 63.800 119.005 ;
        RECT 62.645 118.405 63.135 118.605 ;
        RECT 63.325 118.395 63.800 118.605 ;
        RECT 64.045 118.605 64.255 119.005 ;
        RECT 64.510 118.940 65.265 119.065 ;
        RECT 64.510 118.895 65.355 118.940 ;
        RECT 65.085 118.775 65.355 118.895 ;
        RECT 64.045 118.395 64.375 118.605 ;
        RECT 64.545 118.335 64.955 118.640 ;
        RECT 62.650 118.165 63.825 118.225 ;
        RECT 65.185 118.200 65.355 118.775 ;
        RECT 65.155 118.165 65.355 118.200 ;
        RECT 61.245 117.215 61.500 118.120 ;
        RECT 61.670 117.975 62.385 118.145 ;
        RECT 61.670 117.045 62.000 117.805 ;
        RECT 62.215 117.215 62.385 117.975 ;
        RECT 62.650 118.055 65.355 118.165 ;
        RECT 62.650 117.435 62.905 118.055 ;
        RECT 63.495 117.995 65.295 118.055 ;
        RECT 63.495 117.965 63.825 117.995 ;
        RECT 65.525 117.895 65.695 119.085 ;
        RECT 65.955 119.045 66.125 119.335 ;
        RECT 66.295 119.215 66.625 119.595 ;
        RECT 65.955 118.875 66.620 119.045 ;
        RECT 65.870 118.055 66.220 118.705 ;
        RECT 63.155 117.795 63.340 117.885 ;
        RECT 63.930 117.795 64.765 117.805 ;
        RECT 63.155 117.595 64.765 117.795 ;
        RECT 63.155 117.555 63.385 117.595 ;
        RECT 62.650 117.215 62.985 117.435 ;
        RECT 63.990 117.045 64.345 117.425 ;
        RECT 64.515 117.215 64.765 117.595 ;
        RECT 65.015 117.045 65.265 117.825 ;
        RECT 65.435 117.215 65.695 117.895 ;
        RECT 66.390 117.885 66.620 118.875 ;
        RECT 65.955 117.715 66.620 117.885 ;
        RECT 65.955 117.215 66.125 117.715 ;
        RECT 66.295 117.045 66.625 117.545 ;
        RECT 66.795 117.215 66.980 119.335 ;
        RECT 67.235 119.135 67.485 119.595 ;
        RECT 67.655 119.145 67.990 119.315 ;
        RECT 68.185 119.145 68.860 119.315 ;
        RECT 67.655 119.005 67.825 119.145 ;
        RECT 67.150 118.015 67.430 118.965 ;
        RECT 67.600 118.875 67.825 119.005 ;
        RECT 67.600 117.770 67.770 118.875 ;
        RECT 67.995 118.725 68.520 118.945 ;
        RECT 67.940 117.960 68.180 118.555 ;
        RECT 68.350 118.025 68.520 118.725 ;
        RECT 68.690 118.365 68.860 119.145 ;
        RECT 69.180 119.095 69.550 119.595 ;
        RECT 69.730 119.145 70.135 119.315 ;
        RECT 70.305 119.145 71.090 119.315 ;
        RECT 69.730 118.915 69.900 119.145 ;
        RECT 69.070 118.615 69.900 118.915 ;
        RECT 70.285 118.645 70.750 118.975 ;
        RECT 69.070 118.585 69.270 118.615 ;
        RECT 69.390 118.365 69.560 118.435 ;
        RECT 68.690 118.195 69.560 118.365 ;
        RECT 69.050 118.105 69.560 118.195 ;
        RECT 67.600 117.640 67.905 117.770 ;
        RECT 68.350 117.660 68.880 118.025 ;
        RECT 67.220 117.045 67.485 117.505 ;
        RECT 67.655 117.215 67.905 117.640 ;
        RECT 69.050 117.490 69.220 118.105 ;
        RECT 68.115 117.320 69.220 117.490 ;
        RECT 69.390 117.045 69.560 117.845 ;
        RECT 69.730 117.545 69.900 118.615 ;
        RECT 70.070 117.715 70.260 118.435 ;
        RECT 70.430 117.685 70.750 118.645 ;
        RECT 70.920 118.685 71.090 119.145 ;
        RECT 71.365 119.065 71.575 119.595 ;
        RECT 71.835 118.855 72.165 119.380 ;
        RECT 72.335 118.985 72.505 119.595 ;
        RECT 72.675 118.940 73.005 119.375 ;
        RECT 73.390 119.085 73.630 119.595 ;
        RECT 73.810 119.085 74.090 119.415 ;
        RECT 74.320 119.085 74.535 119.595 ;
        RECT 72.675 118.855 73.055 118.940 ;
        RECT 71.965 118.685 72.165 118.855 ;
        RECT 72.830 118.815 73.055 118.855 ;
        RECT 70.920 118.355 71.795 118.685 ;
        RECT 71.965 118.355 72.715 118.685 ;
        RECT 69.730 117.215 69.980 117.545 ;
        RECT 70.920 117.515 71.090 118.355 ;
        RECT 71.965 118.150 72.155 118.355 ;
        RECT 72.885 118.235 73.055 118.815 ;
        RECT 73.285 118.355 73.640 118.915 ;
        RECT 72.840 118.185 73.055 118.235 ;
        RECT 73.810 118.185 73.980 119.085 ;
        RECT 74.150 118.355 74.415 118.915 ;
        RECT 74.705 118.855 75.320 119.425 ;
        RECT 74.665 118.185 74.835 118.685 ;
        RECT 71.260 117.775 72.155 118.150 ;
        RECT 72.665 118.105 73.055 118.185 ;
        RECT 70.205 117.345 71.090 117.515 ;
        RECT 71.270 117.045 71.585 117.545 ;
        RECT 71.815 117.215 72.155 117.775 ;
        RECT 72.325 117.045 72.495 118.055 ;
        RECT 72.665 117.260 72.995 118.105 ;
        RECT 73.410 118.015 74.835 118.185 ;
        RECT 73.410 117.840 73.800 118.015 ;
        RECT 74.285 117.045 74.615 117.845 ;
        RECT 75.005 117.835 75.320 118.855 ;
        RECT 75.530 118.830 75.985 119.595 ;
        RECT 76.260 119.215 77.560 119.425 ;
        RECT 77.815 119.235 78.145 119.595 ;
        RECT 77.390 119.065 77.560 119.215 ;
        RECT 78.315 119.095 78.575 119.425 ;
        RECT 76.460 118.605 76.680 119.005 ;
        RECT 75.525 118.405 76.015 118.605 ;
        RECT 76.205 118.395 76.680 118.605 ;
        RECT 76.925 118.605 77.135 119.005 ;
        RECT 77.390 118.940 78.145 119.065 ;
        RECT 77.390 118.895 78.235 118.940 ;
        RECT 77.965 118.775 78.235 118.895 ;
        RECT 76.925 118.395 77.255 118.605 ;
        RECT 77.425 118.335 77.835 118.640 ;
        RECT 74.785 117.215 75.320 117.835 ;
        RECT 75.530 118.165 76.705 118.225 ;
        RECT 78.065 118.200 78.235 118.775 ;
        RECT 78.035 118.165 78.235 118.200 ;
        RECT 75.530 118.055 78.235 118.165 ;
        RECT 75.530 117.435 75.785 118.055 ;
        RECT 76.375 117.995 78.175 118.055 ;
        RECT 76.375 117.965 76.705 117.995 ;
        RECT 78.405 117.895 78.575 119.095 ;
        RECT 76.035 117.795 76.220 117.885 ;
        RECT 76.810 117.795 77.645 117.805 ;
        RECT 76.035 117.595 77.645 117.795 ;
        RECT 76.035 117.555 76.265 117.595 ;
        RECT 75.530 117.215 75.865 117.435 ;
        RECT 76.870 117.045 77.225 117.425 ;
        RECT 77.395 117.215 77.645 117.595 ;
        RECT 77.895 117.045 78.145 117.825 ;
        RECT 78.315 117.215 78.575 117.895 ;
        RECT 78.780 118.855 79.395 119.425 ;
        RECT 79.565 119.085 79.780 119.595 ;
        RECT 80.010 119.085 80.290 119.415 ;
        RECT 80.470 119.085 80.710 119.595 ;
        RECT 78.780 117.835 79.095 118.855 ;
        RECT 79.265 118.185 79.435 118.685 ;
        RECT 79.685 118.355 79.950 118.915 ;
        RECT 80.120 118.185 80.290 119.085 ;
        RECT 80.460 118.355 80.815 118.915 ;
        RECT 81.965 118.845 83.175 119.595 ;
        RECT 79.265 118.015 80.690 118.185 ;
        RECT 78.780 117.215 79.315 117.835 ;
        RECT 79.485 117.045 79.815 117.845 ;
        RECT 80.300 117.840 80.690 118.015 ;
        RECT 81.965 118.135 82.485 118.675 ;
        RECT 82.655 118.305 83.175 118.845 ;
        RECT 81.965 117.045 83.175 118.135 ;
        RECT 5.520 116.875 83.260 117.045 ;
        RECT 5.605 115.785 6.815 116.875 ;
        RECT 5.605 115.075 6.125 115.615 ;
        RECT 6.295 115.245 6.815 115.785 ;
        RECT 7.905 115.735 8.165 116.705 ;
        RECT 8.360 116.465 8.690 116.875 ;
        RECT 8.890 116.285 9.060 116.705 ;
        RECT 9.275 116.465 9.945 116.875 ;
        RECT 10.180 116.285 10.350 116.705 ;
        RECT 10.655 116.435 10.985 116.875 ;
        RECT 8.335 116.115 10.350 116.285 ;
        RECT 11.155 116.255 11.330 116.705 ;
        RECT 5.605 114.325 6.815 115.075 ;
        RECT 7.905 115.045 8.075 115.735 ;
        RECT 8.335 115.565 8.505 116.115 ;
        RECT 8.245 115.235 8.505 115.565 ;
        RECT 7.905 114.580 8.245 115.045 ;
        RECT 8.675 114.905 9.015 115.935 ;
        RECT 9.205 115.515 9.475 115.935 ;
        RECT 9.205 115.345 9.515 115.515 ;
        RECT 7.910 114.535 8.245 114.580 ;
        RECT 8.415 114.325 8.745 114.705 ;
        RECT 9.205 114.660 9.475 115.345 ;
        RECT 9.700 114.660 9.980 115.935 ;
        RECT 10.180 114.825 10.350 116.115 ;
        RECT 10.700 116.085 11.330 116.255 ;
        RECT 10.700 115.565 10.870 116.085 ;
        RECT 10.520 115.235 10.870 115.565 ;
        RECT 11.050 115.235 11.415 115.915 ;
        RECT 11.595 115.905 11.925 116.690 ;
        RECT 11.595 115.735 12.275 115.905 ;
        RECT 12.455 115.735 12.785 116.875 ;
        RECT 12.965 116.445 13.305 116.705 ;
        RECT 11.585 115.315 11.935 115.565 ;
        RECT 10.700 115.065 10.870 115.235 ;
        RECT 12.105 115.135 12.275 115.735 ;
        RECT 12.445 115.315 12.795 115.565 ;
        RECT 10.700 114.895 11.330 115.065 ;
        RECT 10.180 114.495 10.410 114.825 ;
        RECT 10.655 114.325 10.985 114.705 ;
        RECT 11.155 114.495 11.330 114.895 ;
        RECT 11.605 114.325 11.845 115.135 ;
        RECT 12.015 114.495 12.345 115.135 ;
        RECT 12.515 114.325 12.785 115.135 ;
        RECT 12.965 115.045 13.225 116.445 ;
        RECT 13.475 116.075 13.805 116.875 ;
        RECT 14.270 115.905 14.520 116.705 ;
        RECT 14.705 116.155 15.035 116.875 ;
        RECT 15.255 115.905 15.505 116.705 ;
        RECT 15.675 116.495 16.010 116.875 ;
        RECT 16.185 116.365 17.375 116.655 ;
        RECT 13.415 115.735 15.605 115.905 ;
        RECT 13.415 115.565 13.730 115.735 ;
        RECT 13.400 115.315 13.730 115.565 ;
        RECT 12.965 114.535 13.305 115.045 ;
        RECT 13.475 114.325 13.745 115.125 ;
        RECT 13.925 114.595 14.205 115.565 ;
        RECT 14.385 114.595 14.685 115.565 ;
        RECT 14.865 114.600 15.215 115.565 ;
        RECT 15.435 114.825 15.605 115.735 ;
        RECT 15.775 115.005 16.015 116.315 ;
        RECT 16.205 116.025 17.375 116.195 ;
        RECT 17.545 116.075 17.825 116.875 ;
        RECT 16.205 115.735 16.530 116.025 ;
        RECT 17.205 115.905 17.375 116.025 ;
        RECT 16.700 115.565 16.895 115.855 ;
        RECT 17.205 115.735 17.865 115.905 ;
        RECT 18.035 115.735 18.310 116.705 ;
        RECT 17.695 115.565 17.865 115.735 ;
        RECT 16.185 115.235 16.530 115.565 ;
        RECT 16.700 115.235 17.525 115.565 ;
        RECT 17.695 115.235 17.970 115.565 ;
        RECT 17.695 115.065 17.865 115.235 ;
        RECT 16.200 114.895 17.865 115.065 ;
        RECT 18.140 115.000 18.310 115.735 ;
        RECT 18.485 115.710 18.775 116.875 ;
        RECT 19.150 115.905 19.480 116.705 ;
        RECT 19.650 116.075 19.980 116.875 ;
        RECT 20.280 115.905 20.610 116.705 ;
        RECT 21.255 116.075 21.505 116.875 ;
        RECT 19.150 115.735 21.585 115.905 ;
        RECT 21.775 115.735 21.945 116.875 ;
        RECT 22.115 115.735 22.455 116.705 ;
        RECT 22.810 115.905 23.200 116.080 ;
        RECT 23.685 116.075 24.015 116.875 ;
        RECT 24.185 116.085 24.720 116.705 ;
        RECT 22.810 115.735 24.235 115.905 ;
        RECT 18.945 115.315 19.295 115.565 ;
        RECT 19.480 115.105 19.650 115.735 ;
        RECT 19.820 115.315 20.150 115.515 ;
        RECT 20.320 115.315 20.650 115.515 ;
        RECT 20.820 115.315 21.240 115.515 ;
        RECT 21.415 115.485 21.585 115.735 ;
        RECT 21.415 115.315 22.110 115.485 ;
        RECT 15.435 114.495 15.930 114.825 ;
        RECT 16.200 114.545 16.455 114.895 ;
        RECT 16.625 114.325 16.955 114.725 ;
        RECT 17.125 114.545 17.295 114.895 ;
        RECT 17.465 114.325 17.845 114.725 ;
        RECT 18.035 114.655 18.310 115.000 ;
        RECT 18.485 114.325 18.775 115.050 ;
        RECT 19.150 114.495 19.650 115.105 ;
        RECT 20.280 114.975 21.505 115.145 ;
        RECT 22.280 115.125 22.455 115.735 ;
        RECT 20.280 114.495 20.610 114.975 ;
        RECT 20.780 114.325 21.005 114.785 ;
        RECT 21.175 114.495 21.505 114.975 ;
        RECT 21.695 114.325 21.945 115.125 ;
        RECT 22.115 114.495 22.455 115.125 ;
        RECT 22.685 115.005 23.040 115.565 ;
        RECT 23.210 114.835 23.380 115.735 ;
        RECT 23.550 115.005 23.815 115.565 ;
        RECT 24.065 115.235 24.235 115.735 ;
        RECT 24.405 115.065 24.720 116.085 ;
        RECT 25.445 115.815 25.775 116.660 ;
        RECT 25.945 115.865 26.115 116.875 ;
        RECT 26.285 116.145 26.625 116.705 ;
        RECT 26.855 116.375 27.170 116.875 ;
        RECT 27.350 116.405 28.235 116.575 ;
        RECT 22.790 114.325 23.030 114.835 ;
        RECT 23.210 114.505 23.490 114.835 ;
        RECT 23.720 114.325 23.935 114.835 ;
        RECT 24.105 114.495 24.720 115.065 ;
        RECT 25.385 115.735 25.775 115.815 ;
        RECT 26.285 115.770 27.180 116.145 ;
        RECT 25.385 115.685 25.600 115.735 ;
        RECT 25.385 115.105 25.555 115.685 ;
        RECT 26.285 115.565 26.475 115.770 ;
        RECT 27.350 115.565 27.520 116.405 ;
        RECT 28.460 116.375 28.710 116.705 ;
        RECT 25.725 115.235 26.475 115.565 ;
        RECT 26.645 115.235 27.520 115.565 ;
        RECT 25.385 115.065 25.610 115.105 ;
        RECT 26.275 115.065 26.475 115.235 ;
        RECT 25.385 114.980 25.765 115.065 ;
        RECT 25.435 114.545 25.765 114.980 ;
        RECT 25.935 114.325 26.105 114.935 ;
        RECT 26.275 114.540 26.605 115.065 ;
        RECT 26.865 114.325 27.075 114.855 ;
        RECT 27.350 114.775 27.520 115.235 ;
        RECT 27.690 115.275 28.010 116.235 ;
        RECT 28.180 115.485 28.370 116.205 ;
        RECT 28.540 115.305 28.710 116.375 ;
        RECT 28.880 116.075 29.050 116.875 ;
        RECT 29.220 116.430 30.325 116.600 ;
        RECT 29.220 115.815 29.390 116.430 ;
        RECT 30.535 116.280 30.785 116.705 ;
        RECT 30.955 116.415 31.220 116.875 ;
        RECT 29.560 115.895 30.090 116.260 ;
        RECT 30.535 116.150 30.840 116.280 ;
        RECT 28.880 115.725 29.390 115.815 ;
        RECT 28.880 115.555 29.750 115.725 ;
        RECT 28.880 115.485 29.050 115.555 ;
        RECT 29.170 115.305 29.370 115.335 ;
        RECT 27.690 114.945 28.155 115.275 ;
        RECT 28.540 115.005 29.370 115.305 ;
        RECT 28.540 114.775 28.710 115.005 ;
        RECT 27.350 114.605 28.135 114.775 ;
        RECT 28.305 114.605 28.710 114.775 ;
        RECT 28.890 114.325 29.260 114.825 ;
        RECT 29.580 114.775 29.750 115.555 ;
        RECT 29.920 115.195 30.090 115.895 ;
        RECT 30.260 115.365 30.500 115.960 ;
        RECT 29.920 114.975 30.445 115.195 ;
        RECT 30.670 115.045 30.840 116.150 ;
        RECT 30.615 114.915 30.840 115.045 ;
        RECT 31.010 114.955 31.290 115.905 ;
        RECT 30.615 114.775 30.785 114.915 ;
        RECT 29.580 114.605 30.255 114.775 ;
        RECT 30.450 114.605 30.785 114.775 ;
        RECT 30.955 114.325 31.205 114.785 ;
        RECT 31.460 114.585 31.645 116.705 ;
        RECT 31.815 116.375 32.145 116.875 ;
        RECT 32.315 116.205 32.485 116.705 ;
        RECT 31.820 116.035 32.485 116.205 ;
        RECT 31.820 115.045 32.050 116.035 ;
        RECT 32.220 115.215 32.570 115.865 ;
        RECT 32.805 115.815 33.135 116.660 ;
        RECT 33.305 115.865 33.475 116.875 ;
        RECT 33.645 116.145 33.985 116.705 ;
        RECT 34.215 116.375 34.530 116.875 ;
        RECT 34.710 116.405 35.595 116.575 ;
        RECT 32.745 115.735 33.135 115.815 ;
        RECT 33.645 115.770 34.540 116.145 ;
        RECT 32.745 115.685 32.960 115.735 ;
        RECT 32.745 115.105 32.915 115.685 ;
        RECT 33.645 115.565 33.835 115.770 ;
        RECT 34.710 115.565 34.880 116.405 ;
        RECT 35.820 116.375 36.070 116.705 ;
        RECT 33.085 115.235 33.835 115.565 ;
        RECT 34.005 115.235 34.880 115.565 ;
        RECT 32.745 115.065 32.970 115.105 ;
        RECT 33.635 115.065 33.835 115.235 ;
        RECT 31.820 114.875 32.485 115.045 ;
        RECT 32.745 114.980 33.125 115.065 ;
        RECT 31.815 114.325 32.145 114.705 ;
        RECT 32.315 114.585 32.485 114.875 ;
        RECT 32.795 114.545 33.125 114.980 ;
        RECT 33.295 114.325 33.465 114.935 ;
        RECT 33.635 114.540 33.965 115.065 ;
        RECT 34.225 114.325 34.435 114.855 ;
        RECT 34.710 114.775 34.880 115.235 ;
        RECT 35.050 115.275 35.370 116.235 ;
        RECT 35.540 115.485 35.730 116.205 ;
        RECT 35.900 115.305 36.070 116.375 ;
        RECT 36.240 116.075 36.410 116.875 ;
        RECT 36.580 116.430 37.685 116.600 ;
        RECT 36.580 115.815 36.750 116.430 ;
        RECT 37.895 116.280 38.145 116.705 ;
        RECT 38.315 116.415 38.580 116.875 ;
        RECT 36.920 115.895 37.450 116.260 ;
        RECT 37.895 116.150 38.200 116.280 ;
        RECT 36.240 115.725 36.750 115.815 ;
        RECT 36.240 115.555 37.110 115.725 ;
        RECT 36.240 115.485 36.410 115.555 ;
        RECT 36.530 115.305 36.730 115.335 ;
        RECT 35.050 114.945 35.515 115.275 ;
        RECT 35.900 115.005 36.730 115.305 ;
        RECT 35.900 114.775 36.070 115.005 ;
        RECT 34.710 114.605 35.495 114.775 ;
        RECT 35.665 114.605 36.070 114.775 ;
        RECT 36.250 114.325 36.620 114.825 ;
        RECT 36.940 114.775 37.110 115.555 ;
        RECT 37.280 115.195 37.450 115.895 ;
        RECT 37.620 115.365 37.860 115.960 ;
        RECT 37.280 114.975 37.805 115.195 ;
        RECT 38.030 115.045 38.200 116.150 ;
        RECT 37.975 114.915 38.200 115.045 ;
        RECT 38.370 114.955 38.650 115.905 ;
        RECT 37.975 114.775 38.145 114.915 ;
        RECT 36.940 114.605 37.615 114.775 ;
        RECT 37.810 114.605 38.145 114.775 ;
        RECT 38.315 114.325 38.565 114.785 ;
        RECT 38.820 114.585 39.005 116.705 ;
        RECT 39.175 116.375 39.505 116.875 ;
        RECT 39.675 116.205 39.845 116.705 ;
        RECT 39.180 116.035 39.845 116.205 ;
        RECT 39.180 115.045 39.410 116.035 ;
        RECT 40.115 115.905 40.445 116.690 ;
        RECT 39.580 115.215 39.930 115.865 ;
        RECT 40.115 115.735 40.795 115.905 ;
        RECT 40.975 115.735 41.305 116.875 ;
        RECT 41.485 115.785 44.075 116.875 ;
        RECT 40.105 115.315 40.455 115.565 ;
        RECT 40.625 115.135 40.795 115.735 ;
        RECT 40.965 115.315 41.315 115.565 ;
        RECT 39.180 114.875 39.845 115.045 ;
        RECT 39.175 114.325 39.505 114.705 ;
        RECT 39.675 114.585 39.845 114.875 ;
        RECT 40.125 114.325 40.365 115.135 ;
        RECT 40.535 114.495 40.865 115.135 ;
        RECT 41.035 114.325 41.305 115.135 ;
        RECT 41.485 115.095 42.695 115.615 ;
        RECT 42.865 115.265 44.075 115.785 ;
        RECT 44.245 115.710 44.535 116.875 ;
        RECT 45.630 115.735 45.965 116.705 ;
        RECT 46.135 115.735 46.305 116.875 ;
        RECT 46.475 116.535 48.505 116.705 ;
        RECT 41.485 114.325 44.075 115.095 ;
        RECT 45.630 115.065 45.800 115.735 ;
        RECT 46.475 115.565 46.645 116.535 ;
        RECT 45.970 115.235 46.225 115.565 ;
        RECT 46.450 115.235 46.645 115.565 ;
        RECT 46.815 116.195 47.940 116.365 ;
        RECT 46.055 115.065 46.225 115.235 ;
        RECT 46.815 115.065 46.985 116.195 ;
        RECT 44.245 114.325 44.535 115.050 ;
        RECT 45.630 114.495 45.885 115.065 ;
        RECT 46.055 114.895 46.985 115.065 ;
        RECT 47.155 115.855 48.165 116.025 ;
        RECT 47.155 115.055 47.325 115.855 ;
        RECT 46.810 114.860 46.985 114.895 ;
        RECT 46.055 114.325 46.385 114.725 ;
        RECT 46.810 114.495 47.340 114.860 ;
        RECT 47.530 114.835 47.805 115.655 ;
        RECT 47.525 114.665 47.805 114.835 ;
        RECT 47.530 114.495 47.805 114.665 ;
        RECT 47.975 114.495 48.165 115.855 ;
        RECT 48.335 115.870 48.505 116.535 ;
        RECT 48.675 116.115 48.845 116.875 ;
        RECT 49.080 116.115 49.595 116.525 ;
        RECT 48.335 115.680 49.085 115.870 ;
        RECT 49.255 115.305 49.595 116.115 ;
        RECT 49.880 116.245 50.165 116.705 ;
        RECT 50.335 116.415 50.605 116.875 ;
        RECT 49.880 116.025 50.835 116.245 ;
        RECT 48.365 115.135 49.595 115.305 ;
        RECT 49.765 115.295 50.455 115.855 ;
        RECT 48.345 114.325 48.855 114.860 ;
        RECT 49.075 114.530 49.320 115.135 ;
        RECT 50.625 115.125 50.835 116.025 ;
        RECT 49.880 114.955 50.835 115.125 ;
        RECT 51.005 115.855 51.405 116.705 ;
        RECT 51.595 116.245 51.875 116.705 ;
        RECT 52.395 116.415 52.720 116.875 ;
        RECT 51.595 116.025 52.720 116.245 ;
        RECT 51.005 115.295 52.100 115.855 ;
        RECT 52.270 115.565 52.720 116.025 ;
        RECT 52.890 115.735 53.275 116.705 ;
        RECT 49.880 114.495 50.165 114.955 ;
        RECT 50.335 114.325 50.605 114.785 ;
        RECT 51.005 114.495 51.405 115.295 ;
        RECT 52.270 115.235 52.825 115.565 ;
        RECT 52.270 115.125 52.720 115.235 ;
        RECT 51.595 114.955 52.720 115.125 ;
        RECT 52.995 115.065 53.275 115.735 ;
        RECT 51.595 114.495 51.875 114.955 ;
        RECT 52.395 114.325 52.720 114.785 ;
        RECT 52.890 114.495 53.275 115.065 ;
        RECT 53.445 114.605 53.725 116.705 ;
        RECT 53.915 116.115 54.700 116.875 ;
        RECT 55.095 116.045 55.480 116.705 ;
        RECT 55.095 115.945 55.505 116.045 ;
        RECT 53.895 115.735 55.505 115.945 ;
        RECT 55.805 115.855 56.005 116.645 ;
        RECT 53.895 115.135 54.170 115.735 ;
        RECT 55.675 115.685 56.005 115.855 ;
        RECT 56.175 115.695 56.495 116.875 ;
        RECT 56.670 115.735 56.990 116.875 ;
        RECT 55.675 115.565 55.855 115.685 ;
        RECT 57.170 115.565 57.365 116.615 ;
        RECT 57.545 116.025 57.875 116.705 ;
        RECT 58.075 116.075 58.330 116.875 ;
        RECT 58.510 116.075 58.765 116.875 ;
        RECT 58.965 116.025 59.295 116.705 ;
        RECT 57.545 115.745 57.895 116.025 ;
        RECT 54.340 115.315 54.695 115.565 ;
        RECT 54.890 115.515 55.355 115.565 ;
        RECT 54.885 115.345 55.355 115.515 ;
        RECT 54.890 115.315 55.355 115.345 ;
        RECT 55.525 115.315 55.855 115.565 ;
        RECT 56.730 115.515 56.990 115.565 ;
        RECT 56.030 115.315 56.495 115.515 ;
        RECT 56.725 115.345 56.990 115.515 ;
        RECT 56.730 115.235 56.990 115.345 ;
        RECT 57.170 115.235 57.555 115.565 ;
        RECT 57.725 115.365 57.895 115.745 ;
        RECT 58.085 115.535 58.330 115.895 ;
        RECT 58.510 115.535 58.755 115.895 ;
        RECT 58.945 115.745 59.295 116.025 ;
        RECT 58.945 115.365 59.115 115.745 ;
        RECT 59.475 115.565 59.670 116.615 ;
        RECT 59.850 115.735 60.170 116.875 ;
        RECT 60.345 116.025 60.605 116.705 ;
        RECT 60.775 116.095 61.025 116.875 ;
        RECT 61.275 116.325 61.525 116.705 ;
        RECT 61.695 116.495 62.050 116.875 ;
        RECT 63.055 116.485 63.390 116.705 ;
        RECT 62.655 116.325 62.885 116.365 ;
        RECT 61.275 116.125 62.885 116.325 ;
        RECT 61.275 116.115 62.110 116.125 ;
        RECT 62.700 116.035 62.885 116.125 ;
        RECT 57.725 115.195 58.245 115.365 ;
        RECT 53.895 114.955 55.145 115.135 ;
        RECT 54.780 114.885 55.145 114.955 ;
        RECT 55.315 114.935 56.495 115.105 ;
        RECT 53.955 114.325 54.125 114.785 ;
        RECT 55.315 114.715 55.645 114.935 ;
        RECT 54.395 114.535 55.645 114.715 ;
        RECT 55.815 114.325 55.985 114.765 ;
        RECT 56.155 114.520 56.495 114.935 ;
        RECT 56.670 114.855 57.885 115.025 ;
        RECT 56.670 114.505 56.960 114.855 ;
        RECT 57.155 114.325 57.485 114.685 ;
        RECT 57.655 114.550 57.885 114.855 ;
        RECT 58.075 114.630 58.245 115.195 ;
        RECT 58.595 115.195 59.115 115.365 ;
        RECT 59.285 115.235 59.670 115.565 ;
        RECT 59.850 115.515 60.110 115.565 ;
        RECT 59.850 115.345 60.115 115.515 ;
        RECT 59.850 115.235 60.110 115.345 ;
        RECT 58.595 114.630 58.765 115.195 ;
        RECT 58.955 114.855 60.170 115.025 ;
        RECT 58.955 114.550 59.185 114.855 ;
        RECT 59.355 114.325 59.685 114.685 ;
        RECT 59.880 114.505 60.170 114.855 ;
        RECT 60.345 114.835 60.515 116.025 ;
        RECT 62.215 115.925 62.545 115.955 ;
        RECT 60.745 115.865 62.545 115.925 ;
        RECT 63.135 115.865 63.390 116.485 ;
        RECT 63.680 116.245 63.965 116.705 ;
        RECT 64.135 116.415 64.405 116.875 ;
        RECT 63.680 116.025 64.635 116.245 ;
        RECT 60.685 115.755 63.390 115.865 ;
        RECT 60.685 115.720 60.885 115.755 ;
        RECT 60.685 115.145 60.855 115.720 ;
        RECT 62.215 115.695 63.390 115.755 ;
        RECT 61.085 115.280 61.495 115.585 ;
        RECT 61.665 115.315 61.995 115.525 ;
        RECT 60.685 115.025 60.955 115.145 ;
        RECT 60.685 114.980 61.530 115.025 ;
        RECT 60.775 114.855 61.530 114.980 ;
        RECT 61.785 114.915 61.995 115.315 ;
        RECT 62.240 115.315 62.715 115.525 ;
        RECT 62.905 115.315 63.395 115.515 ;
        RECT 62.240 114.915 62.460 115.315 ;
        RECT 63.565 115.295 64.255 115.855 ;
        RECT 64.425 115.125 64.635 116.025 ;
        RECT 60.345 114.825 60.575 114.835 ;
        RECT 60.345 114.495 60.605 114.825 ;
        RECT 61.360 114.705 61.530 114.855 ;
        RECT 60.775 114.325 61.105 114.685 ;
        RECT 61.360 114.495 62.660 114.705 ;
        RECT 62.935 114.325 63.390 115.090 ;
        RECT 63.680 114.955 64.635 115.125 ;
        RECT 64.805 115.855 65.205 116.705 ;
        RECT 65.395 116.245 65.675 116.705 ;
        RECT 66.195 116.415 66.520 116.875 ;
        RECT 65.395 116.025 66.520 116.245 ;
        RECT 64.805 115.295 65.900 115.855 ;
        RECT 66.070 115.565 66.520 116.025 ;
        RECT 66.690 115.735 67.075 116.705 ;
        RECT 67.255 115.735 67.585 116.875 ;
        RECT 63.680 114.495 63.965 114.955 ;
        RECT 64.135 114.325 64.405 114.785 ;
        RECT 64.805 114.495 65.205 115.295 ;
        RECT 66.070 115.235 66.625 115.565 ;
        RECT 66.070 115.125 66.520 115.235 ;
        RECT 65.395 114.955 66.520 115.125 ;
        RECT 66.795 115.065 67.075 115.735 ;
        RECT 65.395 114.495 65.675 114.955 ;
        RECT 66.195 114.325 66.520 114.785 ;
        RECT 66.690 114.495 67.075 115.065 ;
        RECT 67.245 114.985 67.585 115.565 ;
        RECT 67.755 115.535 68.115 116.705 ;
        RECT 68.315 115.705 68.645 116.875 ;
        RECT 68.845 115.535 69.175 116.705 ;
        RECT 69.375 115.705 69.705 116.875 ;
        RECT 70.005 115.710 70.295 116.875 ;
        RECT 70.670 115.905 71.000 116.705 ;
        RECT 71.170 116.075 71.500 116.875 ;
        RECT 71.800 115.905 72.130 116.705 ;
        RECT 72.775 116.075 73.025 116.875 ;
        RECT 70.670 115.735 73.105 115.905 ;
        RECT 73.295 115.735 73.465 116.875 ;
        RECT 73.635 115.735 73.975 116.705 ;
        RECT 74.235 116.205 74.405 116.705 ;
        RECT 74.575 116.375 74.905 116.875 ;
        RECT 74.235 116.035 74.900 116.205 ;
        RECT 67.755 115.255 69.175 115.535 ;
        RECT 70.465 115.315 70.815 115.565 ;
        RECT 67.755 114.920 68.115 115.255 ;
        RECT 71.000 115.105 71.170 115.735 ;
        RECT 71.340 115.315 71.670 115.515 ;
        RECT 71.840 115.315 72.170 115.515 ;
        RECT 72.340 115.315 72.760 115.515 ;
        RECT 72.935 115.485 73.105 115.735 ;
        RECT 72.935 115.315 73.630 115.485 ;
        RECT 73.800 115.175 73.975 115.735 ;
        RECT 74.150 115.215 74.500 115.865 ;
        RECT 67.255 114.325 67.585 114.815 ;
        RECT 67.755 114.495 68.375 114.920 ;
        RECT 68.835 114.325 69.165 115.015 ;
        RECT 70.005 114.325 70.295 115.050 ;
        RECT 70.670 114.495 71.170 115.105 ;
        RECT 71.800 114.975 73.025 115.145 ;
        RECT 73.745 115.125 73.975 115.175 ;
        RECT 71.800 114.495 72.130 114.975 ;
        RECT 72.300 114.325 72.525 114.785 ;
        RECT 72.695 114.495 73.025 114.975 ;
        RECT 73.215 114.325 73.465 115.125 ;
        RECT 73.635 114.495 73.975 115.125 ;
        RECT 74.670 115.045 74.900 116.035 ;
        RECT 74.235 114.875 74.900 115.045 ;
        RECT 74.235 114.585 74.405 114.875 ;
        RECT 74.575 114.325 74.905 114.705 ;
        RECT 75.075 114.585 75.260 116.705 ;
        RECT 75.500 116.415 75.765 116.875 ;
        RECT 75.935 116.280 76.185 116.705 ;
        RECT 76.395 116.430 77.500 116.600 ;
        RECT 75.880 116.150 76.185 116.280 ;
        RECT 75.430 114.955 75.710 115.905 ;
        RECT 75.880 115.045 76.050 116.150 ;
        RECT 76.220 115.365 76.460 115.960 ;
        RECT 76.630 115.895 77.160 116.260 ;
        RECT 76.630 115.195 76.800 115.895 ;
        RECT 77.330 115.815 77.500 116.430 ;
        RECT 77.670 116.075 77.840 116.875 ;
        RECT 78.010 116.375 78.260 116.705 ;
        RECT 78.485 116.405 79.370 116.575 ;
        RECT 77.330 115.725 77.840 115.815 ;
        RECT 75.880 114.915 76.105 115.045 ;
        RECT 76.275 114.975 76.800 115.195 ;
        RECT 76.970 115.555 77.840 115.725 ;
        RECT 75.515 114.325 75.765 114.785 ;
        RECT 75.935 114.775 76.105 114.915 ;
        RECT 76.970 114.775 77.140 115.555 ;
        RECT 77.670 115.485 77.840 115.555 ;
        RECT 77.350 115.305 77.550 115.335 ;
        RECT 78.010 115.305 78.180 116.375 ;
        RECT 78.350 115.485 78.540 116.205 ;
        RECT 77.350 115.005 78.180 115.305 ;
        RECT 78.710 115.275 79.030 116.235 ;
        RECT 75.935 114.605 76.270 114.775 ;
        RECT 76.465 114.605 77.140 114.775 ;
        RECT 77.460 114.325 77.830 114.825 ;
        RECT 78.010 114.775 78.180 115.005 ;
        RECT 78.565 114.945 79.030 115.275 ;
        RECT 79.200 115.565 79.370 116.405 ;
        RECT 79.550 116.375 79.865 116.875 ;
        RECT 80.095 116.145 80.435 116.705 ;
        RECT 79.540 115.770 80.435 116.145 ;
        RECT 80.605 115.865 80.775 116.875 ;
        RECT 80.245 115.565 80.435 115.770 ;
        RECT 80.945 115.815 81.275 116.660 ;
        RECT 80.945 115.735 81.335 115.815 ;
        RECT 81.120 115.685 81.335 115.735 ;
        RECT 79.200 115.235 80.075 115.565 ;
        RECT 80.245 115.235 80.995 115.565 ;
        RECT 79.200 114.775 79.370 115.235 ;
        RECT 80.245 115.065 80.445 115.235 ;
        RECT 81.165 115.105 81.335 115.685 ;
        RECT 81.965 115.785 83.175 116.875 ;
        RECT 81.965 115.245 82.485 115.785 ;
        RECT 81.110 115.065 81.335 115.105 ;
        RECT 82.655 115.075 83.175 115.615 ;
        RECT 78.010 114.605 78.415 114.775 ;
        RECT 78.585 114.605 79.370 114.775 ;
        RECT 79.645 114.325 79.855 114.855 ;
        RECT 80.115 114.540 80.445 115.065 ;
        RECT 80.955 114.980 81.335 115.065 ;
        RECT 80.615 114.325 80.785 114.935 ;
        RECT 80.955 114.545 81.285 114.980 ;
        RECT 81.965 114.325 83.175 115.075 ;
        RECT 5.520 114.155 83.260 114.325 ;
        RECT 5.605 113.405 6.815 114.155 ;
        RECT 5.605 112.865 6.125 113.405 ;
        RECT 6.985 113.385 9.575 114.155 ;
        RECT 9.755 113.425 10.055 114.155 ;
        RECT 6.295 112.695 6.815 113.235 ;
        RECT 6.985 112.865 8.195 113.385 ;
        RECT 10.235 113.245 10.465 113.865 ;
        RECT 10.665 113.595 10.890 113.975 ;
        RECT 11.060 113.765 11.390 114.155 ;
        RECT 11.585 113.775 12.475 113.945 ;
        RECT 10.665 113.415 10.995 113.595 ;
        RECT 8.365 112.695 9.575 113.215 ;
        RECT 9.760 112.915 10.055 113.245 ;
        RECT 10.235 112.915 10.650 113.245 ;
        RECT 10.820 112.745 10.995 113.415 ;
        RECT 11.165 112.915 11.405 113.565 ;
        RECT 11.585 113.220 12.135 113.605 ;
        RECT 12.305 113.050 12.475 113.775 ;
        RECT 11.585 112.980 12.475 113.050 ;
        RECT 12.645 113.450 12.865 113.935 ;
        RECT 13.035 113.615 13.285 114.155 ;
        RECT 13.455 113.505 13.715 113.985 ;
        RECT 12.645 113.025 12.975 113.450 ;
        RECT 11.585 112.955 12.480 112.980 ;
        RECT 11.585 112.940 12.490 112.955 ;
        RECT 11.585 112.925 12.495 112.940 ;
        RECT 11.585 112.920 12.505 112.925 ;
        RECT 11.585 112.910 12.510 112.920 ;
        RECT 11.585 112.900 12.515 112.910 ;
        RECT 11.585 112.895 12.525 112.900 ;
        RECT 11.585 112.885 12.535 112.895 ;
        RECT 11.585 112.880 12.545 112.885 ;
        RECT 5.605 111.605 6.815 112.695 ;
        RECT 6.985 111.605 9.575 112.695 ;
        RECT 9.755 112.385 10.650 112.715 ;
        RECT 10.820 112.555 11.405 112.745 ;
        RECT 9.755 112.215 10.960 112.385 ;
        RECT 9.755 111.785 10.085 112.215 ;
        RECT 10.265 111.605 10.460 112.045 ;
        RECT 10.630 111.785 10.960 112.215 ;
        RECT 11.130 111.785 11.405 112.555 ;
        RECT 11.585 112.430 11.845 112.880 ;
        RECT 12.210 112.875 12.545 112.880 ;
        RECT 12.210 112.870 12.560 112.875 ;
        RECT 12.210 112.860 12.575 112.870 ;
        RECT 12.210 112.855 12.600 112.860 ;
        RECT 13.145 112.855 13.375 113.250 ;
        RECT 12.210 112.850 13.375 112.855 ;
        RECT 12.240 112.815 13.375 112.850 ;
        RECT 12.275 112.790 13.375 112.815 ;
        RECT 12.305 112.760 13.375 112.790 ;
        RECT 12.325 112.730 13.375 112.760 ;
        RECT 12.345 112.700 13.375 112.730 ;
        RECT 12.415 112.690 13.375 112.700 ;
        RECT 12.440 112.680 13.375 112.690 ;
        RECT 12.460 112.665 13.375 112.680 ;
        RECT 12.480 112.650 13.375 112.665 ;
        RECT 12.485 112.640 13.270 112.650 ;
        RECT 12.500 112.605 13.270 112.640 ;
        RECT 12.015 112.285 12.345 112.530 ;
        RECT 12.515 112.355 13.270 112.605 ;
        RECT 13.545 112.475 13.715 113.505 ;
        RECT 12.015 112.260 12.200 112.285 ;
        RECT 11.585 112.160 12.200 112.260 ;
        RECT 11.585 111.605 12.190 112.160 ;
        RECT 12.365 111.775 12.845 112.115 ;
        RECT 13.015 111.605 13.270 112.150 ;
        RECT 13.440 111.775 13.715 112.475 ;
        RECT 14.345 113.415 14.810 113.960 ;
        RECT 14.345 112.455 14.515 113.415 ;
        RECT 15.315 113.335 15.485 114.155 ;
        RECT 15.655 113.505 15.985 113.985 ;
        RECT 16.155 113.765 16.505 114.155 ;
        RECT 16.675 113.585 16.905 113.985 ;
        RECT 16.395 113.505 16.905 113.585 ;
        RECT 15.655 113.415 16.905 113.505 ;
        RECT 17.075 113.415 17.395 113.895 ;
        RECT 15.655 113.335 16.565 113.415 ;
        RECT 14.685 112.795 14.930 113.245 ;
        RECT 15.190 112.965 15.885 113.165 ;
        RECT 16.055 112.995 16.655 113.165 ;
        RECT 16.055 112.795 16.225 112.995 ;
        RECT 16.885 112.825 17.055 113.245 ;
        RECT 14.685 112.625 16.225 112.795 ;
        RECT 16.395 112.655 17.055 112.825 ;
        RECT 16.395 112.455 16.565 112.655 ;
        RECT 17.225 112.485 17.395 113.415 ;
        RECT 17.565 113.385 19.235 114.155 ;
        RECT 17.565 112.865 18.315 113.385 ;
        RECT 19.405 113.335 19.665 114.155 ;
        RECT 19.835 113.335 20.165 113.755 ;
        RECT 20.345 113.585 20.605 113.985 ;
        RECT 20.775 113.755 21.105 114.155 ;
        RECT 21.275 113.585 21.445 113.935 ;
        RECT 21.615 113.755 21.990 114.155 ;
        RECT 20.345 113.415 22.010 113.585 ;
        RECT 22.180 113.480 22.455 113.825 ;
        RECT 19.915 113.245 20.165 113.335 ;
        RECT 21.840 113.245 22.010 113.415 ;
        RECT 18.485 112.695 19.235 113.215 ;
        RECT 19.410 112.915 19.745 113.165 ;
        RECT 19.915 112.915 20.630 113.245 ;
        RECT 20.845 112.915 21.670 113.245 ;
        RECT 21.840 112.915 22.115 113.245 ;
        RECT 14.345 112.285 16.565 112.455 ;
        RECT 16.735 112.285 17.395 112.485 ;
        RECT 14.345 111.605 14.645 112.115 ;
        RECT 14.815 111.775 15.145 112.285 ;
        RECT 16.735 112.115 16.905 112.285 ;
        RECT 15.315 111.605 15.945 112.115 ;
        RECT 16.525 111.945 16.905 112.115 ;
        RECT 17.075 111.605 17.375 112.115 ;
        RECT 17.565 111.605 19.235 112.695 ;
        RECT 19.405 111.605 19.665 112.745 ;
        RECT 19.915 112.355 20.085 112.915 ;
        RECT 20.345 112.455 20.675 112.745 ;
        RECT 20.845 112.625 21.090 112.915 ;
        RECT 21.840 112.745 22.010 112.915 ;
        RECT 22.285 112.745 22.455 113.480 ;
        RECT 22.640 113.585 22.895 113.935 ;
        RECT 23.065 113.755 23.395 114.155 ;
        RECT 23.565 113.585 23.735 113.935 ;
        RECT 23.905 113.755 24.285 114.155 ;
        RECT 22.640 113.415 24.305 113.585 ;
        RECT 24.475 113.480 24.750 113.825 ;
        RECT 24.975 113.765 25.305 114.155 ;
        RECT 25.475 113.585 25.645 113.905 ;
        RECT 25.815 113.765 26.145 114.155 ;
        RECT 26.560 113.755 27.515 113.925 ;
        RECT 24.135 113.245 24.305 113.415 ;
        RECT 22.625 112.915 22.970 113.245 ;
        RECT 23.140 112.915 23.965 113.245 ;
        RECT 24.135 112.915 24.410 113.245 ;
        RECT 21.350 112.575 22.010 112.745 ;
        RECT 21.350 112.455 21.520 112.575 ;
        RECT 20.345 112.285 21.520 112.455 ;
        RECT 19.905 111.785 21.520 112.115 ;
        RECT 21.690 111.605 21.970 112.405 ;
        RECT 22.180 111.775 22.455 112.745 ;
        RECT 22.645 112.455 22.970 112.745 ;
        RECT 23.140 112.625 23.335 112.915 ;
        RECT 24.135 112.745 24.305 112.915 ;
        RECT 24.580 112.745 24.750 113.480 ;
        RECT 23.645 112.575 24.305 112.745 ;
        RECT 23.645 112.455 23.815 112.575 ;
        RECT 22.645 112.285 23.815 112.455 ;
        RECT 22.625 111.825 23.815 112.115 ;
        RECT 23.985 111.605 24.265 112.405 ;
        RECT 24.475 111.775 24.750 112.745 ;
        RECT 24.925 113.415 27.175 113.585 ;
        RECT 24.925 112.455 25.095 113.415 ;
        RECT 25.265 112.795 25.510 113.245 ;
        RECT 25.680 112.965 26.230 113.165 ;
        RECT 26.400 112.995 26.775 113.165 ;
        RECT 26.400 112.795 26.570 112.995 ;
        RECT 26.945 112.915 27.175 113.415 ;
        RECT 25.265 112.625 26.570 112.795 ;
        RECT 27.345 112.875 27.515 113.755 ;
        RECT 27.685 113.320 27.975 114.155 ;
        RECT 28.155 113.430 28.485 113.940 ;
        RECT 28.655 113.755 28.985 114.155 ;
        RECT 30.035 113.585 30.365 113.925 ;
        RECT 30.535 113.755 30.865 114.155 ;
        RECT 27.345 112.705 27.975 112.875 ;
        RECT 24.925 111.775 25.305 112.455 ;
        RECT 25.895 111.605 26.065 112.455 ;
        RECT 26.235 112.285 27.475 112.455 ;
        RECT 26.235 111.775 26.565 112.285 ;
        RECT 26.735 111.605 26.905 112.115 ;
        RECT 27.075 111.775 27.475 112.285 ;
        RECT 27.655 111.775 27.975 112.705 ;
        RECT 28.155 112.665 28.345 113.430 ;
        RECT 28.655 113.415 31.020 113.585 ;
        RECT 31.365 113.430 31.655 114.155 ;
        RECT 31.830 113.755 32.165 114.155 ;
        RECT 32.335 113.585 32.540 113.985 ;
        RECT 32.750 113.675 33.025 114.155 ;
        RECT 33.235 113.655 33.495 113.985 ;
        RECT 28.655 113.245 28.825 113.415 ;
        RECT 28.515 112.915 28.825 113.245 ;
        RECT 28.995 112.915 29.300 113.245 ;
        RECT 28.155 111.815 28.485 112.665 ;
        RECT 28.655 111.605 28.905 112.745 ;
        RECT 29.085 112.585 29.300 112.915 ;
        RECT 29.475 112.585 29.760 113.245 ;
        RECT 29.955 112.585 30.220 113.245 ;
        RECT 30.435 112.585 30.680 113.245 ;
        RECT 30.850 112.415 31.020 113.415 ;
        RECT 31.855 113.415 32.540 113.585 ;
        RECT 29.095 112.245 30.385 112.415 ;
        RECT 29.095 111.825 29.345 112.245 ;
        RECT 29.575 111.605 29.905 112.075 ;
        RECT 30.135 111.825 30.385 112.245 ;
        RECT 30.565 112.245 31.020 112.415 ;
        RECT 30.565 111.815 30.895 112.245 ;
        RECT 31.365 111.605 31.655 112.770 ;
        RECT 31.855 112.385 32.195 113.415 ;
        RECT 32.365 112.745 32.615 113.245 ;
        RECT 32.795 112.915 33.155 113.495 ;
        RECT 33.325 112.745 33.495 113.655 ;
        RECT 34.675 113.605 34.845 113.895 ;
        RECT 35.015 113.775 35.345 114.155 ;
        RECT 34.675 113.435 35.340 113.605 ;
        RECT 32.365 112.575 33.495 112.745 ;
        RECT 34.590 112.615 34.940 113.265 ;
        RECT 31.855 112.210 32.520 112.385 ;
        RECT 31.830 111.605 32.165 112.030 ;
        RECT 32.335 111.805 32.520 112.210 ;
        RECT 32.725 111.605 33.055 112.385 ;
        RECT 33.225 111.805 33.495 112.575 ;
        RECT 35.110 112.445 35.340 113.435 ;
        RECT 34.675 112.275 35.340 112.445 ;
        RECT 34.675 111.775 34.845 112.275 ;
        RECT 35.015 111.605 35.345 112.105 ;
        RECT 35.515 111.775 35.700 113.895 ;
        RECT 35.955 113.695 36.205 114.155 ;
        RECT 36.375 113.705 36.710 113.875 ;
        RECT 36.905 113.705 37.580 113.875 ;
        RECT 36.375 113.565 36.545 113.705 ;
        RECT 35.870 112.575 36.150 113.525 ;
        RECT 36.320 113.435 36.545 113.565 ;
        RECT 36.320 112.330 36.490 113.435 ;
        RECT 36.715 113.285 37.240 113.505 ;
        RECT 36.660 112.520 36.900 113.115 ;
        RECT 37.070 112.585 37.240 113.285 ;
        RECT 37.410 112.925 37.580 113.705 ;
        RECT 37.900 113.655 38.270 114.155 ;
        RECT 38.450 113.705 38.855 113.875 ;
        RECT 39.025 113.705 39.810 113.875 ;
        RECT 38.450 113.475 38.620 113.705 ;
        RECT 37.790 113.175 38.620 113.475 ;
        RECT 39.005 113.205 39.470 113.535 ;
        RECT 37.790 113.145 37.990 113.175 ;
        RECT 38.110 112.925 38.280 112.995 ;
        RECT 37.410 112.755 38.280 112.925 ;
        RECT 37.770 112.665 38.280 112.755 ;
        RECT 36.320 112.200 36.625 112.330 ;
        RECT 37.070 112.220 37.600 112.585 ;
        RECT 35.940 111.605 36.205 112.065 ;
        RECT 36.375 111.775 36.625 112.200 ;
        RECT 37.770 112.050 37.940 112.665 ;
        RECT 36.835 111.880 37.940 112.050 ;
        RECT 38.110 111.605 38.280 112.405 ;
        RECT 38.450 112.105 38.620 113.175 ;
        RECT 38.790 112.275 38.980 112.995 ;
        RECT 39.150 112.245 39.470 113.205 ;
        RECT 39.640 113.245 39.810 113.705 ;
        RECT 40.085 113.625 40.295 114.155 ;
        RECT 40.555 113.415 40.885 113.940 ;
        RECT 41.055 113.545 41.225 114.155 ;
        RECT 41.395 113.500 41.725 113.935 ;
        RECT 42.035 113.605 42.205 113.895 ;
        RECT 42.375 113.775 42.705 114.155 ;
        RECT 41.395 113.415 41.775 113.500 ;
        RECT 42.035 113.435 42.700 113.605 ;
        RECT 40.685 113.245 40.885 113.415 ;
        RECT 41.550 113.375 41.775 113.415 ;
        RECT 39.640 112.915 40.515 113.245 ;
        RECT 40.685 112.915 41.435 113.245 ;
        RECT 38.450 111.775 38.700 112.105 ;
        RECT 39.640 112.075 39.810 112.915 ;
        RECT 40.685 112.710 40.875 112.915 ;
        RECT 41.605 112.795 41.775 113.375 ;
        RECT 41.560 112.745 41.775 112.795 ;
        RECT 39.980 112.335 40.875 112.710 ;
        RECT 41.385 112.665 41.775 112.745 ;
        RECT 38.925 111.905 39.810 112.075 ;
        RECT 39.990 111.605 40.305 112.105 ;
        RECT 40.535 111.775 40.875 112.335 ;
        RECT 41.045 111.605 41.215 112.615 ;
        RECT 41.385 111.820 41.715 112.665 ;
        RECT 41.950 112.615 42.300 113.265 ;
        RECT 42.470 112.445 42.700 113.435 ;
        RECT 42.035 112.275 42.700 112.445 ;
        RECT 42.035 111.775 42.205 112.275 ;
        RECT 42.375 111.605 42.705 112.105 ;
        RECT 42.875 111.775 43.060 113.895 ;
        RECT 43.315 113.695 43.565 114.155 ;
        RECT 43.735 113.705 44.070 113.875 ;
        RECT 44.265 113.705 44.940 113.875 ;
        RECT 43.735 113.565 43.905 113.705 ;
        RECT 43.230 112.575 43.510 113.525 ;
        RECT 43.680 113.435 43.905 113.565 ;
        RECT 43.680 112.330 43.850 113.435 ;
        RECT 44.075 113.285 44.600 113.505 ;
        RECT 44.020 112.520 44.260 113.115 ;
        RECT 44.430 112.585 44.600 113.285 ;
        RECT 44.770 112.925 44.940 113.705 ;
        RECT 45.260 113.655 45.630 114.155 ;
        RECT 45.810 113.705 46.215 113.875 ;
        RECT 46.385 113.705 47.170 113.875 ;
        RECT 45.810 113.475 45.980 113.705 ;
        RECT 45.150 113.175 45.980 113.475 ;
        RECT 46.365 113.205 46.830 113.535 ;
        RECT 45.150 113.145 45.350 113.175 ;
        RECT 45.470 112.925 45.640 112.995 ;
        RECT 44.770 112.755 45.640 112.925 ;
        RECT 45.130 112.665 45.640 112.755 ;
        RECT 43.680 112.200 43.985 112.330 ;
        RECT 44.430 112.220 44.960 112.585 ;
        RECT 43.300 111.605 43.565 112.065 ;
        RECT 43.735 111.775 43.985 112.200 ;
        RECT 45.130 112.050 45.300 112.665 ;
        RECT 44.195 111.880 45.300 112.050 ;
        RECT 45.470 111.605 45.640 112.405 ;
        RECT 45.810 112.105 45.980 113.175 ;
        RECT 46.150 112.275 46.340 112.995 ;
        RECT 46.510 112.245 46.830 113.205 ;
        RECT 47.000 113.245 47.170 113.705 ;
        RECT 47.445 113.625 47.655 114.155 ;
        RECT 47.915 113.415 48.245 113.940 ;
        RECT 48.415 113.545 48.585 114.155 ;
        RECT 48.755 113.500 49.085 113.935 ;
        RECT 48.755 113.415 49.135 113.500 ;
        RECT 48.045 113.245 48.245 113.415 ;
        RECT 48.910 113.375 49.135 113.415 ;
        RECT 47.000 112.915 47.875 113.245 ;
        RECT 48.045 112.915 48.795 113.245 ;
        RECT 45.810 111.775 46.060 112.105 ;
        RECT 47.000 112.075 47.170 112.915 ;
        RECT 48.045 112.710 48.235 112.915 ;
        RECT 48.965 112.795 49.135 113.375 ;
        RECT 48.920 112.745 49.135 112.795 ;
        RECT 47.340 112.335 48.235 112.710 ;
        RECT 48.745 112.665 49.135 112.745 ;
        RECT 49.305 113.415 49.690 113.985 ;
        RECT 49.860 113.695 50.185 114.155 ;
        RECT 50.705 113.525 50.985 113.985 ;
        RECT 49.305 112.745 49.585 113.415 ;
        RECT 49.860 113.355 50.985 113.525 ;
        RECT 49.860 113.245 50.310 113.355 ;
        RECT 49.755 112.915 50.310 113.245 ;
        RECT 51.175 113.185 51.575 113.985 ;
        RECT 51.975 113.695 52.245 114.155 ;
        RECT 52.415 113.525 52.700 113.985 ;
        RECT 46.285 111.905 47.170 112.075 ;
        RECT 47.350 111.605 47.665 112.105 ;
        RECT 47.895 111.775 48.235 112.335 ;
        RECT 48.405 111.605 48.575 112.615 ;
        RECT 48.745 111.820 49.075 112.665 ;
        RECT 49.305 111.775 49.690 112.745 ;
        RECT 49.860 112.455 50.310 112.915 ;
        RECT 50.480 112.625 51.575 113.185 ;
        RECT 49.860 112.235 50.985 112.455 ;
        RECT 49.860 111.605 50.185 112.065 ;
        RECT 50.705 111.775 50.985 112.235 ;
        RECT 51.175 111.775 51.575 112.625 ;
        RECT 51.745 113.355 52.700 113.525 ;
        RECT 52.990 113.390 53.445 114.155 ;
        RECT 53.720 113.775 55.020 113.985 ;
        RECT 55.275 113.795 55.605 114.155 ;
        RECT 54.850 113.625 55.020 113.775 ;
        RECT 55.775 113.655 56.035 113.985 ;
        RECT 55.805 113.645 56.035 113.655 ;
        RECT 51.745 112.455 51.955 113.355 ;
        RECT 52.125 112.625 52.815 113.185 ;
        RECT 53.920 113.165 54.140 113.565 ;
        RECT 52.985 112.965 53.475 113.165 ;
        RECT 53.665 112.955 54.140 113.165 ;
        RECT 54.385 113.165 54.595 113.565 ;
        RECT 54.850 113.500 55.605 113.625 ;
        RECT 54.850 113.455 55.695 113.500 ;
        RECT 55.425 113.335 55.695 113.455 ;
        RECT 54.385 112.955 54.715 113.165 ;
        RECT 54.885 112.895 55.295 113.200 ;
        RECT 52.990 112.725 54.165 112.785 ;
        RECT 55.525 112.760 55.695 113.335 ;
        RECT 55.495 112.725 55.695 112.760 ;
        RECT 52.990 112.615 55.695 112.725 ;
        RECT 51.745 112.235 52.700 112.455 ;
        RECT 51.975 111.605 52.245 112.065 ;
        RECT 52.415 111.775 52.700 112.235 ;
        RECT 52.990 111.995 53.245 112.615 ;
        RECT 53.835 112.555 55.635 112.615 ;
        RECT 53.835 112.525 54.165 112.555 ;
        RECT 55.865 112.455 56.035 113.645 ;
        RECT 57.125 113.430 57.415 114.155 ;
        RECT 57.630 113.695 57.895 114.155 ;
        RECT 58.265 113.515 58.435 113.985 ;
        RECT 58.685 113.695 58.855 114.155 ;
        RECT 59.105 113.515 59.275 113.985 ;
        RECT 59.525 113.695 59.695 114.155 ;
        RECT 59.945 113.515 60.115 113.985 ;
        RECT 60.285 113.690 60.535 114.155 ;
        RECT 58.265 113.335 60.635 113.515 ;
        RECT 60.855 113.500 61.185 113.935 ;
        RECT 61.355 113.545 61.525 114.155 ;
        RECT 57.605 112.915 60.115 113.165 ;
        RECT 53.495 112.355 53.680 112.445 ;
        RECT 54.270 112.355 55.105 112.365 ;
        RECT 53.495 112.155 55.105 112.355 ;
        RECT 53.495 112.115 53.725 112.155 ;
        RECT 52.990 111.775 53.325 111.995 ;
        RECT 54.330 111.605 54.685 111.985 ;
        RECT 54.855 111.775 55.105 112.155 ;
        RECT 55.355 111.605 55.605 112.385 ;
        RECT 55.775 111.775 56.035 112.455 ;
        RECT 57.125 111.605 57.415 112.770 ;
        RECT 60.285 112.745 60.635 113.335 ;
        RECT 57.630 111.605 57.925 112.745 ;
        RECT 58.185 112.575 60.635 112.745 ;
        RECT 60.805 113.415 61.185 113.500 ;
        RECT 61.695 113.415 62.025 113.940 ;
        RECT 62.285 113.625 62.495 114.155 ;
        RECT 62.770 113.705 63.555 113.875 ;
        RECT 63.725 113.705 64.130 113.875 ;
        RECT 60.805 113.375 61.030 113.415 ;
        RECT 60.805 112.795 60.975 113.375 ;
        RECT 61.695 113.245 61.895 113.415 ;
        RECT 62.770 113.245 62.940 113.705 ;
        RECT 61.145 112.915 61.895 113.245 ;
        RECT 62.065 112.915 62.940 113.245 ;
        RECT 60.805 112.745 61.020 112.795 ;
        RECT 60.805 112.665 61.195 112.745 ;
        RECT 58.185 111.775 58.515 112.575 ;
        RECT 58.685 111.605 58.855 112.405 ;
        RECT 59.025 111.775 59.355 112.575 ;
        RECT 59.865 112.555 60.635 112.575 ;
        RECT 59.525 111.605 59.695 112.405 ;
        RECT 59.865 111.775 60.195 112.555 ;
        RECT 60.365 111.605 60.535 112.065 ;
        RECT 60.865 111.820 61.195 112.665 ;
        RECT 61.705 112.710 61.895 112.915 ;
        RECT 61.365 111.605 61.535 112.615 ;
        RECT 61.705 112.335 62.600 112.710 ;
        RECT 61.705 111.775 62.045 112.335 ;
        RECT 62.275 111.605 62.590 112.105 ;
        RECT 62.770 112.075 62.940 112.915 ;
        RECT 63.110 113.205 63.575 113.535 ;
        RECT 63.960 113.475 64.130 113.705 ;
        RECT 64.310 113.655 64.680 114.155 ;
        RECT 65.000 113.705 65.675 113.875 ;
        RECT 65.870 113.705 66.205 113.875 ;
        RECT 63.110 112.245 63.430 113.205 ;
        RECT 63.960 113.175 64.790 113.475 ;
        RECT 63.600 112.275 63.790 112.995 ;
        RECT 63.960 112.105 64.130 113.175 ;
        RECT 64.590 113.145 64.790 113.175 ;
        RECT 64.300 112.925 64.470 112.995 ;
        RECT 65.000 112.925 65.170 113.705 ;
        RECT 66.035 113.565 66.205 113.705 ;
        RECT 66.375 113.695 66.625 114.155 ;
        RECT 64.300 112.755 65.170 112.925 ;
        RECT 65.340 113.285 65.865 113.505 ;
        RECT 66.035 113.435 66.260 113.565 ;
        RECT 64.300 112.665 64.810 112.755 ;
        RECT 62.770 111.905 63.655 112.075 ;
        RECT 63.880 111.775 64.130 112.105 ;
        RECT 64.300 111.605 64.470 112.405 ;
        RECT 64.640 112.050 64.810 112.665 ;
        RECT 65.340 112.585 65.510 113.285 ;
        RECT 64.980 112.220 65.510 112.585 ;
        RECT 65.680 112.520 65.920 113.115 ;
        RECT 66.090 112.330 66.260 113.435 ;
        RECT 66.430 112.575 66.710 113.525 ;
        RECT 65.955 112.200 66.260 112.330 ;
        RECT 64.640 111.880 65.745 112.050 ;
        RECT 65.955 111.775 66.205 112.200 ;
        RECT 66.375 111.605 66.640 112.065 ;
        RECT 66.880 111.775 67.065 113.895 ;
        RECT 67.235 113.775 67.565 114.155 ;
        RECT 67.735 113.605 67.905 113.895 ;
        RECT 67.240 113.435 67.905 113.605 ;
        RECT 67.240 112.445 67.470 113.435 ;
        RECT 68.165 113.355 68.860 113.985 ;
        RECT 69.065 113.355 69.375 114.155 ;
        RECT 69.635 113.605 69.805 113.895 ;
        RECT 69.975 113.775 70.305 114.155 ;
        RECT 69.635 113.435 70.300 113.605 ;
        RECT 68.685 113.305 68.860 113.355 ;
        RECT 67.640 112.615 67.990 113.265 ;
        RECT 68.185 112.915 68.520 113.165 ;
        RECT 68.690 112.755 68.860 113.305 ;
        RECT 69.030 112.915 69.365 113.185 ;
        RECT 67.240 112.275 67.905 112.445 ;
        RECT 67.235 111.605 67.565 112.105 ;
        RECT 67.735 111.775 67.905 112.275 ;
        RECT 68.165 111.605 68.425 112.745 ;
        RECT 68.595 111.775 68.925 112.755 ;
        RECT 69.095 111.605 69.375 112.745 ;
        RECT 69.550 112.615 69.900 113.265 ;
        RECT 70.070 112.445 70.300 113.435 ;
        RECT 69.635 112.275 70.300 112.445 ;
        RECT 69.635 111.775 69.805 112.275 ;
        RECT 69.975 111.605 70.305 112.105 ;
        RECT 70.475 111.775 70.660 113.895 ;
        RECT 70.915 113.695 71.165 114.155 ;
        RECT 71.335 113.705 71.670 113.875 ;
        RECT 71.865 113.705 72.540 113.875 ;
        RECT 71.335 113.565 71.505 113.705 ;
        RECT 70.830 112.575 71.110 113.525 ;
        RECT 71.280 113.435 71.505 113.565 ;
        RECT 71.280 112.330 71.450 113.435 ;
        RECT 71.675 113.285 72.200 113.505 ;
        RECT 71.620 112.520 71.860 113.115 ;
        RECT 72.030 112.585 72.200 113.285 ;
        RECT 72.370 112.925 72.540 113.705 ;
        RECT 72.860 113.655 73.230 114.155 ;
        RECT 73.410 113.705 73.815 113.875 ;
        RECT 73.985 113.705 74.770 113.875 ;
        RECT 73.410 113.475 73.580 113.705 ;
        RECT 72.750 113.175 73.580 113.475 ;
        RECT 73.965 113.205 74.430 113.535 ;
        RECT 72.750 113.145 72.950 113.175 ;
        RECT 73.070 112.925 73.240 112.995 ;
        RECT 72.370 112.755 73.240 112.925 ;
        RECT 72.730 112.665 73.240 112.755 ;
        RECT 71.280 112.200 71.585 112.330 ;
        RECT 72.030 112.220 72.560 112.585 ;
        RECT 70.900 111.605 71.165 112.065 ;
        RECT 71.335 111.775 71.585 112.200 ;
        RECT 72.730 112.050 72.900 112.665 ;
        RECT 71.795 111.880 72.900 112.050 ;
        RECT 73.070 111.605 73.240 112.405 ;
        RECT 73.410 112.105 73.580 113.175 ;
        RECT 73.750 112.275 73.940 112.995 ;
        RECT 74.110 112.245 74.430 113.205 ;
        RECT 74.600 113.245 74.770 113.705 ;
        RECT 75.045 113.625 75.255 114.155 ;
        RECT 75.515 113.415 75.845 113.940 ;
        RECT 76.015 113.545 76.185 114.155 ;
        RECT 76.355 113.500 76.685 113.935 ;
        RECT 76.355 113.415 76.735 113.500 ;
        RECT 75.645 113.245 75.845 113.415 ;
        RECT 76.510 113.375 76.735 113.415 ;
        RECT 74.600 112.915 75.475 113.245 ;
        RECT 75.645 112.915 76.395 113.245 ;
        RECT 73.410 111.775 73.660 112.105 ;
        RECT 74.600 112.075 74.770 112.915 ;
        RECT 75.645 112.710 75.835 112.915 ;
        RECT 76.565 112.795 76.735 113.375 ;
        RECT 76.520 112.745 76.735 112.795 ;
        RECT 74.940 112.335 75.835 112.710 ;
        RECT 76.345 112.665 76.735 112.745 ;
        RECT 76.940 113.415 77.555 113.985 ;
        RECT 77.725 113.645 77.940 114.155 ;
        RECT 78.170 113.645 78.450 113.975 ;
        RECT 78.630 113.645 78.870 114.155 ;
        RECT 79.370 113.645 79.610 114.155 ;
        RECT 79.790 113.645 80.070 113.975 ;
        RECT 80.300 113.645 80.515 114.155 ;
        RECT 73.885 111.905 74.770 112.075 ;
        RECT 74.950 111.605 75.265 112.105 ;
        RECT 75.495 111.775 75.835 112.335 ;
        RECT 76.005 111.605 76.175 112.615 ;
        RECT 76.345 111.820 76.675 112.665 ;
        RECT 76.940 112.395 77.255 113.415 ;
        RECT 77.425 112.745 77.595 113.245 ;
        RECT 77.845 112.915 78.110 113.475 ;
        RECT 78.280 112.745 78.450 113.645 ;
        RECT 78.620 112.915 78.975 113.475 ;
        RECT 79.265 112.915 79.620 113.475 ;
        RECT 79.790 112.745 79.960 113.645 ;
        RECT 80.130 112.915 80.395 113.475 ;
        RECT 80.685 113.415 81.300 113.985 ;
        RECT 80.645 112.745 80.815 113.245 ;
        RECT 77.425 112.575 78.850 112.745 ;
        RECT 76.940 111.775 77.475 112.395 ;
        RECT 77.645 111.605 77.975 112.405 ;
        RECT 78.460 112.400 78.850 112.575 ;
        RECT 79.390 112.575 80.815 112.745 ;
        RECT 79.390 112.400 79.780 112.575 ;
        RECT 80.265 111.605 80.595 112.405 ;
        RECT 80.985 112.395 81.300 113.415 ;
        RECT 81.965 113.405 83.175 114.155 ;
        RECT 80.765 111.775 81.300 112.395 ;
        RECT 81.965 112.695 82.485 113.235 ;
        RECT 82.655 112.865 83.175 113.405 ;
        RECT 81.965 111.605 83.175 112.695 ;
        RECT 5.520 111.435 83.260 111.605 ;
        RECT 5.605 110.345 6.815 111.435 ;
        RECT 6.985 111.000 12.330 111.435 ;
        RECT 5.605 109.635 6.125 110.175 ;
        RECT 6.295 109.805 6.815 110.345 ;
        RECT 5.605 108.885 6.815 109.635 ;
        RECT 8.570 109.430 8.910 110.260 ;
        RECT 10.390 109.750 10.740 111.000 ;
        RECT 12.505 110.345 15.095 111.435 ;
        RECT 15.265 110.925 15.565 111.435 ;
        RECT 15.735 110.755 16.065 111.265 ;
        RECT 16.235 110.925 16.865 111.435 ;
        RECT 17.445 110.925 17.825 111.095 ;
        RECT 17.995 110.925 18.295 111.435 ;
        RECT 17.655 110.755 17.825 110.925 ;
        RECT 12.505 109.655 13.715 110.175 ;
        RECT 13.885 109.825 15.095 110.345 ;
        RECT 15.265 110.585 17.485 110.755 ;
        RECT 6.985 108.885 12.330 109.430 ;
        RECT 12.505 108.885 15.095 109.655 ;
        RECT 15.265 109.625 15.435 110.585 ;
        RECT 15.605 110.245 17.145 110.415 ;
        RECT 15.605 109.795 15.850 110.245 ;
        RECT 16.110 109.875 16.805 110.075 ;
        RECT 16.975 110.045 17.145 110.245 ;
        RECT 17.315 110.385 17.485 110.585 ;
        RECT 17.655 110.555 18.315 110.755 ;
        RECT 17.315 110.215 17.975 110.385 ;
        RECT 16.975 109.875 17.575 110.045 ;
        RECT 17.805 109.795 17.975 110.215 ;
        RECT 15.265 109.080 15.730 109.625 ;
        RECT 16.235 108.885 16.405 109.705 ;
        RECT 16.575 109.625 17.485 109.705 ;
        RECT 18.145 109.625 18.315 110.555 ;
        RECT 18.485 110.270 18.775 111.435 ;
        RECT 19.955 110.425 20.125 111.265 ;
        RECT 20.295 111.095 21.465 111.265 ;
        RECT 20.295 110.595 20.625 111.095 ;
        RECT 21.135 111.055 21.465 111.095 ;
        RECT 21.655 111.015 22.010 111.435 ;
        RECT 20.795 110.835 21.025 110.925 ;
        RECT 22.180 110.835 22.430 111.265 ;
        RECT 20.795 110.595 22.430 110.835 ;
        RECT 22.600 110.675 22.930 111.435 ;
        RECT 23.100 110.595 23.355 111.265 ;
        RECT 24.175 110.635 24.430 111.435 ;
        RECT 19.955 110.255 23.015 110.425 ;
        RECT 19.870 109.875 20.220 110.085 ;
        RECT 20.390 109.875 20.835 110.075 ;
        RECT 21.005 109.875 21.480 110.075 ;
        RECT 16.575 109.535 17.825 109.625 ;
        RECT 16.575 109.055 16.905 109.535 ;
        RECT 17.315 109.455 17.825 109.535 ;
        RECT 17.075 108.885 17.425 109.275 ;
        RECT 17.595 109.055 17.825 109.455 ;
        RECT 17.995 109.145 18.315 109.625 ;
        RECT 18.485 108.885 18.775 109.610 ;
        RECT 19.955 109.535 21.020 109.705 ;
        RECT 19.955 109.055 20.125 109.535 ;
        RECT 20.295 108.885 20.625 109.365 ;
        RECT 20.850 109.305 21.020 109.535 ;
        RECT 21.200 109.475 21.480 109.875 ;
        RECT 21.750 109.875 22.080 110.075 ;
        RECT 22.250 109.905 22.625 110.075 ;
        RECT 22.250 109.875 22.615 109.905 ;
        RECT 21.750 109.475 22.035 109.875 ;
        RECT 22.845 109.705 23.015 110.255 ;
        RECT 22.215 109.535 23.015 109.705 ;
        RECT 22.215 109.305 22.385 109.535 ;
        RECT 23.185 109.465 23.355 110.595 ;
        RECT 24.600 110.465 24.930 111.265 ;
        RECT 25.100 110.635 25.270 111.435 ;
        RECT 25.440 110.465 25.770 111.265 ;
        RECT 25.940 110.635 26.110 111.435 ;
        RECT 26.280 110.465 26.610 111.265 ;
        RECT 26.780 110.635 26.950 111.435 ;
        RECT 27.120 110.465 27.450 111.265 ;
        RECT 27.620 110.635 27.920 111.435 ;
        RECT 24.005 110.295 27.975 110.465 ;
        RECT 28.155 110.325 28.450 111.435 ;
        RECT 24.005 109.705 24.350 110.295 ;
        RECT 24.600 109.875 27.455 110.125 ;
        RECT 27.655 109.705 27.975 110.295 ;
        RECT 28.630 110.125 28.880 111.260 ;
        RECT 29.050 110.325 29.310 111.435 ;
        RECT 29.480 110.535 29.740 111.260 ;
        RECT 29.910 110.705 30.170 111.435 ;
        RECT 30.340 110.535 30.600 111.260 ;
        RECT 30.770 110.705 31.030 111.435 ;
        RECT 31.200 110.535 31.460 111.260 ;
        RECT 31.630 110.705 31.890 111.435 ;
        RECT 32.060 110.535 32.320 111.260 ;
        RECT 32.490 110.705 32.785 111.435 ;
        RECT 29.480 110.295 32.790 110.535 ;
        RECT 33.205 110.295 33.485 111.435 ;
        RECT 24.005 109.515 27.975 109.705 ;
        RECT 28.145 109.515 28.460 110.125 ;
        RECT 28.630 109.875 31.650 110.125 ;
        RECT 23.170 109.395 23.355 109.465 ;
        RECT 23.145 109.385 23.355 109.395 ;
        RECT 20.850 109.055 22.385 109.305 ;
        RECT 22.555 108.885 22.885 109.365 ;
        RECT 23.100 109.055 23.355 109.385 ;
        RECT 24.175 108.885 24.430 109.345 ;
        RECT 24.600 109.055 24.930 109.515 ;
        RECT 25.100 108.885 25.270 109.345 ;
        RECT 25.440 109.055 25.770 109.515 ;
        RECT 25.940 108.885 26.110 109.345 ;
        RECT 26.280 109.055 26.610 109.515 ;
        RECT 26.780 108.885 26.950 109.345 ;
        RECT 27.120 109.055 27.450 109.515 ;
        RECT 27.620 108.885 27.925 109.345 ;
        RECT 28.205 108.885 28.450 109.345 ;
        RECT 28.630 109.065 28.880 109.875 ;
        RECT 31.820 109.705 32.790 110.295 ;
        RECT 33.655 110.285 33.985 111.265 ;
        RECT 34.155 110.295 34.415 111.435 ;
        RECT 34.675 110.765 34.845 111.265 ;
        RECT 35.015 110.935 35.345 111.435 ;
        RECT 34.675 110.595 35.340 110.765 ;
        RECT 33.215 109.855 33.550 110.125 ;
        RECT 29.480 109.535 32.790 109.705 ;
        RECT 33.720 109.685 33.890 110.285 ;
        RECT 34.060 109.875 34.395 110.125 ;
        RECT 34.590 109.775 34.940 110.425 ;
        RECT 29.050 108.885 29.310 109.410 ;
        RECT 29.480 109.080 29.740 109.535 ;
        RECT 29.910 108.885 30.170 109.365 ;
        RECT 30.340 109.080 30.600 109.535 ;
        RECT 30.770 108.885 31.030 109.365 ;
        RECT 31.200 109.080 31.460 109.535 ;
        RECT 31.630 108.885 31.890 109.365 ;
        RECT 32.060 109.080 32.320 109.535 ;
        RECT 32.490 108.885 32.790 109.365 ;
        RECT 33.205 108.885 33.515 109.685 ;
        RECT 33.720 109.055 34.415 109.685 ;
        RECT 35.110 109.605 35.340 110.595 ;
        RECT 34.675 109.435 35.340 109.605 ;
        RECT 34.675 109.145 34.845 109.435 ;
        RECT 35.015 108.885 35.345 109.265 ;
        RECT 35.515 109.145 35.700 111.265 ;
        RECT 35.940 110.975 36.205 111.435 ;
        RECT 36.375 110.840 36.625 111.265 ;
        RECT 36.835 110.990 37.940 111.160 ;
        RECT 36.320 110.710 36.625 110.840 ;
        RECT 35.870 109.515 36.150 110.465 ;
        RECT 36.320 109.605 36.490 110.710 ;
        RECT 36.660 109.925 36.900 110.520 ;
        RECT 37.070 110.455 37.600 110.820 ;
        RECT 37.070 109.755 37.240 110.455 ;
        RECT 37.770 110.375 37.940 110.990 ;
        RECT 38.110 110.635 38.280 111.435 ;
        RECT 38.450 110.935 38.700 111.265 ;
        RECT 38.925 110.965 39.810 111.135 ;
        RECT 37.770 110.285 38.280 110.375 ;
        RECT 36.320 109.475 36.545 109.605 ;
        RECT 36.715 109.535 37.240 109.755 ;
        RECT 37.410 110.115 38.280 110.285 ;
        RECT 35.955 108.885 36.205 109.345 ;
        RECT 36.375 109.335 36.545 109.475 ;
        RECT 37.410 109.335 37.580 110.115 ;
        RECT 38.110 110.045 38.280 110.115 ;
        RECT 37.790 109.865 37.990 109.895 ;
        RECT 38.450 109.865 38.620 110.935 ;
        RECT 38.790 110.045 38.980 110.765 ;
        RECT 37.790 109.565 38.620 109.865 ;
        RECT 39.150 109.835 39.470 110.795 ;
        RECT 36.375 109.165 36.710 109.335 ;
        RECT 36.905 109.165 37.580 109.335 ;
        RECT 37.900 108.885 38.270 109.385 ;
        RECT 38.450 109.335 38.620 109.565 ;
        RECT 39.005 109.505 39.470 109.835 ;
        RECT 39.640 110.125 39.810 110.965 ;
        RECT 39.990 110.935 40.305 111.435 ;
        RECT 40.535 110.705 40.875 111.265 ;
        RECT 39.980 110.330 40.875 110.705 ;
        RECT 41.045 110.425 41.215 111.435 ;
        RECT 40.685 110.125 40.875 110.330 ;
        RECT 41.385 110.375 41.715 111.220 ;
        RECT 41.385 110.295 41.775 110.375 ;
        RECT 41.945 110.345 43.615 111.435 ;
        RECT 41.560 110.245 41.775 110.295 ;
        RECT 39.640 109.795 40.515 110.125 ;
        RECT 40.685 109.795 41.435 110.125 ;
        RECT 39.640 109.335 39.810 109.795 ;
        RECT 40.685 109.625 40.885 109.795 ;
        RECT 41.605 109.665 41.775 110.245 ;
        RECT 41.550 109.625 41.775 109.665 ;
        RECT 38.450 109.165 38.855 109.335 ;
        RECT 39.025 109.165 39.810 109.335 ;
        RECT 40.085 108.885 40.295 109.415 ;
        RECT 40.555 109.100 40.885 109.625 ;
        RECT 41.395 109.540 41.775 109.625 ;
        RECT 41.945 109.655 42.695 110.175 ;
        RECT 42.865 109.825 43.615 110.345 ;
        RECT 44.245 110.270 44.535 111.435 ;
        RECT 44.710 110.295 45.045 111.265 ;
        RECT 45.215 110.295 45.385 111.435 ;
        RECT 45.555 111.095 47.585 111.265 ;
        RECT 41.055 108.885 41.225 109.495 ;
        RECT 41.395 109.105 41.725 109.540 ;
        RECT 41.945 108.885 43.615 109.655 ;
        RECT 44.710 109.625 44.880 110.295 ;
        RECT 45.555 110.125 45.725 111.095 ;
        RECT 45.050 109.795 45.305 110.125 ;
        RECT 45.530 109.795 45.725 110.125 ;
        RECT 45.895 110.755 47.020 110.925 ;
        RECT 45.135 109.625 45.305 109.795 ;
        RECT 45.895 109.625 46.065 110.755 ;
        RECT 44.245 108.885 44.535 109.610 ;
        RECT 44.710 109.055 44.965 109.625 ;
        RECT 45.135 109.455 46.065 109.625 ;
        RECT 46.235 110.415 47.245 110.585 ;
        RECT 46.235 109.615 46.405 110.415 ;
        RECT 45.890 109.420 46.065 109.455 ;
        RECT 45.135 108.885 45.465 109.285 ;
        RECT 45.890 109.055 46.420 109.420 ;
        RECT 46.610 109.395 46.885 110.215 ;
        RECT 46.605 109.225 46.885 109.395 ;
        RECT 46.610 109.055 46.885 109.225 ;
        RECT 47.055 109.055 47.245 110.415 ;
        RECT 47.415 110.430 47.585 111.095 ;
        RECT 47.755 110.675 47.925 111.435 ;
        RECT 48.160 110.675 48.675 111.085 ;
        RECT 47.415 110.240 48.165 110.430 ;
        RECT 48.335 109.865 48.675 110.675 ;
        RECT 48.885 110.485 49.175 111.255 ;
        RECT 49.745 110.895 50.005 111.255 ;
        RECT 50.175 111.065 50.505 111.435 ;
        RECT 50.675 110.895 50.935 111.255 ;
        RECT 49.745 110.665 50.935 110.895 ;
        RECT 51.125 110.715 51.455 111.435 ;
        RECT 51.625 110.485 51.890 111.255 ;
        RECT 52.725 110.765 53.005 111.435 ;
        RECT 53.175 110.545 53.475 111.095 ;
        RECT 53.675 110.715 54.005 111.435 ;
        RECT 54.195 110.715 54.655 111.265 ;
        RECT 48.885 110.305 51.380 110.485 ;
        RECT 47.445 109.695 48.675 109.865 ;
        RECT 48.855 109.795 49.125 110.125 ;
        RECT 49.305 109.795 49.740 110.125 ;
        RECT 49.920 109.795 50.495 110.125 ;
        RECT 50.675 109.795 50.955 110.125 ;
        RECT 47.425 108.885 47.935 109.420 ;
        RECT 48.155 109.090 48.400 109.695 ;
        RECT 51.155 109.615 51.380 110.305 ;
        RECT 48.895 109.425 51.380 109.615 ;
        RECT 48.895 109.065 49.120 109.425 ;
        RECT 49.300 108.885 49.630 109.255 ;
        RECT 49.810 109.065 50.065 109.425 ;
        RECT 50.630 108.885 51.375 109.255 ;
        RECT 51.555 109.065 51.890 110.485 ;
        RECT 52.540 110.125 52.805 110.485 ;
        RECT 53.175 110.375 54.115 110.545 ;
        RECT 53.945 110.125 54.115 110.375 ;
        RECT 52.540 109.875 53.215 110.125 ;
        RECT 53.435 109.875 53.775 110.125 ;
        RECT 53.945 109.795 54.235 110.125 ;
        RECT 53.945 109.705 54.115 109.795 ;
        RECT 52.725 109.515 54.115 109.705 ;
        RECT 52.725 109.155 53.055 109.515 ;
        RECT 54.405 109.345 54.655 110.715 ;
        RECT 54.835 110.325 55.130 111.435 ;
        RECT 55.310 110.125 55.560 111.260 ;
        RECT 55.730 110.325 55.990 111.435 ;
        RECT 56.160 110.535 56.420 111.260 ;
        RECT 56.590 110.705 56.850 111.435 ;
        RECT 57.020 110.535 57.280 111.260 ;
        RECT 57.450 110.705 57.710 111.435 ;
        RECT 57.880 110.535 58.140 111.260 ;
        RECT 58.310 110.705 58.570 111.435 ;
        RECT 58.740 110.535 59.000 111.260 ;
        RECT 59.170 110.705 59.465 111.435 ;
        RECT 56.160 110.295 59.470 110.535 ;
        RECT 54.825 109.515 55.140 110.125 ;
        RECT 55.310 109.875 58.330 110.125 ;
        RECT 53.675 108.885 53.925 109.345 ;
        RECT 54.095 109.055 54.655 109.345 ;
        RECT 54.885 108.885 55.130 109.345 ;
        RECT 55.310 109.065 55.560 109.875 ;
        RECT 58.500 109.705 59.470 110.295 ;
        RECT 56.160 109.535 59.470 109.705 ;
        RECT 59.895 110.375 60.225 111.225 ;
        RECT 59.895 109.610 60.085 110.375 ;
        RECT 60.395 110.295 60.645 111.435 ;
        RECT 60.835 110.795 61.085 111.215 ;
        RECT 61.315 110.965 61.645 111.435 ;
        RECT 61.875 110.795 62.125 111.215 ;
        RECT 60.835 110.625 62.125 110.795 ;
        RECT 62.305 110.795 62.635 111.225 ;
        RECT 62.305 110.625 62.760 110.795 ;
        RECT 60.825 110.125 61.040 110.455 ;
        RECT 60.255 109.795 60.565 110.125 ;
        RECT 60.735 109.795 61.040 110.125 ;
        RECT 61.215 109.795 61.500 110.455 ;
        RECT 61.695 109.795 61.960 110.455 ;
        RECT 62.175 109.795 62.420 110.455 ;
        RECT 60.395 109.625 60.565 109.795 ;
        RECT 62.590 109.625 62.760 110.625 ;
        RECT 64.025 110.675 64.540 111.085 ;
        RECT 64.775 110.675 64.945 111.435 ;
        RECT 65.115 111.095 67.145 111.265 ;
        RECT 64.025 109.865 64.365 110.675 ;
        RECT 65.115 110.430 65.285 111.095 ;
        RECT 65.680 110.755 66.805 110.925 ;
        RECT 64.535 110.240 65.285 110.430 ;
        RECT 65.455 110.415 66.465 110.585 ;
        RECT 64.025 109.695 65.255 109.865 ;
        RECT 55.730 108.885 55.990 109.410 ;
        RECT 56.160 109.080 56.420 109.535 ;
        RECT 56.590 108.885 56.850 109.365 ;
        RECT 57.020 109.080 57.280 109.535 ;
        RECT 57.450 108.885 57.710 109.365 ;
        RECT 57.880 109.080 58.140 109.535 ;
        RECT 58.310 108.885 58.570 109.365 ;
        RECT 58.740 109.080 59.000 109.535 ;
        RECT 59.170 108.885 59.470 109.365 ;
        RECT 59.895 109.100 60.225 109.610 ;
        RECT 60.395 109.455 62.760 109.625 ;
        RECT 60.395 108.885 60.725 109.285 ;
        RECT 61.775 109.115 62.105 109.455 ;
        RECT 62.275 108.885 62.605 109.285 ;
        RECT 64.300 109.090 64.545 109.695 ;
        RECT 64.765 108.885 65.275 109.420 ;
        RECT 65.455 109.055 65.645 110.415 ;
        RECT 65.815 110.075 66.090 110.215 ;
        RECT 65.815 109.905 66.095 110.075 ;
        RECT 65.815 109.055 66.090 109.905 ;
        RECT 66.295 109.615 66.465 110.415 ;
        RECT 66.635 109.625 66.805 110.755 ;
        RECT 66.975 110.125 67.145 111.095 ;
        RECT 67.315 110.295 67.485 111.435 ;
        RECT 67.655 110.295 67.990 111.265 ;
        RECT 66.975 109.795 67.170 110.125 ;
        RECT 67.395 109.795 67.650 110.125 ;
        RECT 67.395 109.625 67.565 109.795 ;
        RECT 67.820 109.625 67.990 110.295 ;
        RECT 68.170 110.285 68.430 111.435 ;
        RECT 68.605 110.360 68.860 111.265 ;
        RECT 69.030 110.675 69.360 111.435 ;
        RECT 69.575 110.505 69.745 111.265 ;
        RECT 66.635 109.455 67.565 109.625 ;
        RECT 66.635 109.420 66.810 109.455 ;
        RECT 66.280 109.055 66.810 109.420 ;
        RECT 67.235 108.885 67.565 109.285 ;
        RECT 67.735 109.055 67.990 109.625 ;
        RECT 68.170 108.885 68.430 109.725 ;
        RECT 68.605 109.630 68.775 110.360 ;
        RECT 69.030 110.335 69.745 110.505 ;
        RECT 69.030 110.125 69.200 110.335 ;
        RECT 70.005 110.270 70.295 111.435 ;
        RECT 70.475 110.325 70.770 111.435 ;
        RECT 68.945 109.795 69.200 110.125 ;
        RECT 68.605 109.055 68.860 109.630 ;
        RECT 69.030 109.605 69.200 109.795 ;
        RECT 69.480 109.785 69.835 110.155 ;
        RECT 70.950 110.125 71.200 111.260 ;
        RECT 71.370 110.325 71.630 111.435 ;
        RECT 71.800 110.535 72.060 111.260 ;
        RECT 72.230 110.705 72.490 111.435 ;
        RECT 72.660 110.535 72.920 111.260 ;
        RECT 73.090 110.705 73.350 111.435 ;
        RECT 73.520 110.535 73.780 111.260 ;
        RECT 73.950 110.705 74.210 111.435 ;
        RECT 74.380 110.535 74.640 111.260 ;
        RECT 74.810 110.705 75.105 111.435 ;
        RECT 71.800 110.295 75.110 110.535 ;
        RECT 69.030 109.435 69.745 109.605 ;
        RECT 69.030 108.885 69.360 109.265 ;
        RECT 69.575 109.055 69.745 109.435 ;
        RECT 70.005 108.885 70.295 109.610 ;
        RECT 70.465 109.515 70.780 110.125 ;
        RECT 70.950 109.875 73.970 110.125 ;
        RECT 70.525 108.885 70.770 109.345 ;
        RECT 70.950 109.065 71.200 109.875 ;
        RECT 74.140 109.705 75.110 110.295 ;
        RECT 75.530 110.285 75.790 111.435 ;
        RECT 75.965 110.360 76.220 111.265 ;
        RECT 76.390 110.675 76.720 111.435 ;
        RECT 76.935 110.505 77.105 111.265 ;
        RECT 71.800 109.535 75.110 109.705 ;
        RECT 71.370 108.885 71.630 109.410 ;
        RECT 71.800 109.080 72.060 109.535 ;
        RECT 72.230 108.885 72.490 109.365 ;
        RECT 72.660 109.080 72.920 109.535 ;
        RECT 73.090 108.885 73.350 109.365 ;
        RECT 73.520 109.080 73.780 109.535 ;
        RECT 73.950 108.885 74.210 109.365 ;
        RECT 74.380 109.080 74.640 109.535 ;
        RECT 74.810 108.885 75.110 109.365 ;
        RECT 75.530 108.885 75.790 109.725 ;
        RECT 75.965 109.630 76.135 110.360 ;
        RECT 76.390 110.335 77.105 110.505 ;
        RECT 78.375 110.505 78.545 111.265 ;
        RECT 78.760 110.675 79.090 111.435 ;
        RECT 78.375 110.335 79.090 110.505 ;
        RECT 79.260 110.360 79.515 111.265 ;
        RECT 76.390 110.125 76.560 110.335 ;
        RECT 76.305 109.795 76.560 110.125 ;
        RECT 75.965 109.055 76.220 109.630 ;
        RECT 76.390 109.605 76.560 109.795 ;
        RECT 76.840 109.785 77.195 110.155 ;
        RECT 78.285 109.785 78.640 110.155 ;
        RECT 78.920 110.125 79.090 110.335 ;
        RECT 78.920 109.795 79.175 110.125 ;
        RECT 78.920 109.605 79.090 109.795 ;
        RECT 79.345 109.630 79.515 110.360 ;
        RECT 79.690 110.285 79.950 111.435 ;
        RECT 80.215 110.505 80.385 111.265 ;
        RECT 80.600 110.675 80.930 111.435 ;
        RECT 80.215 110.335 80.930 110.505 ;
        RECT 81.100 110.360 81.355 111.265 ;
        RECT 80.125 109.785 80.480 110.155 ;
        RECT 80.760 110.125 80.930 110.335 ;
        RECT 80.760 109.795 81.015 110.125 ;
        RECT 76.390 109.435 77.105 109.605 ;
        RECT 76.390 108.885 76.720 109.265 ;
        RECT 76.935 109.055 77.105 109.435 ;
        RECT 78.375 109.435 79.090 109.605 ;
        RECT 78.375 109.055 78.545 109.435 ;
        RECT 78.760 108.885 79.090 109.265 ;
        RECT 79.260 109.055 79.515 109.630 ;
        RECT 79.690 108.885 79.950 109.725 ;
        RECT 80.760 109.605 80.930 109.795 ;
        RECT 81.185 109.630 81.355 110.360 ;
        RECT 81.530 110.285 81.790 111.435 ;
        RECT 81.965 110.345 83.175 111.435 ;
        RECT 81.965 109.805 82.485 110.345 ;
        RECT 80.215 109.435 80.930 109.605 ;
        RECT 80.215 109.055 80.385 109.435 ;
        RECT 80.600 108.885 80.930 109.265 ;
        RECT 81.100 109.055 81.355 109.630 ;
        RECT 81.530 108.885 81.790 109.725 ;
        RECT 82.655 109.635 83.175 110.175 ;
        RECT 81.965 108.885 83.175 109.635 ;
        RECT 5.520 108.715 83.260 108.885 ;
        RECT 5.605 107.965 6.815 108.715 ;
        RECT 7.075 108.165 7.245 108.545 ;
        RECT 7.425 108.335 7.755 108.715 ;
        RECT 7.075 107.995 7.740 108.165 ;
        RECT 7.935 108.040 8.195 108.545 ;
        RECT 8.365 108.170 13.710 108.715 ;
        RECT 5.605 107.425 6.125 107.965 ;
        RECT 6.295 107.255 6.815 107.795 ;
        RECT 7.005 107.445 7.345 107.815 ;
        RECT 7.570 107.740 7.740 107.995 ;
        RECT 7.570 107.410 7.845 107.740 ;
        RECT 7.570 107.265 7.740 107.410 ;
        RECT 5.605 106.165 6.815 107.255 ;
        RECT 7.065 107.095 7.740 107.265 ;
        RECT 8.015 107.240 8.195 108.040 ;
        RECT 9.950 107.340 10.290 108.170 ;
        RECT 14.355 107.905 14.625 108.715 ;
        RECT 14.795 107.905 15.125 108.545 ;
        RECT 15.295 107.905 15.535 108.715 ;
        RECT 16.190 107.950 16.645 108.715 ;
        RECT 16.920 108.335 18.220 108.545 ;
        RECT 18.475 108.355 18.805 108.715 ;
        RECT 18.050 108.185 18.220 108.335 ;
        RECT 18.975 108.215 19.235 108.545 ;
        RECT 7.065 106.335 7.245 107.095 ;
        RECT 7.425 106.165 7.755 106.925 ;
        RECT 7.925 106.335 8.195 107.240 ;
        RECT 11.770 106.600 12.120 107.850 ;
        RECT 14.345 107.475 14.695 107.725 ;
        RECT 14.865 107.305 15.035 107.905 ;
        RECT 17.120 107.725 17.340 108.125 ;
        RECT 15.205 107.475 15.555 107.725 ;
        RECT 16.185 107.525 16.675 107.725 ;
        RECT 16.865 107.515 17.340 107.725 ;
        RECT 17.585 107.725 17.795 108.125 ;
        RECT 18.050 108.060 18.805 108.185 ;
        RECT 18.050 108.015 18.895 108.060 ;
        RECT 18.625 107.895 18.895 108.015 ;
        RECT 17.585 107.515 17.915 107.725 ;
        RECT 18.085 107.455 18.495 107.760 ;
        RECT 8.365 106.165 13.710 106.600 ;
        RECT 14.355 106.165 14.685 107.305 ;
        RECT 14.865 107.135 15.545 107.305 ;
        RECT 15.215 106.350 15.545 107.135 ;
        RECT 16.190 107.285 17.365 107.345 ;
        RECT 18.725 107.320 18.895 107.895 ;
        RECT 18.695 107.285 18.895 107.320 ;
        RECT 16.190 107.175 18.895 107.285 ;
        RECT 16.190 106.555 16.445 107.175 ;
        RECT 17.035 107.115 18.835 107.175 ;
        RECT 17.035 107.085 17.365 107.115 ;
        RECT 19.065 107.015 19.235 108.215 ;
        RECT 16.695 106.915 16.880 107.005 ;
        RECT 17.470 106.915 18.305 106.925 ;
        RECT 16.695 106.715 18.305 106.915 ;
        RECT 16.695 106.675 16.925 106.715 ;
        RECT 16.190 106.335 16.525 106.555 ;
        RECT 17.530 106.165 17.885 106.545 ;
        RECT 18.055 106.335 18.305 106.715 ;
        RECT 18.555 106.165 18.805 106.945 ;
        RECT 18.975 106.335 19.235 107.015 ;
        RECT 19.410 107.115 19.745 108.535 ;
        RECT 19.925 108.345 20.670 108.715 ;
        RECT 21.235 108.175 21.490 108.535 ;
        RECT 21.670 108.345 22.000 108.715 ;
        RECT 22.180 108.175 22.405 108.535 ;
        RECT 19.920 107.985 22.405 108.175 ;
        RECT 19.920 107.295 20.145 107.985 ;
        RECT 22.660 107.975 23.275 108.545 ;
        RECT 23.445 108.205 23.660 108.715 ;
        RECT 23.890 108.205 24.170 108.535 ;
        RECT 24.350 108.205 24.590 108.715 ;
        RECT 20.345 107.475 20.625 107.805 ;
        RECT 20.805 107.475 21.380 107.805 ;
        RECT 21.560 107.475 21.995 107.805 ;
        RECT 22.175 107.475 22.445 107.805 ;
        RECT 19.920 107.115 22.415 107.295 ;
        RECT 19.410 106.345 19.675 107.115 ;
        RECT 19.845 106.165 20.175 106.885 ;
        RECT 20.365 106.705 21.555 106.935 ;
        RECT 20.365 106.345 20.625 106.705 ;
        RECT 20.795 106.165 21.125 106.535 ;
        RECT 21.295 106.345 21.555 106.705 ;
        RECT 22.125 106.345 22.415 107.115 ;
        RECT 22.660 106.955 22.975 107.975 ;
        RECT 23.145 107.305 23.315 107.805 ;
        RECT 23.565 107.475 23.830 108.035 ;
        RECT 24.000 107.305 24.170 108.205 ;
        RECT 25.010 108.145 25.185 108.545 ;
        RECT 25.355 108.335 25.685 108.715 ;
        RECT 25.930 108.215 26.160 108.545 ;
        RECT 24.340 107.475 24.695 108.035 ;
        RECT 25.010 107.975 25.640 108.145 ;
        RECT 25.470 107.805 25.640 107.975 ;
        RECT 23.145 107.135 24.570 107.305 ;
        RECT 22.660 106.335 23.195 106.955 ;
        RECT 23.365 106.165 23.695 106.965 ;
        RECT 24.180 106.960 24.570 107.135 ;
        RECT 24.925 107.125 25.290 107.805 ;
        RECT 25.470 107.475 25.820 107.805 ;
        RECT 25.470 106.955 25.640 107.475 ;
        RECT 25.010 106.785 25.640 106.955 ;
        RECT 25.990 106.925 26.160 108.215 ;
        RECT 26.360 107.105 26.640 108.380 ;
        RECT 26.865 108.375 27.135 108.380 ;
        RECT 26.825 108.205 27.135 108.375 ;
        RECT 27.595 108.335 27.925 108.715 ;
        RECT 28.095 108.460 28.430 108.505 ;
        RECT 26.865 107.105 27.135 108.205 ;
        RECT 27.325 107.105 27.665 108.135 ;
        RECT 28.095 107.995 28.435 108.460 ;
        RECT 27.835 107.475 28.095 107.805 ;
        RECT 27.835 106.925 28.005 107.475 ;
        RECT 28.265 107.305 28.435 107.995 ;
        RECT 25.010 106.335 25.185 106.785 ;
        RECT 25.990 106.755 28.005 106.925 ;
        RECT 25.355 106.165 25.685 106.605 ;
        RECT 25.990 106.335 26.160 106.755 ;
        RECT 26.395 106.165 27.065 106.575 ;
        RECT 27.280 106.335 27.450 106.755 ;
        RECT 27.650 106.165 27.980 106.575 ;
        RECT 28.175 106.335 28.435 107.305 ;
        RECT 28.615 106.345 28.875 108.535 ;
        RECT 29.135 108.345 29.805 108.715 ;
        RECT 29.985 108.165 30.295 108.535 ;
        RECT 29.065 107.965 30.295 108.165 ;
        RECT 29.065 107.295 29.355 107.965 ;
        RECT 30.475 107.785 30.705 108.425 ;
        RECT 30.885 107.985 31.175 108.715 ;
        RECT 31.365 107.990 31.655 108.715 ;
        RECT 31.830 108.315 32.165 108.715 ;
        RECT 32.335 108.145 32.540 108.545 ;
        RECT 32.750 108.235 33.025 108.715 ;
        RECT 33.235 108.215 33.495 108.545 ;
        RECT 31.855 107.975 32.540 108.145 ;
        RECT 29.535 107.475 30.000 107.785 ;
        RECT 30.180 107.475 30.705 107.785 ;
        RECT 30.885 107.475 31.185 107.805 ;
        RECT 29.065 107.075 29.835 107.295 ;
        RECT 29.045 106.165 29.385 106.895 ;
        RECT 29.565 106.345 29.835 107.075 ;
        RECT 30.015 107.055 31.175 107.295 ;
        RECT 30.015 106.345 30.245 107.055 ;
        RECT 30.415 106.165 30.745 106.875 ;
        RECT 30.915 106.345 31.175 107.055 ;
        RECT 31.365 106.165 31.655 107.330 ;
        RECT 31.855 106.945 32.195 107.975 ;
        RECT 32.365 107.305 32.615 107.805 ;
        RECT 32.795 107.475 33.155 108.055 ;
        RECT 33.325 107.305 33.495 108.215 ;
        RECT 34.700 108.085 34.985 108.545 ;
        RECT 35.155 108.255 35.425 108.715 ;
        RECT 34.700 107.915 35.655 108.085 ;
        RECT 32.365 107.135 33.495 107.305 ;
        RECT 34.585 107.185 35.275 107.745 ;
        RECT 31.855 106.770 32.520 106.945 ;
        RECT 31.830 106.165 32.165 106.590 ;
        RECT 32.335 106.365 32.520 106.770 ;
        RECT 32.725 106.165 33.055 106.945 ;
        RECT 33.225 106.365 33.495 107.135 ;
        RECT 35.445 107.015 35.655 107.915 ;
        RECT 34.700 106.795 35.655 107.015 ;
        RECT 35.825 107.745 36.225 108.545 ;
        RECT 36.415 108.085 36.695 108.545 ;
        RECT 37.215 108.255 37.540 108.715 ;
        RECT 36.415 107.915 37.540 108.085 ;
        RECT 37.710 107.975 38.095 108.545 ;
        RECT 37.090 107.805 37.540 107.915 ;
        RECT 35.825 107.185 36.920 107.745 ;
        RECT 37.090 107.475 37.645 107.805 ;
        RECT 34.700 106.335 34.985 106.795 ;
        RECT 35.155 106.165 35.425 106.625 ;
        RECT 35.825 106.335 36.225 107.185 ;
        RECT 37.090 107.015 37.540 107.475 ;
        RECT 37.815 107.305 38.095 107.975 ;
        RECT 38.285 107.905 38.525 108.715 ;
        RECT 38.695 107.905 39.025 108.545 ;
        RECT 39.195 107.905 39.465 108.715 ;
        RECT 39.645 107.965 40.855 108.715 ;
        RECT 41.085 108.255 41.330 108.715 ;
        RECT 38.265 107.475 38.615 107.725 ;
        RECT 38.785 107.305 38.955 107.905 ;
        RECT 39.125 107.475 39.475 107.725 ;
        RECT 39.645 107.425 40.165 107.965 ;
        RECT 36.415 106.795 37.540 107.015 ;
        RECT 36.415 106.335 36.695 106.795 ;
        RECT 37.215 106.165 37.540 106.625 ;
        RECT 37.710 106.335 38.095 107.305 ;
        RECT 38.275 107.135 38.955 107.305 ;
        RECT 38.275 106.350 38.605 107.135 ;
        RECT 39.135 106.165 39.465 107.305 ;
        RECT 40.335 107.255 40.855 107.795 ;
        RECT 41.025 107.475 41.340 108.085 ;
        RECT 41.510 107.725 41.760 108.535 ;
        RECT 41.930 108.190 42.190 108.715 ;
        RECT 42.360 108.065 42.620 108.520 ;
        RECT 42.790 108.235 43.050 108.715 ;
        RECT 43.220 108.065 43.480 108.520 ;
        RECT 43.650 108.235 43.910 108.715 ;
        RECT 44.080 108.065 44.340 108.520 ;
        RECT 44.510 108.235 44.770 108.715 ;
        RECT 44.940 108.065 45.200 108.520 ;
        RECT 45.370 108.235 45.670 108.715 ;
        RECT 42.360 107.895 45.670 108.065 ;
        RECT 41.510 107.475 44.530 107.725 ;
        RECT 39.645 106.165 40.855 107.255 ;
        RECT 41.035 106.165 41.330 107.275 ;
        RECT 41.510 106.340 41.760 107.475 ;
        RECT 44.700 107.305 45.670 107.895 ;
        RECT 46.085 107.965 47.295 108.715 ;
        RECT 47.555 108.165 47.725 108.455 ;
        RECT 47.895 108.335 48.225 108.715 ;
        RECT 47.555 107.995 48.220 108.165 ;
        RECT 46.085 107.425 46.605 107.965 ;
        RECT 41.930 106.165 42.190 107.275 ;
        RECT 42.360 107.065 45.670 107.305 ;
        RECT 46.775 107.255 47.295 107.795 ;
        RECT 42.360 106.340 42.620 107.065 ;
        RECT 42.790 106.165 43.050 106.895 ;
        RECT 43.220 106.340 43.480 107.065 ;
        RECT 43.650 106.165 43.910 106.895 ;
        RECT 44.080 106.340 44.340 107.065 ;
        RECT 44.510 106.165 44.770 106.895 ;
        RECT 44.940 106.340 45.200 107.065 ;
        RECT 45.370 106.165 45.665 106.895 ;
        RECT 46.085 106.165 47.295 107.255 ;
        RECT 47.470 107.175 47.820 107.825 ;
        RECT 47.990 107.005 48.220 107.995 ;
        RECT 47.555 106.835 48.220 107.005 ;
        RECT 47.555 106.335 47.725 106.835 ;
        RECT 47.895 106.165 48.225 106.665 ;
        RECT 48.395 106.335 48.580 108.455 ;
        RECT 48.835 108.255 49.085 108.715 ;
        RECT 49.255 108.265 49.590 108.435 ;
        RECT 49.785 108.265 50.460 108.435 ;
        RECT 49.255 108.125 49.425 108.265 ;
        RECT 48.750 107.135 49.030 108.085 ;
        RECT 49.200 107.995 49.425 108.125 ;
        RECT 49.200 106.890 49.370 107.995 ;
        RECT 49.595 107.845 50.120 108.065 ;
        RECT 49.540 107.080 49.780 107.675 ;
        RECT 49.950 107.145 50.120 107.845 ;
        RECT 50.290 107.485 50.460 108.265 ;
        RECT 50.780 108.215 51.150 108.715 ;
        RECT 51.330 108.265 51.735 108.435 ;
        RECT 51.905 108.265 52.690 108.435 ;
        RECT 51.330 108.035 51.500 108.265 ;
        RECT 50.670 107.735 51.500 108.035 ;
        RECT 51.885 107.765 52.350 108.095 ;
        RECT 50.670 107.705 50.870 107.735 ;
        RECT 50.990 107.485 51.160 107.555 ;
        RECT 50.290 107.315 51.160 107.485 ;
        RECT 50.650 107.225 51.160 107.315 ;
        RECT 49.200 106.760 49.505 106.890 ;
        RECT 49.950 106.780 50.480 107.145 ;
        RECT 48.820 106.165 49.085 106.625 ;
        RECT 49.255 106.335 49.505 106.760 ;
        RECT 50.650 106.610 50.820 107.225 ;
        RECT 49.715 106.440 50.820 106.610 ;
        RECT 50.990 106.165 51.160 106.965 ;
        RECT 51.330 106.665 51.500 107.735 ;
        RECT 51.670 106.835 51.860 107.555 ;
        RECT 52.030 106.805 52.350 107.765 ;
        RECT 52.520 107.805 52.690 108.265 ;
        RECT 52.965 108.185 53.175 108.715 ;
        RECT 53.435 107.975 53.765 108.500 ;
        RECT 53.935 108.105 54.105 108.715 ;
        RECT 54.275 108.060 54.605 108.495 ;
        RECT 54.840 108.145 55.095 108.495 ;
        RECT 55.265 108.315 55.595 108.715 ;
        RECT 55.765 108.145 55.935 108.495 ;
        RECT 56.105 108.315 56.485 108.715 ;
        RECT 54.275 107.975 54.655 108.060 ;
        RECT 54.840 107.975 56.505 108.145 ;
        RECT 56.675 108.040 56.950 108.385 ;
        RECT 53.565 107.805 53.765 107.975 ;
        RECT 54.430 107.935 54.655 107.975 ;
        RECT 52.520 107.475 53.395 107.805 ;
        RECT 53.565 107.475 54.315 107.805 ;
        RECT 51.330 106.335 51.580 106.665 ;
        RECT 52.520 106.635 52.690 107.475 ;
        RECT 53.565 107.270 53.755 107.475 ;
        RECT 54.485 107.355 54.655 107.935 ;
        RECT 56.335 107.805 56.505 107.975 ;
        RECT 54.825 107.475 55.170 107.805 ;
        RECT 55.340 107.475 56.165 107.805 ;
        RECT 56.335 107.475 56.610 107.805 ;
        RECT 54.440 107.305 54.655 107.355 ;
        RECT 52.860 106.895 53.755 107.270 ;
        RECT 54.265 107.225 54.655 107.305 ;
        RECT 51.805 106.465 52.690 106.635 ;
        RECT 52.870 106.165 53.185 106.665 ;
        RECT 53.415 106.335 53.755 106.895 ;
        RECT 53.925 106.165 54.095 107.175 ;
        RECT 54.265 106.380 54.595 107.225 ;
        RECT 54.845 107.015 55.170 107.305 ;
        RECT 55.340 107.185 55.535 107.475 ;
        RECT 56.335 107.305 56.505 107.475 ;
        RECT 56.780 107.305 56.950 108.040 ;
        RECT 57.125 107.990 57.415 108.715 ;
        RECT 57.745 108.155 58.075 108.545 ;
        RECT 58.245 108.325 59.430 108.495 ;
        RECT 59.690 108.245 59.860 108.715 ;
        RECT 57.745 107.975 58.255 108.155 ;
        RECT 57.585 107.515 57.915 107.805 ;
        RECT 58.085 107.345 58.255 107.975 ;
        RECT 58.660 108.065 59.045 108.155 ;
        RECT 60.030 108.065 60.360 108.530 ;
        RECT 58.660 107.895 60.360 108.065 ;
        RECT 60.530 107.895 60.700 108.715 ;
        RECT 60.870 107.895 61.555 108.535 ;
        RECT 61.815 108.165 61.985 108.455 ;
        RECT 62.155 108.335 62.485 108.715 ;
        RECT 61.815 107.995 62.480 108.165 ;
        RECT 58.425 107.515 58.755 107.725 ;
        RECT 58.935 107.475 59.315 107.725 ;
        RECT 55.845 107.135 56.505 107.305 ;
        RECT 55.845 107.015 56.015 107.135 ;
        RECT 54.845 106.845 56.015 107.015 ;
        RECT 54.825 106.385 56.015 106.675 ;
        RECT 56.185 106.165 56.465 106.965 ;
        RECT 56.675 106.335 56.950 107.305 ;
        RECT 57.125 106.165 57.415 107.330 ;
        RECT 57.740 107.175 58.825 107.345 ;
        RECT 57.740 106.335 58.040 107.175 ;
        RECT 58.235 106.165 58.485 107.005 ;
        RECT 58.655 106.925 58.825 107.175 ;
        RECT 58.995 107.095 59.315 107.475 ;
        RECT 59.505 107.515 59.990 107.725 ;
        RECT 60.180 107.515 60.630 107.725 ;
        RECT 60.800 107.515 61.135 107.725 ;
        RECT 59.505 107.355 59.880 107.515 ;
        RECT 59.485 107.185 59.880 107.355 ;
        RECT 60.800 107.345 60.970 107.515 ;
        RECT 59.505 107.095 59.880 107.185 ;
        RECT 60.050 107.175 60.970 107.345 ;
        RECT 60.050 106.925 60.220 107.175 ;
        RECT 58.655 106.755 60.220 106.925 ;
        RECT 59.075 106.335 59.880 106.755 ;
        RECT 60.390 106.165 60.720 107.005 ;
        RECT 61.305 106.925 61.555 107.895 ;
        RECT 61.730 107.175 62.080 107.825 ;
        RECT 62.250 107.005 62.480 107.995 ;
        RECT 60.890 106.335 61.555 106.925 ;
        RECT 61.815 106.835 62.480 107.005 ;
        RECT 61.815 106.335 61.985 106.835 ;
        RECT 62.155 106.165 62.485 106.665 ;
        RECT 62.655 106.335 62.840 108.455 ;
        RECT 63.095 108.255 63.345 108.715 ;
        RECT 63.515 108.265 63.850 108.435 ;
        RECT 64.045 108.265 64.720 108.435 ;
        RECT 63.515 108.125 63.685 108.265 ;
        RECT 63.010 107.135 63.290 108.085 ;
        RECT 63.460 107.995 63.685 108.125 ;
        RECT 63.460 106.890 63.630 107.995 ;
        RECT 63.855 107.845 64.380 108.065 ;
        RECT 63.800 107.080 64.040 107.675 ;
        RECT 64.210 107.145 64.380 107.845 ;
        RECT 64.550 107.485 64.720 108.265 ;
        RECT 65.040 108.215 65.410 108.715 ;
        RECT 65.590 108.265 65.995 108.435 ;
        RECT 66.165 108.265 66.950 108.435 ;
        RECT 65.590 108.035 65.760 108.265 ;
        RECT 64.930 107.735 65.760 108.035 ;
        RECT 66.145 107.765 66.610 108.095 ;
        RECT 64.930 107.705 65.130 107.735 ;
        RECT 65.250 107.485 65.420 107.555 ;
        RECT 64.550 107.315 65.420 107.485 ;
        RECT 64.910 107.225 65.420 107.315 ;
        RECT 63.460 106.760 63.765 106.890 ;
        RECT 64.210 106.780 64.740 107.145 ;
        RECT 63.080 106.165 63.345 106.625 ;
        RECT 63.515 106.335 63.765 106.760 ;
        RECT 64.910 106.610 65.080 107.225 ;
        RECT 63.975 106.440 65.080 106.610 ;
        RECT 65.250 106.165 65.420 106.965 ;
        RECT 65.590 106.665 65.760 107.735 ;
        RECT 65.930 106.835 66.120 107.555 ;
        RECT 66.290 106.805 66.610 107.765 ;
        RECT 66.780 107.805 66.950 108.265 ;
        RECT 67.225 108.185 67.435 108.715 ;
        RECT 67.695 107.975 68.025 108.500 ;
        RECT 68.195 108.105 68.365 108.715 ;
        RECT 68.535 108.060 68.865 108.495 ;
        RECT 68.535 107.975 68.915 108.060 ;
        RECT 67.825 107.805 68.025 107.975 ;
        RECT 68.690 107.935 68.915 107.975 ;
        RECT 66.780 107.475 67.655 107.805 ;
        RECT 67.825 107.475 68.575 107.805 ;
        RECT 65.590 106.335 65.840 106.665 ;
        RECT 66.780 106.635 66.950 107.475 ;
        RECT 67.825 107.270 68.015 107.475 ;
        RECT 68.745 107.355 68.915 107.935 ;
        RECT 68.700 107.305 68.915 107.355 ;
        RECT 67.120 106.895 68.015 107.270 ;
        RECT 68.525 107.225 68.915 107.305 ;
        RECT 69.085 107.975 69.470 108.545 ;
        RECT 69.640 108.255 69.965 108.715 ;
        RECT 70.485 108.085 70.765 108.545 ;
        RECT 69.085 107.305 69.365 107.975 ;
        RECT 69.640 107.915 70.765 108.085 ;
        RECT 69.640 107.805 70.090 107.915 ;
        RECT 69.535 107.475 70.090 107.805 ;
        RECT 70.955 107.745 71.355 108.545 ;
        RECT 71.755 108.255 72.025 108.715 ;
        RECT 72.195 108.085 72.480 108.545 ;
        RECT 66.065 106.465 66.950 106.635 ;
        RECT 67.130 106.165 67.445 106.665 ;
        RECT 67.675 106.335 68.015 106.895 ;
        RECT 68.185 106.165 68.355 107.175 ;
        RECT 68.525 106.380 68.855 107.225 ;
        RECT 69.085 106.335 69.470 107.305 ;
        RECT 69.640 107.015 70.090 107.475 ;
        RECT 70.260 107.185 71.355 107.745 ;
        RECT 69.640 106.795 70.765 107.015 ;
        RECT 69.640 106.165 69.965 106.625 ;
        RECT 70.485 106.335 70.765 106.795 ;
        RECT 70.955 106.335 71.355 107.185 ;
        RECT 71.525 107.915 72.480 108.085 ;
        RECT 72.765 107.915 73.105 108.545 ;
        RECT 73.275 107.915 73.525 108.715 ;
        RECT 73.715 108.065 74.045 108.545 ;
        RECT 74.215 108.255 74.440 108.715 ;
        RECT 74.610 108.065 74.940 108.545 ;
        RECT 71.525 107.015 71.735 107.915 ;
        RECT 71.905 107.185 72.595 107.745 ;
        RECT 72.765 107.305 72.940 107.915 ;
        RECT 73.715 107.895 74.940 108.065 ;
        RECT 75.570 107.935 76.070 108.545 ;
        RECT 76.535 108.165 76.705 108.545 ;
        RECT 76.885 108.335 77.215 108.715 ;
        RECT 76.535 107.995 77.200 108.165 ;
        RECT 77.395 108.040 77.655 108.545 ;
        RECT 73.110 107.555 73.805 107.725 ;
        RECT 73.635 107.305 73.805 107.555 ;
        RECT 73.980 107.525 74.400 107.725 ;
        RECT 74.570 107.525 74.900 107.725 ;
        RECT 75.070 107.525 75.400 107.725 ;
        RECT 75.570 107.305 75.740 107.935 ;
        RECT 75.925 107.475 76.275 107.725 ;
        RECT 76.465 107.445 76.795 107.815 ;
        RECT 77.030 107.740 77.200 107.995 ;
        RECT 77.030 107.410 77.315 107.740 ;
        RECT 71.525 106.795 72.480 107.015 ;
        RECT 71.755 106.165 72.025 106.625 ;
        RECT 72.195 106.335 72.480 106.795 ;
        RECT 72.765 106.335 73.105 107.305 ;
        RECT 73.275 106.165 73.445 107.305 ;
        RECT 73.635 107.135 76.070 107.305 ;
        RECT 77.030 107.265 77.200 107.410 ;
        RECT 73.715 106.165 73.965 106.965 ;
        RECT 74.610 106.335 74.940 107.135 ;
        RECT 75.240 106.165 75.570 106.965 ;
        RECT 75.740 106.335 76.070 107.135 ;
        RECT 76.535 107.095 77.200 107.265 ;
        RECT 77.485 107.240 77.655 108.040 ;
        RECT 76.535 106.335 76.705 107.095 ;
        RECT 76.885 106.165 77.215 106.925 ;
        RECT 77.385 106.335 77.655 107.240 ;
        RECT 77.860 107.975 78.475 108.545 ;
        RECT 78.645 108.205 78.860 108.715 ;
        RECT 79.090 108.205 79.370 108.535 ;
        RECT 79.550 108.205 79.790 108.715 ;
        RECT 77.860 106.955 78.175 107.975 ;
        RECT 78.345 107.305 78.515 107.805 ;
        RECT 78.765 107.475 79.030 108.035 ;
        RECT 79.200 107.305 79.370 108.205 ;
        RECT 80.215 108.165 80.385 108.545 ;
        RECT 80.600 108.335 80.930 108.715 ;
        RECT 79.540 107.475 79.895 108.035 ;
        RECT 80.215 107.995 80.930 108.165 ;
        RECT 80.125 107.445 80.480 107.815 ;
        RECT 80.760 107.805 80.930 107.995 ;
        RECT 81.100 107.970 81.355 108.545 ;
        RECT 80.760 107.475 81.015 107.805 ;
        RECT 78.345 107.135 79.770 107.305 ;
        RECT 80.760 107.265 80.930 107.475 ;
        RECT 77.860 106.335 78.395 106.955 ;
        RECT 78.565 106.165 78.895 106.965 ;
        RECT 79.380 106.960 79.770 107.135 ;
        RECT 80.215 107.095 80.930 107.265 ;
        RECT 81.185 107.240 81.355 107.970 ;
        RECT 81.530 107.875 81.790 108.715 ;
        RECT 81.965 107.965 83.175 108.715 ;
        RECT 80.215 106.335 80.385 107.095 ;
        RECT 80.600 106.165 80.930 106.925 ;
        RECT 81.100 106.335 81.355 107.240 ;
        RECT 81.530 106.165 81.790 107.315 ;
        RECT 81.965 107.255 82.485 107.795 ;
        RECT 82.655 107.425 83.175 107.965 ;
        RECT 81.965 106.165 83.175 107.255 ;
        RECT 5.520 105.995 83.260 106.165 ;
        RECT 5.605 104.905 6.815 105.995 ;
        RECT 5.605 104.195 6.125 104.735 ;
        RECT 6.295 104.365 6.815 104.905 ;
        RECT 5.605 103.445 6.815 104.195 ;
        RECT 7.445 103.615 7.705 105.825 ;
        RECT 7.875 105.615 8.205 105.995 ;
        RECT 8.630 105.445 8.800 105.825 ;
        RECT 9.060 105.615 9.390 105.995 ;
        RECT 9.585 105.445 9.755 105.825 ;
        RECT 9.965 105.615 10.295 105.995 ;
        RECT 10.545 105.445 10.735 105.825 ;
        RECT 10.975 105.615 11.305 105.995 ;
        RECT 11.615 105.495 11.875 105.825 ;
        RECT 7.875 105.275 9.825 105.445 ;
        RECT 7.875 104.355 8.045 105.275 ;
        RECT 8.415 104.685 8.610 104.995 ;
        RECT 8.880 104.685 9.065 104.995 ;
        RECT 8.355 104.355 8.610 104.685 ;
        RECT 8.835 104.355 9.065 104.685 ;
        RECT 7.875 103.445 8.205 103.825 ;
        RECT 8.415 103.780 8.610 104.355 ;
        RECT 8.880 103.775 9.065 104.355 ;
        RECT 9.315 103.785 9.485 104.685 ;
        RECT 9.655 104.285 9.825 105.275 ;
        RECT 9.995 105.275 10.735 105.445 ;
        RECT 9.995 104.765 10.165 105.275 ;
        RECT 10.335 104.935 10.915 105.105 ;
        RECT 11.185 104.985 11.535 105.315 ;
        RECT 10.745 104.815 10.915 104.935 ;
        RECT 11.705 104.815 11.875 105.495 ;
        RECT 9.995 104.595 10.565 104.765 ;
        RECT 10.745 104.645 11.875 104.815 ;
        RECT 9.655 103.955 10.205 104.285 ;
        RECT 10.395 104.115 10.565 104.595 ;
        RECT 10.735 104.305 11.355 104.475 ;
        RECT 11.145 104.125 11.355 104.305 ;
        RECT 10.395 103.785 10.795 104.115 ;
        RECT 11.705 103.945 11.875 104.645 ;
        RECT 9.315 103.615 10.795 103.785 ;
        RECT 10.975 103.445 11.305 103.825 ;
        RECT 11.615 103.615 11.875 103.945 ;
        RECT 12.045 104.855 12.305 105.825 ;
        RECT 12.500 105.585 12.830 105.995 ;
        RECT 13.030 105.405 13.200 105.825 ;
        RECT 13.415 105.585 14.085 105.995 ;
        RECT 14.320 105.405 14.490 105.825 ;
        RECT 14.795 105.555 15.125 105.995 ;
        RECT 12.475 105.235 14.490 105.405 ;
        RECT 15.295 105.375 15.470 105.825 ;
        RECT 12.045 104.165 12.215 104.855 ;
        RECT 12.475 104.685 12.645 105.235 ;
        RECT 12.385 104.355 12.645 104.685 ;
        RECT 12.045 103.700 12.385 104.165 ;
        RECT 12.815 104.025 13.155 105.055 ;
        RECT 13.345 104.975 13.615 105.055 ;
        RECT 13.345 104.805 13.655 104.975 ;
        RECT 12.050 103.655 12.385 103.700 ;
        RECT 12.555 103.445 12.885 103.825 ;
        RECT 13.345 103.780 13.615 104.805 ;
        RECT 13.840 103.780 14.120 105.055 ;
        RECT 14.320 103.945 14.490 105.235 ;
        RECT 14.840 105.205 15.470 105.375 ;
        RECT 14.840 104.685 15.010 105.205 ;
        RECT 16.220 105.195 16.470 105.995 ;
        RECT 16.640 105.365 16.970 105.825 ;
        RECT 17.140 105.535 17.355 105.995 ;
        RECT 16.640 105.195 17.810 105.365 ;
        RECT 14.660 104.355 15.010 104.685 ;
        RECT 15.190 104.355 15.555 105.035 ;
        RECT 15.730 105.025 16.010 105.185 ;
        RECT 15.730 104.855 17.065 105.025 ;
        RECT 16.895 104.685 17.065 104.855 ;
        RECT 15.730 104.435 16.080 104.675 ;
        RECT 16.250 104.435 16.725 104.675 ;
        RECT 16.895 104.435 17.270 104.685 ;
        RECT 14.840 104.185 15.010 104.355 ;
        RECT 16.895 104.265 17.065 104.435 ;
        RECT 14.840 104.015 15.470 104.185 ;
        RECT 14.320 103.615 14.550 103.945 ;
        RECT 14.795 103.445 15.125 103.825 ;
        RECT 15.295 103.615 15.470 104.015 ;
        RECT 15.730 104.095 17.065 104.265 ;
        RECT 15.730 103.885 16.000 104.095 ;
        RECT 17.440 103.905 17.810 105.195 ;
        RECT 18.485 104.830 18.775 105.995 ;
        RECT 18.945 105.155 19.205 105.825 ;
        RECT 19.375 105.595 19.705 105.995 ;
        RECT 20.575 105.595 20.975 105.995 ;
        RECT 21.265 105.415 21.595 105.650 ;
        RECT 19.515 105.245 21.595 105.415 ;
        RECT 18.945 104.185 19.120 105.155 ;
        RECT 19.515 104.975 19.685 105.245 ;
        RECT 19.290 104.805 19.685 104.975 ;
        RECT 19.855 104.855 20.870 105.075 ;
        RECT 19.290 104.355 19.460 104.805 ;
        RECT 20.595 104.715 20.870 104.855 ;
        RECT 21.040 104.855 21.595 105.245 ;
        RECT 19.630 104.435 20.080 104.635 ;
        RECT 20.250 104.265 20.425 104.460 ;
        RECT 16.220 103.445 16.550 103.905 ;
        RECT 17.060 103.615 17.810 103.905 ;
        RECT 18.485 103.445 18.775 104.170 ;
        RECT 18.945 103.615 19.285 104.185 ;
        RECT 19.480 103.445 19.650 104.110 ;
        RECT 19.930 104.095 20.425 104.265 ;
        RECT 19.930 103.955 20.150 104.095 ;
        RECT 19.925 103.785 20.150 103.955 ;
        RECT 20.595 103.925 20.765 104.715 ;
        RECT 21.040 104.605 21.210 104.855 ;
        RECT 21.765 104.685 21.940 105.785 ;
        RECT 22.110 105.175 22.455 105.995 ;
        RECT 22.625 105.400 23.060 105.825 ;
        RECT 23.230 105.570 23.615 105.995 ;
        RECT 22.625 105.230 23.615 105.400 ;
        RECT 21.015 104.435 21.210 104.605 ;
        RECT 21.380 104.435 21.940 104.685 ;
        RECT 22.110 104.435 22.455 105.005 ;
        RECT 21.015 104.050 21.185 104.435 ;
        RECT 22.625 104.355 23.110 105.060 ;
        RECT 23.280 104.685 23.615 105.230 ;
        RECT 23.785 105.035 24.210 105.825 ;
        RECT 24.380 105.400 24.655 105.825 ;
        RECT 24.825 105.570 25.210 105.995 ;
        RECT 24.380 105.205 25.210 105.400 ;
        RECT 23.785 104.855 24.690 105.035 ;
        RECT 23.280 104.355 23.690 104.685 ;
        RECT 23.860 104.355 24.690 104.855 ;
        RECT 24.860 104.685 25.210 105.205 ;
        RECT 25.380 105.035 25.625 105.825 ;
        RECT 25.815 105.400 26.070 105.825 ;
        RECT 26.240 105.570 26.625 105.995 ;
        RECT 25.815 105.205 26.625 105.400 ;
        RECT 25.380 104.855 26.105 105.035 ;
        RECT 24.860 104.355 25.285 104.685 ;
        RECT 25.455 104.355 26.105 104.855 ;
        RECT 26.275 104.685 26.625 105.205 ;
        RECT 26.795 104.855 27.055 105.825 ;
        RECT 27.770 105.375 27.945 105.825 ;
        RECT 28.115 105.555 28.445 105.995 ;
        RECT 28.750 105.405 28.920 105.825 ;
        RECT 29.155 105.585 29.825 105.995 ;
        RECT 30.040 105.405 30.210 105.825 ;
        RECT 30.410 105.585 30.740 105.995 ;
        RECT 27.770 105.205 28.400 105.375 ;
        RECT 26.275 104.355 26.700 104.685 ;
        RECT 19.930 103.740 20.150 103.785 ;
        RECT 20.320 103.755 20.765 103.925 ;
        RECT 20.935 103.680 21.185 104.050 ;
        RECT 21.355 104.085 22.455 104.265 ;
        RECT 23.280 104.185 23.615 104.355 ;
        RECT 23.860 104.185 24.210 104.355 ;
        RECT 24.860 104.185 25.210 104.355 ;
        RECT 25.455 104.185 25.625 104.355 ;
        RECT 26.275 104.185 26.625 104.355 ;
        RECT 26.870 104.185 27.055 104.855 ;
        RECT 27.685 104.355 28.050 105.035 ;
        RECT 28.230 104.685 28.400 105.205 ;
        RECT 28.750 105.235 30.765 105.405 ;
        RECT 28.230 104.355 28.580 104.685 ;
        RECT 28.230 104.185 28.400 104.355 ;
        RECT 21.355 103.680 21.605 104.085 ;
        RECT 21.775 103.445 21.945 103.915 ;
        RECT 22.115 103.680 22.455 104.085 ;
        RECT 22.625 104.015 23.615 104.185 ;
        RECT 22.625 103.615 23.060 104.015 ;
        RECT 23.230 103.445 23.615 103.845 ;
        RECT 23.785 103.615 24.210 104.185 ;
        RECT 24.400 104.015 25.210 104.185 ;
        RECT 24.400 103.615 24.655 104.015 ;
        RECT 24.825 103.445 25.210 103.845 ;
        RECT 25.380 103.615 25.625 104.185 ;
        RECT 25.815 104.015 26.625 104.185 ;
        RECT 25.815 103.615 26.070 104.015 ;
        RECT 26.240 103.445 26.625 103.845 ;
        RECT 26.795 103.615 27.055 104.185 ;
        RECT 27.770 104.015 28.400 104.185 ;
        RECT 27.770 103.615 27.945 104.015 ;
        RECT 28.750 103.945 28.920 105.235 ;
        RECT 28.115 103.445 28.445 103.825 ;
        RECT 28.690 103.615 28.920 103.945 ;
        RECT 29.120 103.780 29.400 105.055 ;
        RECT 29.625 104.295 29.895 105.055 ;
        RECT 29.585 104.125 29.895 104.295 ;
        RECT 29.625 103.780 29.895 104.125 ;
        RECT 30.085 104.025 30.425 105.055 ;
        RECT 30.595 104.685 30.765 105.235 ;
        RECT 30.935 104.855 31.195 105.825 ;
        RECT 31.385 105.485 31.685 105.995 ;
        RECT 31.855 105.485 32.235 105.655 ;
        RECT 32.815 105.485 33.445 105.995 ;
        RECT 31.855 105.315 32.025 105.485 ;
        RECT 33.615 105.315 33.945 105.825 ;
        RECT 34.115 105.485 34.415 105.995 ;
        RECT 34.675 105.325 34.845 105.825 ;
        RECT 35.015 105.495 35.345 105.995 ;
        RECT 30.595 104.355 30.855 104.685 ;
        RECT 31.025 104.165 31.195 104.855 ;
        RECT 30.355 103.445 30.685 103.825 ;
        RECT 30.855 103.700 31.195 104.165 ;
        RECT 31.365 105.115 32.025 105.315 ;
        RECT 32.195 105.145 34.415 105.315 ;
        RECT 34.675 105.155 35.340 105.325 ;
        RECT 31.365 104.185 31.535 105.115 ;
        RECT 32.195 104.945 32.365 105.145 ;
        RECT 31.705 104.775 32.365 104.945 ;
        RECT 32.535 104.805 34.075 104.975 ;
        RECT 31.705 104.355 31.875 104.775 ;
        RECT 32.535 104.605 32.705 104.805 ;
        RECT 32.105 104.435 32.705 104.605 ;
        RECT 32.875 104.435 33.570 104.635 ;
        RECT 33.830 104.355 34.075 104.805 ;
        RECT 32.195 104.185 33.105 104.265 ;
        RECT 31.365 103.705 31.685 104.185 ;
        RECT 31.855 104.095 33.105 104.185 ;
        RECT 31.855 104.015 32.365 104.095 ;
        RECT 30.855 103.655 31.190 103.700 ;
        RECT 31.855 103.615 32.085 104.015 ;
        RECT 32.255 103.445 32.605 103.835 ;
        RECT 32.775 103.615 33.105 104.095 ;
        RECT 33.275 103.445 33.445 104.265 ;
        RECT 34.245 104.185 34.415 105.145 ;
        RECT 34.590 104.335 34.940 104.985 ;
        RECT 33.950 103.640 34.415 104.185 ;
        RECT 35.110 104.165 35.340 105.155 ;
        RECT 34.675 103.995 35.340 104.165 ;
        RECT 34.675 103.705 34.845 103.995 ;
        RECT 35.015 103.445 35.345 103.825 ;
        RECT 35.515 103.705 35.700 105.825 ;
        RECT 35.940 105.535 36.205 105.995 ;
        RECT 36.375 105.400 36.625 105.825 ;
        RECT 36.835 105.550 37.940 105.720 ;
        RECT 36.320 105.270 36.625 105.400 ;
        RECT 35.870 104.075 36.150 105.025 ;
        RECT 36.320 104.165 36.490 105.270 ;
        RECT 36.660 104.485 36.900 105.080 ;
        RECT 37.070 105.015 37.600 105.380 ;
        RECT 37.070 104.315 37.240 105.015 ;
        RECT 37.770 104.935 37.940 105.550 ;
        RECT 38.110 105.195 38.280 105.995 ;
        RECT 38.450 105.495 38.700 105.825 ;
        RECT 38.925 105.525 39.810 105.695 ;
        RECT 37.770 104.845 38.280 104.935 ;
        RECT 36.320 104.035 36.545 104.165 ;
        RECT 36.715 104.095 37.240 104.315 ;
        RECT 37.410 104.675 38.280 104.845 ;
        RECT 35.955 103.445 36.205 103.905 ;
        RECT 36.375 103.895 36.545 104.035 ;
        RECT 37.410 103.895 37.580 104.675 ;
        RECT 38.110 104.605 38.280 104.675 ;
        RECT 37.790 104.425 37.990 104.455 ;
        RECT 38.450 104.425 38.620 105.495 ;
        RECT 38.790 104.605 38.980 105.325 ;
        RECT 37.790 104.125 38.620 104.425 ;
        RECT 39.150 104.395 39.470 105.355 ;
        RECT 36.375 103.725 36.710 103.895 ;
        RECT 36.905 103.725 37.580 103.895 ;
        RECT 37.900 103.445 38.270 103.945 ;
        RECT 38.450 103.895 38.620 104.125 ;
        RECT 39.005 104.065 39.470 104.395 ;
        RECT 39.640 104.685 39.810 105.525 ;
        RECT 39.990 105.495 40.305 105.995 ;
        RECT 40.535 105.265 40.875 105.825 ;
        RECT 39.980 104.890 40.875 105.265 ;
        RECT 41.045 104.985 41.215 105.995 ;
        RECT 40.685 104.685 40.875 104.890 ;
        RECT 41.385 104.935 41.715 105.780 ;
        RECT 41.385 104.855 41.775 104.935 ;
        RECT 41.945 104.905 43.615 105.995 ;
        RECT 41.560 104.805 41.775 104.855 ;
        RECT 39.640 104.355 40.515 104.685 ;
        RECT 40.685 104.355 41.435 104.685 ;
        RECT 39.640 103.895 39.810 104.355 ;
        RECT 40.685 104.185 40.885 104.355 ;
        RECT 41.605 104.225 41.775 104.805 ;
        RECT 41.550 104.185 41.775 104.225 ;
        RECT 38.450 103.725 38.855 103.895 ;
        RECT 39.025 103.725 39.810 103.895 ;
        RECT 40.085 103.445 40.295 103.975 ;
        RECT 40.555 103.660 40.885 104.185 ;
        RECT 41.395 104.100 41.775 104.185 ;
        RECT 41.945 104.215 42.695 104.735 ;
        RECT 42.865 104.385 43.615 104.905 ;
        RECT 44.245 104.830 44.535 105.995 ;
        RECT 44.750 104.855 45.045 105.995 ;
        RECT 45.305 105.025 45.635 105.825 ;
        RECT 45.805 105.195 45.975 105.995 ;
        RECT 46.145 105.025 46.475 105.825 ;
        RECT 46.645 105.195 46.815 105.995 ;
        RECT 46.985 105.045 47.315 105.825 ;
        RECT 47.485 105.535 47.655 105.995 ;
        RECT 48.845 105.195 49.285 105.825 ;
        RECT 46.985 105.025 47.755 105.045 ;
        RECT 45.305 104.855 47.755 105.025 ;
        RECT 44.725 104.435 47.235 104.685 ;
        RECT 47.405 104.265 47.755 104.855 ;
        RECT 41.055 103.445 41.225 104.055 ;
        RECT 41.395 103.665 41.725 104.100 ;
        RECT 41.945 103.445 43.615 104.215 ;
        RECT 44.245 103.445 44.535 104.170 ;
        RECT 45.385 104.085 47.755 104.265 ;
        RECT 48.845 104.185 49.155 105.195 ;
        RECT 49.460 105.145 49.775 105.995 ;
        RECT 49.945 105.655 51.375 105.825 ;
        RECT 49.945 104.975 50.115 105.655 ;
        RECT 49.325 104.805 50.115 104.975 ;
        RECT 49.325 104.355 49.495 104.805 ;
        RECT 50.285 104.685 50.485 105.485 ;
        RECT 49.665 104.355 50.055 104.635 ;
        RECT 50.240 104.355 50.485 104.685 ;
        RECT 50.685 104.355 50.935 105.485 ;
        RECT 51.125 105.025 51.375 105.655 ;
        RECT 51.555 105.195 51.885 105.995 ;
        RECT 52.075 105.025 52.405 105.810 ;
        RECT 51.125 104.855 51.895 105.025 ;
        RECT 52.075 104.855 52.755 105.025 ;
        RECT 52.935 104.855 53.265 105.995 ;
        RECT 53.445 104.855 53.705 105.995 ;
        RECT 51.150 104.355 51.555 104.685 ;
        RECT 51.725 104.185 51.895 104.855 ;
        RECT 52.065 104.435 52.415 104.685 ;
        RECT 52.585 104.255 52.755 104.855 ;
        RECT 53.875 104.845 54.205 105.825 ;
        RECT 54.375 104.855 54.655 105.995 ;
        RECT 54.940 105.365 55.225 105.825 ;
        RECT 55.395 105.535 55.665 105.995 ;
        RECT 54.940 105.145 55.895 105.365 ;
        RECT 52.925 104.435 53.275 104.685 ;
        RECT 53.465 104.435 53.800 104.685 ;
        RECT 44.750 103.445 45.015 103.905 ;
        RECT 45.385 103.615 45.555 104.085 ;
        RECT 45.805 103.445 45.975 103.905 ;
        RECT 46.225 103.615 46.395 104.085 ;
        RECT 46.645 103.445 46.815 103.905 ;
        RECT 47.065 103.615 47.235 104.085 ;
        RECT 47.405 103.445 47.655 103.910 ;
        RECT 48.845 103.625 49.285 104.185 ;
        RECT 49.455 103.445 49.905 104.185 ;
        RECT 50.075 104.015 51.235 104.185 ;
        RECT 50.075 103.615 50.245 104.015 ;
        RECT 50.415 103.445 50.835 103.845 ;
        RECT 51.005 103.615 51.235 104.015 ;
        RECT 51.405 103.615 51.895 104.185 ;
        RECT 52.085 103.445 52.325 104.255 ;
        RECT 52.495 103.615 52.825 104.255 ;
        RECT 52.995 103.445 53.265 104.255 ;
        RECT 53.970 104.245 54.140 104.845 ;
        RECT 54.310 104.415 54.645 104.685 ;
        RECT 54.825 104.415 55.515 104.975 ;
        RECT 55.685 104.245 55.895 105.145 ;
        RECT 53.445 103.615 54.140 104.245 ;
        RECT 54.345 103.445 54.655 104.245 ;
        RECT 54.940 104.075 55.895 104.245 ;
        RECT 56.065 104.975 56.465 105.825 ;
        RECT 56.655 105.365 56.935 105.825 ;
        RECT 57.455 105.535 57.780 105.995 ;
        RECT 56.655 105.145 57.780 105.365 ;
        RECT 56.065 104.415 57.160 104.975 ;
        RECT 57.330 104.685 57.780 105.145 ;
        RECT 57.950 104.855 58.335 105.825 ;
        RECT 58.710 105.025 59.040 105.825 ;
        RECT 59.210 105.195 59.540 105.995 ;
        RECT 59.840 105.025 60.170 105.825 ;
        RECT 60.815 105.195 61.065 105.995 ;
        RECT 58.710 104.855 61.145 105.025 ;
        RECT 61.335 104.855 61.505 105.995 ;
        RECT 61.675 104.855 62.015 105.825 ;
        RECT 62.185 104.855 62.465 105.995 ;
        RECT 54.940 103.615 55.225 104.075 ;
        RECT 55.395 103.445 55.665 103.905 ;
        RECT 56.065 103.615 56.465 104.415 ;
        RECT 57.330 104.355 57.885 104.685 ;
        RECT 57.330 104.245 57.780 104.355 ;
        RECT 56.655 104.075 57.780 104.245 ;
        RECT 58.055 104.185 58.335 104.855 ;
        RECT 58.505 104.435 58.855 104.685 ;
        RECT 59.040 104.225 59.210 104.855 ;
        RECT 59.380 104.435 59.710 104.635 ;
        RECT 59.880 104.435 60.210 104.635 ;
        RECT 60.380 104.435 60.800 104.635 ;
        RECT 60.975 104.605 61.145 104.855 ;
        RECT 60.975 104.435 61.670 104.605 ;
        RECT 56.655 103.615 56.935 104.075 ;
        RECT 57.455 103.445 57.780 103.905 ;
        RECT 57.950 103.615 58.335 104.185 ;
        RECT 58.710 103.615 59.210 104.225 ;
        RECT 59.840 104.095 61.065 104.265 ;
        RECT 61.840 104.245 62.015 104.855 ;
        RECT 62.635 104.845 62.965 105.825 ;
        RECT 63.135 104.855 63.395 105.995 ;
        RECT 63.570 104.855 63.905 105.825 ;
        RECT 64.075 104.855 64.245 105.995 ;
        RECT 64.415 105.655 66.445 105.825 ;
        RECT 62.195 104.415 62.530 104.685 ;
        RECT 62.700 104.245 62.870 104.845 ;
        RECT 63.040 104.435 63.375 104.685 ;
        RECT 59.840 103.615 60.170 104.095 ;
        RECT 60.340 103.445 60.565 103.905 ;
        RECT 60.735 103.615 61.065 104.095 ;
        RECT 61.255 103.445 61.505 104.245 ;
        RECT 61.675 103.615 62.015 104.245 ;
        RECT 62.185 103.445 62.495 104.245 ;
        RECT 62.700 103.615 63.395 104.245 ;
        RECT 63.570 104.185 63.740 104.855 ;
        RECT 64.415 104.685 64.585 105.655 ;
        RECT 63.910 104.355 64.165 104.685 ;
        RECT 64.390 104.355 64.585 104.685 ;
        RECT 64.755 105.315 65.880 105.485 ;
        RECT 63.995 104.185 64.165 104.355 ;
        RECT 64.755 104.185 64.925 105.315 ;
        RECT 63.570 103.615 63.825 104.185 ;
        RECT 63.995 104.015 64.925 104.185 ;
        RECT 65.095 104.975 66.105 105.145 ;
        RECT 65.095 104.175 65.265 104.975 ;
        RECT 65.470 104.635 65.745 104.775 ;
        RECT 65.465 104.465 65.745 104.635 ;
        RECT 64.750 103.980 64.925 104.015 ;
        RECT 63.995 103.445 64.325 103.845 ;
        RECT 64.750 103.615 65.280 103.980 ;
        RECT 65.470 103.615 65.745 104.465 ;
        RECT 65.915 103.615 66.105 104.975 ;
        RECT 66.275 104.990 66.445 105.655 ;
        RECT 66.615 105.235 66.785 105.995 ;
        RECT 67.020 105.235 67.535 105.645 ;
        RECT 66.275 104.800 67.025 104.990 ;
        RECT 67.195 104.425 67.535 105.235 ;
        RECT 67.705 104.905 69.375 105.995 ;
        RECT 66.305 104.255 67.535 104.425 ;
        RECT 66.285 103.445 66.795 103.980 ;
        RECT 67.015 103.650 67.260 104.255 ;
        RECT 67.705 104.215 68.455 104.735 ;
        RECT 68.625 104.385 69.375 104.905 ;
        RECT 70.005 104.830 70.295 105.995 ;
        RECT 70.960 105.205 71.495 105.825 ;
        RECT 67.705 103.445 69.375 104.215 ;
        RECT 70.960 104.185 71.275 105.205 ;
        RECT 71.665 105.195 71.995 105.995 ;
        RECT 72.480 105.025 72.870 105.200 ;
        RECT 71.445 104.855 72.870 105.025 ;
        RECT 73.225 104.905 74.435 105.995 ;
        RECT 74.695 105.325 74.865 105.825 ;
        RECT 75.035 105.495 75.365 105.995 ;
        RECT 74.695 105.155 75.360 105.325 ;
        RECT 71.445 104.355 71.615 104.855 ;
        RECT 70.005 103.445 70.295 104.170 ;
        RECT 70.960 103.615 71.575 104.185 ;
        RECT 71.865 104.125 72.130 104.685 ;
        RECT 72.300 103.955 72.470 104.855 ;
        RECT 72.640 104.125 72.995 104.685 ;
        RECT 73.225 104.195 73.745 104.735 ;
        RECT 73.915 104.365 74.435 104.905 ;
        RECT 74.610 104.335 74.960 104.985 ;
        RECT 71.745 103.445 71.960 103.955 ;
        RECT 72.190 103.625 72.470 103.955 ;
        RECT 72.650 103.445 72.890 103.955 ;
        RECT 73.225 103.445 74.435 104.195 ;
        RECT 75.130 104.165 75.360 105.155 ;
        RECT 74.695 103.995 75.360 104.165 ;
        RECT 74.695 103.705 74.865 103.995 ;
        RECT 75.035 103.445 75.365 103.825 ;
        RECT 75.535 103.705 75.720 105.825 ;
        RECT 75.960 105.535 76.225 105.995 ;
        RECT 76.395 105.400 76.645 105.825 ;
        RECT 76.855 105.550 77.960 105.720 ;
        RECT 76.340 105.270 76.645 105.400 ;
        RECT 75.890 104.075 76.170 105.025 ;
        RECT 76.340 104.165 76.510 105.270 ;
        RECT 76.680 104.485 76.920 105.080 ;
        RECT 77.090 105.015 77.620 105.380 ;
        RECT 77.090 104.315 77.260 105.015 ;
        RECT 77.790 104.935 77.960 105.550 ;
        RECT 78.130 105.195 78.300 105.995 ;
        RECT 78.470 105.495 78.720 105.825 ;
        RECT 78.945 105.525 79.830 105.695 ;
        RECT 77.790 104.845 78.300 104.935 ;
        RECT 76.340 104.035 76.565 104.165 ;
        RECT 76.735 104.095 77.260 104.315 ;
        RECT 77.430 104.675 78.300 104.845 ;
        RECT 75.975 103.445 76.225 103.905 ;
        RECT 76.395 103.895 76.565 104.035 ;
        RECT 77.430 103.895 77.600 104.675 ;
        RECT 78.130 104.605 78.300 104.675 ;
        RECT 77.810 104.425 78.010 104.455 ;
        RECT 78.470 104.425 78.640 105.495 ;
        RECT 78.810 104.605 79.000 105.325 ;
        RECT 77.810 104.125 78.640 104.425 ;
        RECT 79.170 104.395 79.490 105.355 ;
        RECT 76.395 103.725 76.730 103.895 ;
        RECT 76.925 103.725 77.600 103.895 ;
        RECT 77.920 103.445 78.290 103.945 ;
        RECT 78.470 103.895 78.640 104.125 ;
        RECT 79.025 104.065 79.490 104.395 ;
        RECT 79.660 104.685 79.830 105.525 ;
        RECT 80.010 105.495 80.325 105.995 ;
        RECT 80.555 105.265 80.895 105.825 ;
        RECT 80.000 104.890 80.895 105.265 ;
        RECT 81.065 104.985 81.235 105.995 ;
        RECT 80.705 104.685 80.895 104.890 ;
        RECT 81.405 104.935 81.735 105.780 ;
        RECT 81.405 104.855 81.795 104.935 ;
        RECT 81.580 104.805 81.795 104.855 ;
        RECT 79.660 104.355 80.535 104.685 ;
        RECT 80.705 104.355 81.455 104.685 ;
        RECT 79.660 103.895 79.830 104.355 ;
        RECT 80.705 104.185 80.905 104.355 ;
        RECT 81.625 104.225 81.795 104.805 ;
        RECT 81.965 104.905 83.175 105.995 ;
        RECT 81.965 104.365 82.485 104.905 ;
        RECT 81.570 104.185 81.795 104.225 ;
        RECT 82.655 104.195 83.175 104.735 ;
        RECT 78.470 103.725 78.875 103.895 ;
        RECT 79.045 103.725 79.830 103.895 ;
        RECT 80.105 103.445 80.315 103.975 ;
        RECT 80.575 103.660 80.905 104.185 ;
        RECT 81.415 104.100 81.795 104.185 ;
        RECT 81.075 103.445 81.245 104.055 ;
        RECT 81.415 103.665 81.745 104.100 ;
        RECT 81.965 103.445 83.175 104.195 ;
        RECT 5.520 103.275 83.260 103.445 ;
        RECT 5.605 102.525 6.815 103.275 ;
        RECT 7.535 102.725 7.705 103.015 ;
        RECT 7.875 102.895 8.205 103.275 ;
        RECT 7.535 102.555 8.200 102.725 ;
        RECT 5.605 101.985 6.125 102.525 ;
        RECT 6.295 101.815 6.815 102.355 ;
        RECT 5.605 100.725 6.815 101.815 ;
        RECT 7.450 101.735 7.800 102.385 ;
        RECT 7.970 101.565 8.200 102.555 ;
        RECT 7.535 101.395 8.200 101.565 ;
        RECT 7.535 100.895 7.705 101.395 ;
        RECT 7.875 100.725 8.205 101.225 ;
        RECT 8.375 100.895 8.560 103.015 ;
        RECT 8.815 102.815 9.065 103.275 ;
        RECT 9.235 102.825 9.570 102.995 ;
        RECT 9.765 102.825 10.440 102.995 ;
        RECT 9.235 102.685 9.405 102.825 ;
        RECT 8.730 101.695 9.010 102.645 ;
        RECT 9.180 102.555 9.405 102.685 ;
        RECT 9.180 101.450 9.350 102.555 ;
        RECT 9.575 102.405 10.100 102.625 ;
        RECT 9.520 101.640 9.760 102.235 ;
        RECT 9.930 101.705 10.100 102.405 ;
        RECT 10.270 102.045 10.440 102.825 ;
        RECT 10.760 102.775 11.130 103.275 ;
        RECT 11.310 102.825 11.715 102.995 ;
        RECT 11.885 102.825 12.670 102.995 ;
        RECT 11.310 102.595 11.480 102.825 ;
        RECT 10.650 102.295 11.480 102.595 ;
        RECT 11.865 102.325 12.330 102.655 ;
        RECT 10.650 102.265 10.850 102.295 ;
        RECT 10.970 102.045 11.140 102.115 ;
        RECT 10.270 101.875 11.140 102.045 ;
        RECT 10.630 101.785 11.140 101.875 ;
        RECT 9.180 101.320 9.485 101.450 ;
        RECT 9.930 101.340 10.460 101.705 ;
        RECT 8.800 100.725 9.065 101.185 ;
        RECT 9.235 100.895 9.485 101.320 ;
        RECT 10.630 101.170 10.800 101.785 ;
        RECT 9.695 101.000 10.800 101.170 ;
        RECT 10.970 100.725 11.140 101.525 ;
        RECT 11.310 101.225 11.480 102.295 ;
        RECT 11.650 101.395 11.840 102.115 ;
        RECT 12.010 101.365 12.330 102.325 ;
        RECT 12.500 102.365 12.670 102.825 ;
        RECT 12.945 102.745 13.155 103.275 ;
        RECT 13.415 102.535 13.745 103.060 ;
        RECT 13.915 102.665 14.085 103.275 ;
        RECT 14.255 102.620 14.585 103.055 ;
        RECT 14.255 102.535 14.635 102.620 ;
        RECT 13.545 102.365 13.745 102.535 ;
        RECT 14.410 102.495 14.635 102.535 ;
        RECT 12.500 102.035 13.375 102.365 ;
        RECT 13.545 102.035 14.295 102.365 ;
        RECT 11.310 100.895 11.560 101.225 ;
        RECT 12.500 101.195 12.670 102.035 ;
        RECT 13.545 101.830 13.735 102.035 ;
        RECT 14.465 101.915 14.635 102.495 ;
        RECT 14.805 102.440 15.095 103.275 ;
        RECT 15.265 102.875 16.220 103.045 ;
        RECT 16.635 102.885 16.965 103.275 ;
        RECT 15.265 101.995 15.435 102.875 ;
        RECT 17.135 102.705 17.305 103.025 ;
        RECT 17.475 102.885 17.805 103.275 ;
        RECT 18.945 102.775 19.285 103.275 ;
        RECT 15.605 102.535 17.855 102.705 ;
        RECT 15.605 102.035 15.835 102.535 ;
        RECT 16.005 102.115 16.380 102.285 ;
        RECT 14.420 101.865 14.635 101.915 ;
        RECT 12.840 101.455 13.735 101.830 ;
        RECT 14.245 101.785 14.635 101.865 ;
        RECT 14.805 101.825 15.435 101.995 ;
        RECT 16.210 101.915 16.380 102.115 ;
        RECT 16.550 102.085 17.100 102.285 ;
        RECT 17.270 101.915 17.515 102.365 ;
        RECT 11.785 101.025 12.670 101.195 ;
        RECT 12.850 100.725 13.165 101.225 ;
        RECT 13.395 100.895 13.735 101.455 ;
        RECT 13.905 100.725 14.075 101.735 ;
        RECT 14.245 100.940 14.575 101.785 ;
        RECT 14.805 100.895 15.125 101.825 ;
        RECT 16.210 101.745 17.515 101.915 ;
        RECT 17.685 101.575 17.855 102.535 ;
        RECT 18.945 102.035 19.285 102.605 ;
        RECT 19.455 102.365 19.700 103.055 ;
        RECT 19.895 102.775 20.225 103.275 ;
        RECT 20.425 102.705 20.595 103.055 ;
        RECT 20.770 102.875 21.100 103.275 ;
        RECT 21.270 102.705 21.440 103.055 ;
        RECT 21.610 102.875 21.990 103.275 ;
        RECT 20.425 102.535 22.010 102.705 ;
        RECT 22.180 102.600 22.455 102.945 ;
        RECT 23.600 102.880 24.300 103.050 ;
        RECT 24.545 102.910 26.000 103.090 ;
        RECT 23.600 102.765 23.770 102.880 ;
        RECT 24.545 102.705 24.715 102.910 ;
        RECT 26.360 102.905 27.675 103.105 ;
        RECT 27.845 102.915 28.175 103.275 ;
        RECT 28.705 102.915 29.035 103.275 ;
        RECT 27.445 102.735 27.675 102.905 ;
        RECT 29.645 102.835 29.815 103.275 ;
        RECT 30.040 102.735 30.255 102.935 ;
        RECT 30.425 102.915 30.755 103.275 ;
        RECT 30.925 102.735 31.125 102.825 ;
        RECT 21.840 102.365 22.010 102.535 ;
        RECT 19.455 102.035 20.110 102.365 ;
        RECT 15.305 101.405 16.545 101.575 ;
        RECT 15.305 100.895 15.705 101.405 ;
        RECT 15.875 100.725 16.045 101.235 ;
        RECT 16.215 100.895 16.545 101.405 ;
        RECT 16.715 100.725 16.885 101.575 ;
        RECT 17.475 100.895 17.855 101.575 ;
        RECT 18.945 100.725 19.285 101.800 ;
        RECT 19.455 101.440 19.695 102.035 ;
        RECT 19.890 101.575 20.210 101.865 ;
        RECT 20.380 101.745 21.120 102.365 ;
        RECT 21.290 102.035 21.670 102.365 ;
        RECT 21.840 102.035 22.115 102.365 ;
        RECT 21.840 101.865 22.010 102.035 ;
        RECT 22.285 101.865 22.455 102.600 ;
        RECT 23.930 102.535 24.715 102.705 ;
        RECT 25.110 102.545 27.275 102.725 ;
        RECT 27.445 102.665 29.505 102.735 ;
        RECT 30.040 102.665 31.125 102.735 ;
        RECT 27.445 102.565 31.125 102.665 ;
        RECT 23.930 102.020 24.110 102.535 ;
        RECT 28.150 102.495 31.125 102.565 ;
        RECT 31.365 102.550 31.655 103.275 ;
        RECT 31.875 102.620 32.205 103.055 ;
        RECT 32.375 102.665 32.545 103.275 ;
        RECT 29.485 102.455 31.125 102.495 ;
        RECT 31.825 102.535 32.205 102.620 ;
        RECT 32.715 102.535 33.045 103.060 ;
        RECT 33.305 102.745 33.515 103.275 ;
        RECT 33.790 102.825 34.575 102.995 ;
        RECT 34.745 102.825 35.150 102.995 ;
        RECT 31.825 102.495 32.050 102.535 ;
        RECT 21.350 101.695 22.010 101.865 ;
        RECT 21.350 101.575 21.520 101.695 ;
        RECT 19.890 101.405 21.520 101.575 ;
        RECT 19.465 101.065 21.520 101.235 ;
        RECT 19.470 100.945 21.520 101.065 ;
        RECT 21.690 100.725 21.970 101.525 ;
        RECT 22.180 100.895 22.455 101.865 ;
        RECT 23.600 101.505 24.110 102.020 ;
        RECT 24.280 101.845 24.450 102.365 ;
        RECT 24.840 102.015 25.910 102.285 ;
        RECT 26.305 101.950 27.480 102.365 ;
        RECT 26.305 101.845 27.020 101.950 ;
        RECT 24.280 101.675 27.020 101.845 ;
        RECT 27.650 101.845 27.930 102.365 ;
        RECT 28.100 102.015 29.575 102.285 ;
        RECT 29.870 102.030 30.880 102.285 ;
        RECT 29.870 101.845 30.315 102.030 ;
        RECT 31.825 101.915 31.995 102.495 ;
        RECT 32.715 102.365 32.915 102.535 ;
        RECT 33.790 102.365 33.960 102.825 ;
        RECT 32.165 102.035 32.915 102.365 ;
        RECT 33.085 102.035 33.960 102.365 ;
        RECT 27.650 101.675 30.315 101.845 ;
        RECT 27.285 101.505 27.455 101.575 ;
        RECT 23.600 101.335 29.475 101.505 ;
        RECT 30.505 101.425 30.725 101.500 ;
        RECT 23.600 101.255 27.235 101.335 ;
        RECT 27.810 101.255 29.475 101.335 ;
        RECT 29.645 101.255 30.725 101.425 ;
        RECT 23.595 100.725 23.925 101.085 ;
        RECT 24.825 100.725 25.160 101.085 ;
        RECT 25.670 100.725 26.000 101.085 ;
        RECT 26.515 100.725 26.845 101.085 ;
        RECT 27.395 100.725 27.665 101.165 ;
        RECT 29.645 101.085 29.825 101.255 ;
        RECT 30.505 101.170 30.725 101.255 ;
        RECT 27.845 100.895 29.825 101.085 ;
        RECT 29.995 100.725 30.325 101.085 ;
        RECT 30.895 100.725 31.190 101.695 ;
        RECT 31.365 100.725 31.655 101.890 ;
        RECT 31.825 101.865 32.040 101.915 ;
        RECT 31.825 101.785 32.215 101.865 ;
        RECT 31.885 100.940 32.215 101.785 ;
        RECT 32.725 101.830 32.915 102.035 ;
        RECT 32.385 100.725 32.555 101.735 ;
        RECT 32.725 101.455 33.620 101.830 ;
        RECT 32.725 100.895 33.065 101.455 ;
        RECT 33.295 100.725 33.610 101.225 ;
        RECT 33.790 101.195 33.960 102.035 ;
        RECT 34.130 102.325 34.595 102.655 ;
        RECT 34.980 102.595 35.150 102.825 ;
        RECT 35.330 102.775 35.700 103.275 ;
        RECT 36.020 102.825 36.695 102.995 ;
        RECT 36.890 102.825 37.225 102.995 ;
        RECT 34.130 101.365 34.450 102.325 ;
        RECT 34.980 102.295 35.810 102.595 ;
        RECT 34.620 101.395 34.810 102.115 ;
        RECT 34.980 101.225 35.150 102.295 ;
        RECT 35.610 102.265 35.810 102.295 ;
        RECT 35.320 102.045 35.490 102.115 ;
        RECT 36.020 102.045 36.190 102.825 ;
        RECT 37.055 102.685 37.225 102.825 ;
        RECT 37.395 102.815 37.645 103.275 ;
        RECT 35.320 101.875 36.190 102.045 ;
        RECT 36.360 102.405 36.885 102.625 ;
        RECT 37.055 102.555 37.280 102.685 ;
        RECT 35.320 101.785 35.830 101.875 ;
        RECT 33.790 101.025 34.675 101.195 ;
        RECT 34.900 100.895 35.150 101.225 ;
        RECT 35.320 100.725 35.490 101.525 ;
        RECT 35.660 101.170 35.830 101.785 ;
        RECT 36.360 101.705 36.530 102.405 ;
        RECT 36.000 101.340 36.530 101.705 ;
        RECT 36.700 101.640 36.940 102.235 ;
        RECT 37.110 101.450 37.280 102.555 ;
        RECT 37.450 101.695 37.730 102.645 ;
        RECT 36.975 101.320 37.280 101.450 ;
        RECT 35.660 101.000 36.765 101.170 ;
        RECT 36.975 100.895 37.225 101.320 ;
        RECT 37.395 100.725 37.660 101.185 ;
        RECT 37.900 100.895 38.085 103.015 ;
        RECT 38.255 102.895 38.585 103.275 ;
        RECT 38.755 102.725 38.925 103.015 ;
        RECT 38.260 102.555 38.925 102.725 ;
        RECT 38.260 101.565 38.490 102.555 ;
        RECT 39.185 102.525 40.395 103.275 ;
        RECT 40.565 102.535 40.950 103.105 ;
        RECT 41.120 102.815 41.445 103.275 ;
        RECT 41.965 102.645 42.245 103.105 ;
        RECT 38.660 101.735 39.010 102.385 ;
        RECT 39.185 101.985 39.705 102.525 ;
        RECT 39.875 101.815 40.395 102.355 ;
        RECT 38.260 101.395 38.925 101.565 ;
        RECT 38.255 100.725 38.585 101.225 ;
        RECT 38.755 100.895 38.925 101.395 ;
        RECT 39.185 100.725 40.395 101.815 ;
        RECT 40.565 101.865 40.845 102.535 ;
        RECT 41.120 102.475 42.245 102.645 ;
        RECT 41.120 102.365 41.570 102.475 ;
        RECT 41.015 102.035 41.570 102.365 ;
        RECT 42.435 102.305 42.835 103.105 ;
        RECT 43.235 102.815 43.505 103.275 ;
        RECT 43.675 102.645 43.960 103.105 ;
        RECT 40.565 100.895 40.950 101.865 ;
        RECT 41.120 101.575 41.570 102.035 ;
        RECT 41.740 101.745 42.835 102.305 ;
        RECT 41.120 101.355 42.245 101.575 ;
        RECT 41.120 100.725 41.445 101.185 ;
        RECT 41.965 100.895 42.245 101.355 ;
        RECT 42.435 100.895 42.835 101.745 ;
        RECT 43.005 102.475 43.960 102.645 ;
        RECT 44.245 102.535 44.630 103.105 ;
        RECT 44.800 102.815 45.125 103.275 ;
        RECT 45.645 102.645 45.925 103.105 ;
        RECT 43.005 101.575 43.215 102.475 ;
        RECT 43.385 101.745 44.075 102.305 ;
        RECT 44.245 101.865 44.525 102.535 ;
        RECT 44.800 102.475 45.925 102.645 ;
        RECT 44.800 102.365 45.250 102.475 ;
        RECT 44.695 102.035 45.250 102.365 ;
        RECT 46.115 102.305 46.515 103.105 ;
        RECT 46.915 102.815 47.185 103.275 ;
        RECT 47.355 102.645 47.640 103.105 ;
        RECT 43.005 101.355 43.960 101.575 ;
        RECT 43.235 100.725 43.505 101.185 ;
        RECT 43.675 100.895 43.960 101.355 ;
        RECT 44.245 100.895 44.630 101.865 ;
        RECT 44.800 101.575 45.250 102.035 ;
        RECT 45.420 101.745 46.515 102.305 ;
        RECT 44.800 101.355 45.925 101.575 ;
        RECT 44.800 100.725 45.125 101.185 ;
        RECT 45.645 100.895 45.925 101.355 ;
        RECT 46.115 100.895 46.515 101.745 ;
        RECT 46.685 102.475 47.640 102.645 ;
        RECT 47.925 102.505 51.435 103.275 ;
        RECT 51.605 102.525 52.815 103.275 ;
        RECT 52.995 102.550 53.325 103.060 ;
        RECT 53.495 102.875 53.825 103.275 ;
        RECT 54.875 102.705 55.205 103.045 ;
        RECT 55.375 102.875 55.705 103.275 ;
        RECT 46.685 101.575 46.895 102.475 ;
        RECT 47.065 101.745 47.755 102.305 ;
        RECT 47.925 101.985 49.575 102.505 ;
        RECT 49.745 101.815 51.435 102.335 ;
        RECT 51.605 101.985 52.125 102.525 ;
        RECT 52.295 101.815 52.815 102.355 ;
        RECT 46.685 101.355 47.640 101.575 ;
        RECT 46.915 100.725 47.185 101.185 ;
        RECT 47.355 100.895 47.640 101.355 ;
        RECT 47.925 100.725 51.435 101.815 ;
        RECT 51.605 100.725 52.815 101.815 ;
        RECT 52.995 101.785 53.185 102.550 ;
        RECT 53.495 102.535 55.860 102.705 ;
        RECT 57.125 102.550 57.415 103.275 ;
        RECT 53.495 102.365 53.665 102.535 ;
        RECT 53.355 102.035 53.665 102.365 ;
        RECT 53.835 102.035 54.140 102.365 ;
        RECT 52.995 100.935 53.325 101.785 ;
        RECT 53.495 100.725 53.745 101.865 ;
        RECT 53.925 101.705 54.140 102.035 ;
        RECT 54.315 101.705 54.600 102.365 ;
        RECT 54.795 101.705 55.060 102.365 ;
        RECT 55.275 101.705 55.520 102.365 ;
        RECT 55.690 101.535 55.860 102.535 ;
        RECT 57.625 102.455 57.855 103.275 ;
        RECT 58.025 102.475 58.355 103.105 ;
        RECT 57.605 102.035 57.935 102.285 ;
        RECT 53.935 101.365 55.225 101.535 ;
        RECT 53.935 100.945 54.185 101.365 ;
        RECT 54.415 100.725 54.745 101.195 ;
        RECT 54.975 100.945 55.225 101.365 ;
        RECT 55.405 101.365 55.860 101.535 ;
        RECT 55.405 100.935 55.735 101.365 ;
        RECT 57.125 100.725 57.415 101.890 ;
        RECT 58.105 101.875 58.355 102.475 ;
        RECT 58.525 102.455 58.735 103.275 ;
        RECT 58.965 102.505 62.475 103.275 ;
        RECT 58.965 101.985 60.615 102.505 ;
        RECT 63.770 102.495 64.270 103.105 ;
        RECT 57.625 100.725 57.855 101.865 ;
        RECT 58.025 100.895 58.355 101.875 ;
        RECT 58.525 100.725 58.735 101.865 ;
        RECT 60.785 101.815 62.475 102.335 ;
        RECT 63.565 102.035 63.915 102.285 ;
        RECT 64.100 101.865 64.270 102.495 ;
        RECT 64.900 102.625 65.230 103.105 ;
        RECT 65.400 102.815 65.625 103.275 ;
        RECT 65.795 102.625 66.125 103.105 ;
        RECT 64.900 102.455 66.125 102.625 ;
        RECT 66.315 102.475 66.565 103.275 ;
        RECT 66.735 102.475 67.075 103.105 ;
        RECT 67.335 102.725 67.505 103.015 ;
        RECT 67.675 102.895 68.005 103.275 ;
        RECT 67.335 102.555 68.000 102.725 ;
        RECT 66.845 102.425 67.075 102.475 ;
        RECT 64.440 102.085 64.770 102.285 ;
        RECT 64.940 102.085 65.270 102.285 ;
        RECT 65.440 102.085 65.860 102.285 ;
        RECT 66.035 102.115 66.730 102.285 ;
        RECT 66.035 101.865 66.205 102.115 ;
        RECT 66.900 101.865 67.075 102.425 ;
        RECT 58.965 100.725 62.475 101.815 ;
        RECT 63.770 101.695 66.205 101.865 ;
        RECT 63.770 100.895 64.100 101.695 ;
        RECT 64.270 100.725 64.600 101.525 ;
        RECT 64.900 100.895 65.230 101.695 ;
        RECT 65.875 100.725 66.125 101.525 ;
        RECT 66.395 100.725 66.565 101.865 ;
        RECT 66.735 100.895 67.075 101.865 ;
        RECT 67.250 101.735 67.600 102.385 ;
        RECT 67.770 101.565 68.000 102.555 ;
        RECT 67.335 101.395 68.000 101.565 ;
        RECT 67.335 100.895 67.505 101.395 ;
        RECT 67.675 100.725 68.005 101.225 ;
        RECT 68.175 100.895 68.360 103.015 ;
        RECT 68.615 102.815 68.865 103.275 ;
        RECT 69.035 102.825 69.370 102.995 ;
        RECT 69.565 102.825 70.240 102.995 ;
        RECT 69.035 102.685 69.205 102.825 ;
        RECT 68.530 101.695 68.810 102.645 ;
        RECT 68.980 102.555 69.205 102.685 ;
        RECT 68.980 101.450 69.150 102.555 ;
        RECT 69.375 102.405 69.900 102.625 ;
        RECT 69.320 101.640 69.560 102.235 ;
        RECT 69.730 101.705 69.900 102.405 ;
        RECT 70.070 102.045 70.240 102.825 ;
        RECT 70.560 102.775 70.930 103.275 ;
        RECT 71.110 102.825 71.515 102.995 ;
        RECT 71.685 102.825 72.470 102.995 ;
        RECT 71.110 102.595 71.280 102.825 ;
        RECT 70.450 102.295 71.280 102.595 ;
        RECT 71.665 102.325 72.130 102.655 ;
        RECT 70.450 102.265 70.650 102.295 ;
        RECT 70.770 102.045 70.940 102.115 ;
        RECT 70.070 101.875 70.940 102.045 ;
        RECT 70.430 101.785 70.940 101.875 ;
        RECT 68.980 101.320 69.285 101.450 ;
        RECT 69.730 101.340 70.260 101.705 ;
        RECT 68.600 100.725 68.865 101.185 ;
        RECT 69.035 100.895 69.285 101.320 ;
        RECT 70.430 101.170 70.600 101.785 ;
        RECT 69.495 101.000 70.600 101.170 ;
        RECT 70.770 100.725 70.940 101.525 ;
        RECT 71.110 101.225 71.280 102.295 ;
        RECT 71.450 101.395 71.640 102.115 ;
        RECT 71.810 101.365 72.130 102.325 ;
        RECT 72.300 102.365 72.470 102.825 ;
        RECT 72.745 102.745 72.955 103.275 ;
        RECT 73.215 102.535 73.545 103.060 ;
        RECT 73.715 102.665 73.885 103.275 ;
        RECT 74.055 102.620 74.385 103.055 ;
        RECT 74.055 102.535 74.435 102.620 ;
        RECT 73.345 102.365 73.545 102.535 ;
        RECT 74.210 102.495 74.435 102.535 ;
        RECT 72.300 102.035 73.175 102.365 ;
        RECT 73.345 102.035 74.095 102.365 ;
        RECT 71.110 100.895 71.360 101.225 ;
        RECT 72.300 101.195 72.470 102.035 ;
        RECT 73.345 101.830 73.535 102.035 ;
        RECT 74.265 101.915 74.435 102.495 ;
        RECT 74.220 101.865 74.435 101.915 ;
        RECT 72.640 101.455 73.535 101.830 ;
        RECT 74.045 101.785 74.435 101.865 ;
        RECT 74.605 102.475 74.945 103.105 ;
        RECT 75.115 102.475 75.365 103.275 ;
        RECT 75.555 102.625 75.885 103.105 ;
        RECT 76.055 102.815 76.280 103.275 ;
        RECT 76.450 102.625 76.780 103.105 ;
        RECT 74.605 101.865 74.780 102.475 ;
        RECT 75.555 102.455 76.780 102.625 ;
        RECT 77.410 102.495 77.910 103.105 ;
        RECT 74.950 102.115 75.645 102.285 ;
        RECT 75.475 101.865 75.645 102.115 ;
        RECT 75.820 102.085 76.240 102.285 ;
        RECT 76.410 102.085 76.740 102.285 ;
        RECT 76.910 102.085 77.240 102.285 ;
        RECT 77.410 101.865 77.580 102.495 ;
        RECT 77.765 102.035 78.115 102.285 ;
        RECT 71.585 101.025 72.470 101.195 ;
        RECT 72.650 100.725 72.965 101.225 ;
        RECT 73.195 100.895 73.535 101.455 ;
        RECT 73.705 100.725 73.875 101.735 ;
        RECT 74.045 100.940 74.375 101.785 ;
        RECT 74.605 100.895 74.945 101.865 ;
        RECT 75.115 100.725 75.285 101.865 ;
        RECT 75.475 101.695 77.910 101.865 ;
        RECT 75.555 100.725 75.805 101.525 ;
        RECT 76.450 100.895 76.780 101.695 ;
        RECT 77.080 100.725 77.410 101.525 ;
        RECT 77.580 100.895 77.910 101.695 ;
        RECT 78.290 101.675 78.625 103.095 ;
        RECT 78.805 102.905 79.550 103.275 ;
        RECT 80.115 102.735 80.370 103.095 ;
        RECT 80.550 102.905 80.880 103.275 ;
        RECT 81.060 102.735 81.285 103.095 ;
        RECT 78.800 102.545 81.285 102.735 ;
        RECT 78.800 101.855 79.025 102.545 ;
        RECT 81.965 102.525 83.175 103.275 ;
        RECT 79.225 102.035 79.505 102.365 ;
        RECT 79.685 102.035 80.260 102.365 ;
        RECT 80.440 102.035 80.875 102.365 ;
        RECT 81.055 102.035 81.325 102.365 ;
        RECT 78.800 101.675 81.295 101.855 ;
        RECT 78.290 100.905 78.555 101.675 ;
        RECT 78.725 100.725 79.055 101.445 ;
        RECT 79.245 101.265 80.435 101.495 ;
        RECT 79.245 100.905 79.505 101.265 ;
        RECT 79.675 100.725 80.005 101.095 ;
        RECT 80.175 100.905 80.435 101.265 ;
        RECT 81.005 100.905 81.295 101.675 ;
        RECT 81.965 101.815 82.485 102.355 ;
        RECT 82.655 101.985 83.175 102.525 ;
        RECT 81.965 100.725 83.175 101.815 ;
        RECT 5.520 100.555 83.260 100.725 ;
        RECT 5.605 99.465 6.815 100.555 ;
        RECT 7.075 99.885 7.245 100.385 ;
        RECT 7.415 100.055 7.745 100.555 ;
        RECT 7.075 99.715 7.740 99.885 ;
        RECT 5.605 98.755 6.125 99.295 ;
        RECT 6.295 98.925 6.815 99.465 ;
        RECT 6.990 98.895 7.340 99.545 ;
        RECT 5.605 98.005 6.815 98.755 ;
        RECT 7.510 98.725 7.740 99.715 ;
        RECT 7.075 98.555 7.740 98.725 ;
        RECT 7.075 98.265 7.245 98.555 ;
        RECT 7.415 98.005 7.745 98.385 ;
        RECT 7.915 98.265 8.100 100.385 ;
        RECT 8.340 100.095 8.605 100.555 ;
        RECT 8.775 99.960 9.025 100.385 ;
        RECT 9.235 100.110 10.340 100.280 ;
        RECT 8.720 99.830 9.025 99.960 ;
        RECT 8.270 98.635 8.550 99.585 ;
        RECT 8.720 98.725 8.890 99.830 ;
        RECT 9.060 99.045 9.300 99.640 ;
        RECT 9.470 99.575 10.000 99.940 ;
        RECT 9.470 98.875 9.640 99.575 ;
        RECT 10.170 99.495 10.340 100.110 ;
        RECT 10.510 99.755 10.680 100.555 ;
        RECT 10.850 100.055 11.100 100.385 ;
        RECT 11.325 100.085 12.210 100.255 ;
        RECT 10.170 99.405 10.680 99.495 ;
        RECT 8.720 98.595 8.945 98.725 ;
        RECT 9.115 98.655 9.640 98.875 ;
        RECT 9.810 99.235 10.680 99.405 ;
        RECT 8.355 98.005 8.605 98.465 ;
        RECT 8.775 98.455 8.945 98.595 ;
        RECT 9.810 98.455 9.980 99.235 ;
        RECT 10.510 99.165 10.680 99.235 ;
        RECT 10.190 98.985 10.390 99.015 ;
        RECT 10.850 98.985 11.020 100.055 ;
        RECT 11.190 99.165 11.380 99.885 ;
        RECT 10.190 98.685 11.020 98.985 ;
        RECT 11.550 98.955 11.870 99.915 ;
        RECT 8.775 98.285 9.110 98.455 ;
        RECT 9.305 98.285 9.980 98.455 ;
        RECT 10.300 98.005 10.670 98.505 ;
        RECT 10.850 98.455 11.020 98.685 ;
        RECT 11.405 98.625 11.870 98.955 ;
        RECT 12.040 99.245 12.210 100.085 ;
        RECT 12.390 100.055 12.705 100.555 ;
        RECT 12.935 99.825 13.275 100.385 ;
        RECT 12.380 99.450 13.275 99.825 ;
        RECT 13.445 99.545 13.615 100.555 ;
        RECT 13.085 99.245 13.275 99.450 ;
        RECT 13.785 99.495 14.115 100.340 ;
        RECT 13.785 99.415 14.175 99.495 ;
        RECT 14.345 99.465 15.555 100.555 ;
        RECT 15.735 99.835 16.065 100.555 ;
        RECT 13.960 99.365 14.175 99.415 ;
        RECT 12.040 98.915 12.915 99.245 ;
        RECT 13.085 98.915 13.835 99.245 ;
        RECT 12.040 98.455 12.210 98.915 ;
        RECT 13.085 98.745 13.285 98.915 ;
        RECT 14.005 98.785 14.175 99.365 ;
        RECT 13.950 98.745 14.175 98.785 ;
        RECT 10.850 98.285 11.255 98.455 ;
        RECT 11.425 98.285 12.210 98.455 ;
        RECT 12.485 98.005 12.695 98.535 ;
        RECT 12.955 98.220 13.285 98.745 ;
        RECT 13.795 98.660 14.175 98.745 ;
        RECT 14.345 98.755 14.865 99.295 ;
        RECT 15.035 98.925 15.555 99.465 ;
        RECT 15.725 99.195 15.955 99.535 ;
        RECT 16.245 99.195 16.460 100.310 ;
        RECT 16.655 99.610 16.985 100.385 ;
        RECT 17.155 99.780 17.865 100.555 ;
        RECT 16.655 99.395 17.805 99.610 ;
        RECT 15.725 98.995 16.055 99.195 ;
        RECT 16.245 99.015 16.695 99.195 ;
        RECT 16.365 98.995 16.695 99.015 ;
        RECT 16.865 98.995 17.335 99.225 ;
        RECT 17.520 98.825 17.805 99.395 ;
        RECT 18.035 98.950 18.315 100.385 ;
        RECT 18.485 99.390 18.775 100.555 ;
        RECT 18.945 99.465 20.615 100.555 ;
        RECT 13.455 98.005 13.625 98.615 ;
        RECT 13.795 98.225 14.125 98.660 ;
        RECT 14.345 98.005 15.555 98.755 ;
        RECT 15.725 98.635 16.905 98.825 ;
        RECT 15.725 98.175 16.065 98.635 ;
        RECT 16.575 98.555 16.905 98.635 ;
        RECT 17.095 98.635 17.805 98.825 ;
        RECT 17.095 98.495 17.395 98.635 ;
        RECT 17.080 98.485 17.395 98.495 ;
        RECT 17.070 98.475 17.395 98.485 ;
        RECT 17.060 98.470 17.395 98.475 ;
        RECT 16.235 98.005 16.405 98.465 ;
        RECT 17.055 98.460 17.395 98.470 ;
        RECT 17.050 98.455 17.395 98.460 ;
        RECT 17.045 98.445 17.395 98.455 ;
        RECT 17.040 98.440 17.395 98.445 ;
        RECT 17.035 98.175 17.395 98.440 ;
        RECT 17.635 98.005 17.805 98.465 ;
        RECT 17.975 98.175 18.315 98.950 ;
        RECT 18.945 98.775 19.695 99.295 ;
        RECT 19.865 98.945 20.615 99.465 ;
        RECT 20.785 99.415 21.055 100.385 ;
        RECT 21.265 99.755 21.545 100.555 ;
        RECT 21.715 100.045 23.370 100.335 ;
        RECT 23.545 100.045 23.845 100.555 ;
        RECT 24.015 99.875 24.345 100.385 ;
        RECT 24.515 100.045 25.145 100.555 ;
        RECT 25.725 100.045 26.105 100.215 ;
        RECT 26.275 100.045 26.575 100.555 ;
        RECT 25.935 99.875 26.105 100.045 ;
        RECT 26.855 99.885 27.025 100.385 ;
        RECT 27.195 100.055 27.525 100.555 ;
        RECT 21.780 99.705 23.370 99.875 ;
        RECT 21.780 99.585 21.950 99.705 ;
        RECT 21.225 99.415 21.950 99.585 ;
        RECT 18.485 98.005 18.775 98.730 ;
        RECT 18.945 98.005 20.615 98.775 ;
        RECT 20.785 98.680 20.955 99.415 ;
        RECT 21.225 99.245 21.395 99.415 ;
        RECT 21.125 98.915 21.395 99.245 ;
        RECT 21.565 98.915 21.970 99.245 ;
        RECT 22.140 98.915 22.850 99.535 ;
        RECT 23.050 99.415 23.370 99.705 ;
        RECT 23.545 99.705 25.765 99.875 ;
        RECT 21.225 98.745 21.395 98.915 ;
        RECT 20.785 98.335 21.055 98.680 ;
        RECT 21.225 98.575 22.835 98.745 ;
        RECT 23.020 98.675 23.370 99.245 ;
        RECT 23.545 98.745 23.715 99.705 ;
        RECT 23.885 99.365 25.425 99.535 ;
        RECT 23.885 98.915 24.130 99.365 ;
        RECT 24.390 98.995 25.085 99.195 ;
        RECT 25.255 99.165 25.425 99.365 ;
        RECT 25.595 99.505 25.765 99.705 ;
        RECT 25.935 99.675 26.595 99.875 ;
        RECT 26.855 99.715 27.520 99.885 ;
        RECT 25.595 99.335 26.255 99.505 ;
        RECT 25.255 98.995 25.855 99.165 ;
        RECT 26.085 98.915 26.255 99.335 ;
        RECT 21.245 98.005 21.625 98.405 ;
        RECT 21.795 98.225 21.965 98.575 ;
        RECT 22.135 98.005 22.465 98.405 ;
        RECT 22.665 98.225 22.835 98.575 ;
        RECT 23.035 98.005 23.365 98.505 ;
        RECT 23.545 98.200 24.010 98.745 ;
        RECT 24.515 98.005 24.685 98.825 ;
        RECT 24.855 98.745 25.765 98.825 ;
        RECT 26.425 98.745 26.595 99.675 ;
        RECT 26.770 98.895 27.120 99.545 ;
        RECT 24.855 98.655 26.105 98.745 ;
        RECT 24.855 98.175 25.185 98.655 ;
        RECT 25.595 98.575 26.105 98.655 ;
        RECT 25.355 98.005 25.705 98.395 ;
        RECT 25.875 98.175 26.105 98.575 ;
        RECT 26.275 98.265 26.595 98.745 ;
        RECT 27.290 98.725 27.520 99.715 ;
        RECT 26.855 98.555 27.520 98.725 ;
        RECT 26.855 98.265 27.025 98.555 ;
        RECT 27.195 98.005 27.525 98.385 ;
        RECT 27.695 98.265 27.880 100.385 ;
        RECT 28.120 100.095 28.385 100.555 ;
        RECT 28.555 99.960 28.805 100.385 ;
        RECT 29.015 100.110 30.120 100.280 ;
        RECT 28.500 99.830 28.805 99.960 ;
        RECT 28.050 98.635 28.330 99.585 ;
        RECT 28.500 98.725 28.670 99.830 ;
        RECT 28.840 99.045 29.080 99.640 ;
        RECT 29.250 99.575 29.780 99.940 ;
        RECT 29.250 98.875 29.420 99.575 ;
        RECT 29.950 99.495 30.120 100.110 ;
        RECT 30.290 99.755 30.460 100.555 ;
        RECT 30.630 100.055 30.880 100.385 ;
        RECT 31.105 100.085 31.990 100.255 ;
        RECT 29.950 99.405 30.460 99.495 ;
        RECT 28.500 98.595 28.725 98.725 ;
        RECT 28.895 98.655 29.420 98.875 ;
        RECT 29.590 99.235 30.460 99.405 ;
        RECT 28.135 98.005 28.385 98.465 ;
        RECT 28.555 98.455 28.725 98.595 ;
        RECT 29.590 98.455 29.760 99.235 ;
        RECT 30.290 99.165 30.460 99.235 ;
        RECT 29.970 98.985 30.170 99.015 ;
        RECT 30.630 98.985 30.800 100.055 ;
        RECT 30.970 99.165 31.160 99.885 ;
        RECT 29.970 98.685 30.800 98.985 ;
        RECT 31.330 98.955 31.650 99.915 ;
        RECT 28.555 98.285 28.890 98.455 ;
        RECT 29.085 98.285 29.760 98.455 ;
        RECT 30.080 98.005 30.450 98.505 ;
        RECT 30.630 98.455 30.800 98.685 ;
        RECT 31.185 98.625 31.650 98.955 ;
        RECT 31.820 99.245 31.990 100.085 ;
        RECT 32.170 100.055 32.485 100.555 ;
        RECT 32.715 99.825 33.055 100.385 ;
        RECT 32.160 99.450 33.055 99.825 ;
        RECT 33.225 99.545 33.395 100.555 ;
        RECT 32.865 99.245 33.055 99.450 ;
        RECT 33.565 99.495 33.895 100.340 ;
        RECT 33.565 99.415 33.955 99.495 ;
        RECT 34.125 99.465 37.635 100.555 ;
        RECT 33.740 99.365 33.955 99.415 ;
        RECT 31.820 98.915 32.695 99.245 ;
        RECT 32.865 98.915 33.615 99.245 ;
        RECT 31.820 98.455 31.990 98.915 ;
        RECT 32.865 98.745 33.065 98.915 ;
        RECT 33.785 98.785 33.955 99.365 ;
        RECT 33.730 98.745 33.955 98.785 ;
        RECT 30.630 98.285 31.035 98.455 ;
        RECT 31.205 98.285 31.990 98.455 ;
        RECT 32.265 98.005 32.475 98.535 ;
        RECT 32.735 98.220 33.065 98.745 ;
        RECT 33.575 98.660 33.955 98.745 ;
        RECT 34.125 98.775 35.775 99.295 ;
        RECT 35.945 98.945 37.635 99.465 ;
        RECT 38.010 99.585 38.340 100.385 ;
        RECT 38.510 99.755 38.840 100.555 ;
        RECT 39.140 99.585 39.470 100.385 ;
        RECT 40.115 99.755 40.365 100.555 ;
        RECT 38.010 99.415 40.445 99.585 ;
        RECT 40.635 99.415 40.805 100.555 ;
        RECT 40.975 99.415 41.315 100.385 ;
        RECT 41.535 100.095 41.745 100.555 ;
        RECT 42.235 99.965 42.735 100.385 ;
        RECT 37.805 98.995 38.155 99.245 ;
        RECT 38.340 98.785 38.510 99.415 ;
        RECT 38.680 98.995 39.010 99.195 ;
        RECT 39.180 98.995 39.510 99.195 ;
        RECT 39.680 98.995 40.100 99.195 ;
        RECT 40.275 99.165 40.445 99.415 ;
        RECT 41.085 99.365 41.315 99.415 ;
        RECT 40.275 98.995 40.970 99.165 ;
        RECT 33.235 98.005 33.405 98.615 ;
        RECT 33.575 98.225 33.905 98.660 ;
        RECT 34.125 98.005 37.635 98.775 ;
        RECT 38.010 98.175 38.510 98.785 ;
        RECT 39.140 98.655 40.365 98.825 ;
        RECT 41.140 98.805 41.315 99.365 ;
        RECT 39.140 98.175 39.470 98.655 ;
        RECT 39.640 98.005 39.865 98.465 ;
        RECT 40.035 98.175 40.365 98.655 ;
        RECT 40.555 98.005 40.805 98.805 ;
        RECT 40.975 98.175 41.315 98.805 ;
        RECT 41.485 98.585 41.725 99.910 ;
        RECT 41.895 99.755 42.735 99.965 ;
        RECT 41.895 98.745 42.065 99.755 ;
        RECT 42.235 99.335 42.635 99.585 ;
        RECT 42.925 99.535 43.125 100.325 ;
        RECT 42.805 99.365 43.125 99.535 ;
        RECT 43.295 99.375 43.615 100.555 ;
        RECT 44.245 99.390 44.535 100.555 ;
        RECT 44.710 99.415 45.030 100.555 ;
        RECT 42.235 98.915 42.405 99.335 ;
        RECT 42.805 99.165 42.985 99.365 ;
        RECT 45.210 99.245 45.405 100.295 ;
        RECT 45.585 99.705 45.915 100.385 ;
        RECT 46.115 99.755 46.370 100.555 ;
        RECT 45.585 99.425 45.935 99.705 ;
        RECT 47.470 99.605 47.735 100.375 ;
        RECT 47.905 99.835 48.235 100.555 ;
        RECT 48.425 100.015 48.685 100.375 ;
        RECT 48.855 100.185 49.185 100.555 ;
        RECT 49.355 100.015 49.615 100.375 ;
        RECT 48.425 99.785 49.615 100.015 ;
        RECT 50.185 99.605 50.475 100.375 ;
        RECT 44.770 99.195 45.030 99.245 ;
        RECT 42.620 98.995 42.985 99.165 ;
        RECT 43.155 98.995 43.615 99.195 ;
        RECT 44.765 99.025 45.030 99.195 ;
        RECT 44.770 98.915 45.030 99.025 ;
        RECT 45.210 98.915 45.595 99.245 ;
        RECT 45.765 99.045 45.935 99.425 ;
        RECT 46.125 99.215 46.370 99.575 ;
        RECT 45.765 98.875 46.285 99.045 ;
        RECT 46.115 98.855 46.285 98.875 ;
        RECT 42.585 98.745 43.615 98.785 ;
        RECT 41.895 98.565 42.245 98.745 ;
        RECT 42.415 98.615 43.615 98.745 ;
        RECT 42.415 98.395 42.745 98.615 ;
        RECT 41.485 98.215 42.745 98.395 ;
        RECT 42.935 98.005 43.105 98.445 ;
        RECT 43.275 98.200 43.615 98.615 ;
        RECT 44.245 98.005 44.535 98.730 ;
        RECT 44.710 98.535 45.925 98.705 ;
        RECT 44.710 98.185 45.000 98.535 ;
        RECT 45.195 98.005 45.525 98.365 ;
        RECT 45.695 98.230 45.925 98.535 ;
        RECT 46.115 98.685 46.315 98.855 ;
        RECT 46.115 98.310 46.285 98.685 ;
        RECT 47.470 98.185 47.805 99.605 ;
        RECT 47.980 99.425 50.475 99.605 ;
        RECT 50.685 99.465 54.195 100.555 ;
        RECT 55.365 99.925 55.545 100.385 ;
        RECT 55.715 100.095 55.965 100.555 ;
        RECT 56.135 100.175 56.465 100.345 ;
        RECT 56.635 100.290 56.890 100.385 ;
        RECT 56.135 99.925 56.305 100.175 ;
        RECT 56.635 100.120 57.775 100.290 ;
        RECT 58.035 100.155 58.365 100.555 ;
        RECT 56.635 99.985 56.890 100.120 ;
        RECT 55.365 99.755 56.305 99.925 ;
        RECT 56.480 99.815 56.890 99.985 ;
        RECT 57.605 99.895 57.775 100.120 ;
        RECT 47.980 98.735 48.205 99.425 ;
        RECT 48.405 98.915 48.685 99.245 ;
        RECT 48.865 98.915 49.440 99.245 ;
        RECT 49.620 98.915 50.055 99.245 ;
        RECT 50.235 98.915 50.505 99.245 ;
        RECT 50.685 98.775 52.335 99.295 ;
        RECT 52.505 98.945 54.195 99.465 ;
        RECT 47.980 98.545 50.465 98.735 ;
        RECT 47.985 98.005 48.730 98.375 ;
        RECT 49.295 98.185 49.550 98.545 ;
        RECT 49.730 98.005 50.060 98.375 ;
        RECT 50.240 98.185 50.465 98.545 ;
        RECT 50.685 98.005 54.195 98.775 ;
        RECT 55.340 98.685 55.600 99.575 ;
        RECT 55.800 99.275 56.280 99.575 ;
        RECT 55.800 98.685 56.060 99.275 ;
        RECT 56.480 98.790 56.650 99.815 ;
        RECT 57.170 99.635 57.340 99.825 ;
        RECT 57.605 99.725 58.365 99.895 ;
        RECT 56.300 98.620 56.650 98.790 ;
        RECT 56.820 99.465 57.340 99.635 ;
        RECT 56.820 98.745 56.990 99.465 ;
        RECT 57.180 98.915 57.470 99.295 ;
        RECT 57.640 98.915 57.970 99.535 ;
        RECT 58.195 99.245 58.365 99.725 ;
        RECT 58.535 99.445 58.795 100.385 ;
        RECT 59.055 99.645 59.225 100.375 ;
        RECT 59.405 99.825 59.735 100.555 ;
        RECT 59.905 99.645 60.095 100.375 ;
        RECT 59.055 99.445 60.095 99.645 ;
        RECT 58.195 98.915 58.450 99.245 ;
        RECT 55.325 98.005 55.725 98.515 ;
        RECT 56.300 98.175 56.470 98.620 ;
        RECT 56.820 98.575 57.700 98.745 ;
        RECT 58.620 98.730 58.795 99.445 ;
        RECT 60.265 99.265 60.595 100.375 ;
        RECT 60.785 100.145 61.115 100.555 ;
        RECT 61.285 99.965 61.545 100.355 ;
        RECT 61.725 100.120 67.070 100.555 ;
        RECT 59.000 98.915 59.290 99.265 ;
        RECT 59.485 98.915 59.880 99.265 ;
        RECT 60.060 98.965 60.595 99.265 ;
        RECT 60.785 99.765 61.545 99.965 ;
        RECT 60.785 99.085 61.125 99.765 ;
        RECT 56.640 98.005 57.360 98.405 ;
        RECT 57.530 98.175 57.700 98.575 ;
        RECT 57.935 98.005 58.365 98.450 ;
        RECT 58.535 98.175 58.795 98.730 ;
        RECT 58.985 98.005 59.315 98.735 ;
        RECT 59.485 98.295 59.695 98.915 ;
        RECT 60.060 98.715 60.305 98.965 ;
        RECT 59.875 98.185 60.305 98.715 ;
        RECT 60.485 98.005 60.715 98.785 ;
        RECT 60.895 98.635 61.125 99.085 ;
        RECT 61.305 98.895 61.535 99.585 ;
        RECT 60.895 98.185 61.275 98.635 ;
        RECT 63.310 98.550 63.650 99.380 ;
        RECT 65.130 98.870 65.480 100.120 ;
        RECT 68.170 99.405 68.430 100.555 ;
        RECT 68.605 99.480 68.860 100.385 ;
        RECT 69.030 99.795 69.360 100.555 ;
        RECT 69.575 99.625 69.745 100.385 ;
        RECT 61.725 98.005 67.070 98.550 ;
        RECT 68.170 98.005 68.430 98.845 ;
        RECT 68.605 98.750 68.775 99.480 ;
        RECT 69.030 99.455 69.745 99.625 ;
        RECT 69.030 99.245 69.200 99.455 ;
        RECT 70.005 99.390 70.295 100.555 ;
        RECT 70.555 99.885 70.725 100.385 ;
        RECT 70.895 100.055 71.225 100.555 ;
        RECT 70.555 99.715 71.220 99.885 ;
        RECT 68.945 98.915 69.200 99.245 ;
        RECT 68.605 98.175 68.860 98.750 ;
        RECT 69.030 98.725 69.200 98.915 ;
        RECT 69.480 98.905 69.835 99.275 ;
        RECT 70.470 98.895 70.820 99.545 ;
        RECT 69.030 98.555 69.745 98.725 ;
        RECT 69.030 98.005 69.360 98.385 ;
        RECT 69.575 98.175 69.745 98.555 ;
        RECT 70.005 98.005 70.295 98.730 ;
        RECT 70.990 98.725 71.220 99.715 ;
        RECT 70.555 98.555 71.220 98.725 ;
        RECT 70.555 98.265 70.725 98.555 ;
        RECT 70.895 98.005 71.225 98.385 ;
        RECT 71.395 98.265 71.580 100.385 ;
        RECT 71.820 100.095 72.085 100.555 ;
        RECT 72.255 99.960 72.505 100.385 ;
        RECT 72.715 100.110 73.820 100.280 ;
        RECT 72.200 99.830 72.505 99.960 ;
        RECT 71.750 98.635 72.030 99.585 ;
        RECT 72.200 98.725 72.370 99.830 ;
        RECT 72.540 99.045 72.780 99.640 ;
        RECT 72.950 99.575 73.480 99.940 ;
        RECT 72.950 98.875 73.120 99.575 ;
        RECT 73.650 99.495 73.820 100.110 ;
        RECT 73.990 99.755 74.160 100.555 ;
        RECT 74.330 100.055 74.580 100.385 ;
        RECT 74.805 100.085 75.690 100.255 ;
        RECT 73.650 99.405 74.160 99.495 ;
        RECT 72.200 98.595 72.425 98.725 ;
        RECT 72.595 98.655 73.120 98.875 ;
        RECT 73.290 99.235 74.160 99.405 ;
        RECT 71.835 98.005 72.085 98.465 ;
        RECT 72.255 98.455 72.425 98.595 ;
        RECT 73.290 98.455 73.460 99.235 ;
        RECT 73.990 99.165 74.160 99.235 ;
        RECT 73.670 98.985 73.870 99.015 ;
        RECT 74.330 98.985 74.500 100.055 ;
        RECT 74.670 99.165 74.860 99.885 ;
        RECT 73.670 98.685 74.500 98.985 ;
        RECT 75.030 98.955 75.350 99.915 ;
        RECT 72.255 98.285 72.590 98.455 ;
        RECT 72.785 98.285 73.460 98.455 ;
        RECT 73.780 98.005 74.150 98.505 ;
        RECT 74.330 98.455 74.500 98.685 ;
        RECT 74.885 98.625 75.350 98.955 ;
        RECT 75.520 99.245 75.690 100.085 ;
        RECT 75.870 100.055 76.185 100.555 ;
        RECT 76.415 99.825 76.755 100.385 ;
        RECT 75.860 99.450 76.755 99.825 ;
        RECT 76.925 99.545 77.095 100.555 ;
        RECT 76.565 99.245 76.755 99.450 ;
        RECT 77.265 99.495 77.595 100.340 ;
        RECT 78.290 100.165 78.625 100.385 ;
        RECT 79.630 100.175 79.985 100.555 ;
        RECT 78.290 99.545 78.545 100.165 ;
        RECT 78.795 100.005 79.025 100.045 ;
        RECT 80.155 100.005 80.405 100.385 ;
        RECT 78.795 99.805 80.405 100.005 ;
        RECT 78.795 99.715 78.980 99.805 ;
        RECT 79.570 99.795 80.405 99.805 ;
        RECT 80.655 99.775 80.905 100.555 ;
        RECT 81.075 99.705 81.335 100.385 ;
        RECT 79.135 99.605 79.465 99.635 ;
        RECT 79.135 99.545 80.935 99.605 ;
        RECT 77.265 99.415 77.655 99.495 ;
        RECT 77.440 99.365 77.655 99.415 ;
        RECT 78.290 99.435 80.995 99.545 ;
        RECT 78.290 99.375 79.465 99.435 ;
        RECT 80.795 99.400 80.995 99.435 ;
        RECT 75.520 98.915 76.395 99.245 ;
        RECT 76.565 98.915 77.315 99.245 ;
        RECT 75.520 98.455 75.690 98.915 ;
        RECT 76.565 98.745 76.765 98.915 ;
        RECT 77.485 98.785 77.655 99.365 ;
        RECT 78.285 98.995 78.775 99.195 ;
        RECT 78.965 98.995 79.440 99.205 ;
        RECT 77.430 98.745 77.655 98.785 ;
        RECT 74.330 98.285 74.735 98.455 ;
        RECT 74.905 98.285 75.690 98.455 ;
        RECT 75.965 98.005 76.175 98.535 ;
        RECT 76.435 98.220 76.765 98.745 ;
        RECT 77.275 98.660 77.655 98.745 ;
        RECT 76.935 98.005 77.105 98.615 ;
        RECT 77.275 98.225 77.605 98.660 ;
        RECT 78.290 98.005 78.745 98.770 ;
        RECT 79.220 98.595 79.440 98.995 ;
        RECT 79.685 98.995 80.015 99.205 ;
        RECT 79.685 98.595 79.895 98.995 ;
        RECT 80.185 98.960 80.595 99.265 ;
        RECT 80.825 98.825 80.995 99.400 ;
        RECT 80.725 98.705 80.995 98.825 ;
        RECT 80.150 98.660 80.995 98.705 ;
        RECT 80.150 98.535 80.905 98.660 ;
        RECT 80.150 98.385 80.320 98.535 ;
        RECT 81.165 98.505 81.335 99.705 ;
        RECT 81.965 99.465 83.175 100.555 ;
        RECT 81.965 98.925 82.485 99.465 ;
        RECT 82.655 98.755 83.175 99.295 ;
        RECT 79.020 98.175 80.320 98.385 ;
        RECT 80.575 98.005 80.905 98.365 ;
        RECT 81.075 98.175 81.335 98.505 ;
        RECT 81.965 98.005 83.175 98.755 ;
        RECT 5.520 97.835 83.260 98.005 ;
        RECT 5.605 97.085 6.815 97.835 ;
        RECT 5.605 96.545 6.125 97.085 ;
        RECT 6.985 97.065 8.655 97.835 ;
        RECT 8.875 97.445 9.205 97.835 ;
        RECT 9.375 97.265 9.545 97.585 ;
        RECT 9.715 97.445 10.045 97.835 ;
        RECT 10.460 97.435 11.415 97.605 ;
        RECT 8.825 97.095 11.075 97.265 ;
        RECT 6.295 96.375 6.815 96.915 ;
        RECT 6.985 96.545 7.735 97.065 ;
        RECT 7.905 96.375 8.655 96.895 ;
        RECT 5.605 95.285 6.815 96.375 ;
        RECT 6.985 95.285 8.655 96.375 ;
        RECT 8.825 96.135 8.995 97.095 ;
        RECT 9.165 96.475 9.410 96.925 ;
        RECT 9.580 96.645 10.130 96.845 ;
        RECT 10.300 96.675 10.675 96.845 ;
        RECT 10.300 96.475 10.470 96.675 ;
        RECT 10.845 96.595 11.075 97.095 ;
        RECT 9.165 96.305 10.470 96.475 ;
        RECT 11.245 96.555 11.415 97.435 ;
        RECT 11.585 97.000 11.875 97.835 ;
        RECT 12.045 97.335 12.345 97.665 ;
        RECT 12.515 97.355 12.790 97.835 ;
        RECT 11.245 96.385 11.875 96.555 ;
        RECT 8.825 95.455 9.205 96.135 ;
        RECT 9.795 95.285 9.965 96.135 ;
        RECT 10.135 95.965 11.375 96.135 ;
        RECT 10.135 95.455 10.465 95.965 ;
        RECT 10.635 95.285 10.805 95.795 ;
        RECT 10.975 95.455 11.375 95.965 ;
        RECT 11.555 95.455 11.875 96.385 ;
        RECT 12.045 96.425 12.215 97.335 ;
        RECT 12.970 97.185 13.265 97.575 ;
        RECT 13.435 97.355 13.690 97.835 ;
        RECT 13.865 97.185 14.125 97.575 ;
        RECT 14.295 97.355 14.575 97.835 ;
        RECT 15.310 97.375 16.060 97.665 ;
        RECT 16.570 97.375 16.900 97.835 ;
        RECT 12.385 96.595 12.735 97.165 ;
        RECT 12.970 97.015 14.620 97.185 ;
        RECT 12.905 96.675 14.045 96.845 ;
        RECT 12.905 96.425 13.075 96.675 ;
        RECT 14.215 96.505 14.620 97.015 ;
        RECT 12.045 96.255 13.075 96.425 ;
        RECT 13.865 96.335 14.620 96.505 ;
        RECT 12.045 95.455 12.355 96.255 ;
        RECT 13.865 96.085 14.125 96.335 ;
        RECT 12.525 95.285 12.835 96.085 ;
        RECT 13.005 95.915 14.125 96.085 ;
        RECT 13.005 95.455 13.265 95.915 ;
        RECT 13.435 95.285 13.690 95.745 ;
        RECT 13.865 95.455 14.125 95.915 ;
        RECT 14.295 95.285 14.580 96.155 ;
        RECT 15.310 96.085 15.680 97.375 ;
        RECT 17.120 97.185 17.390 97.395 ;
        RECT 18.030 97.330 18.365 97.835 ;
        RECT 18.535 97.265 18.775 97.640 ;
        RECT 19.055 97.505 19.225 97.650 ;
        RECT 19.055 97.310 19.430 97.505 ;
        RECT 19.790 97.340 20.185 97.835 ;
        RECT 16.055 97.015 17.390 97.185 ;
        RECT 16.055 96.845 16.225 97.015 ;
        RECT 15.850 96.595 16.225 96.845 ;
        RECT 16.395 96.605 16.870 96.845 ;
        RECT 17.040 96.605 17.390 96.845 ;
        RECT 16.055 96.425 16.225 96.595 ;
        RECT 16.055 96.255 17.390 96.425 ;
        RECT 18.085 96.305 18.385 97.155 ;
        RECT 18.555 97.115 18.775 97.265 ;
        RECT 18.555 96.785 19.090 97.115 ;
        RECT 19.260 96.975 19.430 97.310 ;
        RECT 20.355 97.145 20.595 97.665 ;
        RECT 17.110 96.095 17.390 96.255 ;
        RECT 18.555 96.135 18.790 96.785 ;
        RECT 19.260 96.615 20.245 96.975 ;
        RECT 15.310 95.915 16.480 96.085 ;
        RECT 15.765 95.285 15.980 95.745 ;
        RECT 16.150 95.455 16.480 95.915 ;
        RECT 16.650 95.285 16.900 96.085 ;
        RECT 18.115 95.905 18.790 96.135 ;
        RECT 18.960 96.595 20.245 96.615 ;
        RECT 18.960 96.445 19.820 96.595 ;
        RECT 18.115 95.475 18.285 95.905 ;
        RECT 18.455 95.285 18.785 95.735 ;
        RECT 18.960 95.500 19.245 96.445 ;
        RECT 20.420 96.340 20.595 97.145 ;
        RECT 20.825 97.015 21.055 97.835 ;
        RECT 21.225 97.035 21.555 97.665 ;
        RECT 20.805 96.595 21.135 96.845 ;
        RECT 21.305 96.435 21.555 97.035 ;
        RECT 21.725 97.015 21.935 97.835 ;
        RECT 22.165 97.065 23.835 97.835 ;
        RECT 24.005 97.095 24.495 97.665 ;
        RECT 24.665 97.265 24.895 97.665 ;
        RECT 25.065 97.435 25.485 97.835 ;
        RECT 25.655 97.265 25.825 97.665 ;
        RECT 24.665 97.095 25.825 97.265 ;
        RECT 25.995 97.095 26.445 97.835 ;
        RECT 26.615 97.095 27.055 97.655 ;
        RECT 22.165 96.545 22.915 97.065 ;
        RECT 19.420 95.965 20.115 96.275 ;
        RECT 19.425 95.285 20.110 95.755 ;
        RECT 20.290 95.555 20.595 96.340 ;
        RECT 20.825 95.285 21.055 96.425 ;
        RECT 21.225 95.455 21.555 96.435 ;
        RECT 21.725 95.285 21.935 96.425 ;
        RECT 23.085 96.375 23.835 96.895 ;
        RECT 22.165 95.285 23.835 96.375 ;
        RECT 24.005 96.425 24.175 97.095 ;
        RECT 24.345 96.595 24.750 96.925 ;
        RECT 24.005 96.255 24.775 96.425 ;
        RECT 24.015 95.285 24.345 96.085 ;
        RECT 24.525 95.625 24.775 96.255 ;
        RECT 24.965 95.795 25.215 96.925 ;
        RECT 25.415 96.595 25.660 96.925 ;
        RECT 25.845 96.645 26.235 96.925 ;
        RECT 25.415 95.795 25.615 96.595 ;
        RECT 26.405 96.475 26.575 96.925 ;
        RECT 25.785 96.305 26.575 96.475 ;
        RECT 25.785 95.625 25.955 96.305 ;
        RECT 24.525 95.455 25.955 95.625 ;
        RECT 26.125 95.285 26.440 96.135 ;
        RECT 26.745 96.085 27.055 97.095 ;
        RECT 26.615 95.455 27.055 96.085 ;
        RECT 27.225 97.160 27.495 97.505 ;
        RECT 27.685 97.435 28.065 97.835 ;
        RECT 28.235 97.265 28.405 97.615 ;
        RECT 28.575 97.435 28.905 97.835 ;
        RECT 29.105 97.265 29.275 97.615 ;
        RECT 29.475 97.335 29.805 97.835 ;
        RECT 27.225 96.425 27.395 97.160 ;
        RECT 27.665 97.095 29.275 97.265 ;
        RECT 27.665 96.925 27.835 97.095 ;
        RECT 27.565 96.595 27.835 96.925 ;
        RECT 28.005 96.595 28.410 96.925 ;
        RECT 27.665 96.425 27.835 96.595 ;
        RECT 27.225 95.455 27.495 96.425 ;
        RECT 27.665 96.255 28.390 96.425 ;
        RECT 28.580 96.305 29.290 96.925 ;
        RECT 29.460 96.595 29.810 97.165 ;
        RECT 29.985 97.085 31.195 97.835 ;
        RECT 31.365 97.110 31.655 97.835 ;
        RECT 29.985 96.545 30.505 97.085 ;
        RECT 31.825 97.065 34.415 97.835 ;
        RECT 34.675 97.285 34.845 97.575 ;
        RECT 35.015 97.455 35.345 97.835 ;
        RECT 34.675 97.115 35.340 97.285 ;
        RECT 28.220 96.135 28.390 96.255 ;
        RECT 29.490 96.135 29.810 96.425 ;
        RECT 30.675 96.375 31.195 96.915 ;
        RECT 31.825 96.545 33.035 97.065 ;
        RECT 27.705 95.285 27.985 96.085 ;
        RECT 28.220 95.965 29.810 96.135 ;
        RECT 28.155 95.505 29.810 95.795 ;
        RECT 29.985 95.285 31.195 96.375 ;
        RECT 31.365 95.285 31.655 96.450 ;
        RECT 33.205 96.375 34.415 96.895 ;
        RECT 31.825 95.285 34.415 96.375 ;
        RECT 34.590 96.295 34.940 96.945 ;
        RECT 35.110 96.125 35.340 97.115 ;
        RECT 34.675 95.955 35.340 96.125 ;
        RECT 34.675 95.455 34.845 95.955 ;
        RECT 35.015 95.285 35.345 95.785 ;
        RECT 35.515 95.455 35.700 97.575 ;
        RECT 35.955 97.375 36.205 97.835 ;
        RECT 36.375 97.385 36.710 97.555 ;
        RECT 36.905 97.385 37.580 97.555 ;
        RECT 36.375 97.245 36.545 97.385 ;
        RECT 35.870 96.255 36.150 97.205 ;
        RECT 36.320 97.115 36.545 97.245 ;
        RECT 36.320 96.010 36.490 97.115 ;
        RECT 36.715 96.965 37.240 97.185 ;
        RECT 36.660 96.200 36.900 96.795 ;
        RECT 37.070 96.265 37.240 96.965 ;
        RECT 37.410 96.605 37.580 97.385 ;
        RECT 37.900 97.335 38.270 97.835 ;
        RECT 38.450 97.385 38.855 97.555 ;
        RECT 39.025 97.385 39.810 97.555 ;
        RECT 38.450 97.155 38.620 97.385 ;
        RECT 37.790 96.855 38.620 97.155 ;
        RECT 39.005 96.885 39.470 97.215 ;
        RECT 37.790 96.825 37.990 96.855 ;
        RECT 38.110 96.605 38.280 96.675 ;
        RECT 37.410 96.435 38.280 96.605 ;
        RECT 37.770 96.345 38.280 96.435 ;
        RECT 36.320 95.880 36.625 96.010 ;
        RECT 37.070 95.900 37.600 96.265 ;
        RECT 35.940 95.285 36.205 95.745 ;
        RECT 36.375 95.455 36.625 95.880 ;
        RECT 37.770 95.730 37.940 96.345 ;
        RECT 36.835 95.560 37.940 95.730 ;
        RECT 38.110 95.285 38.280 96.085 ;
        RECT 38.450 95.785 38.620 96.855 ;
        RECT 38.790 95.955 38.980 96.675 ;
        RECT 39.150 95.925 39.470 96.885 ;
        RECT 39.640 96.925 39.810 97.385 ;
        RECT 40.085 97.305 40.295 97.835 ;
        RECT 40.555 97.095 40.885 97.620 ;
        RECT 41.055 97.225 41.225 97.835 ;
        RECT 41.395 97.180 41.725 97.615 ;
        RECT 41.395 97.095 41.775 97.180 ;
        RECT 40.685 96.925 40.885 97.095 ;
        RECT 41.550 97.055 41.775 97.095 ;
        RECT 39.640 96.595 40.515 96.925 ;
        RECT 40.685 96.595 41.435 96.925 ;
        RECT 38.450 95.455 38.700 95.785 ;
        RECT 39.640 95.755 39.810 96.595 ;
        RECT 40.685 96.390 40.875 96.595 ;
        RECT 41.605 96.475 41.775 97.055 ;
        RECT 41.945 97.015 42.205 97.835 ;
        RECT 42.375 97.015 42.705 97.435 ;
        RECT 42.885 97.350 43.675 97.615 ;
        RECT 42.455 96.925 42.705 97.015 ;
        RECT 41.560 96.425 41.775 96.475 ;
        RECT 39.980 96.015 40.875 96.390 ;
        RECT 41.385 96.345 41.775 96.425 ;
        RECT 38.925 95.585 39.810 95.755 ;
        RECT 39.990 95.285 40.305 95.785 ;
        RECT 40.535 95.455 40.875 96.015 ;
        RECT 41.045 95.285 41.215 96.295 ;
        RECT 41.385 95.500 41.715 96.345 ;
        RECT 41.945 95.965 42.285 96.845 ;
        RECT 42.455 96.675 43.250 96.925 ;
        RECT 41.945 95.285 42.205 95.795 ;
        RECT 42.455 95.455 42.625 96.675 ;
        RECT 43.420 96.495 43.675 97.350 ;
        RECT 43.845 97.195 44.045 97.615 ;
        RECT 44.235 97.375 44.565 97.835 ;
        RECT 43.845 96.675 44.255 97.195 ;
        RECT 44.735 97.185 44.995 97.665 ;
        RECT 44.425 96.495 44.655 96.925 ;
        RECT 42.865 96.325 44.655 96.495 ;
        RECT 42.865 95.960 43.115 96.325 ;
        RECT 43.285 95.965 43.615 96.155 ;
        RECT 43.835 96.030 44.550 96.325 ;
        RECT 44.825 96.155 44.995 97.185 ;
        RECT 45.255 97.285 45.425 97.575 ;
        RECT 45.595 97.455 45.925 97.835 ;
        RECT 45.255 97.115 45.920 97.285 ;
        RECT 45.170 96.295 45.520 96.945 ;
        RECT 43.285 95.790 43.480 95.965 ;
        RECT 42.865 95.285 43.480 95.790 ;
        RECT 43.650 95.455 44.125 95.795 ;
        RECT 44.295 95.285 44.510 95.830 ;
        RECT 44.720 95.455 44.995 96.155 ;
        RECT 45.690 96.125 45.920 97.115 ;
        RECT 45.255 95.955 45.920 96.125 ;
        RECT 45.255 95.455 45.425 95.955 ;
        RECT 45.595 95.285 45.925 95.785 ;
        RECT 46.095 95.455 46.280 97.575 ;
        RECT 46.535 97.375 46.785 97.835 ;
        RECT 46.955 97.385 47.290 97.555 ;
        RECT 47.485 97.385 48.160 97.555 ;
        RECT 46.955 97.245 47.125 97.385 ;
        RECT 46.450 96.255 46.730 97.205 ;
        RECT 46.900 97.115 47.125 97.245 ;
        RECT 46.900 96.010 47.070 97.115 ;
        RECT 47.295 96.965 47.820 97.185 ;
        RECT 47.240 96.200 47.480 96.795 ;
        RECT 47.650 96.265 47.820 96.965 ;
        RECT 47.990 96.605 48.160 97.385 ;
        RECT 48.480 97.335 48.850 97.835 ;
        RECT 49.030 97.385 49.435 97.555 ;
        RECT 49.605 97.385 50.390 97.555 ;
        RECT 49.030 97.155 49.200 97.385 ;
        RECT 48.370 96.855 49.200 97.155 ;
        RECT 49.585 96.885 50.050 97.215 ;
        RECT 48.370 96.825 48.570 96.855 ;
        RECT 48.690 96.605 48.860 96.675 ;
        RECT 47.990 96.435 48.860 96.605 ;
        RECT 48.350 96.345 48.860 96.435 ;
        RECT 46.900 95.880 47.205 96.010 ;
        RECT 47.650 95.900 48.180 96.265 ;
        RECT 46.520 95.285 46.785 95.745 ;
        RECT 46.955 95.455 47.205 95.880 ;
        RECT 48.350 95.730 48.520 96.345 ;
        RECT 47.415 95.560 48.520 95.730 ;
        RECT 48.690 95.285 48.860 96.085 ;
        RECT 49.030 95.785 49.200 96.855 ;
        RECT 49.370 95.955 49.560 96.675 ;
        RECT 49.730 95.925 50.050 96.885 ;
        RECT 50.220 96.925 50.390 97.385 ;
        RECT 50.665 97.305 50.875 97.835 ;
        RECT 51.135 97.095 51.465 97.620 ;
        RECT 51.635 97.225 51.805 97.835 ;
        RECT 51.975 97.180 52.305 97.615 ;
        RECT 51.975 97.095 52.355 97.180 ;
        RECT 51.265 96.925 51.465 97.095 ;
        RECT 52.130 97.055 52.355 97.095 ;
        RECT 50.220 96.595 51.095 96.925 ;
        RECT 51.265 96.595 52.015 96.925 ;
        RECT 49.030 95.455 49.280 95.785 ;
        RECT 50.220 95.755 50.390 96.595 ;
        RECT 51.265 96.390 51.455 96.595 ;
        RECT 52.185 96.475 52.355 97.055 ;
        RECT 52.995 97.025 53.265 97.835 ;
        RECT 53.435 97.025 53.765 97.665 ;
        RECT 53.935 97.025 54.175 97.835 ;
        RECT 52.985 96.595 53.335 96.845 ;
        RECT 52.140 96.425 52.355 96.475 ;
        RECT 53.505 96.425 53.675 97.025 ;
        RECT 53.845 96.595 54.195 96.845 ;
        RECT 50.560 96.015 51.455 96.390 ;
        RECT 51.965 96.345 52.355 96.425 ;
        RECT 49.505 95.585 50.390 95.755 ;
        RECT 50.570 95.285 50.885 95.785 ;
        RECT 51.115 95.455 51.455 96.015 ;
        RECT 51.625 95.285 51.795 96.295 ;
        RECT 51.965 95.500 52.295 96.345 ;
        RECT 52.995 95.285 53.325 96.425 ;
        RECT 53.505 96.255 54.185 96.425 ;
        RECT 53.855 95.470 54.185 96.255 ;
        RECT 54.375 95.465 54.635 97.655 ;
        RECT 54.895 97.465 55.565 97.835 ;
        RECT 55.745 97.285 56.055 97.655 ;
        RECT 54.825 97.085 56.055 97.285 ;
        RECT 54.825 96.415 55.115 97.085 ;
        RECT 56.235 96.905 56.465 97.545 ;
        RECT 56.645 97.105 56.935 97.835 ;
        RECT 57.125 97.110 57.415 97.835 ;
        RECT 57.585 97.035 58.280 97.665 ;
        RECT 58.485 97.035 58.795 97.835 ;
        RECT 59.430 97.070 59.885 97.835 ;
        RECT 60.160 97.455 61.460 97.665 ;
        RECT 61.715 97.475 62.045 97.835 ;
        RECT 61.290 97.305 61.460 97.455 ;
        RECT 62.215 97.335 62.475 97.665 ;
        RECT 62.245 97.325 62.475 97.335 ;
        RECT 55.295 96.595 55.760 96.905 ;
        RECT 55.940 96.595 56.465 96.905 ;
        RECT 56.645 96.595 56.945 96.925 ;
        RECT 57.605 96.595 57.940 96.845 ;
        RECT 54.825 96.195 55.595 96.415 ;
        RECT 54.805 95.285 55.145 96.015 ;
        RECT 55.325 95.465 55.595 96.195 ;
        RECT 55.775 96.175 56.935 96.415 ;
        RECT 55.775 95.465 56.005 96.175 ;
        RECT 56.175 95.285 56.505 95.995 ;
        RECT 56.675 95.465 56.935 96.175 ;
        RECT 57.125 95.285 57.415 96.450 ;
        RECT 58.110 96.435 58.280 97.035 ;
        RECT 58.450 96.595 58.785 96.865 ;
        RECT 60.360 96.845 60.580 97.245 ;
        RECT 59.425 96.645 59.915 96.845 ;
        RECT 60.105 96.635 60.580 96.845 ;
        RECT 60.825 96.845 61.035 97.245 ;
        RECT 61.290 97.180 62.045 97.305 ;
        RECT 61.290 97.135 62.135 97.180 ;
        RECT 61.865 97.015 62.135 97.135 ;
        RECT 60.825 96.635 61.155 96.845 ;
        RECT 61.325 96.575 61.735 96.880 ;
        RECT 57.585 95.285 57.845 96.425 ;
        RECT 58.015 95.455 58.345 96.435 ;
        RECT 58.515 95.285 58.795 96.425 ;
        RECT 59.430 96.405 60.605 96.465 ;
        RECT 61.965 96.440 62.135 97.015 ;
        RECT 61.935 96.405 62.135 96.440 ;
        RECT 59.430 96.295 62.135 96.405 ;
        RECT 59.430 95.675 59.685 96.295 ;
        RECT 60.275 96.235 62.075 96.295 ;
        RECT 60.275 96.205 60.605 96.235 ;
        RECT 62.305 96.135 62.475 97.325 ;
        RECT 59.935 96.035 60.120 96.125 ;
        RECT 60.710 96.035 61.545 96.045 ;
        RECT 59.935 95.835 61.545 96.035 ;
        RECT 59.935 95.795 60.165 95.835 ;
        RECT 59.430 95.455 59.765 95.675 ;
        RECT 60.770 95.285 61.125 95.665 ;
        RECT 61.295 95.455 61.545 95.835 ;
        RECT 61.795 95.285 62.045 96.065 ;
        RECT 62.215 95.455 62.475 96.135 ;
        RECT 62.650 97.095 62.905 97.665 ;
        RECT 63.075 97.435 63.405 97.835 ;
        RECT 63.830 97.300 64.360 97.665 ;
        RECT 63.830 97.265 64.005 97.300 ;
        RECT 63.075 97.095 64.005 97.265 ;
        RECT 62.650 96.425 62.820 97.095 ;
        RECT 63.075 96.925 63.245 97.095 ;
        RECT 62.990 96.595 63.245 96.925 ;
        RECT 63.470 96.595 63.665 96.925 ;
        RECT 62.650 95.455 62.985 96.425 ;
        RECT 63.155 95.285 63.325 96.425 ;
        RECT 63.495 95.625 63.665 96.595 ;
        RECT 63.835 95.965 64.005 97.095 ;
        RECT 64.175 96.305 64.345 97.105 ;
        RECT 64.550 96.815 64.825 97.665 ;
        RECT 64.545 96.645 64.825 96.815 ;
        RECT 64.550 96.505 64.825 96.645 ;
        RECT 64.995 96.305 65.185 97.665 ;
        RECT 65.365 97.300 65.875 97.835 ;
        RECT 66.095 97.025 66.340 97.630 ;
        RECT 66.785 97.095 67.170 97.665 ;
        RECT 67.340 97.375 67.665 97.835 ;
        RECT 68.185 97.205 68.465 97.665 ;
        RECT 65.385 96.855 66.615 97.025 ;
        RECT 64.175 96.135 65.185 96.305 ;
        RECT 65.355 96.290 66.105 96.480 ;
        RECT 63.835 95.795 64.960 95.965 ;
        RECT 65.355 95.625 65.525 96.290 ;
        RECT 66.275 96.045 66.615 96.855 ;
        RECT 63.495 95.455 65.525 95.625 ;
        RECT 65.695 95.285 65.865 96.045 ;
        RECT 66.100 95.635 66.615 96.045 ;
        RECT 66.785 96.425 67.065 97.095 ;
        RECT 67.340 97.035 68.465 97.205 ;
        RECT 67.340 96.925 67.790 97.035 ;
        RECT 67.235 96.595 67.790 96.925 ;
        RECT 68.655 96.865 69.055 97.665 ;
        RECT 69.455 97.375 69.725 97.835 ;
        RECT 69.895 97.205 70.180 97.665 ;
        RECT 66.785 95.455 67.170 96.425 ;
        RECT 67.340 96.135 67.790 96.595 ;
        RECT 67.960 96.305 69.055 96.865 ;
        RECT 67.340 95.915 68.465 96.135 ;
        RECT 67.340 95.285 67.665 95.745 ;
        RECT 68.185 95.455 68.465 95.915 ;
        RECT 68.655 95.455 69.055 96.305 ;
        RECT 69.225 97.035 70.180 97.205 ;
        RECT 70.465 97.035 70.805 97.665 ;
        RECT 70.975 97.035 71.225 97.835 ;
        RECT 71.415 97.185 71.745 97.665 ;
        RECT 71.915 97.375 72.140 97.835 ;
        RECT 72.310 97.185 72.640 97.665 ;
        RECT 69.225 96.135 69.435 97.035 ;
        RECT 69.605 96.305 70.295 96.865 ;
        RECT 70.465 96.425 70.640 97.035 ;
        RECT 71.415 97.015 72.640 97.185 ;
        RECT 73.270 97.055 73.770 97.665 ;
        RECT 74.695 97.285 74.865 97.575 ;
        RECT 75.035 97.455 75.365 97.835 ;
        RECT 74.695 97.115 75.360 97.285 ;
        RECT 70.810 96.675 71.505 96.845 ;
        RECT 71.335 96.425 71.505 96.675 ;
        RECT 71.680 96.645 72.100 96.845 ;
        RECT 72.270 96.645 72.600 96.845 ;
        RECT 72.770 96.645 73.100 96.845 ;
        RECT 73.270 96.425 73.440 97.055 ;
        RECT 73.625 96.595 73.975 96.845 ;
        RECT 69.225 95.915 70.180 96.135 ;
        RECT 69.455 95.285 69.725 95.745 ;
        RECT 69.895 95.455 70.180 95.915 ;
        RECT 70.465 95.455 70.805 96.425 ;
        RECT 70.975 95.285 71.145 96.425 ;
        RECT 71.335 96.255 73.770 96.425 ;
        RECT 74.610 96.295 74.960 96.945 ;
        RECT 71.415 95.285 71.665 96.085 ;
        RECT 72.310 95.455 72.640 96.255 ;
        RECT 72.940 95.285 73.270 96.085 ;
        RECT 73.440 95.455 73.770 96.255 ;
        RECT 75.130 96.125 75.360 97.115 ;
        RECT 74.695 95.955 75.360 96.125 ;
        RECT 74.695 95.455 74.865 95.955 ;
        RECT 75.035 95.285 75.365 95.785 ;
        RECT 75.535 95.455 75.720 97.575 ;
        RECT 75.975 97.375 76.225 97.835 ;
        RECT 76.395 97.385 76.730 97.555 ;
        RECT 76.925 97.385 77.600 97.555 ;
        RECT 76.395 97.245 76.565 97.385 ;
        RECT 75.890 96.255 76.170 97.205 ;
        RECT 76.340 97.115 76.565 97.245 ;
        RECT 76.340 96.010 76.510 97.115 ;
        RECT 76.735 96.965 77.260 97.185 ;
        RECT 76.680 96.200 76.920 96.795 ;
        RECT 77.090 96.265 77.260 96.965 ;
        RECT 77.430 96.605 77.600 97.385 ;
        RECT 77.920 97.335 78.290 97.835 ;
        RECT 78.470 97.385 78.875 97.555 ;
        RECT 79.045 97.385 79.830 97.555 ;
        RECT 78.470 97.155 78.640 97.385 ;
        RECT 77.810 96.855 78.640 97.155 ;
        RECT 79.025 96.885 79.490 97.215 ;
        RECT 77.810 96.825 78.010 96.855 ;
        RECT 78.130 96.605 78.300 96.675 ;
        RECT 77.430 96.435 78.300 96.605 ;
        RECT 77.790 96.345 78.300 96.435 ;
        RECT 76.340 95.880 76.645 96.010 ;
        RECT 77.090 95.900 77.620 96.265 ;
        RECT 75.960 95.285 76.225 95.745 ;
        RECT 76.395 95.455 76.645 95.880 ;
        RECT 77.790 95.730 77.960 96.345 ;
        RECT 76.855 95.560 77.960 95.730 ;
        RECT 78.130 95.285 78.300 96.085 ;
        RECT 78.470 95.785 78.640 96.855 ;
        RECT 78.810 95.955 79.000 96.675 ;
        RECT 79.170 95.925 79.490 96.885 ;
        RECT 79.660 96.925 79.830 97.385 ;
        RECT 80.105 97.305 80.315 97.835 ;
        RECT 80.575 97.095 80.905 97.620 ;
        RECT 81.075 97.225 81.245 97.835 ;
        RECT 81.415 97.180 81.745 97.615 ;
        RECT 81.415 97.095 81.795 97.180 ;
        RECT 80.705 96.925 80.905 97.095 ;
        RECT 81.570 97.055 81.795 97.095 ;
        RECT 81.965 97.085 83.175 97.835 ;
        RECT 79.660 96.595 80.535 96.925 ;
        RECT 80.705 96.595 81.455 96.925 ;
        RECT 78.470 95.455 78.720 95.785 ;
        RECT 79.660 95.755 79.830 96.595 ;
        RECT 80.705 96.390 80.895 96.595 ;
        RECT 81.625 96.475 81.795 97.055 ;
        RECT 81.580 96.425 81.795 96.475 ;
        RECT 80.000 96.015 80.895 96.390 ;
        RECT 81.405 96.345 81.795 96.425 ;
        RECT 81.965 96.375 82.485 96.915 ;
        RECT 82.655 96.545 83.175 97.085 ;
        RECT 78.945 95.585 79.830 95.755 ;
        RECT 80.010 95.285 80.325 95.785 ;
        RECT 80.555 95.455 80.895 96.015 ;
        RECT 81.065 95.285 81.235 96.295 ;
        RECT 81.405 95.500 81.735 96.345 ;
        RECT 81.965 95.285 83.175 96.375 ;
        RECT 5.520 95.115 83.260 95.285 ;
        RECT 5.605 94.025 6.815 95.115 ;
        RECT 6.985 94.680 12.330 95.115 ;
        RECT 12.505 94.680 17.850 95.115 ;
        RECT 5.605 93.315 6.125 93.855 ;
        RECT 6.295 93.485 6.815 94.025 ;
        RECT 5.605 92.565 6.815 93.315 ;
        RECT 8.570 93.110 8.910 93.940 ;
        RECT 10.390 93.430 10.740 94.680 ;
        RECT 14.090 93.110 14.430 93.940 ;
        RECT 15.910 93.430 16.260 94.680 ;
        RECT 18.485 93.950 18.775 95.115 ;
        RECT 18.945 94.680 24.290 95.115 ;
        RECT 6.985 92.565 12.330 93.110 ;
        RECT 12.505 92.565 17.850 93.110 ;
        RECT 18.485 92.565 18.775 93.290 ;
        RECT 20.530 93.110 20.870 93.940 ;
        RECT 22.350 93.430 22.700 94.680 ;
        RECT 24.465 94.025 27.975 95.115 ;
        RECT 28.145 94.025 29.355 95.115 ;
        RECT 24.465 93.335 26.115 93.855 ;
        RECT 26.285 93.505 27.975 94.025 ;
        RECT 18.945 92.565 24.290 93.110 ;
        RECT 24.465 92.565 27.975 93.335 ;
        RECT 28.145 93.315 28.665 93.855 ;
        RECT 28.835 93.485 29.355 94.025 ;
        RECT 29.535 93.975 29.865 95.115 ;
        RECT 30.395 94.145 30.725 94.930 ;
        RECT 31.020 94.485 31.305 94.945 ;
        RECT 31.475 94.655 31.745 95.115 ;
        RECT 31.020 94.265 31.975 94.485 ;
        RECT 30.045 93.975 30.725 94.145 ;
        RECT 29.525 93.555 29.875 93.805 ;
        RECT 30.045 93.375 30.215 93.975 ;
        RECT 30.385 93.555 30.735 93.805 ;
        RECT 30.905 93.535 31.595 94.095 ;
        RECT 28.145 92.565 29.355 93.315 ;
        RECT 29.535 92.565 29.805 93.375 ;
        RECT 29.975 92.735 30.305 93.375 ;
        RECT 30.475 92.565 30.715 93.375 ;
        RECT 31.765 93.365 31.975 94.265 ;
        RECT 31.020 93.195 31.975 93.365 ;
        RECT 32.145 94.095 32.545 94.945 ;
        RECT 32.735 94.485 33.015 94.945 ;
        RECT 33.535 94.655 33.860 95.115 ;
        RECT 32.735 94.265 33.860 94.485 ;
        RECT 32.145 93.535 33.240 94.095 ;
        RECT 33.410 93.805 33.860 94.265 ;
        RECT 34.030 93.975 34.415 94.945 ;
        RECT 34.645 94.055 34.975 94.900 ;
        RECT 35.145 94.105 35.315 95.115 ;
        RECT 35.485 94.385 35.825 94.945 ;
        RECT 36.055 94.615 36.370 95.115 ;
        RECT 36.550 94.645 37.435 94.815 ;
        RECT 31.020 92.735 31.305 93.195 ;
        RECT 31.475 92.565 31.745 93.025 ;
        RECT 32.145 92.735 32.545 93.535 ;
        RECT 33.410 93.475 33.965 93.805 ;
        RECT 33.410 93.365 33.860 93.475 ;
        RECT 32.735 93.195 33.860 93.365 ;
        RECT 34.135 93.305 34.415 93.975 ;
        RECT 32.735 92.735 33.015 93.195 ;
        RECT 33.535 92.565 33.860 93.025 ;
        RECT 34.030 92.735 34.415 93.305 ;
        RECT 34.585 93.975 34.975 94.055 ;
        RECT 35.485 94.010 36.380 94.385 ;
        RECT 34.585 93.925 34.800 93.975 ;
        RECT 34.585 93.345 34.755 93.925 ;
        RECT 35.485 93.805 35.675 94.010 ;
        RECT 36.550 93.805 36.720 94.645 ;
        RECT 37.660 94.615 37.910 94.945 ;
        RECT 34.925 93.475 35.675 93.805 ;
        RECT 35.845 93.475 36.720 93.805 ;
        RECT 34.585 93.305 34.810 93.345 ;
        RECT 35.475 93.305 35.675 93.475 ;
        RECT 34.585 93.220 34.965 93.305 ;
        RECT 34.635 92.785 34.965 93.220 ;
        RECT 35.135 92.565 35.305 93.175 ;
        RECT 35.475 92.780 35.805 93.305 ;
        RECT 36.065 92.565 36.275 93.095 ;
        RECT 36.550 93.015 36.720 93.475 ;
        RECT 36.890 93.515 37.210 94.475 ;
        RECT 37.380 93.725 37.570 94.445 ;
        RECT 37.740 93.545 37.910 94.615 ;
        RECT 38.080 94.315 38.250 95.115 ;
        RECT 38.420 94.670 39.525 94.840 ;
        RECT 38.420 94.055 38.590 94.670 ;
        RECT 39.735 94.520 39.985 94.945 ;
        RECT 40.155 94.655 40.420 95.115 ;
        RECT 38.760 94.135 39.290 94.500 ;
        RECT 39.735 94.390 40.040 94.520 ;
        RECT 38.080 93.965 38.590 94.055 ;
        RECT 38.080 93.795 38.950 93.965 ;
        RECT 38.080 93.725 38.250 93.795 ;
        RECT 38.370 93.545 38.570 93.575 ;
        RECT 36.890 93.185 37.355 93.515 ;
        RECT 37.740 93.245 38.570 93.545 ;
        RECT 37.740 93.015 37.910 93.245 ;
        RECT 36.550 92.845 37.335 93.015 ;
        RECT 37.505 92.845 37.910 93.015 ;
        RECT 38.090 92.565 38.460 93.065 ;
        RECT 38.780 93.015 38.950 93.795 ;
        RECT 39.120 93.435 39.290 94.135 ;
        RECT 39.460 93.605 39.700 94.200 ;
        RECT 39.120 93.215 39.645 93.435 ;
        RECT 39.870 93.285 40.040 94.390 ;
        RECT 39.815 93.155 40.040 93.285 ;
        RECT 40.210 93.195 40.490 94.145 ;
        RECT 39.815 93.015 39.985 93.155 ;
        RECT 38.780 92.845 39.455 93.015 ;
        RECT 39.650 92.845 39.985 93.015 ;
        RECT 40.155 92.565 40.405 93.025 ;
        RECT 40.660 92.825 40.845 94.945 ;
        RECT 41.015 94.615 41.345 95.115 ;
        RECT 41.515 94.445 41.685 94.945 ;
        RECT 41.020 94.275 41.685 94.445 ;
        RECT 42.050 94.315 42.305 95.115 ;
        RECT 41.020 93.285 41.250 94.275 ;
        RECT 42.475 94.145 42.805 94.945 ;
        RECT 42.975 94.315 43.145 95.115 ;
        RECT 43.315 94.145 43.645 94.945 ;
        RECT 41.420 93.455 41.770 94.105 ;
        RECT 41.945 93.975 43.645 94.145 ;
        RECT 43.815 93.975 44.075 95.115 ;
        RECT 41.945 93.385 42.225 93.975 ;
        RECT 44.245 93.950 44.535 95.115 ;
        RECT 44.705 93.975 44.965 94.945 ;
        RECT 45.160 94.705 45.490 95.115 ;
        RECT 45.690 94.525 45.860 94.945 ;
        RECT 46.075 94.705 46.745 95.115 ;
        RECT 46.980 94.525 47.150 94.945 ;
        RECT 47.455 94.675 47.785 95.115 ;
        RECT 45.135 94.355 47.150 94.525 ;
        RECT 47.955 94.495 48.130 94.945 ;
        RECT 42.395 93.555 43.145 93.805 ;
        RECT 43.315 93.555 44.075 93.805 ;
        RECT 41.020 93.115 41.685 93.285 ;
        RECT 41.945 93.135 42.805 93.385 ;
        RECT 42.975 93.195 44.075 93.365 ;
        RECT 41.015 92.565 41.345 92.945 ;
        RECT 41.515 92.825 41.685 93.115 ;
        RECT 42.055 92.945 42.385 92.965 ;
        RECT 42.975 92.945 43.225 93.195 ;
        RECT 42.055 92.735 43.225 92.945 ;
        RECT 43.395 92.565 43.565 93.025 ;
        RECT 43.735 92.735 44.075 93.195 ;
        RECT 44.245 92.565 44.535 93.290 ;
        RECT 44.705 93.285 44.875 93.975 ;
        RECT 45.135 93.805 45.305 94.355 ;
        RECT 45.045 93.475 45.305 93.805 ;
        RECT 44.705 92.820 45.045 93.285 ;
        RECT 45.475 93.145 45.815 94.175 ;
        RECT 46.005 93.075 46.275 94.175 ;
        RECT 44.710 92.775 45.045 92.820 ;
        RECT 45.215 92.565 45.545 92.945 ;
        RECT 46.005 92.905 46.315 93.075 ;
        RECT 46.005 92.900 46.275 92.905 ;
        RECT 46.500 92.900 46.780 94.175 ;
        RECT 46.980 93.065 47.150 94.355 ;
        RECT 47.500 94.325 48.130 94.495 ;
        RECT 48.475 94.495 48.645 94.925 ;
        RECT 48.815 94.665 49.145 95.115 ;
        RECT 47.500 93.805 47.670 94.325 ;
        RECT 48.475 94.265 49.150 94.495 ;
        RECT 47.320 93.475 47.670 93.805 ;
        RECT 47.850 93.475 48.215 94.155 ;
        RECT 47.500 93.305 47.670 93.475 ;
        RECT 47.500 93.135 48.130 93.305 ;
        RECT 48.445 93.245 48.745 94.095 ;
        RECT 48.915 93.615 49.150 94.265 ;
        RECT 49.320 93.955 49.605 94.900 ;
        RECT 49.785 94.645 50.470 95.115 ;
        RECT 49.780 94.125 50.475 94.435 ;
        RECT 50.650 94.060 50.955 94.845 ;
        RECT 51.235 94.495 51.405 94.925 ;
        RECT 51.575 94.665 51.905 95.115 ;
        RECT 51.235 94.265 51.910 94.495 ;
        RECT 49.320 93.805 50.180 93.955 ;
        RECT 49.320 93.785 50.605 93.805 ;
        RECT 48.915 93.285 49.450 93.615 ;
        RECT 49.620 93.425 50.605 93.785 ;
        RECT 48.915 93.135 49.135 93.285 ;
        RECT 46.980 92.735 47.210 93.065 ;
        RECT 47.455 92.565 47.785 92.945 ;
        RECT 47.955 92.735 48.130 93.135 ;
        RECT 48.390 92.565 48.725 93.070 ;
        RECT 48.895 92.760 49.135 93.135 ;
        RECT 49.620 93.090 49.790 93.425 ;
        RECT 50.780 93.255 50.955 94.060 ;
        RECT 49.415 92.895 49.790 93.090 ;
        RECT 49.415 92.750 49.585 92.895 ;
        RECT 50.150 92.565 50.545 93.060 ;
        RECT 50.715 92.735 50.955 93.255 ;
        RECT 51.205 93.245 51.505 94.095 ;
        RECT 51.675 93.615 51.910 94.265 ;
        RECT 52.080 93.955 52.365 94.900 ;
        RECT 52.545 94.645 53.230 95.115 ;
        RECT 52.540 94.125 53.235 94.435 ;
        RECT 53.410 94.060 53.715 94.845 ;
        RECT 52.080 93.805 52.940 93.955 ;
        RECT 52.080 93.785 53.365 93.805 ;
        RECT 51.675 93.285 52.210 93.615 ;
        RECT 52.380 93.425 53.365 93.785 ;
        RECT 51.675 93.135 51.895 93.285 ;
        RECT 51.150 92.565 51.485 93.070 ;
        RECT 51.655 92.760 51.895 93.135 ;
        RECT 52.380 93.090 52.550 93.425 ;
        RECT 53.540 93.255 53.715 94.060 ;
        RECT 54.980 94.105 55.280 94.945 ;
        RECT 55.475 94.275 55.725 95.115 ;
        RECT 56.315 94.525 57.120 94.945 ;
        RECT 55.895 94.355 57.460 94.525 ;
        RECT 55.895 94.105 56.065 94.355 ;
        RECT 54.980 93.935 56.065 94.105 ;
        RECT 54.825 93.475 55.155 93.765 ;
        RECT 55.325 93.305 55.495 93.935 ;
        RECT 56.235 93.805 56.555 94.185 ;
        RECT 56.745 94.095 57.120 94.185 ;
        RECT 56.725 93.925 57.120 94.095 ;
        RECT 57.290 94.105 57.460 94.355 ;
        RECT 57.630 94.275 57.960 95.115 ;
        RECT 58.130 94.355 58.795 94.945 ;
        RECT 57.290 93.935 58.210 94.105 ;
        RECT 55.665 93.555 55.995 93.765 ;
        RECT 56.175 93.555 56.555 93.805 ;
        RECT 56.745 93.765 57.120 93.925 ;
        RECT 58.040 93.765 58.210 93.935 ;
        RECT 56.745 93.555 57.230 93.765 ;
        RECT 57.420 93.555 57.870 93.765 ;
        RECT 58.040 93.555 58.375 93.765 ;
        RECT 58.545 93.385 58.795 94.355 ;
        RECT 58.965 93.975 59.245 95.115 ;
        RECT 59.415 93.965 59.745 94.945 ;
        RECT 59.915 93.975 60.175 95.115 ;
        RECT 61.355 94.445 61.525 94.945 ;
        RECT 61.695 94.615 62.025 95.115 ;
        RECT 61.355 94.275 62.020 94.445 ;
        RECT 58.975 93.535 59.310 93.805 ;
        RECT 52.175 92.895 52.550 93.090 ;
        RECT 52.175 92.750 52.345 92.895 ;
        RECT 52.910 92.565 53.305 93.060 ;
        RECT 53.475 92.735 53.715 93.255 ;
        RECT 54.985 93.125 55.495 93.305 ;
        RECT 55.900 93.215 57.600 93.385 ;
        RECT 55.900 93.125 56.285 93.215 ;
        RECT 54.985 92.735 55.315 93.125 ;
        RECT 55.485 92.785 56.670 92.955 ;
        RECT 56.930 92.565 57.100 93.035 ;
        RECT 57.270 92.750 57.600 93.215 ;
        RECT 57.770 92.565 57.940 93.385 ;
        RECT 58.110 92.745 58.795 93.385 ;
        RECT 59.480 93.365 59.650 93.965 ;
        RECT 59.820 93.555 60.155 93.805 ;
        RECT 61.270 93.455 61.620 94.105 ;
        RECT 58.965 92.565 59.275 93.365 ;
        RECT 59.480 92.735 60.175 93.365 ;
        RECT 61.790 93.285 62.020 94.275 ;
        RECT 61.355 93.115 62.020 93.285 ;
        RECT 61.355 92.825 61.525 93.115 ;
        RECT 61.695 92.565 62.025 92.945 ;
        RECT 62.195 92.825 62.380 94.945 ;
        RECT 62.620 94.655 62.885 95.115 ;
        RECT 63.055 94.520 63.305 94.945 ;
        RECT 63.515 94.670 64.620 94.840 ;
        RECT 63.000 94.390 63.305 94.520 ;
        RECT 62.550 93.195 62.830 94.145 ;
        RECT 63.000 93.285 63.170 94.390 ;
        RECT 63.340 93.605 63.580 94.200 ;
        RECT 63.750 94.135 64.280 94.500 ;
        RECT 63.750 93.435 63.920 94.135 ;
        RECT 64.450 94.055 64.620 94.670 ;
        RECT 64.790 94.315 64.960 95.115 ;
        RECT 65.130 94.615 65.380 94.945 ;
        RECT 65.605 94.645 66.490 94.815 ;
        RECT 64.450 93.965 64.960 94.055 ;
        RECT 63.000 93.155 63.225 93.285 ;
        RECT 63.395 93.215 63.920 93.435 ;
        RECT 64.090 93.795 64.960 93.965 ;
        RECT 62.635 92.565 62.885 93.025 ;
        RECT 63.055 93.015 63.225 93.155 ;
        RECT 64.090 93.015 64.260 93.795 ;
        RECT 64.790 93.725 64.960 93.795 ;
        RECT 64.470 93.545 64.670 93.575 ;
        RECT 65.130 93.545 65.300 94.615 ;
        RECT 65.470 93.725 65.660 94.445 ;
        RECT 64.470 93.245 65.300 93.545 ;
        RECT 65.830 93.515 66.150 94.475 ;
        RECT 63.055 92.845 63.390 93.015 ;
        RECT 63.585 92.845 64.260 93.015 ;
        RECT 64.580 92.565 64.950 93.065 ;
        RECT 65.130 93.015 65.300 93.245 ;
        RECT 65.685 93.185 66.150 93.515 ;
        RECT 66.320 93.805 66.490 94.645 ;
        RECT 66.670 94.615 66.985 95.115 ;
        RECT 67.215 94.385 67.555 94.945 ;
        RECT 66.660 94.010 67.555 94.385 ;
        RECT 67.725 94.105 67.895 95.115 ;
        RECT 67.365 93.805 67.555 94.010 ;
        RECT 68.065 94.055 68.395 94.900 ;
        RECT 68.065 93.975 68.455 94.055 ;
        RECT 68.240 93.925 68.455 93.975 ;
        RECT 66.320 93.475 67.195 93.805 ;
        RECT 67.365 93.475 68.115 93.805 ;
        RECT 66.320 93.015 66.490 93.475 ;
        RECT 67.365 93.305 67.565 93.475 ;
        RECT 68.285 93.345 68.455 93.925 ;
        RECT 68.230 93.305 68.455 93.345 ;
        RECT 65.130 92.845 65.535 93.015 ;
        RECT 65.705 92.845 66.490 93.015 ;
        RECT 66.765 92.565 66.975 93.095 ;
        RECT 67.235 92.780 67.565 93.305 ;
        RECT 68.075 93.220 68.455 93.305 ;
        RECT 68.625 94.040 68.895 94.945 ;
        RECT 69.065 94.355 69.395 95.115 ;
        RECT 69.575 94.185 69.745 94.945 ;
        RECT 68.625 93.240 68.795 94.040 ;
        RECT 69.080 94.015 69.745 94.185 ;
        RECT 69.080 93.870 69.250 94.015 ;
        RECT 70.005 93.950 70.295 95.115 ;
        RECT 71.390 94.165 71.655 94.935 ;
        RECT 71.825 94.395 72.155 95.115 ;
        RECT 72.345 94.575 72.605 94.935 ;
        RECT 72.775 94.745 73.105 95.115 ;
        RECT 73.275 94.575 73.535 94.935 ;
        RECT 72.345 94.345 73.535 94.575 ;
        RECT 74.105 94.165 74.395 94.935 ;
        RECT 68.965 93.540 69.250 93.870 ;
        RECT 69.080 93.285 69.250 93.540 ;
        RECT 69.485 93.465 69.815 93.835 ;
        RECT 67.735 92.565 67.905 93.175 ;
        RECT 68.075 92.785 68.405 93.220 ;
        RECT 68.625 92.735 68.885 93.240 ;
        RECT 69.080 93.115 69.745 93.285 ;
        RECT 69.065 92.565 69.395 92.945 ;
        RECT 69.575 92.735 69.745 93.115 ;
        RECT 70.005 92.565 70.295 93.290 ;
        RECT 71.390 92.745 71.725 94.165 ;
        RECT 71.900 93.985 74.395 94.165 ;
        RECT 71.900 93.295 72.125 93.985 ;
        RECT 74.605 93.975 74.945 94.945 ;
        RECT 75.115 93.975 75.285 95.115 ;
        RECT 75.555 94.315 75.805 95.115 ;
        RECT 76.450 94.145 76.780 94.945 ;
        RECT 77.080 94.315 77.410 95.115 ;
        RECT 77.580 94.145 77.910 94.945 ;
        RECT 75.475 93.975 77.910 94.145 ;
        RECT 78.285 94.265 78.545 94.945 ;
        RECT 78.715 94.335 78.965 95.115 ;
        RECT 79.215 94.565 79.465 94.945 ;
        RECT 79.635 94.735 79.990 95.115 ;
        RECT 80.995 94.725 81.330 94.945 ;
        RECT 80.595 94.565 80.825 94.605 ;
        RECT 79.215 94.365 80.825 94.565 ;
        RECT 79.215 94.355 80.050 94.365 ;
        RECT 80.640 94.275 80.825 94.365 ;
        RECT 72.325 93.475 72.605 93.805 ;
        RECT 72.785 93.475 73.360 93.805 ;
        RECT 73.540 93.475 73.975 93.805 ;
        RECT 74.155 93.475 74.425 93.805 ;
        RECT 74.605 93.365 74.780 93.975 ;
        RECT 75.475 93.725 75.645 93.975 ;
        RECT 74.950 93.555 75.645 93.725 ;
        RECT 75.820 93.555 76.240 93.755 ;
        RECT 76.410 93.555 76.740 93.755 ;
        RECT 76.910 93.555 77.240 93.755 ;
        RECT 71.900 93.105 74.385 93.295 ;
        RECT 71.905 92.565 72.650 92.935 ;
        RECT 73.215 92.745 73.470 93.105 ;
        RECT 73.650 92.565 73.980 92.935 ;
        RECT 74.160 92.745 74.385 93.105 ;
        RECT 74.605 92.735 74.945 93.365 ;
        RECT 75.115 92.565 75.365 93.365 ;
        RECT 75.555 93.215 76.780 93.385 ;
        RECT 75.555 92.735 75.885 93.215 ;
        RECT 76.055 92.565 76.280 93.025 ;
        RECT 76.450 92.735 76.780 93.215 ;
        RECT 77.410 93.345 77.580 93.975 ;
        RECT 77.765 93.555 78.115 93.805 ;
        RECT 77.410 92.735 77.910 93.345 ;
        RECT 78.285 93.075 78.455 94.265 ;
        RECT 80.155 94.165 80.485 94.195 ;
        RECT 78.685 94.105 80.485 94.165 ;
        RECT 81.075 94.105 81.330 94.725 ;
        RECT 78.625 93.995 81.330 94.105 ;
        RECT 78.625 93.960 78.825 93.995 ;
        RECT 78.625 93.385 78.795 93.960 ;
        RECT 80.155 93.935 81.330 93.995 ;
        RECT 81.965 94.025 83.175 95.115 ;
        RECT 79.025 93.520 79.435 93.825 ;
        RECT 79.605 93.555 79.935 93.765 ;
        RECT 78.625 93.265 78.895 93.385 ;
        RECT 78.625 93.220 79.470 93.265 ;
        RECT 78.715 93.095 79.470 93.220 ;
        RECT 79.725 93.155 79.935 93.555 ;
        RECT 80.180 93.555 80.655 93.765 ;
        RECT 80.845 93.555 81.335 93.755 ;
        RECT 80.180 93.155 80.400 93.555 ;
        RECT 81.965 93.485 82.485 94.025 ;
        RECT 78.285 93.065 78.515 93.075 ;
        RECT 78.285 92.735 78.545 93.065 ;
        RECT 79.300 92.945 79.470 93.095 ;
        RECT 78.715 92.565 79.045 92.925 ;
        RECT 79.300 92.735 80.600 92.945 ;
        RECT 80.875 92.565 81.330 93.330 ;
        RECT 82.655 93.315 83.175 93.855 ;
        RECT 81.965 92.565 83.175 93.315 ;
        RECT 5.520 92.395 83.260 92.565 ;
        RECT 5.605 91.645 6.815 92.395 ;
        RECT 5.605 91.105 6.125 91.645 ;
        RECT 6.985 91.625 10.495 92.395 ;
        RECT 6.295 90.935 6.815 91.475 ;
        RECT 6.985 91.105 8.635 91.625 ;
        RECT 11.605 91.585 11.845 92.395 ;
        RECT 12.015 91.585 12.345 92.225 ;
        RECT 12.515 91.585 12.785 92.395 ;
        RECT 12.965 91.850 18.310 92.395 ;
        RECT 19.470 92.005 21.480 92.175 ;
        RECT 8.805 90.935 10.495 91.455 ;
        RECT 11.585 91.155 11.935 91.405 ;
        RECT 12.105 90.985 12.275 91.585 ;
        RECT 12.445 91.155 12.795 91.405 ;
        RECT 14.550 91.020 14.890 91.850 ;
        RECT 19.405 91.575 21.060 91.835 ;
        RECT 21.230 91.745 21.480 92.005 ;
        RECT 21.670 91.925 21.940 92.395 ;
        RECT 22.110 91.755 22.440 92.225 ;
        RECT 22.610 91.925 22.780 92.395 ;
        RECT 22.950 91.755 23.280 92.225 ;
        RECT 23.450 91.925 23.620 92.395 ;
        RECT 23.790 91.755 24.120 92.225 ;
        RECT 24.290 91.925 24.460 92.395 ;
        RECT 24.630 91.755 24.960 92.225 ;
        RECT 22.010 91.745 24.960 91.755 ;
        RECT 21.230 91.575 24.960 91.745 ;
        RECT 25.130 91.575 25.405 92.395 ;
        RECT 25.580 91.755 25.910 92.225 ;
        RECT 26.080 91.925 26.250 92.395 ;
        RECT 26.420 91.755 26.750 92.225 ;
        RECT 26.920 91.925 27.090 92.395 ;
        RECT 27.260 92.005 29.270 92.225 ;
        RECT 27.260 91.755 27.510 92.005 ;
        RECT 25.580 91.575 27.510 91.755 ;
        RECT 27.680 91.575 29.355 91.835 ;
        RECT 19.405 91.545 19.635 91.575 ;
        RECT 5.605 89.845 6.815 90.935 ;
        RECT 6.985 89.845 10.495 90.935 ;
        RECT 11.595 90.815 12.275 90.985 ;
        RECT 11.595 90.030 11.925 90.815 ;
        RECT 12.455 89.845 12.785 90.985 ;
        RECT 16.370 90.280 16.720 91.530 ;
        RECT 19.405 91.035 19.625 91.545 ;
        RECT 19.795 91.205 21.840 91.405 ;
        RECT 22.010 91.205 23.880 91.405 ;
        RECT 24.050 91.205 27.265 91.405 ;
        RECT 27.585 91.205 28.950 91.405 ;
        RECT 21.670 91.035 21.840 91.205 ;
        RECT 23.710 91.035 23.880 91.205 ;
        RECT 27.585 91.035 27.755 91.205 ;
        RECT 29.120 91.035 29.355 91.575 ;
        RECT 29.525 91.625 31.195 92.395 ;
        RECT 31.365 91.670 31.655 92.395 ;
        RECT 29.525 91.105 30.275 91.625 ;
        RECT 31.825 91.595 32.135 92.395 ;
        RECT 32.340 91.595 33.035 92.225 ;
        RECT 19.405 90.815 21.480 91.035 ;
        RECT 21.670 90.865 23.540 91.035 ;
        RECT 23.710 90.865 27.755 91.035 ;
        RECT 28.140 90.865 29.355 91.035 ;
        RECT 30.445 90.935 31.195 91.455 ;
        RECT 31.835 91.155 32.170 91.425 ;
        RECT 12.965 89.845 18.310 90.280 ;
        RECT 19.405 90.015 19.760 90.815 ;
        RECT 19.930 89.845 20.180 90.645 ;
        RECT 20.350 90.015 20.600 90.815 ;
        RECT 21.190 90.695 21.480 90.815 ;
        RECT 28.140 90.695 28.390 90.865 ;
        RECT 20.770 89.845 21.020 90.645 ;
        RECT 21.190 90.435 23.280 90.695 ;
        RECT 23.450 90.475 25.405 90.695 ;
        RECT 21.190 90.015 21.480 90.435 ;
        RECT 23.450 90.265 23.660 90.475 ;
        RECT 21.690 90.015 23.660 90.265 ;
        RECT 23.830 89.845 24.080 90.305 ;
        RECT 24.250 90.015 24.500 90.475 ;
        RECT 24.670 89.845 24.920 90.305 ;
        RECT 25.090 90.015 25.405 90.475 ;
        RECT 25.620 90.475 28.390 90.695 ;
        RECT 25.620 90.015 25.870 90.475 ;
        RECT 26.040 89.845 26.290 90.305 ;
        RECT 26.460 90.015 26.710 90.475 ;
        RECT 26.880 89.845 27.130 90.305 ;
        RECT 27.300 90.015 27.550 90.475 ;
        RECT 27.720 89.845 27.970 90.305 ;
        RECT 28.140 90.015 28.390 90.475 ;
        RECT 28.560 89.845 28.810 90.645 ;
        RECT 28.980 90.015 29.355 90.865 ;
        RECT 29.525 89.845 31.195 90.935 ;
        RECT 31.365 89.845 31.655 91.010 ;
        RECT 32.340 90.995 32.510 91.595 ;
        RECT 33.265 91.575 33.475 92.395 ;
        RECT 33.645 91.595 33.975 92.225 ;
        RECT 32.680 91.155 33.015 91.405 ;
        RECT 33.645 90.995 33.895 91.595 ;
        RECT 34.145 91.575 34.375 92.395 ;
        RECT 35.595 91.845 35.765 92.135 ;
        RECT 35.935 92.015 36.265 92.395 ;
        RECT 35.595 91.675 36.260 91.845 ;
        RECT 34.065 91.155 34.395 91.405 ;
        RECT 31.825 89.845 32.105 90.985 ;
        RECT 32.275 90.015 32.605 90.995 ;
        RECT 32.775 89.845 33.035 90.985 ;
        RECT 33.265 89.845 33.475 90.985 ;
        RECT 33.645 90.015 33.975 90.995 ;
        RECT 34.145 89.845 34.375 90.985 ;
        RECT 35.510 90.855 35.860 91.505 ;
        RECT 36.030 90.685 36.260 91.675 ;
        RECT 35.595 90.515 36.260 90.685 ;
        RECT 35.595 90.015 35.765 90.515 ;
        RECT 35.935 89.845 36.265 90.345 ;
        RECT 36.435 90.015 36.620 92.135 ;
        RECT 36.875 91.935 37.125 92.395 ;
        RECT 37.295 91.945 37.630 92.115 ;
        RECT 37.825 91.945 38.500 92.115 ;
        RECT 37.295 91.805 37.465 91.945 ;
        RECT 36.790 90.815 37.070 91.765 ;
        RECT 37.240 91.675 37.465 91.805 ;
        RECT 37.240 90.570 37.410 91.675 ;
        RECT 37.635 91.525 38.160 91.745 ;
        RECT 37.580 90.760 37.820 91.355 ;
        RECT 37.990 90.825 38.160 91.525 ;
        RECT 38.330 91.165 38.500 91.945 ;
        RECT 38.820 91.895 39.190 92.395 ;
        RECT 39.370 91.945 39.775 92.115 ;
        RECT 39.945 91.945 40.730 92.115 ;
        RECT 39.370 91.715 39.540 91.945 ;
        RECT 38.710 91.415 39.540 91.715 ;
        RECT 39.925 91.445 40.390 91.775 ;
        RECT 38.710 91.385 38.910 91.415 ;
        RECT 39.030 91.165 39.200 91.235 ;
        RECT 38.330 90.995 39.200 91.165 ;
        RECT 38.690 90.905 39.200 90.995 ;
        RECT 37.240 90.440 37.545 90.570 ;
        RECT 37.990 90.460 38.520 90.825 ;
        RECT 36.860 89.845 37.125 90.305 ;
        RECT 37.295 90.015 37.545 90.440 ;
        RECT 38.690 90.290 38.860 90.905 ;
        RECT 37.755 90.120 38.860 90.290 ;
        RECT 39.030 89.845 39.200 90.645 ;
        RECT 39.370 90.345 39.540 91.415 ;
        RECT 39.710 90.515 39.900 91.235 ;
        RECT 40.070 90.485 40.390 91.445 ;
        RECT 40.560 91.485 40.730 91.945 ;
        RECT 41.005 91.865 41.215 92.395 ;
        RECT 41.475 91.655 41.805 92.180 ;
        RECT 41.975 91.785 42.145 92.395 ;
        RECT 42.315 91.740 42.645 92.175 ;
        RECT 42.870 91.890 43.205 92.395 ;
        RECT 43.375 91.825 43.615 92.200 ;
        RECT 43.895 92.065 44.065 92.210 ;
        RECT 43.895 91.870 44.270 92.065 ;
        RECT 44.630 91.900 45.025 92.395 ;
        RECT 42.315 91.655 42.695 91.740 ;
        RECT 41.605 91.485 41.805 91.655 ;
        RECT 42.470 91.615 42.695 91.655 ;
        RECT 40.560 91.155 41.435 91.485 ;
        RECT 41.605 91.155 42.355 91.485 ;
        RECT 39.370 90.015 39.620 90.345 ;
        RECT 40.560 90.315 40.730 91.155 ;
        RECT 41.605 90.950 41.795 91.155 ;
        RECT 42.525 91.035 42.695 91.615 ;
        RECT 42.480 90.985 42.695 91.035 ;
        RECT 40.900 90.575 41.795 90.950 ;
        RECT 42.305 90.905 42.695 90.985 ;
        RECT 39.845 90.145 40.730 90.315 ;
        RECT 40.910 89.845 41.225 90.345 ;
        RECT 41.455 90.015 41.795 90.575 ;
        RECT 41.965 89.845 42.135 90.855 ;
        RECT 42.305 90.060 42.635 90.905 ;
        RECT 42.925 90.865 43.225 91.715 ;
        RECT 43.395 91.675 43.615 91.825 ;
        RECT 43.395 91.345 43.930 91.675 ;
        RECT 44.100 91.535 44.270 91.870 ;
        RECT 45.195 91.705 45.435 92.225 ;
        RECT 43.395 90.695 43.630 91.345 ;
        RECT 44.100 91.175 45.085 91.535 ;
        RECT 42.955 90.465 43.630 90.695 ;
        RECT 43.800 91.155 45.085 91.175 ;
        RECT 43.800 91.005 44.660 91.155 ;
        RECT 42.955 90.035 43.125 90.465 ;
        RECT 43.295 89.845 43.625 90.295 ;
        RECT 43.800 90.060 44.085 91.005 ;
        RECT 45.260 90.900 45.435 91.705 ;
        RECT 46.545 91.765 46.885 92.225 ;
        RECT 47.055 91.935 47.225 92.395 ;
        RECT 47.395 92.015 48.565 92.225 ;
        RECT 48.845 92.015 49.735 92.185 ;
        RECT 47.395 91.765 47.645 92.015 ;
        RECT 48.235 91.995 48.565 92.015 ;
        RECT 46.545 91.595 47.645 91.765 ;
        RECT 47.815 91.575 48.675 91.825 ;
        RECT 46.545 91.155 47.305 91.405 ;
        RECT 47.475 91.155 48.225 91.405 ;
        RECT 48.395 90.985 48.675 91.575 ;
        RECT 48.845 91.460 49.395 91.845 ;
        RECT 49.565 91.290 49.735 92.015 ;
        RECT 44.260 90.525 44.955 90.835 ;
        RECT 44.265 89.845 44.950 90.315 ;
        RECT 45.130 90.115 45.435 90.900 ;
        RECT 46.545 89.845 46.805 90.985 ;
        RECT 46.975 90.815 48.675 90.985 ;
        RECT 48.845 91.220 49.735 91.290 ;
        RECT 49.905 91.715 50.125 92.175 ;
        RECT 50.295 91.855 50.545 92.395 ;
        RECT 50.715 91.745 50.975 92.225 ;
        RECT 51.165 91.885 51.405 92.395 ;
        RECT 51.575 91.885 51.865 92.225 ;
        RECT 52.095 91.885 52.410 92.395 ;
        RECT 49.905 91.690 50.155 91.715 ;
        RECT 49.905 91.265 50.235 91.690 ;
        RECT 48.845 91.195 49.740 91.220 ;
        RECT 48.845 91.180 49.750 91.195 ;
        RECT 48.845 91.165 49.755 91.180 ;
        RECT 48.845 91.160 49.765 91.165 ;
        RECT 48.845 91.150 49.770 91.160 ;
        RECT 48.845 91.140 49.775 91.150 ;
        RECT 48.845 91.135 49.785 91.140 ;
        RECT 48.845 91.125 49.795 91.135 ;
        RECT 48.845 91.120 49.805 91.125 ;
        RECT 46.975 90.015 47.305 90.815 ;
        RECT 47.475 89.845 47.645 90.645 ;
        RECT 47.815 90.015 48.145 90.815 ;
        RECT 48.845 90.670 49.105 91.120 ;
        RECT 49.470 91.115 49.805 91.120 ;
        RECT 49.470 91.110 49.820 91.115 ;
        RECT 49.470 91.100 49.835 91.110 ;
        RECT 49.470 91.095 49.860 91.100 ;
        RECT 50.405 91.095 50.635 91.490 ;
        RECT 49.470 91.090 50.635 91.095 ;
        RECT 49.500 91.055 50.635 91.090 ;
        RECT 49.535 91.030 50.635 91.055 ;
        RECT 49.565 91.000 50.635 91.030 ;
        RECT 49.585 90.970 50.635 91.000 ;
        RECT 49.605 90.940 50.635 90.970 ;
        RECT 49.675 90.930 50.635 90.940 ;
        RECT 49.700 90.920 50.635 90.930 ;
        RECT 49.720 90.905 50.635 90.920 ;
        RECT 49.740 90.890 50.635 90.905 ;
        RECT 49.745 90.880 50.530 90.890 ;
        RECT 49.760 90.845 50.530 90.880 ;
        RECT 48.315 89.845 48.570 90.645 ;
        RECT 49.275 90.525 49.605 90.770 ;
        RECT 49.775 90.595 50.530 90.845 ;
        RECT 50.805 90.715 50.975 91.745 ;
        RECT 51.210 91.375 51.405 91.715 ;
        RECT 51.205 91.205 51.405 91.375 ;
        RECT 51.210 91.155 51.405 91.205 ;
        RECT 51.575 90.985 51.755 91.885 ;
        RECT 52.580 91.825 52.750 92.095 ;
        RECT 52.920 91.995 53.250 92.395 ;
        RECT 51.925 91.155 52.335 91.715 ;
        RECT 52.580 91.655 53.275 91.825 ;
        RECT 54.385 91.665 54.675 92.395 ;
        RECT 52.505 90.985 52.675 91.485 ;
        RECT 49.275 90.500 49.460 90.525 ;
        RECT 48.845 90.400 49.460 90.500 ;
        RECT 48.845 89.845 49.450 90.400 ;
        RECT 49.625 90.015 50.105 90.355 ;
        RECT 50.275 89.845 50.530 90.390 ;
        RECT 50.700 90.015 50.975 90.715 ;
        RECT 51.215 90.815 52.675 90.985 ;
        RECT 51.215 90.640 51.575 90.815 ;
        RECT 52.845 90.645 53.275 91.655 ;
        RECT 54.375 91.155 54.675 91.485 ;
        RECT 54.855 91.465 55.085 92.105 ;
        RECT 55.265 91.845 55.575 92.215 ;
        RECT 55.755 92.025 56.425 92.395 ;
        RECT 55.265 91.645 56.495 91.845 ;
        RECT 54.855 91.155 55.380 91.465 ;
        RECT 55.560 91.155 56.025 91.465 ;
        RECT 56.205 90.975 56.495 91.645 ;
        RECT 52.160 89.845 52.330 90.645 ;
        RECT 52.500 90.475 53.275 90.645 ;
        RECT 54.385 90.735 55.545 90.975 ;
        RECT 52.500 90.015 52.830 90.475 ;
        RECT 53.000 89.845 53.170 90.305 ;
        RECT 54.385 90.025 54.645 90.735 ;
        RECT 54.815 89.845 55.145 90.555 ;
        RECT 55.315 90.025 55.545 90.735 ;
        RECT 55.725 90.755 56.495 90.975 ;
        RECT 55.725 90.025 55.995 90.755 ;
        RECT 56.175 89.845 56.515 90.575 ;
        RECT 56.685 90.025 56.945 92.215 ;
        RECT 57.125 91.670 57.415 92.395 ;
        RECT 57.585 91.625 59.255 92.395 ;
        RECT 59.515 91.845 59.685 92.135 ;
        RECT 59.855 92.015 60.185 92.395 ;
        RECT 59.515 91.675 60.180 91.845 ;
        RECT 57.585 91.105 58.335 91.625 ;
        RECT 57.125 89.845 57.415 91.010 ;
        RECT 58.505 90.935 59.255 91.455 ;
        RECT 57.585 89.845 59.255 90.935 ;
        RECT 59.430 90.855 59.780 91.505 ;
        RECT 59.950 90.685 60.180 91.675 ;
        RECT 59.515 90.515 60.180 90.685 ;
        RECT 59.515 90.015 59.685 90.515 ;
        RECT 59.855 89.845 60.185 90.345 ;
        RECT 60.355 90.015 60.540 92.135 ;
        RECT 60.795 91.935 61.045 92.395 ;
        RECT 61.215 91.945 61.550 92.115 ;
        RECT 61.745 91.945 62.420 92.115 ;
        RECT 61.215 91.805 61.385 91.945 ;
        RECT 60.710 90.815 60.990 91.765 ;
        RECT 61.160 91.675 61.385 91.805 ;
        RECT 61.160 90.570 61.330 91.675 ;
        RECT 61.555 91.525 62.080 91.745 ;
        RECT 61.500 90.760 61.740 91.355 ;
        RECT 61.910 90.825 62.080 91.525 ;
        RECT 62.250 91.165 62.420 91.945 ;
        RECT 62.740 91.895 63.110 92.395 ;
        RECT 63.290 91.945 63.695 92.115 ;
        RECT 63.865 91.945 64.650 92.115 ;
        RECT 63.290 91.715 63.460 91.945 ;
        RECT 62.630 91.415 63.460 91.715 ;
        RECT 63.845 91.445 64.310 91.775 ;
        RECT 62.630 91.385 62.830 91.415 ;
        RECT 62.950 91.165 63.120 91.235 ;
        RECT 62.250 90.995 63.120 91.165 ;
        RECT 62.610 90.905 63.120 90.995 ;
        RECT 61.160 90.440 61.465 90.570 ;
        RECT 61.910 90.460 62.440 90.825 ;
        RECT 60.780 89.845 61.045 90.305 ;
        RECT 61.215 90.015 61.465 90.440 ;
        RECT 62.610 90.290 62.780 90.905 ;
        RECT 61.675 90.120 62.780 90.290 ;
        RECT 62.950 89.845 63.120 90.645 ;
        RECT 63.290 90.345 63.460 91.415 ;
        RECT 63.630 90.515 63.820 91.235 ;
        RECT 63.990 90.485 64.310 91.445 ;
        RECT 64.480 91.485 64.650 91.945 ;
        RECT 64.925 91.865 65.135 92.395 ;
        RECT 65.395 91.655 65.725 92.180 ;
        RECT 65.895 91.785 66.065 92.395 ;
        RECT 66.235 91.740 66.565 92.175 ;
        RECT 66.235 91.655 66.615 91.740 ;
        RECT 65.525 91.485 65.725 91.655 ;
        RECT 66.390 91.615 66.615 91.655 ;
        RECT 64.480 91.155 65.355 91.485 ;
        RECT 65.525 91.155 66.275 91.485 ;
        RECT 63.290 90.015 63.540 90.345 ;
        RECT 64.480 90.315 64.650 91.155 ;
        RECT 65.525 90.950 65.715 91.155 ;
        RECT 66.445 91.035 66.615 91.615 ;
        RECT 66.400 90.985 66.615 91.035 ;
        RECT 64.820 90.575 65.715 90.950 ;
        RECT 66.225 90.905 66.615 90.985 ;
        RECT 66.785 91.655 67.170 92.225 ;
        RECT 67.340 91.935 67.665 92.395 ;
        RECT 68.185 91.765 68.465 92.225 ;
        RECT 66.785 90.985 67.065 91.655 ;
        RECT 67.340 91.595 68.465 91.765 ;
        RECT 67.340 91.485 67.790 91.595 ;
        RECT 67.235 91.155 67.790 91.485 ;
        RECT 68.655 91.425 69.055 92.225 ;
        RECT 69.455 91.935 69.725 92.395 ;
        RECT 69.895 91.765 70.180 92.225 ;
        RECT 63.765 90.145 64.650 90.315 ;
        RECT 64.830 89.845 65.145 90.345 ;
        RECT 65.375 90.015 65.715 90.575 ;
        RECT 65.885 89.845 66.055 90.855 ;
        RECT 66.225 90.060 66.555 90.905 ;
        RECT 66.785 90.015 67.170 90.985 ;
        RECT 67.340 90.695 67.790 91.155 ;
        RECT 67.960 90.865 69.055 91.425 ;
        RECT 67.340 90.475 68.465 90.695 ;
        RECT 67.340 89.845 67.665 90.305 ;
        RECT 68.185 90.015 68.465 90.475 ;
        RECT 68.655 90.015 69.055 90.865 ;
        RECT 69.225 91.595 70.180 91.765 ;
        RECT 69.225 90.695 69.435 91.595 ;
        RECT 70.470 91.555 70.730 92.395 ;
        RECT 70.905 91.650 71.160 92.225 ;
        RECT 71.330 92.015 71.660 92.395 ;
        RECT 71.875 91.845 72.045 92.225 ;
        RECT 71.330 91.675 72.045 91.845 ;
        RECT 72.395 91.845 72.565 92.135 ;
        RECT 72.735 92.015 73.065 92.395 ;
        RECT 72.395 91.675 73.060 91.845 ;
        RECT 69.605 90.865 70.295 91.425 ;
        RECT 69.225 90.475 70.180 90.695 ;
        RECT 69.455 89.845 69.725 90.305 ;
        RECT 69.895 90.015 70.180 90.475 ;
        RECT 70.470 89.845 70.730 90.995 ;
        RECT 70.905 90.920 71.075 91.650 ;
        RECT 71.330 91.485 71.500 91.675 ;
        RECT 71.245 91.155 71.500 91.485 ;
        RECT 71.330 90.945 71.500 91.155 ;
        RECT 71.780 91.125 72.135 91.495 ;
        RECT 70.905 90.015 71.160 90.920 ;
        RECT 71.330 90.775 72.045 90.945 ;
        RECT 72.310 90.855 72.660 91.505 ;
        RECT 71.330 89.845 71.660 90.605 ;
        RECT 71.875 90.015 72.045 90.775 ;
        RECT 72.830 90.685 73.060 91.675 ;
        RECT 72.395 90.515 73.060 90.685 ;
        RECT 72.395 90.015 72.565 90.515 ;
        RECT 72.735 89.845 73.065 90.345 ;
        RECT 73.235 90.015 73.420 92.135 ;
        RECT 73.675 91.935 73.925 92.395 ;
        RECT 74.095 91.945 74.430 92.115 ;
        RECT 74.625 91.945 75.300 92.115 ;
        RECT 74.095 91.805 74.265 91.945 ;
        RECT 73.590 90.815 73.870 91.765 ;
        RECT 74.040 91.675 74.265 91.805 ;
        RECT 74.040 90.570 74.210 91.675 ;
        RECT 74.435 91.525 74.960 91.745 ;
        RECT 74.380 90.760 74.620 91.355 ;
        RECT 74.790 90.825 74.960 91.525 ;
        RECT 75.130 91.165 75.300 91.945 ;
        RECT 75.620 91.895 75.990 92.395 ;
        RECT 76.170 91.945 76.575 92.115 ;
        RECT 76.745 91.945 77.530 92.115 ;
        RECT 76.170 91.715 76.340 91.945 ;
        RECT 75.510 91.415 76.340 91.715 ;
        RECT 76.725 91.445 77.190 91.775 ;
        RECT 75.510 91.385 75.710 91.415 ;
        RECT 75.830 91.165 76.000 91.235 ;
        RECT 75.130 90.995 76.000 91.165 ;
        RECT 75.490 90.905 76.000 90.995 ;
        RECT 74.040 90.440 74.345 90.570 ;
        RECT 74.790 90.460 75.320 90.825 ;
        RECT 73.660 89.845 73.925 90.305 ;
        RECT 74.095 90.015 74.345 90.440 ;
        RECT 75.490 90.290 75.660 90.905 ;
        RECT 74.555 90.120 75.660 90.290 ;
        RECT 75.830 89.845 76.000 90.645 ;
        RECT 76.170 90.345 76.340 91.415 ;
        RECT 76.510 90.515 76.700 91.235 ;
        RECT 76.870 90.485 77.190 91.445 ;
        RECT 77.360 91.485 77.530 91.945 ;
        RECT 77.805 91.865 78.015 92.395 ;
        RECT 78.275 91.655 78.605 92.180 ;
        RECT 78.775 91.785 78.945 92.395 ;
        RECT 79.115 91.740 79.445 92.175 ;
        RECT 79.830 91.885 80.070 92.395 ;
        RECT 80.250 91.885 80.530 92.215 ;
        RECT 80.760 91.885 80.975 92.395 ;
        RECT 79.115 91.655 79.495 91.740 ;
        RECT 78.405 91.485 78.605 91.655 ;
        RECT 79.270 91.615 79.495 91.655 ;
        RECT 77.360 91.155 78.235 91.485 ;
        RECT 78.405 91.155 79.155 91.485 ;
        RECT 76.170 90.015 76.420 90.345 ;
        RECT 77.360 90.315 77.530 91.155 ;
        RECT 78.405 90.950 78.595 91.155 ;
        RECT 79.325 91.035 79.495 91.615 ;
        RECT 79.725 91.155 80.080 91.715 ;
        RECT 79.280 90.985 79.495 91.035 ;
        RECT 80.250 90.985 80.420 91.885 ;
        RECT 80.590 91.155 80.855 91.715 ;
        RECT 81.145 91.655 81.760 92.225 ;
        RECT 81.105 90.985 81.275 91.485 ;
        RECT 77.700 90.575 78.595 90.950 ;
        RECT 79.105 90.905 79.495 90.985 ;
        RECT 76.645 90.145 77.530 90.315 ;
        RECT 77.710 89.845 78.025 90.345 ;
        RECT 78.255 90.015 78.595 90.575 ;
        RECT 78.765 89.845 78.935 90.855 ;
        RECT 79.105 90.060 79.435 90.905 ;
        RECT 79.850 90.815 81.275 90.985 ;
        RECT 79.850 90.640 80.240 90.815 ;
        RECT 80.725 89.845 81.055 90.645 ;
        RECT 81.445 90.635 81.760 91.655 ;
        RECT 81.965 91.645 83.175 92.395 ;
        RECT 81.225 90.015 81.760 90.635 ;
        RECT 81.965 90.935 82.485 91.475 ;
        RECT 82.655 91.105 83.175 91.645 ;
        RECT 81.965 89.845 83.175 90.935 ;
        RECT 5.520 89.675 83.260 89.845 ;
        RECT 5.605 88.585 6.815 89.675 ;
        RECT 5.605 87.875 6.125 88.415 ;
        RECT 6.295 88.045 6.815 88.585 ;
        RECT 6.985 88.805 7.260 89.505 ;
        RECT 7.430 89.130 7.685 89.675 ;
        RECT 7.855 89.165 8.335 89.505 ;
        RECT 8.510 89.120 9.115 89.675 ;
        RECT 8.500 89.020 9.115 89.120 ;
        RECT 8.500 88.995 8.685 89.020 ;
        RECT 5.605 87.125 6.815 87.875 ;
        RECT 6.985 87.775 7.155 88.805 ;
        RECT 7.430 88.675 8.185 88.925 ;
        RECT 8.355 88.750 8.685 88.995 ;
        RECT 7.430 88.640 8.200 88.675 ;
        RECT 7.430 88.630 8.215 88.640 ;
        RECT 7.325 88.615 8.220 88.630 ;
        RECT 7.325 88.600 8.240 88.615 ;
        RECT 7.325 88.590 8.260 88.600 ;
        RECT 7.325 88.580 8.285 88.590 ;
        RECT 7.325 88.550 8.355 88.580 ;
        RECT 7.325 88.520 8.375 88.550 ;
        RECT 7.325 88.490 8.395 88.520 ;
        RECT 7.325 88.465 8.425 88.490 ;
        RECT 7.325 88.430 8.460 88.465 ;
        RECT 7.325 88.425 8.490 88.430 ;
        RECT 7.325 88.030 7.555 88.425 ;
        RECT 8.100 88.420 8.490 88.425 ;
        RECT 8.125 88.410 8.490 88.420 ;
        RECT 8.140 88.405 8.490 88.410 ;
        RECT 8.155 88.400 8.490 88.405 ;
        RECT 8.855 88.400 9.115 88.850 ;
        RECT 8.155 88.395 9.115 88.400 ;
        RECT 8.165 88.385 9.115 88.395 ;
        RECT 8.175 88.380 9.115 88.385 ;
        RECT 8.185 88.370 9.115 88.380 ;
        RECT 8.190 88.360 9.115 88.370 ;
        RECT 8.195 88.355 9.115 88.360 ;
        RECT 8.205 88.340 9.115 88.355 ;
        RECT 8.210 88.325 9.115 88.340 ;
        RECT 8.220 88.300 9.115 88.325 ;
        RECT 7.725 87.830 8.055 88.255 ;
        RECT 6.985 87.295 7.245 87.775 ;
        RECT 7.415 87.125 7.665 87.665 ;
        RECT 7.835 87.345 8.055 87.830 ;
        RECT 8.225 88.230 9.115 88.300 ;
        RECT 9.285 88.805 9.560 89.505 ;
        RECT 9.730 89.130 9.985 89.675 ;
        RECT 10.155 89.165 10.635 89.505 ;
        RECT 10.810 89.120 11.415 89.675 ;
        RECT 10.800 89.020 11.415 89.120 ;
        RECT 10.800 88.995 10.985 89.020 ;
        RECT 8.225 87.505 8.395 88.230 ;
        RECT 8.565 87.675 9.115 88.060 ;
        RECT 9.285 87.775 9.455 88.805 ;
        RECT 9.730 88.675 10.485 88.925 ;
        RECT 10.655 88.750 10.985 88.995 ;
        RECT 9.730 88.640 10.500 88.675 ;
        RECT 9.730 88.630 10.515 88.640 ;
        RECT 9.625 88.615 10.520 88.630 ;
        RECT 9.625 88.600 10.540 88.615 ;
        RECT 9.625 88.590 10.560 88.600 ;
        RECT 9.625 88.580 10.585 88.590 ;
        RECT 9.625 88.550 10.655 88.580 ;
        RECT 9.625 88.520 10.675 88.550 ;
        RECT 9.625 88.490 10.695 88.520 ;
        RECT 9.625 88.465 10.725 88.490 ;
        RECT 9.625 88.430 10.760 88.465 ;
        RECT 9.625 88.425 10.790 88.430 ;
        RECT 9.625 88.030 9.855 88.425 ;
        RECT 10.400 88.420 10.790 88.425 ;
        RECT 10.425 88.410 10.790 88.420 ;
        RECT 10.440 88.405 10.790 88.410 ;
        RECT 10.455 88.400 10.790 88.405 ;
        RECT 11.155 88.400 11.415 88.850 ;
        RECT 12.055 88.535 12.385 89.675 ;
        RECT 12.915 88.705 13.245 89.490 ;
        RECT 13.425 88.855 13.770 89.675 ;
        RECT 12.565 88.535 13.245 88.705 ;
        RECT 10.455 88.395 11.415 88.400 ;
        RECT 10.465 88.385 11.415 88.395 ;
        RECT 10.475 88.380 11.415 88.385 ;
        RECT 10.485 88.370 11.415 88.380 ;
        RECT 10.490 88.360 11.415 88.370 ;
        RECT 10.495 88.355 11.415 88.360 ;
        RECT 10.505 88.340 11.415 88.355 ;
        RECT 10.510 88.325 11.415 88.340 ;
        RECT 10.520 88.300 11.415 88.325 ;
        RECT 10.025 87.830 10.355 88.255 ;
        RECT 8.225 87.335 9.115 87.505 ;
        RECT 9.285 87.295 9.545 87.775 ;
        RECT 9.715 87.125 9.965 87.665 ;
        RECT 10.135 87.345 10.355 87.830 ;
        RECT 10.525 88.230 11.415 88.300 ;
        RECT 10.525 87.505 10.695 88.230 ;
        RECT 12.045 88.115 12.395 88.365 ;
        RECT 10.865 87.675 11.415 88.060 ;
        RECT 12.565 87.935 12.735 88.535 ;
        RECT 12.905 88.115 13.255 88.365 ;
        RECT 13.425 88.115 13.770 88.685 ;
        RECT 13.940 88.365 14.115 89.465 ;
        RECT 14.285 89.095 14.615 89.330 ;
        RECT 14.905 89.275 15.305 89.675 ;
        RECT 16.175 89.275 16.505 89.675 ;
        RECT 14.285 88.925 16.365 89.095 ;
        RECT 14.285 88.535 14.840 88.925 ;
        RECT 13.940 88.115 14.500 88.365 ;
        RECT 14.670 88.285 14.840 88.535 ;
        RECT 15.010 88.535 16.025 88.755 ;
        RECT 16.195 88.655 16.365 88.925 ;
        RECT 16.675 88.835 16.935 89.505 ;
        RECT 15.010 88.395 15.285 88.535 ;
        RECT 16.195 88.485 16.590 88.655 ;
        RECT 14.670 88.115 14.865 88.285 ;
        RECT 10.525 87.335 11.415 87.505 ;
        RECT 12.055 87.125 12.325 87.935 ;
        RECT 12.495 87.295 12.825 87.935 ;
        RECT 12.995 87.125 13.235 87.935 ;
        RECT 13.425 87.765 14.525 87.945 ;
        RECT 13.425 87.360 13.765 87.765 ;
        RECT 13.935 87.125 14.105 87.595 ;
        RECT 14.275 87.360 14.525 87.765 ;
        RECT 14.695 87.730 14.865 88.115 ;
        RECT 14.695 87.360 14.945 87.730 ;
        RECT 15.115 87.605 15.285 88.395 ;
        RECT 15.455 87.945 15.630 88.140 ;
        RECT 15.800 88.115 16.250 88.315 ;
        RECT 16.420 88.035 16.590 88.485 ;
        RECT 15.455 87.775 15.950 87.945 ;
        RECT 16.760 87.865 16.935 88.835 ;
        RECT 17.105 88.535 17.365 89.675 ;
        RECT 17.535 88.525 17.865 89.505 ;
        RECT 18.035 88.535 18.315 89.675 ;
        RECT 17.125 88.115 17.460 88.365 ;
        RECT 17.630 87.925 17.800 88.525 ;
        RECT 18.485 88.510 18.775 89.675 ;
        RECT 18.985 88.535 19.215 89.675 ;
        RECT 19.385 88.525 19.715 89.505 ;
        RECT 19.885 88.535 20.095 89.675 ;
        RECT 20.325 88.585 21.995 89.675 ;
        RECT 17.970 88.095 18.305 88.365 ;
        RECT 18.965 88.115 19.295 88.365 ;
        RECT 15.730 87.635 15.950 87.775 ;
        RECT 15.115 87.435 15.560 87.605 ;
        RECT 15.730 87.465 15.955 87.635 ;
        RECT 15.730 87.420 15.950 87.465 ;
        RECT 16.230 87.125 16.400 87.790 ;
        RECT 16.595 87.295 16.935 87.865 ;
        RECT 17.105 87.295 17.800 87.925 ;
        RECT 18.005 87.125 18.315 87.925 ;
        RECT 18.485 87.125 18.775 87.850 ;
        RECT 18.985 87.125 19.215 87.945 ;
        RECT 19.465 87.925 19.715 88.525 ;
        RECT 19.385 87.295 19.715 87.925 ;
        RECT 19.885 87.125 20.095 87.945 ;
        RECT 20.325 87.895 21.075 88.415 ;
        RECT 21.245 88.065 21.995 88.585 ;
        RECT 22.660 88.885 23.195 89.505 ;
        RECT 20.325 87.125 21.995 87.895 ;
        RECT 22.660 87.865 22.975 88.885 ;
        RECT 23.365 88.875 23.695 89.675 ;
        RECT 24.180 88.705 24.570 88.880 ;
        RECT 26.340 88.875 26.590 89.675 ;
        RECT 26.760 89.045 27.090 89.505 ;
        RECT 27.260 89.215 27.475 89.675 ;
        RECT 28.145 89.240 33.490 89.675 ;
        RECT 26.760 88.875 27.930 89.045 ;
        RECT 23.145 88.535 24.570 88.705 ;
        RECT 25.850 88.705 26.130 88.865 ;
        RECT 25.850 88.535 27.185 88.705 ;
        RECT 23.145 88.035 23.315 88.535 ;
        RECT 22.660 87.295 23.275 87.865 ;
        RECT 23.565 87.805 23.830 88.365 ;
        RECT 24.000 87.635 24.170 88.535 ;
        RECT 27.015 88.365 27.185 88.535 ;
        RECT 24.340 87.805 24.695 88.365 ;
        RECT 25.850 88.115 26.200 88.355 ;
        RECT 26.370 88.115 26.845 88.355 ;
        RECT 27.015 88.115 27.390 88.365 ;
        RECT 27.015 87.945 27.185 88.115 ;
        RECT 25.850 87.775 27.185 87.945 ;
        RECT 23.445 87.125 23.660 87.635 ;
        RECT 23.890 87.305 24.170 87.635 ;
        RECT 24.350 87.125 24.590 87.635 ;
        RECT 25.850 87.565 26.120 87.775 ;
        RECT 27.560 87.585 27.930 88.875 ;
        RECT 29.730 87.670 30.070 88.500 ;
        RECT 31.550 87.990 31.900 89.240 ;
        RECT 33.665 88.585 36.255 89.675 ;
        RECT 33.665 87.895 34.875 88.415 ;
        RECT 35.045 88.065 36.255 88.585 ;
        RECT 36.435 88.705 36.765 89.490 ;
        RECT 36.435 88.535 37.115 88.705 ;
        RECT 37.295 88.535 37.625 89.675 ;
        RECT 37.805 88.825 38.065 89.505 ;
        RECT 38.235 88.895 38.485 89.675 ;
        RECT 38.735 89.125 38.985 89.505 ;
        RECT 39.155 89.295 39.510 89.675 ;
        RECT 40.515 89.285 40.850 89.505 ;
        RECT 40.115 89.125 40.345 89.165 ;
        RECT 38.735 88.925 40.345 89.125 ;
        RECT 38.735 88.915 39.570 88.925 ;
        RECT 40.160 88.835 40.345 88.925 ;
        RECT 36.425 88.115 36.775 88.365 ;
        RECT 36.945 87.935 37.115 88.535 ;
        RECT 37.285 88.115 37.635 88.365 ;
        RECT 26.340 87.125 26.670 87.585 ;
        RECT 27.180 87.295 27.930 87.585 ;
        RECT 28.145 87.125 33.490 87.670 ;
        RECT 33.665 87.125 36.255 87.895 ;
        RECT 36.445 87.125 36.685 87.935 ;
        RECT 36.855 87.295 37.185 87.935 ;
        RECT 37.355 87.125 37.625 87.935 ;
        RECT 37.805 87.625 37.975 88.825 ;
        RECT 39.675 88.725 40.005 88.755 ;
        RECT 38.205 88.665 40.005 88.725 ;
        RECT 40.595 88.665 40.850 89.285 ;
        RECT 38.145 88.555 40.850 88.665 ;
        RECT 38.145 88.520 38.345 88.555 ;
        RECT 38.145 87.945 38.315 88.520 ;
        RECT 39.675 88.495 40.850 88.555 ;
        RECT 38.545 88.080 38.955 88.385 ;
        RECT 39.125 88.115 39.455 88.325 ;
        RECT 38.145 87.825 38.415 87.945 ;
        RECT 38.145 87.780 38.990 87.825 ;
        RECT 38.235 87.655 38.990 87.780 ;
        RECT 39.245 87.715 39.455 88.115 ;
        RECT 39.700 88.115 40.175 88.325 ;
        RECT 40.365 88.115 40.855 88.315 ;
        RECT 39.700 87.715 39.920 88.115 ;
        RECT 41.025 88.070 41.305 89.505 ;
        RECT 41.475 88.900 42.185 89.675 ;
        RECT 42.355 88.730 42.685 89.505 ;
        RECT 41.535 88.515 42.685 88.730 ;
        RECT 37.805 87.295 38.065 87.625 ;
        RECT 38.820 87.505 38.990 87.655 ;
        RECT 38.235 87.125 38.565 87.485 ;
        RECT 38.820 87.295 40.120 87.505 ;
        RECT 40.395 87.125 40.850 87.890 ;
        RECT 41.025 87.295 41.365 88.070 ;
        RECT 41.535 87.945 41.820 88.515 ;
        RECT 42.005 88.115 42.475 88.345 ;
        RECT 42.880 88.315 43.095 89.430 ;
        RECT 43.275 88.955 43.605 89.675 ;
        RECT 43.385 88.315 43.615 88.655 ;
        RECT 44.245 88.510 44.535 89.675 ;
        RECT 44.715 88.865 45.010 89.675 ;
        RECT 45.190 88.365 45.435 89.505 ;
        RECT 45.610 88.865 45.870 89.675 ;
        RECT 46.470 89.670 52.745 89.675 ;
        RECT 46.050 88.365 46.300 89.500 ;
        RECT 46.470 88.875 46.730 89.670 ;
        RECT 46.900 88.775 47.160 89.500 ;
        RECT 47.330 88.945 47.590 89.670 ;
        RECT 47.760 88.775 48.020 89.500 ;
        RECT 48.190 88.945 48.450 89.670 ;
        RECT 48.620 88.775 48.880 89.500 ;
        RECT 49.050 88.945 49.310 89.670 ;
        RECT 49.480 88.775 49.740 89.500 ;
        RECT 49.910 88.945 50.155 89.670 ;
        RECT 50.325 88.775 50.585 89.500 ;
        RECT 50.770 88.945 51.015 89.670 ;
        RECT 51.185 88.775 51.445 89.500 ;
        RECT 51.630 88.945 51.875 89.670 ;
        RECT 52.045 88.775 52.305 89.500 ;
        RECT 52.490 88.945 52.745 89.670 ;
        RECT 46.900 88.760 52.305 88.775 ;
        RECT 52.915 88.760 53.205 89.500 ;
        RECT 53.375 88.930 53.645 89.675 ;
        RECT 53.905 89.240 59.250 89.675 ;
        RECT 46.900 88.535 53.645 88.760 ;
        RECT 42.645 88.135 43.095 88.315 ;
        RECT 42.645 88.115 42.975 88.135 ;
        RECT 43.285 88.115 43.615 88.315 ;
        RECT 41.535 87.755 42.245 87.945 ;
        RECT 41.945 87.615 42.245 87.755 ;
        RECT 42.435 87.755 43.615 87.945 ;
        RECT 42.435 87.675 42.765 87.755 ;
        RECT 41.945 87.605 42.260 87.615 ;
        RECT 41.945 87.595 42.270 87.605 ;
        RECT 41.945 87.590 42.280 87.595 ;
        RECT 41.535 87.125 41.705 87.585 ;
        RECT 41.945 87.580 42.285 87.590 ;
        RECT 41.945 87.575 42.290 87.580 ;
        RECT 41.945 87.565 42.295 87.575 ;
        RECT 41.945 87.560 42.300 87.565 ;
        RECT 41.945 87.295 42.305 87.560 ;
        RECT 42.935 87.125 43.105 87.585 ;
        RECT 43.275 87.295 43.615 87.755 ;
        RECT 44.245 87.125 44.535 87.850 ;
        RECT 44.705 87.805 45.020 88.365 ;
        RECT 45.190 88.115 52.310 88.365 ;
        RECT 44.705 87.125 45.010 87.635 ;
        RECT 45.190 87.305 45.440 88.115 ;
        RECT 45.610 87.125 45.870 87.650 ;
        RECT 46.050 87.305 46.300 88.115 ;
        RECT 52.480 87.945 53.645 88.535 ;
        RECT 46.900 87.775 53.645 87.945 ;
        RECT 46.470 87.125 46.730 87.685 ;
        RECT 46.900 87.320 47.160 87.775 ;
        RECT 47.330 87.125 47.590 87.605 ;
        RECT 47.760 87.320 48.020 87.775 ;
        RECT 48.190 87.125 48.450 87.605 ;
        RECT 48.620 87.320 48.880 87.775 ;
        RECT 49.050 87.125 49.295 87.605 ;
        RECT 49.465 87.320 49.740 87.775 ;
        RECT 49.910 87.125 50.155 87.605 ;
        RECT 50.325 87.320 50.585 87.775 ;
        RECT 50.765 87.125 51.015 87.605 ;
        RECT 51.185 87.320 51.445 87.775 ;
        RECT 51.625 87.125 51.875 87.605 ;
        RECT 52.045 87.320 52.305 87.775 ;
        RECT 52.485 87.125 52.745 87.605 ;
        RECT 52.915 87.320 53.175 87.775 ;
        RECT 55.490 87.670 55.830 88.500 ;
        RECT 57.310 87.990 57.660 89.240 ;
        RECT 59.425 88.585 61.095 89.675 ;
        RECT 59.425 87.895 60.175 88.415 ;
        RECT 60.345 88.065 61.095 88.585 ;
        RECT 61.270 88.535 61.605 89.505 ;
        RECT 61.775 88.535 61.945 89.675 ;
        RECT 62.115 89.335 64.145 89.505 ;
        RECT 53.345 87.125 53.645 87.605 ;
        RECT 53.905 87.125 59.250 87.670 ;
        RECT 59.425 87.125 61.095 87.895 ;
        RECT 61.270 87.865 61.440 88.535 ;
        RECT 62.115 88.365 62.285 89.335 ;
        RECT 61.610 88.035 61.865 88.365 ;
        RECT 62.090 88.035 62.285 88.365 ;
        RECT 62.455 88.995 63.580 89.165 ;
        RECT 61.695 87.865 61.865 88.035 ;
        RECT 62.455 87.865 62.625 88.995 ;
        RECT 61.270 87.295 61.525 87.865 ;
        RECT 61.695 87.695 62.625 87.865 ;
        RECT 62.795 88.655 63.805 88.825 ;
        RECT 62.795 87.855 62.965 88.655 ;
        RECT 63.170 88.315 63.445 88.455 ;
        RECT 63.165 88.145 63.445 88.315 ;
        RECT 62.450 87.660 62.625 87.695 ;
        RECT 61.695 87.125 62.025 87.525 ;
        RECT 62.450 87.295 62.980 87.660 ;
        RECT 63.170 87.295 63.445 88.145 ;
        RECT 63.615 87.295 63.805 88.655 ;
        RECT 63.975 88.670 64.145 89.335 ;
        RECT 64.315 88.915 64.485 89.675 ;
        RECT 64.720 88.915 65.235 89.325 ;
        RECT 63.975 88.480 64.725 88.670 ;
        RECT 64.895 88.105 65.235 88.915 ;
        RECT 65.405 88.585 66.615 89.675 ;
        RECT 64.005 87.935 65.235 88.105 ;
        RECT 63.985 87.125 64.495 87.660 ;
        RECT 64.715 87.330 64.960 87.935 ;
        RECT 65.405 87.875 65.925 88.415 ;
        RECT 66.095 88.045 66.615 88.585 ;
        RECT 66.785 88.825 67.045 89.505 ;
        RECT 67.215 88.895 67.465 89.675 ;
        RECT 67.715 89.125 67.965 89.505 ;
        RECT 68.135 89.295 68.490 89.675 ;
        RECT 69.495 89.285 69.830 89.505 ;
        RECT 69.095 89.125 69.325 89.165 ;
        RECT 67.715 88.925 69.325 89.125 ;
        RECT 67.715 88.915 68.550 88.925 ;
        RECT 69.140 88.835 69.325 88.925 ;
        RECT 65.405 87.125 66.615 87.875 ;
        RECT 66.785 87.635 66.955 88.825 ;
        RECT 68.655 88.725 68.985 88.755 ;
        RECT 67.185 88.665 68.985 88.725 ;
        RECT 69.575 88.665 69.830 89.285 ;
        RECT 67.125 88.555 69.830 88.665 ;
        RECT 67.125 88.520 67.325 88.555 ;
        RECT 67.125 87.945 67.295 88.520 ;
        RECT 68.655 88.495 69.830 88.555 ;
        RECT 70.005 88.510 70.295 89.675 ;
        RECT 70.555 88.745 70.725 89.505 ;
        RECT 70.905 88.915 71.235 89.675 ;
        RECT 70.555 88.575 71.220 88.745 ;
        RECT 71.405 88.600 71.675 89.505 ;
        RECT 71.050 88.430 71.220 88.575 ;
        RECT 67.525 88.080 67.935 88.385 ;
        RECT 68.105 88.115 68.435 88.325 ;
        RECT 67.125 87.825 67.395 87.945 ;
        RECT 67.125 87.780 67.970 87.825 ;
        RECT 67.215 87.655 67.970 87.780 ;
        RECT 68.225 87.715 68.435 88.115 ;
        RECT 68.680 88.115 69.155 88.325 ;
        RECT 69.345 88.115 69.835 88.315 ;
        RECT 68.680 87.715 68.900 88.115 ;
        RECT 70.485 88.025 70.815 88.395 ;
        RECT 71.050 88.100 71.335 88.430 ;
        RECT 66.785 87.625 67.015 87.635 ;
        RECT 66.785 87.295 67.045 87.625 ;
        RECT 67.800 87.505 67.970 87.655 ;
        RECT 67.215 87.125 67.545 87.485 ;
        RECT 67.800 87.295 69.100 87.505 ;
        RECT 69.375 87.125 69.830 87.890 ;
        RECT 70.005 87.125 70.295 87.850 ;
        RECT 71.050 87.845 71.220 88.100 ;
        RECT 70.555 87.675 71.220 87.845 ;
        RECT 71.505 87.800 71.675 88.600 ;
        RECT 70.555 87.295 70.725 87.675 ;
        RECT 70.905 87.125 71.235 87.505 ;
        RECT 71.415 87.295 71.675 87.800 ;
        RECT 71.845 88.535 72.185 89.505 ;
        RECT 72.355 88.535 72.525 89.675 ;
        RECT 72.795 88.875 73.045 89.675 ;
        RECT 73.690 88.705 74.020 89.505 ;
        RECT 74.320 88.875 74.650 89.675 ;
        RECT 74.820 88.705 75.150 89.505 ;
        RECT 72.715 88.535 75.150 88.705 ;
        RECT 75.560 88.885 76.095 89.505 ;
        RECT 71.845 87.925 72.020 88.535 ;
        RECT 72.715 88.285 72.885 88.535 ;
        RECT 72.190 88.115 72.885 88.285 ;
        RECT 73.060 88.115 73.480 88.315 ;
        RECT 73.650 88.115 73.980 88.315 ;
        RECT 74.150 88.115 74.480 88.315 ;
        RECT 71.845 87.295 72.185 87.925 ;
        RECT 72.355 87.125 72.605 87.925 ;
        RECT 72.795 87.775 74.020 87.945 ;
        RECT 72.795 87.295 73.125 87.775 ;
        RECT 73.295 87.125 73.520 87.585 ;
        RECT 73.690 87.295 74.020 87.775 ;
        RECT 74.650 87.905 74.820 88.535 ;
        RECT 75.005 88.115 75.355 88.365 ;
        RECT 74.650 87.295 75.150 87.905 ;
        RECT 75.560 87.865 75.875 88.885 ;
        RECT 76.265 88.875 76.595 89.675 ;
        RECT 77.080 88.705 77.470 88.880 ;
        RECT 76.045 88.535 77.470 88.705 ;
        RECT 78.010 88.705 78.400 88.880 ;
        RECT 78.885 88.875 79.215 89.675 ;
        RECT 79.385 88.885 79.920 89.505 ;
        RECT 78.010 88.535 79.435 88.705 ;
        RECT 76.045 88.035 76.215 88.535 ;
        RECT 75.560 87.295 76.175 87.865 ;
        RECT 76.465 87.805 76.730 88.365 ;
        RECT 76.900 87.635 77.070 88.535 ;
        RECT 77.240 87.805 77.595 88.365 ;
        RECT 77.885 87.805 78.240 88.365 ;
        RECT 78.410 87.635 78.580 88.535 ;
        RECT 78.750 87.805 79.015 88.365 ;
        RECT 79.265 88.035 79.435 88.535 ;
        RECT 79.605 87.865 79.920 88.885 ;
        RECT 80.130 88.525 80.390 89.675 ;
        RECT 80.565 88.600 80.820 89.505 ;
        RECT 80.990 88.915 81.320 89.675 ;
        RECT 81.535 88.745 81.705 89.505 ;
        RECT 76.345 87.125 76.560 87.635 ;
        RECT 76.790 87.305 77.070 87.635 ;
        RECT 77.250 87.125 77.490 87.635 ;
        RECT 77.990 87.125 78.230 87.635 ;
        RECT 78.410 87.305 78.690 87.635 ;
        RECT 78.920 87.125 79.135 87.635 ;
        RECT 79.305 87.295 79.920 87.865 ;
        RECT 80.130 87.125 80.390 87.965 ;
        RECT 80.565 87.870 80.735 88.600 ;
        RECT 80.990 88.575 81.705 88.745 ;
        RECT 81.965 88.585 83.175 89.675 ;
        RECT 80.990 88.365 81.160 88.575 ;
        RECT 80.905 88.035 81.160 88.365 ;
        RECT 80.565 87.295 80.820 87.870 ;
        RECT 80.990 87.845 81.160 88.035 ;
        RECT 81.440 88.025 81.795 88.395 ;
        RECT 81.965 88.045 82.485 88.585 ;
        RECT 82.655 87.875 83.175 88.415 ;
        RECT 80.990 87.675 81.705 87.845 ;
        RECT 80.990 87.125 81.320 87.505 ;
        RECT 81.535 87.295 81.705 87.675 ;
        RECT 81.965 87.125 83.175 87.875 ;
        RECT 5.520 86.955 83.260 87.125 ;
        RECT 5.605 86.205 6.815 86.955 ;
        RECT 7.995 86.405 8.165 86.695 ;
        RECT 8.335 86.575 8.665 86.955 ;
        RECT 7.995 86.235 8.660 86.405 ;
        RECT 5.605 85.665 6.125 86.205 ;
        RECT 6.295 85.495 6.815 86.035 ;
        RECT 5.605 84.405 6.815 85.495 ;
        RECT 7.910 85.415 8.260 86.065 ;
        RECT 8.430 85.245 8.660 86.235 ;
        RECT 7.995 85.075 8.660 85.245 ;
        RECT 7.995 84.575 8.165 85.075 ;
        RECT 8.335 84.405 8.665 84.905 ;
        RECT 8.835 84.575 9.020 86.695 ;
        RECT 9.275 86.495 9.525 86.955 ;
        RECT 9.695 86.505 10.030 86.675 ;
        RECT 10.225 86.505 10.900 86.675 ;
        RECT 9.695 86.365 9.865 86.505 ;
        RECT 9.190 85.375 9.470 86.325 ;
        RECT 9.640 86.235 9.865 86.365 ;
        RECT 9.640 85.130 9.810 86.235 ;
        RECT 10.035 86.085 10.560 86.305 ;
        RECT 9.980 85.320 10.220 85.915 ;
        RECT 10.390 85.385 10.560 86.085 ;
        RECT 10.730 85.725 10.900 86.505 ;
        RECT 11.220 86.455 11.590 86.955 ;
        RECT 11.770 86.505 12.175 86.675 ;
        RECT 12.345 86.505 13.130 86.675 ;
        RECT 11.770 86.275 11.940 86.505 ;
        RECT 11.110 85.975 11.940 86.275 ;
        RECT 12.325 86.005 12.790 86.335 ;
        RECT 11.110 85.945 11.310 85.975 ;
        RECT 11.430 85.725 11.600 85.795 ;
        RECT 10.730 85.555 11.600 85.725 ;
        RECT 11.090 85.465 11.600 85.555 ;
        RECT 9.640 85.000 9.945 85.130 ;
        RECT 10.390 85.020 10.920 85.385 ;
        RECT 9.260 84.405 9.525 84.865 ;
        RECT 9.695 84.575 9.945 85.000 ;
        RECT 11.090 84.850 11.260 85.465 ;
        RECT 10.155 84.680 11.260 84.850 ;
        RECT 11.430 84.405 11.600 85.205 ;
        RECT 11.770 84.905 11.940 85.975 ;
        RECT 12.110 85.075 12.300 85.795 ;
        RECT 12.470 85.045 12.790 86.005 ;
        RECT 12.960 86.045 13.130 86.505 ;
        RECT 13.405 86.425 13.615 86.955 ;
        RECT 13.875 86.215 14.205 86.740 ;
        RECT 14.375 86.345 14.545 86.955 ;
        RECT 14.715 86.300 15.045 86.735 ;
        RECT 14.715 86.215 15.095 86.300 ;
        RECT 14.005 86.045 14.205 86.215 ;
        RECT 14.870 86.175 15.095 86.215 ;
        RECT 12.960 85.715 13.835 86.045 ;
        RECT 14.005 85.715 14.755 86.045 ;
        RECT 11.770 84.575 12.020 84.905 ;
        RECT 12.960 84.875 13.130 85.715 ;
        RECT 14.005 85.510 14.195 85.715 ;
        RECT 14.925 85.595 15.095 86.175 ;
        RECT 15.735 86.145 16.005 86.955 ;
        RECT 16.175 86.145 16.505 86.785 ;
        RECT 16.675 86.145 16.915 86.955 ;
        RECT 17.195 86.405 17.365 86.695 ;
        RECT 17.535 86.575 17.865 86.955 ;
        RECT 17.195 86.235 17.860 86.405 ;
        RECT 15.725 85.715 16.075 85.965 ;
        RECT 14.880 85.545 15.095 85.595 ;
        RECT 16.245 85.545 16.415 86.145 ;
        RECT 16.585 85.715 16.935 85.965 ;
        RECT 13.300 85.135 14.195 85.510 ;
        RECT 14.705 85.465 15.095 85.545 ;
        RECT 12.245 84.705 13.130 84.875 ;
        RECT 13.310 84.405 13.625 84.905 ;
        RECT 13.855 84.575 14.195 85.135 ;
        RECT 14.365 84.405 14.535 85.415 ;
        RECT 14.705 84.620 15.035 85.465 ;
        RECT 15.735 84.405 16.065 85.545 ;
        RECT 16.245 85.375 16.925 85.545 ;
        RECT 17.110 85.415 17.460 86.065 ;
        RECT 16.595 84.590 16.925 85.375 ;
        RECT 17.630 85.245 17.860 86.235 ;
        RECT 17.195 85.075 17.860 85.245 ;
        RECT 17.195 84.575 17.365 85.075 ;
        RECT 17.535 84.405 17.865 84.905 ;
        RECT 18.035 84.575 18.220 86.695 ;
        RECT 18.475 86.495 18.725 86.955 ;
        RECT 18.895 86.505 19.230 86.675 ;
        RECT 19.425 86.505 20.100 86.675 ;
        RECT 18.895 86.365 19.065 86.505 ;
        RECT 18.390 85.375 18.670 86.325 ;
        RECT 18.840 86.235 19.065 86.365 ;
        RECT 18.840 85.130 19.010 86.235 ;
        RECT 19.235 86.085 19.760 86.305 ;
        RECT 19.180 85.320 19.420 85.915 ;
        RECT 19.590 85.385 19.760 86.085 ;
        RECT 19.930 85.725 20.100 86.505 ;
        RECT 20.420 86.455 20.790 86.955 ;
        RECT 20.970 86.505 21.375 86.675 ;
        RECT 21.545 86.505 22.330 86.675 ;
        RECT 20.970 86.275 21.140 86.505 ;
        RECT 20.310 85.975 21.140 86.275 ;
        RECT 21.525 86.005 21.990 86.335 ;
        RECT 20.310 85.945 20.510 85.975 ;
        RECT 20.630 85.725 20.800 85.795 ;
        RECT 19.930 85.555 20.800 85.725 ;
        RECT 20.290 85.465 20.800 85.555 ;
        RECT 18.840 85.000 19.145 85.130 ;
        RECT 19.590 85.020 20.120 85.385 ;
        RECT 18.460 84.405 18.725 84.865 ;
        RECT 18.895 84.575 19.145 85.000 ;
        RECT 20.290 84.850 20.460 85.465 ;
        RECT 19.355 84.680 20.460 84.850 ;
        RECT 20.630 84.405 20.800 85.205 ;
        RECT 20.970 84.905 21.140 85.975 ;
        RECT 21.310 85.075 21.500 85.795 ;
        RECT 21.670 85.045 21.990 86.005 ;
        RECT 22.160 86.045 22.330 86.505 ;
        RECT 22.605 86.425 22.815 86.955 ;
        RECT 23.075 86.215 23.405 86.740 ;
        RECT 23.575 86.345 23.745 86.955 ;
        RECT 23.915 86.300 24.245 86.735 ;
        RECT 23.915 86.215 24.295 86.300 ;
        RECT 23.205 86.045 23.405 86.215 ;
        RECT 24.070 86.175 24.295 86.215 ;
        RECT 22.160 85.715 23.035 86.045 ;
        RECT 23.205 85.715 23.955 86.045 ;
        RECT 20.970 84.575 21.220 84.905 ;
        RECT 22.160 84.875 22.330 85.715 ;
        RECT 23.205 85.510 23.395 85.715 ;
        RECT 24.125 85.595 24.295 86.175 ;
        RECT 24.465 86.205 25.675 86.955 ;
        RECT 25.845 86.575 26.735 86.745 ;
        RECT 24.465 85.665 24.985 86.205 ;
        RECT 24.080 85.545 24.295 85.595 ;
        RECT 22.500 85.135 23.395 85.510 ;
        RECT 23.905 85.465 24.295 85.545 ;
        RECT 25.155 85.495 25.675 86.035 ;
        RECT 25.845 86.020 26.395 86.405 ;
        RECT 26.565 85.850 26.735 86.575 ;
        RECT 21.445 84.705 22.330 84.875 ;
        RECT 22.510 84.405 22.825 84.905 ;
        RECT 23.055 84.575 23.395 85.135 ;
        RECT 23.565 84.405 23.735 85.415 ;
        RECT 23.905 84.620 24.235 85.465 ;
        RECT 24.465 84.405 25.675 85.495 ;
        RECT 25.845 85.780 26.735 85.850 ;
        RECT 26.905 86.250 27.125 86.735 ;
        RECT 27.295 86.415 27.545 86.955 ;
        RECT 27.715 86.305 27.975 86.785 ;
        RECT 26.905 85.825 27.235 86.250 ;
        RECT 25.845 85.755 26.740 85.780 ;
        RECT 25.845 85.740 26.750 85.755 ;
        RECT 25.845 85.725 26.755 85.740 ;
        RECT 25.845 85.720 26.765 85.725 ;
        RECT 25.845 85.710 26.770 85.720 ;
        RECT 25.845 85.700 26.775 85.710 ;
        RECT 25.845 85.695 26.785 85.700 ;
        RECT 25.845 85.685 26.795 85.695 ;
        RECT 25.845 85.680 26.805 85.685 ;
        RECT 25.845 85.230 26.105 85.680 ;
        RECT 26.470 85.675 26.805 85.680 ;
        RECT 26.470 85.670 26.820 85.675 ;
        RECT 26.470 85.660 26.835 85.670 ;
        RECT 26.470 85.655 26.860 85.660 ;
        RECT 27.405 85.655 27.635 86.050 ;
        RECT 26.470 85.650 27.635 85.655 ;
        RECT 26.500 85.615 27.635 85.650 ;
        RECT 26.535 85.590 27.635 85.615 ;
        RECT 26.565 85.560 27.635 85.590 ;
        RECT 26.585 85.530 27.635 85.560 ;
        RECT 26.605 85.500 27.635 85.530 ;
        RECT 26.675 85.490 27.635 85.500 ;
        RECT 26.700 85.480 27.635 85.490 ;
        RECT 26.720 85.465 27.635 85.480 ;
        RECT 26.740 85.450 27.635 85.465 ;
        RECT 26.745 85.440 27.530 85.450 ;
        RECT 26.760 85.405 27.530 85.440 ;
        RECT 26.275 85.085 26.605 85.330 ;
        RECT 26.775 85.155 27.530 85.405 ;
        RECT 27.805 85.275 27.975 86.305 ;
        RECT 28.165 86.225 28.455 86.955 ;
        RECT 28.155 85.715 28.455 86.045 ;
        RECT 28.635 86.025 28.865 86.665 ;
        RECT 29.045 86.405 29.355 86.775 ;
        RECT 29.535 86.585 30.205 86.955 ;
        RECT 29.045 86.205 30.275 86.405 ;
        RECT 28.635 85.715 29.160 86.025 ;
        RECT 29.340 85.715 29.805 86.025 ;
        RECT 29.985 85.535 30.275 86.205 ;
        RECT 26.275 85.060 26.460 85.085 ;
        RECT 25.845 84.960 26.460 85.060 ;
        RECT 25.845 84.405 26.450 84.960 ;
        RECT 26.625 84.575 27.105 84.915 ;
        RECT 27.275 84.405 27.530 84.950 ;
        RECT 27.700 84.575 27.975 85.275 ;
        RECT 28.165 85.295 29.325 85.535 ;
        RECT 28.165 84.585 28.425 85.295 ;
        RECT 28.595 84.405 28.925 85.115 ;
        RECT 29.095 84.585 29.325 85.295 ;
        RECT 29.505 85.315 30.275 85.535 ;
        RECT 29.505 84.585 29.775 85.315 ;
        RECT 29.955 84.405 30.295 85.135 ;
        RECT 30.465 84.585 30.725 86.775 ;
        RECT 31.365 86.230 31.655 86.955 ;
        RECT 31.825 86.410 37.170 86.955 ;
        RECT 33.410 85.580 33.750 86.410 ;
        RECT 37.345 86.185 40.855 86.955 ;
        RECT 41.025 86.205 42.235 86.955 ;
        RECT 42.420 86.385 42.675 86.735 ;
        RECT 42.845 86.555 43.175 86.955 ;
        RECT 43.345 86.385 43.515 86.735 ;
        RECT 43.685 86.555 44.065 86.955 ;
        RECT 42.420 86.215 44.085 86.385 ;
        RECT 44.255 86.280 44.530 86.625 ;
        RECT 31.365 84.405 31.655 85.570 ;
        RECT 35.230 84.840 35.580 86.090 ;
        RECT 37.345 85.665 38.995 86.185 ;
        RECT 39.165 85.495 40.855 86.015 ;
        RECT 41.025 85.665 41.545 86.205 ;
        RECT 43.915 86.045 44.085 86.215 ;
        RECT 41.715 85.495 42.235 86.035 ;
        RECT 42.405 85.715 42.750 86.045 ;
        RECT 42.920 85.715 43.745 86.045 ;
        RECT 43.915 85.715 44.190 86.045 ;
        RECT 31.825 84.405 37.170 84.840 ;
        RECT 37.345 84.405 40.855 85.495 ;
        RECT 41.025 84.405 42.235 85.495 ;
        RECT 42.425 85.255 42.750 85.545 ;
        RECT 42.920 85.425 43.115 85.715 ;
        RECT 43.915 85.545 44.085 85.715 ;
        RECT 44.360 85.545 44.530 86.280 ;
        RECT 44.765 86.135 44.975 86.955 ;
        RECT 45.145 86.155 45.475 86.785 ;
        RECT 45.145 85.555 45.395 86.155 ;
        RECT 45.645 86.135 45.875 86.955 ;
        RECT 46.130 86.495 46.880 86.785 ;
        RECT 47.390 86.495 47.720 86.955 ;
        RECT 45.565 85.715 45.895 85.965 ;
        RECT 43.425 85.375 44.085 85.545 ;
        RECT 43.425 85.255 43.595 85.375 ;
        RECT 42.425 85.085 43.595 85.255 ;
        RECT 42.405 84.625 43.595 84.915 ;
        RECT 43.765 84.405 44.045 85.205 ;
        RECT 44.255 84.575 44.530 85.545 ;
        RECT 44.765 84.405 44.975 85.545 ;
        RECT 45.145 84.575 45.475 85.555 ;
        RECT 45.645 84.405 45.875 85.545 ;
        RECT 46.130 85.205 46.500 86.495 ;
        RECT 47.940 86.305 48.210 86.515 ;
        RECT 46.875 86.135 48.210 86.305 ;
        RECT 48.385 86.205 49.595 86.955 ;
        RECT 49.785 86.445 50.025 86.955 ;
        RECT 50.195 86.445 50.485 86.785 ;
        RECT 50.715 86.445 51.030 86.955 ;
        RECT 46.875 85.965 47.045 86.135 ;
        RECT 46.670 85.715 47.045 85.965 ;
        RECT 47.215 85.725 47.690 85.965 ;
        RECT 47.860 85.725 48.210 85.965 ;
        RECT 46.875 85.545 47.045 85.715 ;
        RECT 48.385 85.665 48.905 86.205 ;
        RECT 49.825 86.105 50.025 86.275 ;
        RECT 46.875 85.375 48.210 85.545 ;
        RECT 49.075 85.495 49.595 86.035 ;
        RECT 49.830 85.715 50.025 86.105 ;
        RECT 50.195 85.545 50.375 86.445 ;
        RECT 51.200 86.385 51.370 86.655 ;
        RECT 51.540 86.555 51.870 86.955 ;
        RECT 50.545 85.715 50.955 86.275 ;
        RECT 51.200 86.215 51.895 86.385 ;
        RECT 51.125 85.545 51.295 86.045 ;
        RECT 47.930 85.215 48.210 85.375 ;
        RECT 46.130 85.035 47.300 85.205 ;
        RECT 46.585 84.405 46.800 84.865 ;
        RECT 46.970 84.575 47.300 85.035 ;
        RECT 47.470 84.405 47.720 85.205 ;
        RECT 48.385 84.405 49.595 85.495 ;
        RECT 49.835 85.375 51.295 85.545 ;
        RECT 49.835 85.200 50.195 85.375 ;
        RECT 51.465 85.205 51.895 86.215 ;
        RECT 52.070 86.135 52.345 86.955 ;
        RECT 52.515 86.315 52.845 86.785 ;
        RECT 53.015 86.485 53.185 86.955 ;
        RECT 53.355 86.315 53.685 86.785 ;
        RECT 53.855 86.485 54.145 86.955 ;
        RECT 52.515 86.305 53.685 86.315 ;
        RECT 52.515 86.135 54.115 86.305 ;
        RECT 54.370 86.135 54.645 86.955 ;
        RECT 54.815 86.315 55.145 86.785 ;
        RECT 55.315 86.485 55.485 86.955 ;
        RECT 55.655 86.315 55.985 86.785 ;
        RECT 56.155 86.485 56.445 86.955 ;
        RECT 54.815 86.305 55.985 86.315 ;
        RECT 54.815 86.135 56.415 86.305 ;
        RECT 57.125 86.230 57.415 86.955 ;
        RECT 57.585 86.410 62.930 86.955 ;
        RECT 52.070 85.765 52.790 85.965 ;
        RECT 52.960 85.765 53.730 85.965 ;
        RECT 53.900 85.595 54.115 86.135 ;
        RECT 54.370 85.765 55.090 85.965 ;
        RECT 55.260 85.765 56.030 85.965 ;
        RECT 56.200 85.595 56.415 86.135 ;
        RECT 50.780 84.405 50.950 85.205 ;
        RECT 51.120 85.035 51.895 85.205 ;
        RECT 52.070 85.375 53.185 85.585 ;
        RECT 51.120 84.575 51.450 85.035 ;
        RECT 51.620 84.405 51.790 84.865 ;
        RECT 52.070 84.575 52.345 85.375 ;
        RECT 52.515 84.405 52.845 85.205 ;
        RECT 53.015 84.745 53.185 85.375 ;
        RECT 53.355 85.375 54.115 85.595 ;
        RECT 54.370 85.375 55.485 85.585 ;
        RECT 53.355 84.915 53.685 85.375 ;
        RECT 53.855 84.745 54.155 85.205 ;
        RECT 53.015 84.575 54.155 84.745 ;
        RECT 54.370 84.575 54.645 85.375 ;
        RECT 54.815 84.405 55.145 85.205 ;
        RECT 55.315 84.745 55.485 85.375 ;
        RECT 55.655 85.425 56.435 85.595 ;
        RECT 59.170 85.580 59.510 86.410 ;
        RECT 63.105 86.185 64.775 86.955 ;
        RECT 55.655 85.375 56.415 85.425 ;
        RECT 55.655 84.915 55.985 85.375 ;
        RECT 56.155 84.745 56.455 85.205 ;
        RECT 55.315 84.575 56.455 84.745 ;
        RECT 57.125 84.405 57.415 85.570 ;
        RECT 60.990 84.840 61.340 86.090 ;
        RECT 63.105 85.665 63.855 86.185 ;
        RECT 64.950 86.115 65.210 86.955 ;
        RECT 65.385 86.210 65.640 86.785 ;
        RECT 65.810 86.575 66.140 86.955 ;
        RECT 66.355 86.405 66.525 86.785 ;
        RECT 65.810 86.235 66.525 86.405 ;
        RECT 64.025 85.495 64.775 86.015 ;
        RECT 57.585 84.405 62.930 84.840 ;
        RECT 63.105 84.405 64.775 85.495 ;
        RECT 64.950 84.405 65.210 85.555 ;
        RECT 65.385 85.480 65.555 86.210 ;
        RECT 65.810 86.045 65.980 86.235 ;
        RECT 66.790 86.115 67.050 86.955 ;
        RECT 67.225 86.210 67.480 86.785 ;
        RECT 67.650 86.575 67.980 86.955 ;
        RECT 68.195 86.405 68.365 86.785 ;
        RECT 67.650 86.235 68.365 86.405 ;
        RECT 65.725 85.715 65.980 86.045 ;
        RECT 65.810 85.505 65.980 85.715 ;
        RECT 66.260 85.685 66.615 86.055 ;
        RECT 65.385 84.575 65.640 85.480 ;
        RECT 65.810 85.335 66.525 85.505 ;
        RECT 65.810 84.405 66.140 85.165 ;
        RECT 66.355 84.575 66.525 85.335 ;
        RECT 66.790 84.405 67.050 85.555 ;
        RECT 67.225 85.480 67.395 86.210 ;
        RECT 67.650 86.045 67.820 86.235 ;
        RECT 68.630 86.115 68.890 86.955 ;
        RECT 69.065 86.210 69.320 86.785 ;
        RECT 69.490 86.575 69.820 86.955 ;
        RECT 70.035 86.405 70.205 86.785 ;
        RECT 70.630 86.445 70.870 86.955 ;
        RECT 71.050 86.445 71.330 86.775 ;
        RECT 71.560 86.445 71.775 86.955 ;
        RECT 69.490 86.235 70.205 86.405 ;
        RECT 67.565 85.715 67.820 86.045 ;
        RECT 67.650 85.505 67.820 85.715 ;
        RECT 68.100 85.685 68.455 86.055 ;
        RECT 67.225 84.575 67.480 85.480 ;
        RECT 67.650 85.335 68.365 85.505 ;
        RECT 67.650 84.405 67.980 85.165 ;
        RECT 68.195 84.575 68.365 85.335 ;
        RECT 68.630 84.405 68.890 85.555 ;
        RECT 69.065 85.480 69.235 86.210 ;
        RECT 69.490 86.045 69.660 86.235 ;
        RECT 69.405 85.715 69.660 86.045 ;
        RECT 69.490 85.505 69.660 85.715 ;
        RECT 69.940 85.685 70.295 86.055 ;
        RECT 70.525 85.715 70.880 86.275 ;
        RECT 71.050 85.545 71.220 86.445 ;
        RECT 71.390 85.715 71.655 86.275 ;
        RECT 71.945 86.215 72.560 86.785 ;
        RECT 72.875 86.575 74.045 86.785 ;
        RECT 72.875 86.555 73.205 86.575 ;
        RECT 71.905 85.545 72.075 86.045 ;
        RECT 69.065 84.575 69.320 85.480 ;
        RECT 69.490 85.335 70.205 85.505 ;
        RECT 69.490 84.405 69.820 85.165 ;
        RECT 70.035 84.575 70.205 85.335 ;
        RECT 70.650 85.375 72.075 85.545 ;
        RECT 70.650 85.200 71.040 85.375 ;
        RECT 71.525 84.405 71.855 85.205 ;
        RECT 72.245 85.195 72.560 86.215 ;
        RECT 72.765 86.135 73.625 86.385 ;
        RECT 73.795 86.325 74.045 86.575 ;
        RECT 74.215 86.495 74.385 86.955 ;
        RECT 74.555 86.325 74.895 86.785 ;
        RECT 73.795 86.155 74.895 86.325 ;
        RECT 75.155 86.405 75.325 86.785 ;
        RECT 75.540 86.575 75.870 86.955 ;
        RECT 75.155 86.235 75.870 86.405 ;
        RECT 72.765 85.545 73.045 86.135 ;
        RECT 73.215 85.715 73.965 85.965 ;
        RECT 74.135 85.715 74.895 85.965 ;
        RECT 75.065 85.685 75.420 86.055 ;
        RECT 75.700 86.045 75.870 86.235 ;
        RECT 76.040 86.210 76.295 86.785 ;
        RECT 75.700 85.715 75.955 86.045 ;
        RECT 72.765 85.375 74.465 85.545 ;
        RECT 72.025 84.575 72.560 85.195 ;
        RECT 72.870 84.405 73.125 85.205 ;
        RECT 73.295 84.575 73.625 85.375 ;
        RECT 73.795 84.405 73.965 85.205 ;
        RECT 74.135 84.575 74.465 85.375 ;
        RECT 74.635 84.405 74.895 85.545 ;
        RECT 75.700 85.505 75.870 85.715 ;
        RECT 75.155 85.335 75.870 85.505 ;
        RECT 76.125 85.480 76.295 86.210 ;
        RECT 76.470 86.115 76.730 86.955 ;
        RECT 77.365 86.455 77.625 86.785 ;
        RECT 77.795 86.595 78.125 86.955 ;
        RECT 78.380 86.575 79.680 86.785 ;
        RECT 77.365 86.445 77.595 86.455 ;
        RECT 75.155 84.575 75.325 85.335 ;
        RECT 75.540 84.405 75.870 85.165 ;
        RECT 76.040 84.575 76.295 85.480 ;
        RECT 76.470 84.405 76.730 85.555 ;
        RECT 77.365 85.255 77.535 86.445 ;
        RECT 78.380 86.425 78.550 86.575 ;
        RECT 77.795 86.300 78.550 86.425 ;
        RECT 77.705 86.255 78.550 86.300 ;
        RECT 77.705 86.135 77.975 86.255 ;
        RECT 77.705 85.560 77.875 86.135 ;
        RECT 78.105 85.695 78.515 86.000 ;
        RECT 78.805 85.965 79.015 86.365 ;
        RECT 78.685 85.755 79.015 85.965 ;
        RECT 79.260 85.965 79.480 86.365 ;
        RECT 79.955 86.190 80.410 86.955 ;
        RECT 80.585 86.205 81.795 86.955 ;
        RECT 81.965 86.205 83.175 86.955 ;
        RECT 79.260 85.755 79.735 85.965 ;
        RECT 79.925 85.765 80.415 85.965 ;
        RECT 80.585 85.665 81.105 86.205 ;
        RECT 77.705 85.525 77.905 85.560 ;
        RECT 79.235 85.525 80.410 85.585 ;
        RECT 77.705 85.415 80.410 85.525 ;
        RECT 81.275 85.495 81.795 86.035 ;
        RECT 77.765 85.355 79.565 85.415 ;
        RECT 79.235 85.325 79.565 85.355 ;
        RECT 77.365 84.575 77.625 85.255 ;
        RECT 77.795 84.405 78.045 85.185 ;
        RECT 78.295 85.155 79.130 85.165 ;
        RECT 79.720 85.155 79.905 85.245 ;
        RECT 78.295 84.955 79.905 85.155 ;
        RECT 78.295 84.575 78.545 84.955 ;
        RECT 79.675 84.915 79.905 84.955 ;
        RECT 80.155 84.795 80.410 85.415 ;
        RECT 78.715 84.405 79.070 84.785 ;
        RECT 80.075 84.575 80.410 84.795 ;
        RECT 80.585 84.405 81.795 85.495 ;
        RECT 81.965 85.495 82.485 86.035 ;
        RECT 82.655 85.665 83.175 86.205 ;
        RECT 81.965 84.405 83.175 85.495 ;
        RECT 5.520 84.235 83.260 84.405 ;
        RECT 5.605 83.145 6.815 84.235 ;
        RECT 7.075 83.565 7.245 84.065 ;
        RECT 7.415 83.735 7.745 84.235 ;
        RECT 7.075 83.395 7.740 83.565 ;
        RECT 5.605 82.435 6.125 82.975 ;
        RECT 6.295 82.605 6.815 83.145 ;
        RECT 6.990 82.575 7.340 83.225 ;
        RECT 5.605 81.685 6.815 82.435 ;
        RECT 7.510 82.405 7.740 83.395 ;
        RECT 7.075 82.235 7.740 82.405 ;
        RECT 7.075 81.945 7.245 82.235 ;
        RECT 7.415 81.685 7.745 82.065 ;
        RECT 7.915 81.945 8.100 84.065 ;
        RECT 8.340 83.775 8.605 84.235 ;
        RECT 8.775 83.640 9.025 84.065 ;
        RECT 9.235 83.790 10.340 83.960 ;
        RECT 8.720 83.510 9.025 83.640 ;
        RECT 8.270 82.315 8.550 83.265 ;
        RECT 8.720 82.405 8.890 83.510 ;
        RECT 9.060 82.725 9.300 83.320 ;
        RECT 9.470 83.255 10.000 83.620 ;
        RECT 9.470 82.555 9.640 83.255 ;
        RECT 10.170 83.175 10.340 83.790 ;
        RECT 10.510 83.435 10.680 84.235 ;
        RECT 10.850 83.735 11.100 84.065 ;
        RECT 11.325 83.765 12.210 83.935 ;
        RECT 10.170 83.085 10.680 83.175 ;
        RECT 8.720 82.275 8.945 82.405 ;
        RECT 9.115 82.335 9.640 82.555 ;
        RECT 9.810 82.915 10.680 83.085 ;
        RECT 8.355 81.685 8.605 82.145 ;
        RECT 8.775 82.135 8.945 82.275 ;
        RECT 9.810 82.135 9.980 82.915 ;
        RECT 10.510 82.845 10.680 82.915 ;
        RECT 10.190 82.665 10.390 82.695 ;
        RECT 10.850 82.665 11.020 83.735 ;
        RECT 11.190 82.845 11.380 83.565 ;
        RECT 10.190 82.365 11.020 82.665 ;
        RECT 11.550 82.635 11.870 83.595 ;
        RECT 8.775 81.965 9.110 82.135 ;
        RECT 9.305 81.965 9.980 82.135 ;
        RECT 10.300 81.685 10.670 82.185 ;
        RECT 10.850 82.135 11.020 82.365 ;
        RECT 11.405 82.305 11.870 82.635 ;
        RECT 12.040 82.925 12.210 83.765 ;
        RECT 12.390 83.735 12.705 84.235 ;
        RECT 12.935 83.505 13.275 84.065 ;
        RECT 12.380 83.130 13.275 83.505 ;
        RECT 13.445 83.225 13.615 84.235 ;
        RECT 13.085 82.925 13.275 83.130 ;
        RECT 13.785 83.175 14.115 84.020 ;
        RECT 15.270 83.855 15.605 84.235 ;
        RECT 13.785 83.095 14.175 83.175 ;
        RECT 13.960 83.045 14.175 83.095 ;
        RECT 12.040 82.595 12.915 82.925 ;
        RECT 13.085 82.595 13.835 82.925 ;
        RECT 12.040 82.135 12.210 82.595 ;
        RECT 13.085 82.425 13.285 82.595 ;
        RECT 14.005 82.465 14.175 83.045 ;
        RECT 13.950 82.425 14.175 82.465 ;
        RECT 10.850 81.965 11.255 82.135 ;
        RECT 11.425 81.965 12.210 82.135 ;
        RECT 12.485 81.685 12.695 82.215 ;
        RECT 12.955 81.900 13.285 82.425 ;
        RECT 13.795 82.340 14.175 82.425 ;
        RECT 15.265 82.365 15.505 83.675 ;
        RECT 15.775 83.265 16.025 84.065 ;
        RECT 16.245 83.515 16.575 84.235 ;
        RECT 16.760 83.265 17.010 84.065 ;
        RECT 17.475 83.435 17.805 84.235 ;
        RECT 17.975 83.805 18.315 84.065 ;
        RECT 15.675 83.095 17.865 83.265 ;
        RECT 13.455 81.685 13.625 82.295 ;
        RECT 13.795 81.905 14.125 82.340 ;
        RECT 15.675 82.185 15.845 83.095 ;
        RECT 17.550 82.925 17.865 83.095 ;
        RECT 15.350 81.855 15.845 82.185 ;
        RECT 16.065 81.960 16.415 82.925 ;
        RECT 16.595 81.955 16.895 82.925 ;
        RECT 17.075 81.955 17.355 82.925 ;
        RECT 17.550 82.675 17.880 82.925 ;
        RECT 17.535 81.685 17.805 82.485 ;
        RECT 18.055 82.405 18.315 83.805 ;
        RECT 18.485 83.070 18.775 84.235 ;
        RECT 18.950 83.845 19.285 84.065 ;
        RECT 20.290 83.855 20.645 84.235 ;
        RECT 18.950 83.225 19.205 83.845 ;
        RECT 19.455 83.685 19.685 83.725 ;
        RECT 20.815 83.685 21.065 84.065 ;
        RECT 19.455 83.485 21.065 83.685 ;
        RECT 19.455 83.395 19.640 83.485 ;
        RECT 20.230 83.475 21.065 83.485 ;
        RECT 21.315 83.455 21.565 84.235 ;
        RECT 21.735 83.385 21.995 84.065 ;
        RECT 19.795 83.285 20.125 83.315 ;
        RECT 19.795 83.225 21.595 83.285 ;
        RECT 18.950 83.115 21.655 83.225 ;
        RECT 18.950 83.055 20.125 83.115 ;
        RECT 21.455 83.080 21.655 83.115 ;
        RECT 18.945 82.675 19.435 82.875 ;
        RECT 19.625 82.675 20.100 82.885 ;
        RECT 17.975 81.895 18.315 82.405 ;
        RECT 18.485 81.685 18.775 82.410 ;
        RECT 18.950 81.685 19.405 82.450 ;
        RECT 19.880 82.275 20.100 82.675 ;
        RECT 20.345 82.675 20.675 82.885 ;
        RECT 20.345 82.275 20.555 82.675 ;
        RECT 20.845 82.640 21.255 82.945 ;
        RECT 21.485 82.505 21.655 83.080 ;
        RECT 21.385 82.385 21.655 82.505 ;
        RECT 20.810 82.340 21.655 82.385 ;
        RECT 20.810 82.215 21.565 82.340 ;
        RECT 20.810 82.065 20.980 82.215 ;
        RECT 21.825 82.195 21.995 83.385 ;
        RECT 22.220 83.365 22.505 84.235 ;
        RECT 22.675 83.605 22.935 84.065 ;
        RECT 23.110 83.775 23.365 84.235 ;
        RECT 23.535 83.605 23.795 84.065 ;
        RECT 22.675 83.435 23.795 83.605 ;
        RECT 23.965 83.435 24.275 84.235 ;
        RECT 22.675 83.185 22.935 83.435 ;
        RECT 24.445 83.265 24.755 84.065 ;
        RECT 22.180 83.015 22.935 83.185 ;
        RECT 23.725 83.095 24.755 83.265 ;
        RECT 24.925 83.095 25.205 84.235 ;
        RECT 22.180 82.505 22.585 83.015 ;
        RECT 23.725 82.845 23.895 83.095 ;
        RECT 22.755 82.675 23.895 82.845 ;
        RECT 22.180 82.335 23.830 82.505 ;
        RECT 24.065 82.355 24.415 82.925 ;
        RECT 21.765 82.185 21.995 82.195 ;
        RECT 19.680 81.855 20.980 82.065 ;
        RECT 21.235 81.685 21.565 82.045 ;
        RECT 21.735 81.855 21.995 82.185 ;
        RECT 22.225 81.685 22.505 82.165 ;
        RECT 22.675 81.945 22.935 82.335 ;
        RECT 23.110 81.685 23.365 82.165 ;
        RECT 23.535 81.945 23.830 82.335 ;
        RECT 24.585 82.185 24.755 83.095 ;
        RECT 25.375 83.085 25.705 84.065 ;
        RECT 25.875 83.095 26.135 84.235 ;
        RECT 26.395 83.565 26.565 84.065 ;
        RECT 26.735 83.735 27.065 84.235 ;
        RECT 26.395 83.395 27.060 83.565 ;
        RECT 24.935 82.655 25.270 82.925 ;
        RECT 25.440 82.485 25.610 83.085 ;
        RECT 25.780 82.675 26.115 82.925 ;
        RECT 26.310 82.575 26.660 83.225 ;
        RECT 24.010 81.685 24.285 82.165 ;
        RECT 24.455 81.855 24.755 82.185 ;
        RECT 24.925 81.685 25.235 82.485 ;
        RECT 25.440 81.855 26.135 82.485 ;
        RECT 26.830 82.405 27.060 83.395 ;
        RECT 26.395 82.235 27.060 82.405 ;
        RECT 26.395 81.945 26.565 82.235 ;
        RECT 26.735 81.685 27.065 82.065 ;
        RECT 27.235 81.945 27.420 84.065 ;
        RECT 27.660 83.775 27.925 84.235 ;
        RECT 28.095 83.640 28.345 84.065 ;
        RECT 28.555 83.790 29.660 83.960 ;
        RECT 28.040 83.510 28.345 83.640 ;
        RECT 27.590 82.315 27.870 83.265 ;
        RECT 28.040 82.405 28.210 83.510 ;
        RECT 28.380 82.725 28.620 83.320 ;
        RECT 28.790 83.255 29.320 83.620 ;
        RECT 28.790 82.555 28.960 83.255 ;
        RECT 29.490 83.175 29.660 83.790 ;
        RECT 29.830 83.435 30.000 84.235 ;
        RECT 30.170 83.735 30.420 84.065 ;
        RECT 30.645 83.765 31.530 83.935 ;
        RECT 29.490 83.085 30.000 83.175 ;
        RECT 28.040 82.275 28.265 82.405 ;
        RECT 28.435 82.335 28.960 82.555 ;
        RECT 29.130 82.915 30.000 83.085 ;
        RECT 27.675 81.685 27.925 82.145 ;
        RECT 28.095 82.135 28.265 82.275 ;
        RECT 29.130 82.135 29.300 82.915 ;
        RECT 29.830 82.845 30.000 82.915 ;
        RECT 29.510 82.665 29.710 82.695 ;
        RECT 30.170 82.665 30.340 83.735 ;
        RECT 30.510 82.845 30.700 83.565 ;
        RECT 29.510 82.365 30.340 82.665 ;
        RECT 30.870 82.635 31.190 83.595 ;
        RECT 28.095 81.965 28.430 82.135 ;
        RECT 28.625 81.965 29.300 82.135 ;
        RECT 29.620 81.685 29.990 82.185 ;
        RECT 30.170 82.135 30.340 82.365 ;
        RECT 30.725 82.305 31.190 82.635 ;
        RECT 31.360 82.925 31.530 83.765 ;
        RECT 31.710 83.735 32.025 84.235 ;
        RECT 32.255 83.505 32.595 84.065 ;
        RECT 31.700 83.130 32.595 83.505 ;
        RECT 32.765 83.225 32.935 84.235 ;
        RECT 32.405 82.925 32.595 83.130 ;
        RECT 33.105 83.175 33.435 84.020 ;
        RECT 33.725 83.175 34.055 84.020 ;
        RECT 34.225 83.225 34.395 84.235 ;
        RECT 34.565 83.505 34.905 84.065 ;
        RECT 35.135 83.735 35.450 84.235 ;
        RECT 35.630 83.765 36.515 83.935 ;
        RECT 33.105 83.095 33.495 83.175 ;
        RECT 33.280 83.045 33.495 83.095 ;
        RECT 31.360 82.595 32.235 82.925 ;
        RECT 32.405 82.595 33.155 82.925 ;
        RECT 31.360 82.135 31.530 82.595 ;
        RECT 32.405 82.425 32.605 82.595 ;
        RECT 33.325 82.465 33.495 83.045 ;
        RECT 33.270 82.425 33.495 82.465 ;
        RECT 30.170 81.965 30.575 82.135 ;
        RECT 30.745 81.965 31.530 82.135 ;
        RECT 31.805 81.685 32.015 82.215 ;
        RECT 32.275 81.900 32.605 82.425 ;
        RECT 33.115 82.340 33.495 82.425 ;
        RECT 33.665 83.095 34.055 83.175 ;
        RECT 34.565 83.130 35.460 83.505 ;
        RECT 33.665 83.045 33.880 83.095 ;
        RECT 33.665 82.465 33.835 83.045 ;
        RECT 34.565 82.925 34.755 83.130 ;
        RECT 35.630 82.925 35.800 83.765 ;
        RECT 36.740 83.735 36.990 84.065 ;
        RECT 34.005 82.595 34.755 82.925 ;
        RECT 34.925 82.595 35.800 82.925 ;
        RECT 33.665 82.425 33.890 82.465 ;
        RECT 34.555 82.425 34.755 82.595 ;
        RECT 33.665 82.340 34.045 82.425 ;
        RECT 32.775 81.685 32.945 82.295 ;
        RECT 33.115 81.905 33.445 82.340 ;
        RECT 33.715 81.905 34.045 82.340 ;
        RECT 34.215 81.685 34.385 82.295 ;
        RECT 34.555 81.900 34.885 82.425 ;
        RECT 35.145 81.685 35.355 82.215 ;
        RECT 35.630 82.135 35.800 82.595 ;
        RECT 35.970 82.635 36.290 83.595 ;
        RECT 36.460 82.845 36.650 83.565 ;
        RECT 36.820 82.665 36.990 83.735 ;
        RECT 37.160 83.435 37.330 84.235 ;
        RECT 37.500 83.790 38.605 83.960 ;
        RECT 37.500 83.175 37.670 83.790 ;
        RECT 38.815 83.640 39.065 84.065 ;
        RECT 39.235 83.775 39.500 84.235 ;
        RECT 37.840 83.255 38.370 83.620 ;
        RECT 38.815 83.510 39.120 83.640 ;
        RECT 37.160 83.085 37.670 83.175 ;
        RECT 37.160 82.915 38.030 83.085 ;
        RECT 37.160 82.845 37.330 82.915 ;
        RECT 37.450 82.665 37.650 82.695 ;
        RECT 35.970 82.305 36.435 82.635 ;
        RECT 36.820 82.365 37.650 82.665 ;
        RECT 36.820 82.135 36.990 82.365 ;
        RECT 35.630 81.965 36.415 82.135 ;
        RECT 36.585 81.965 36.990 82.135 ;
        RECT 37.170 81.685 37.540 82.185 ;
        RECT 37.860 82.135 38.030 82.915 ;
        RECT 38.200 82.555 38.370 83.255 ;
        RECT 38.540 82.725 38.780 83.320 ;
        RECT 38.200 82.335 38.725 82.555 ;
        RECT 38.950 82.405 39.120 83.510 ;
        RECT 38.895 82.275 39.120 82.405 ;
        RECT 39.290 82.315 39.570 83.265 ;
        RECT 38.895 82.135 39.065 82.275 ;
        RECT 37.860 81.965 38.535 82.135 ;
        RECT 38.730 81.965 39.065 82.135 ;
        RECT 39.235 81.685 39.485 82.145 ;
        RECT 39.740 81.945 39.925 84.065 ;
        RECT 40.095 83.735 40.425 84.235 ;
        RECT 40.595 83.565 40.765 84.065 ;
        RECT 40.100 83.395 40.765 83.565 ;
        RECT 40.100 82.405 40.330 83.395 ;
        RECT 40.500 82.575 40.850 83.225 ;
        RECT 41.025 83.145 43.615 84.235 ;
        RECT 41.025 82.455 42.235 82.975 ;
        RECT 42.405 82.625 43.615 83.145 ;
        RECT 44.245 83.070 44.535 84.235 ;
        RECT 44.705 83.145 46.375 84.235 ;
        RECT 44.705 82.455 45.455 82.975 ;
        RECT 45.625 82.625 46.375 83.145 ;
        RECT 46.545 83.095 46.825 84.235 ;
        RECT 46.995 83.085 47.325 84.065 ;
        RECT 47.495 83.095 47.755 84.235 ;
        RECT 47.925 83.680 48.530 84.235 ;
        RECT 48.705 83.725 49.185 84.065 ;
        RECT 49.355 83.690 49.610 84.235 ;
        RECT 47.925 83.580 48.540 83.680 ;
        RECT 48.355 83.555 48.540 83.580 ;
        RECT 46.555 82.655 46.890 82.925 ;
        RECT 47.060 82.485 47.230 83.085 ;
        RECT 47.925 82.960 48.185 83.410 ;
        RECT 48.355 83.310 48.685 83.555 ;
        RECT 48.855 83.235 49.610 83.485 ;
        RECT 49.780 83.365 50.055 84.065 ;
        RECT 48.840 83.200 49.610 83.235 ;
        RECT 48.825 83.190 49.610 83.200 ;
        RECT 48.820 83.175 49.715 83.190 ;
        RECT 48.800 83.160 49.715 83.175 ;
        RECT 48.780 83.150 49.715 83.160 ;
        RECT 48.755 83.140 49.715 83.150 ;
        RECT 48.685 83.110 49.715 83.140 ;
        RECT 48.665 83.080 49.715 83.110 ;
        RECT 48.645 83.050 49.715 83.080 ;
        RECT 48.615 83.025 49.715 83.050 ;
        RECT 48.580 82.990 49.715 83.025 ;
        RECT 48.550 82.985 49.715 82.990 ;
        RECT 48.550 82.980 48.940 82.985 ;
        RECT 48.550 82.970 48.915 82.980 ;
        RECT 48.550 82.965 48.900 82.970 ;
        RECT 48.550 82.960 48.885 82.965 ;
        RECT 47.925 82.955 48.885 82.960 ;
        RECT 47.925 82.945 48.875 82.955 ;
        RECT 47.925 82.940 48.865 82.945 ;
        RECT 47.925 82.930 48.855 82.940 ;
        RECT 47.400 82.675 47.735 82.925 ;
        RECT 47.925 82.920 48.850 82.930 ;
        RECT 47.925 82.915 48.845 82.920 ;
        RECT 47.925 82.900 48.835 82.915 ;
        RECT 47.925 82.885 48.830 82.900 ;
        RECT 47.925 82.860 48.820 82.885 ;
        RECT 47.925 82.790 48.815 82.860 ;
        RECT 40.100 82.235 40.765 82.405 ;
        RECT 40.095 81.685 40.425 82.065 ;
        RECT 40.595 81.945 40.765 82.235 ;
        RECT 41.025 81.685 43.615 82.455 ;
        RECT 44.245 81.685 44.535 82.410 ;
        RECT 44.705 81.685 46.375 82.455 ;
        RECT 46.545 81.685 46.855 82.485 ;
        RECT 47.060 81.855 47.755 82.485 ;
        RECT 47.925 82.235 48.475 82.620 ;
        RECT 48.645 82.065 48.815 82.790 ;
        RECT 47.925 81.895 48.815 82.065 ;
        RECT 48.985 82.390 49.315 82.815 ;
        RECT 49.485 82.590 49.715 82.985 ;
        RECT 48.985 82.365 49.235 82.390 ;
        RECT 48.985 81.905 49.205 82.365 ;
        RECT 49.885 82.335 50.055 83.365 ;
        RECT 49.375 81.685 49.625 82.225 ;
        RECT 49.795 81.855 50.055 82.335 ;
        RECT 50.690 83.095 50.965 84.065 ;
        RECT 51.175 83.435 51.455 84.235 ;
        RECT 51.625 83.725 52.815 84.015 ;
        RECT 51.625 83.385 52.795 83.555 ;
        RECT 51.625 83.265 51.795 83.385 ;
        RECT 51.135 83.095 51.795 83.265 ;
        RECT 50.690 82.360 50.860 83.095 ;
        RECT 51.135 82.925 51.305 83.095 ;
        RECT 52.105 82.925 52.300 83.215 ;
        RECT 52.470 83.095 52.795 83.385 ;
        RECT 52.990 83.095 53.310 84.235 ;
        RECT 53.490 82.925 53.685 83.975 ;
        RECT 53.865 83.385 54.195 84.065 ;
        RECT 54.395 83.435 54.650 84.235 ;
        RECT 53.865 83.105 54.215 83.385 ;
        RECT 55.010 83.265 55.400 83.440 ;
        RECT 55.885 83.435 56.215 84.235 ;
        RECT 56.385 83.445 56.920 84.065 ;
        RECT 57.125 83.800 62.470 84.235 ;
        RECT 51.030 82.595 51.305 82.925 ;
        RECT 51.475 82.595 52.300 82.925 ;
        RECT 52.470 82.595 52.815 82.925 ;
        RECT 53.050 82.875 53.310 82.925 ;
        RECT 53.045 82.705 53.310 82.875 ;
        RECT 53.050 82.595 53.310 82.705 ;
        RECT 53.490 82.595 53.875 82.925 ;
        RECT 54.045 82.725 54.215 83.105 ;
        RECT 54.405 82.895 54.650 83.255 ;
        RECT 55.010 83.095 56.435 83.265 ;
        RECT 51.135 82.425 51.305 82.595 ;
        RECT 54.045 82.555 54.565 82.725 ;
        RECT 50.690 82.015 50.965 82.360 ;
        RECT 51.135 82.255 52.800 82.425 ;
        RECT 51.155 81.685 51.535 82.085 ;
        RECT 51.705 81.905 51.875 82.255 ;
        RECT 52.045 81.685 52.375 82.085 ;
        RECT 52.545 81.905 52.800 82.255 ;
        RECT 52.990 82.215 54.205 82.385 ;
        RECT 52.990 81.865 53.280 82.215 ;
        RECT 53.475 81.685 53.805 82.045 ;
        RECT 53.975 81.910 54.205 82.215 ;
        RECT 54.395 81.990 54.565 82.555 ;
        RECT 54.885 82.365 55.240 82.925 ;
        RECT 55.410 82.195 55.580 83.095 ;
        RECT 55.750 82.365 56.015 82.925 ;
        RECT 56.265 82.595 56.435 83.095 ;
        RECT 56.605 82.425 56.920 83.445 ;
        RECT 54.990 81.685 55.230 82.195 ;
        RECT 55.410 81.865 55.690 82.195 ;
        RECT 55.920 81.685 56.135 82.195 ;
        RECT 56.305 81.855 56.920 82.425 ;
        RECT 58.710 82.230 59.050 83.060 ;
        RECT 60.530 82.550 60.880 83.800 ;
        RECT 62.645 83.145 64.315 84.235 ;
        RECT 62.645 82.455 63.395 82.975 ;
        RECT 63.565 82.625 64.315 83.145 ;
        RECT 65.005 83.095 65.215 84.235 ;
        RECT 65.385 83.085 65.715 84.065 ;
        RECT 65.885 83.095 66.115 84.235 ;
        RECT 66.530 83.265 66.860 84.065 ;
        RECT 67.030 83.435 67.360 84.235 ;
        RECT 67.660 83.265 67.990 84.065 ;
        RECT 68.635 83.435 68.885 84.235 ;
        RECT 66.530 83.095 68.965 83.265 ;
        RECT 69.155 83.095 69.325 84.235 ;
        RECT 69.495 83.095 69.835 84.065 ;
        RECT 57.125 81.685 62.470 82.230 ;
        RECT 62.645 81.685 64.315 82.455 ;
        RECT 65.005 81.685 65.215 82.505 ;
        RECT 65.385 82.485 65.635 83.085 ;
        RECT 65.805 82.675 66.135 82.925 ;
        RECT 66.325 82.675 66.675 82.925 ;
        RECT 65.385 81.855 65.715 82.485 ;
        RECT 65.885 81.685 66.115 82.505 ;
        RECT 66.860 82.465 67.030 83.095 ;
        RECT 67.200 82.675 67.530 82.875 ;
        RECT 67.700 82.675 68.030 82.875 ;
        RECT 68.200 82.675 68.620 82.875 ;
        RECT 68.795 82.845 68.965 83.095 ;
        RECT 68.795 82.675 69.490 82.845 ;
        RECT 69.660 82.535 69.835 83.095 ;
        RECT 70.005 83.070 70.295 84.235 ;
        RECT 70.555 83.565 70.725 84.065 ;
        RECT 70.895 83.735 71.225 84.235 ;
        RECT 70.555 83.395 71.220 83.565 ;
        RECT 70.470 82.575 70.820 83.225 ;
        RECT 66.530 81.855 67.030 82.465 ;
        RECT 67.660 82.335 68.885 82.505 ;
        RECT 69.605 82.485 69.835 82.535 ;
        RECT 67.660 81.855 67.990 82.335 ;
        RECT 68.160 81.685 68.385 82.145 ;
        RECT 68.555 81.855 68.885 82.335 ;
        RECT 69.075 81.685 69.325 82.485 ;
        RECT 69.495 81.855 69.835 82.485 ;
        RECT 70.005 81.685 70.295 82.410 ;
        RECT 70.990 82.405 71.220 83.395 ;
        RECT 70.555 82.235 71.220 82.405 ;
        RECT 70.555 81.945 70.725 82.235 ;
        RECT 70.895 81.685 71.225 82.065 ;
        RECT 71.395 81.945 71.580 84.065 ;
        RECT 71.820 83.775 72.085 84.235 ;
        RECT 72.255 83.640 72.505 84.065 ;
        RECT 72.715 83.790 73.820 83.960 ;
        RECT 72.200 83.510 72.505 83.640 ;
        RECT 71.750 82.315 72.030 83.265 ;
        RECT 72.200 82.405 72.370 83.510 ;
        RECT 72.540 82.725 72.780 83.320 ;
        RECT 72.950 83.255 73.480 83.620 ;
        RECT 72.950 82.555 73.120 83.255 ;
        RECT 73.650 83.175 73.820 83.790 ;
        RECT 73.990 83.435 74.160 84.235 ;
        RECT 74.330 83.735 74.580 84.065 ;
        RECT 74.805 83.765 75.690 83.935 ;
        RECT 73.650 83.085 74.160 83.175 ;
        RECT 72.200 82.275 72.425 82.405 ;
        RECT 72.595 82.335 73.120 82.555 ;
        RECT 73.290 82.915 74.160 83.085 ;
        RECT 71.835 81.685 72.085 82.145 ;
        RECT 72.255 82.135 72.425 82.275 ;
        RECT 73.290 82.135 73.460 82.915 ;
        RECT 73.990 82.845 74.160 82.915 ;
        RECT 73.670 82.665 73.870 82.695 ;
        RECT 74.330 82.665 74.500 83.735 ;
        RECT 74.670 82.845 74.860 83.565 ;
        RECT 73.670 82.365 74.500 82.665 ;
        RECT 75.030 82.635 75.350 83.595 ;
        RECT 72.255 81.965 72.590 82.135 ;
        RECT 72.785 81.965 73.460 82.135 ;
        RECT 73.780 81.685 74.150 82.185 ;
        RECT 74.330 82.135 74.500 82.365 ;
        RECT 74.885 82.305 75.350 82.635 ;
        RECT 75.520 82.925 75.690 83.765 ;
        RECT 75.870 83.735 76.185 84.235 ;
        RECT 76.415 83.505 76.755 84.065 ;
        RECT 75.860 83.130 76.755 83.505 ;
        RECT 76.925 83.225 77.095 84.235 ;
        RECT 76.565 82.925 76.755 83.130 ;
        RECT 77.265 83.175 77.595 84.020 ;
        RECT 77.265 83.095 77.655 83.175 ;
        RECT 77.440 83.045 77.655 83.095 ;
        RECT 75.520 82.595 76.395 82.925 ;
        RECT 76.565 82.595 77.315 82.925 ;
        RECT 75.520 82.135 75.690 82.595 ;
        RECT 76.565 82.425 76.765 82.595 ;
        RECT 77.485 82.465 77.655 83.045 ;
        RECT 77.430 82.425 77.655 82.465 ;
        RECT 74.330 81.965 74.735 82.135 ;
        RECT 74.905 81.965 75.690 82.135 ;
        RECT 75.965 81.685 76.175 82.215 ;
        RECT 76.435 81.900 76.765 82.425 ;
        RECT 77.275 82.340 77.655 82.425 ;
        RECT 77.825 83.095 78.165 84.065 ;
        RECT 78.335 83.095 78.505 84.235 ;
        RECT 78.775 83.435 79.025 84.235 ;
        RECT 79.670 83.265 80.000 84.065 ;
        RECT 80.300 83.435 80.630 84.235 ;
        RECT 80.800 83.265 81.130 84.065 ;
        RECT 78.695 83.095 81.130 83.265 ;
        RECT 81.965 83.145 83.175 84.235 ;
        RECT 77.825 82.485 78.000 83.095 ;
        RECT 78.695 82.845 78.865 83.095 ;
        RECT 78.170 82.675 78.865 82.845 ;
        RECT 79.040 82.675 79.460 82.875 ;
        RECT 79.630 82.675 79.960 82.875 ;
        RECT 80.130 82.675 80.460 82.875 ;
        RECT 76.935 81.685 77.105 82.295 ;
        RECT 77.275 81.905 77.605 82.340 ;
        RECT 77.825 81.855 78.165 82.485 ;
        RECT 78.335 81.685 78.585 82.485 ;
        RECT 78.775 82.335 80.000 82.505 ;
        RECT 78.775 81.855 79.105 82.335 ;
        RECT 79.275 81.685 79.500 82.145 ;
        RECT 79.670 81.855 80.000 82.335 ;
        RECT 80.630 82.465 80.800 83.095 ;
        RECT 80.985 82.675 81.335 82.925 ;
        RECT 81.965 82.605 82.485 83.145 ;
        RECT 80.630 81.855 81.130 82.465 ;
        RECT 82.655 82.435 83.175 82.975 ;
        RECT 81.965 81.685 83.175 82.435 ;
        RECT 5.520 81.515 83.260 81.685 ;
        RECT 5.605 80.765 6.815 81.515 ;
        RECT 7.075 80.965 7.245 81.255 ;
        RECT 7.415 81.135 7.745 81.515 ;
        RECT 7.075 80.795 7.740 80.965 ;
        RECT 5.605 80.225 6.125 80.765 ;
        RECT 6.295 80.055 6.815 80.595 ;
        RECT 5.605 78.965 6.815 80.055 ;
        RECT 6.990 79.975 7.340 80.625 ;
        RECT 7.510 79.805 7.740 80.795 ;
        RECT 7.075 79.635 7.740 79.805 ;
        RECT 7.075 79.135 7.245 79.635 ;
        RECT 7.415 78.965 7.745 79.465 ;
        RECT 7.915 79.135 8.100 81.255 ;
        RECT 8.355 81.055 8.605 81.515 ;
        RECT 8.775 81.065 9.110 81.235 ;
        RECT 9.305 81.065 9.980 81.235 ;
        RECT 8.775 80.925 8.945 81.065 ;
        RECT 8.270 79.935 8.550 80.885 ;
        RECT 8.720 80.795 8.945 80.925 ;
        RECT 8.720 79.690 8.890 80.795 ;
        RECT 9.115 80.645 9.640 80.865 ;
        RECT 9.060 79.880 9.300 80.475 ;
        RECT 9.470 79.945 9.640 80.645 ;
        RECT 9.810 80.285 9.980 81.065 ;
        RECT 10.300 81.015 10.670 81.515 ;
        RECT 10.850 81.065 11.255 81.235 ;
        RECT 11.425 81.065 12.210 81.235 ;
        RECT 10.850 80.835 11.020 81.065 ;
        RECT 10.190 80.535 11.020 80.835 ;
        RECT 11.405 80.565 11.870 80.895 ;
        RECT 10.190 80.505 10.390 80.535 ;
        RECT 10.510 80.285 10.680 80.355 ;
        RECT 9.810 80.115 10.680 80.285 ;
        RECT 10.170 80.025 10.680 80.115 ;
        RECT 8.720 79.560 9.025 79.690 ;
        RECT 9.470 79.580 10.000 79.945 ;
        RECT 8.340 78.965 8.605 79.425 ;
        RECT 8.775 79.135 9.025 79.560 ;
        RECT 10.170 79.410 10.340 80.025 ;
        RECT 9.235 79.240 10.340 79.410 ;
        RECT 10.510 78.965 10.680 79.765 ;
        RECT 10.850 79.465 11.020 80.535 ;
        RECT 11.190 79.635 11.380 80.355 ;
        RECT 11.550 79.605 11.870 80.565 ;
        RECT 12.040 80.605 12.210 81.065 ;
        RECT 12.485 80.985 12.695 81.515 ;
        RECT 12.955 80.775 13.285 81.300 ;
        RECT 13.455 80.905 13.625 81.515 ;
        RECT 13.795 80.860 14.125 81.295 ;
        RECT 13.795 80.775 14.175 80.860 ;
        RECT 13.085 80.605 13.285 80.775 ;
        RECT 13.950 80.735 14.175 80.775 ;
        RECT 12.040 80.275 12.915 80.605 ;
        RECT 13.085 80.275 13.835 80.605 ;
        RECT 10.850 79.135 11.100 79.465 ;
        RECT 12.040 79.435 12.210 80.275 ;
        RECT 13.085 80.070 13.275 80.275 ;
        RECT 14.005 80.155 14.175 80.735 ;
        RECT 13.960 80.105 14.175 80.155 ;
        RECT 12.380 79.695 13.275 80.070 ;
        RECT 13.785 80.025 14.175 80.105 ;
        RECT 14.345 80.795 14.685 81.305 ;
        RECT 11.325 79.265 12.210 79.435 ;
        RECT 12.390 78.965 12.705 79.465 ;
        RECT 12.935 79.135 13.275 79.695 ;
        RECT 13.445 78.965 13.615 79.975 ;
        RECT 13.785 79.180 14.115 80.025 ;
        RECT 14.345 79.395 14.605 80.795 ;
        RECT 14.855 80.715 15.125 81.515 ;
        RECT 14.780 80.275 15.110 80.525 ;
        RECT 15.305 80.275 15.585 81.245 ;
        RECT 15.765 80.275 16.065 81.245 ;
        RECT 16.245 80.275 16.595 81.240 ;
        RECT 16.815 81.015 17.310 81.345 ;
        RECT 14.795 80.105 15.110 80.275 ;
        RECT 16.815 80.105 16.985 81.015 ;
        RECT 14.795 79.935 16.985 80.105 ;
        RECT 14.345 79.135 14.685 79.395 ;
        RECT 14.855 78.965 15.185 79.765 ;
        RECT 15.650 79.135 15.900 79.935 ;
        RECT 16.085 78.965 16.415 79.685 ;
        RECT 16.635 79.135 16.885 79.935 ;
        RECT 17.155 79.525 17.395 80.835 ;
        RECT 17.600 80.775 18.215 81.345 ;
        RECT 18.385 81.005 18.600 81.515 ;
        RECT 18.830 81.005 19.110 81.335 ;
        RECT 19.290 81.005 19.530 81.515 ;
        RECT 19.910 81.055 20.660 81.345 ;
        RECT 21.170 81.055 21.500 81.515 ;
        RECT 17.600 79.755 17.915 80.775 ;
        RECT 18.085 80.105 18.255 80.605 ;
        RECT 18.505 80.275 18.770 80.835 ;
        RECT 18.940 80.105 19.110 81.005 ;
        RECT 19.280 80.275 19.635 80.835 ;
        RECT 18.085 79.935 19.510 80.105 ;
        RECT 17.055 78.965 17.390 79.345 ;
        RECT 17.600 79.135 18.135 79.755 ;
        RECT 18.305 78.965 18.635 79.765 ;
        RECT 19.120 79.760 19.510 79.935 ;
        RECT 19.910 79.765 20.280 81.055 ;
        RECT 21.720 80.865 21.990 81.075 ;
        RECT 20.655 80.695 21.990 80.865 ;
        RECT 22.165 81.055 22.725 81.345 ;
        RECT 22.895 81.055 23.145 81.515 ;
        RECT 20.655 80.525 20.825 80.695 ;
        RECT 20.450 80.275 20.825 80.525 ;
        RECT 20.995 80.285 21.470 80.525 ;
        RECT 21.640 80.285 21.990 80.525 ;
        RECT 20.655 80.105 20.825 80.275 ;
        RECT 20.655 79.935 21.990 80.105 ;
        RECT 21.710 79.775 21.990 79.935 ;
        RECT 19.910 79.595 21.080 79.765 ;
        RECT 20.365 78.965 20.580 79.425 ;
        RECT 20.750 79.135 21.080 79.595 ;
        RECT 21.250 78.965 21.500 79.765 ;
        RECT 22.165 79.685 22.415 81.055 ;
        RECT 23.765 80.885 24.095 81.245 ;
        RECT 24.925 81.135 25.815 81.305 ;
        RECT 22.705 80.695 24.095 80.885 ;
        RECT 22.705 80.605 22.875 80.695 ;
        RECT 22.585 80.275 22.875 80.605 ;
        RECT 24.925 80.580 25.475 80.965 ;
        RECT 23.045 80.275 23.385 80.525 ;
        RECT 23.605 80.275 24.280 80.525 ;
        RECT 25.645 80.410 25.815 81.135 ;
        RECT 22.705 80.025 22.875 80.275 ;
        RECT 22.705 79.855 23.645 80.025 ;
        RECT 24.015 79.915 24.280 80.275 ;
        RECT 24.925 80.340 25.815 80.410 ;
        RECT 25.985 80.810 26.205 81.295 ;
        RECT 26.375 80.975 26.625 81.515 ;
        RECT 26.795 80.865 27.055 81.345 ;
        RECT 25.985 80.385 26.315 80.810 ;
        RECT 24.925 80.315 25.820 80.340 ;
        RECT 24.925 80.300 25.830 80.315 ;
        RECT 24.925 80.285 25.835 80.300 ;
        RECT 24.925 80.280 25.845 80.285 ;
        RECT 24.925 80.270 25.850 80.280 ;
        RECT 24.925 80.260 25.855 80.270 ;
        RECT 24.925 80.255 25.865 80.260 ;
        RECT 24.925 80.245 25.875 80.255 ;
        RECT 24.925 80.240 25.885 80.245 ;
        RECT 22.165 79.135 22.625 79.685 ;
        RECT 22.815 78.965 23.145 79.685 ;
        RECT 23.345 79.305 23.645 79.855 ;
        RECT 24.925 79.790 25.185 80.240 ;
        RECT 25.550 80.235 25.885 80.240 ;
        RECT 25.550 80.230 25.900 80.235 ;
        RECT 25.550 80.220 25.915 80.230 ;
        RECT 25.550 80.215 25.940 80.220 ;
        RECT 26.485 80.215 26.715 80.610 ;
        RECT 25.550 80.210 26.715 80.215 ;
        RECT 25.580 80.175 26.715 80.210 ;
        RECT 25.615 80.150 26.715 80.175 ;
        RECT 25.645 80.120 26.715 80.150 ;
        RECT 25.665 80.090 26.715 80.120 ;
        RECT 25.685 80.060 26.715 80.090 ;
        RECT 25.755 80.050 26.715 80.060 ;
        RECT 25.780 80.040 26.715 80.050 ;
        RECT 25.800 80.025 26.715 80.040 ;
        RECT 25.820 80.010 26.715 80.025 ;
        RECT 25.825 80.000 26.610 80.010 ;
        RECT 25.840 79.965 26.610 80.000 ;
        RECT 25.355 79.645 25.685 79.890 ;
        RECT 25.855 79.715 26.610 79.965 ;
        RECT 26.885 79.835 27.055 80.865 ;
        RECT 27.225 80.695 27.485 81.515 ;
        RECT 27.655 80.695 27.985 81.115 ;
        RECT 28.165 81.030 28.955 81.295 ;
        RECT 27.735 80.605 27.985 80.695 ;
        RECT 23.815 78.965 24.095 79.635 ;
        RECT 25.355 79.620 25.540 79.645 ;
        RECT 24.925 79.520 25.540 79.620 ;
        RECT 24.925 78.965 25.530 79.520 ;
        RECT 25.705 79.135 26.185 79.475 ;
        RECT 26.355 78.965 26.610 79.510 ;
        RECT 26.780 79.135 27.055 79.835 ;
        RECT 27.225 79.645 27.565 80.525 ;
        RECT 27.735 80.355 28.530 80.605 ;
        RECT 27.225 78.965 27.485 79.475 ;
        RECT 27.735 79.135 27.905 80.355 ;
        RECT 28.700 80.175 28.955 81.030 ;
        RECT 29.125 80.875 29.325 81.295 ;
        RECT 29.515 81.055 29.845 81.515 ;
        RECT 29.125 80.355 29.535 80.875 ;
        RECT 30.015 80.865 30.275 81.345 ;
        RECT 29.705 80.175 29.935 80.605 ;
        RECT 28.145 80.005 29.935 80.175 ;
        RECT 28.145 79.640 28.395 80.005 ;
        RECT 28.565 79.645 28.895 79.835 ;
        RECT 29.115 79.710 29.830 80.005 ;
        RECT 30.105 79.835 30.275 80.865 ;
        RECT 31.365 80.790 31.655 81.515 ;
        RECT 31.825 80.765 33.035 81.515 ;
        RECT 31.825 80.225 32.345 80.765 ;
        RECT 33.205 80.695 33.465 81.515 ;
        RECT 33.635 80.695 33.965 81.115 ;
        RECT 34.145 81.030 34.935 81.295 ;
        RECT 33.715 80.605 33.965 80.695 ;
        RECT 28.565 79.470 28.760 79.645 ;
        RECT 28.145 78.965 28.760 79.470 ;
        RECT 28.930 79.135 29.405 79.475 ;
        RECT 29.575 78.965 29.790 79.510 ;
        RECT 30.000 79.135 30.275 79.835 ;
        RECT 31.365 78.965 31.655 80.130 ;
        RECT 32.515 80.055 33.035 80.595 ;
        RECT 31.825 78.965 33.035 80.055 ;
        RECT 33.205 79.645 33.545 80.525 ;
        RECT 33.715 80.355 34.510 80.605 ;
        RECT 33.205 78.965 33.465 79.475 ;
        RECT 33.715 79.135 33.885 80.355 ;
        RECT 34.680 80.175 34.935 81.030 ;
        RECT 35.105 80.875 35.305 81.295 ;
        RECT 35.495 81.055 35.825 81.515 ;
        RECT 35.105 80.355 35.515 80.875 ;
        RECT 35.995 80.865 36.255 81.345 ;
        RECT 36.590 81.005 36.830 81.515 ;
        RECT 37.010 81.005 37.290 81.335 ;
        RECT 37.520 81.005 37.735 81.515 ;
        RECT 35.685 80.175 35.915 80.605 ;
        RECT 34.125 80.005 35.915 80.175 ;
        RECT 34.125 79.640 34.375 80.005 ;
        RECT 34.545 79.645 34.875 79.835 ;
        RECT 35.095 79.710 35.810 80.005 ;
        RECT 36.085 79.835 36.255 80.865 ;
        RECT 36.485 80.275 36.840 80.835 ;
        RECT 37.010 80.105 37.180 81.005 ;
        RECT 37.350 80.275 37.615 80.835 ;
        RECT 37.905 80.775 38.520 81.345 ;
        RECT 37.865 80.105 38.035 80.605 ;
        RECT 34.545 79.470 34.740 79.645 ;
        RECT 34.125 78.965 34.740 79.470 ;
        RECT 34.910 79.135 35.385 79.475 ;
        RECT 35.555 78.965 35.770 79.510 ;
        RECT 35.980 79.135 36.255 79.835 ;
        RECT 36.610 79.935 38.035 80.105 ;
        RECT 36.610 79.760 37.000 79.935 ;
        RECT 37.485 78.965 37.815 79.765 ;
        RECT 38.205 79.755 38.520 80.775 ;
        RECT 38.725 80.745 42.235 81.515 ;
        RECT 42.405 80.765 43.615 81.515 ;
        RECT 38.725 80.225 40.375 80.745 ;
        RECT 40.545 80.055 42.235 80.575 ;
        RECT 42.405 80.225 42.925 80.765 ;
        RECT 43.795 80.705 44.065 81.515 ;
        RECT 44.235 80.705 44.565 81.345 ;
        RECT 44.735 80.705 44.975 81.515 ;
        RECT 43.095 80.055 43.615 80.595 ;
        RECT 43.785 80.275 44.135 80.525 ;
        RECT 44.305 80.105 44.475 80.705 ;
        RECT 45.170 80.675 45.430 81.515 ;
        RECT 45.605 80.770 45.860 81.345 ;
        RECT 46.030 81.135 46.360 81.515 ;
        RECT 46.575 80.965 46.745 81.345 ;
        RECT 46.030 80.795 46.745 80.965 ;
        RECT 44.645 80.275 44.995 80.525 ;
        RECT 37.985 79.135 38.520 79.755 ;
        RECT 38.725 78.965 42.235 80.055 ;
        RECT 42.405 78.965 43.615 80.055 ;
        RECT 43.795 78.965 44.125 80.105 ;
        RECT 44.305 79.935 44.985 80.105 ;
        RECT 44.655 79.150 44.985 79.935 ;
        RECT 45.170 78.965 45.430 80.115 ;
        RECT 45.605 80.040 45.775 80.770 ;
        RECT 46.030 80.605 46.200 80.795 ;
        RECT 47.005 80.775 47.445 81.335 ;
        RECT 47.615 80.775 48.065 81.515 ;
        RECT 48.235 80.945 48.405 81.345 ;
        RECT 48.575 81.115 48.995 81.515 ;
        RECT 49.165 80.945 49.395 81.345 ;
        RECT 48.235 80.775 49.395 80.945 ;
        RECT 49.565 80.775 50.055 81.345 ;
        RECT 45.945 80.275 46.200 80.605 ;
        RECT 46.030 80.065 46.200 80.275 ;
        RECT 46.480 80.245 46.835 80.615 ;
        RECT 45.605 79.135 45.860 80.040 ;
        RECT 46.030 79.895 46.745 80.065 ;
        RECT 46.030 78.965 46.360 79.725 ;
        RECT 46.575 79.135 46.745 79.895 ;
        RECT 47.005 79.765 47.315 80.775 ;
        RECT 47.485 80.155 47.655 80.605 ;
        RECT 47.825 80.325 48.215 80.605 ;
        RECT 48.400 80.275 48.645 80.605 ;
        RECT 47.485 79.985 48.275 80.155 ;
        RECT 47.005 79.135 47.445 79.765 ;
        RECT 47.620 78.965 47.935 79.815 ;
        RECT 48.105 79.305 48.275 79.985 ;
        RECT 48.445 79.475 48.645 80.275 ;
        RECT 48.845 79.475 49.095 80.605 ;
        RECT 49.310 80.275 49.715 80.605 ;
        RECT 49.885 80.105 50.055 80.775 ;
        RECT 49.285 79.935 50.055 80.105 ;
        RECT 50.230 80.840 50.505 81.185 ;
        RECT 50.695 81.115 51.075 81.515 ;
        RECT 51.245 80.945 51.415 81.295 ;
        RECT 51.585 81.115 51.915 81.515 ;
        RECT 52.085 80.945 52.340 81.295 ;
        RECT 50.230 80.105 50.400 80.840 ;
        RECT 50.675 80.775 52.340 80.945 ;
        RECT 52.540 80.945 52.795 81.295 ;
        RECT 52.965 81.115 53.295 81.515 ;
        RECT 53.465 80.945 53.635 81.295 ;
        RECT 53.805 81.115 54.185 81.515 ;
        RECT 52.540 80.775 54.205 80.945 ;
        RECT 54.375 80.840 54.650 81.185 ;
        RECT 54.825 81.135 55.715 81.305 ;
        RECT 50.675 80.605 50.845 80.775 ;
        RECT 54.035 80.605 54.205 80.775 ;
        RECT 50.570 80.275 50.845 80.605 ;
        RECT 51.015 80.275 51.840 80.605 ;
        RECT 52.010 80.275 52.355 80.605 ;
        RECT 52.525 80.275 52.870 80.605 ;
        RECT 53.040 80.275 53.865 80.605 ;
        RECT 54.035 80.275 54.310 80.605 ;
        RECT 50.675 80.105 50.845 80.275 ;
        RECT 49.285 79.305 49.535 79.935 ;
        RECT 48.105 79.135 49.535 79.305 ;
        RECT 49.715 78.965 50.045 79.765 ;
        RECT 50.230 79.135 50.505 80.105 ;
        RECT 50.675 79.935 51.335 80.105 ;
        RECT 51.645 79.985 51.840 80.275 ;
        RECT 51.165 79.815 51.335 79.935 ;
        RECT 52.010 79.815 52.335 80.105 ;
        RECT 50.715 78.965 50.995 79.765 ;
        RECT 51.165 79.645 52.335 79.815 ;
        RECT 52.545 79.815 52.870 80.105 ;
        RECT 53.040 79.985 53.235 80.275 ;
        RECT 54.035 80.105 54.205 80.275 ;
        RECT 54.480 80.105 54.650 80.840 ;
        RECT 54.825 80.580 55.375 80.965 ;
        RECT 55.545 80.410 55.715 81.135 ;
        RECT 53.545 79.935 54.205 80.105 ;
        RECT 53.545 79.815 53.715 79.935 ;
        RECT 52.545 79.645 53.715 79.815 ;
        RECT 51.165 79.185 52.355 79.475 ;
        RECT 52.525 79.185 53.715 79.475 ;
        RECT 53.885 78.965 54.165 79.765 ;
        RECT 54.375 79.135 54.650 80.105 ;
        RECT 54.825 80.340 55.715 80.410 ;
        RECT 55.885 80.810 56.105 81.295 ;
        RECT 56.275 80.975 56.525 81.515 ;
        RECT 56.695 80.865 56.955 81.345 ;
        RECT 55.885 80.385 56.215 80.810 ;
        RECT 54.825 80.315 55.720 80.340 ;
        RECT 54.825 80.300 55.730 80.315 ;
        RECT 54.825 80.285 55.735 80.300 ;
        RECT 54.825 80.280 55.745 80.285 ;
        RECT 54.825 80.270 55.750 80.280 ;
        RECT 54.825 80.260 55.755 80.270 ;
        RECT 54.825 80.255 55.765 80.260 ;
        RECT 54.825 80.245 55.775 80.255 ;
        RECT 54.825 80.240 55.785 80.245 ;
        RECT 54.825 79.790 55.085 80.240 ;
        RECT 55.450 80.235 55.785 80.240 ;
        RECT 55.450 80.230 55.800 80.235 ;
        RECT 55.450 80.220 55.815 80.230 ;
        RECT 55.450 80.215 55.840 80.220 ;
        RECT 56.385 80.215 56.615 80.610 ;
        RECT 55.450 80.210 56.615 80.215 ;
        RECT 55.480 80.175 56.615 80.210 ;
        RECT 55.515 80.150 56.615 80.175 ;
        RECT 55.545 80.120 56.615 80.150 ;
        RECT 55.565 80.090 56.615 80.120 ;
        RECT 55.585 80.060 56.615 80.090 ;
        RECT 55.655 80.050 56.615 80.060 ;
        RECT 55.680 80.040 56.615 80.050 ;
        RECT 55.700 80.025 56.615 80.040 ;
        RECT 55.720 80.010 56.615 80.025 ;
        RECT 55.725 80.000 56.510 80.010 ;
        RECT 55.740 79.965 56.510 80.000 ;
        RECT 55.255 79.645 55.585 79.890 ;
        RECT 55.755 79.715 56.510 79.965 ;
        RECT 56.785 79.835 56.955 80.865 ;
        RECT 57.125 80.790 57.415 81.515 ;
        RECT 57.585 80.865 57.845 81.345 ;
        RECT 58.015 80.975 58.265 81.515 ;
        RECT 55.255 79.620 55.440 79.645 ;
        RECT 54.825 79.520 55.440 79.620 ;
        RECT 54.825 78.965 55.430 79.520 ;
        RECT 55.605 79.135 56.085 79.475 ;
        RECT 56.255 78.965 56.510 79.510 ;
        RECT 56.680 79.135 56.955 79.835 ;
        RECT 57.125 78.965 57.415 80.130 ;
        RECT 57.585 79.835 57.755 80.865 ;
        RECT 58.435 80.835 58.655 81.295 ;
        RECT 58.405 80.810 58.655 80.835 ;
        RECT 57.925 80.215 58.155 80.610 ;
        RECT 58.325 80.385 58.655 80.810 ;
        RECT 58.825 81.135 59.715 81.305 ;
        RECT 58.825 80.410 58.995 81.135 ;
        RECT 59.165 80.580 59.715 80.965 ;
        RECT 59.885 80.765 61.095 81.515 ;
        RECT 58.825 80.340 59.715 80.410 ;
        RECT 58.820 80.315 59.715 80.340 ;
        RECT 58.810 80.300 59.715 80.315 ;
        RECT 58.805 80.285 59.715 80.300 ;
        RECT 58.795 80.280 59.715 80.285 ;
        RECT 58.790 80.270 59.715 80.280 ;
        RECT 58.785 80.260 59.715 80.270 ;
        RECT 58.775 80.255 59.715 80.260 ;
        RECT 58.765 80.245 59.715 80.255 ;
        RECT 58.755 80.240 59.715 80.245 ;
        RECT 58.755 80.235 59.090 80.240 ;
        RECT 58.740 80.230 59.090 80.235 ;
        RECT 58.725 80.220 59.090 80.230 ;
        RECT 58.700 80.215 59.090 80.220 ;
        RECT 57.925 80.210 59.090 80.215 ;
        RECT 57.925 80.175 59.060 80.210 ;
        RECT 57.925 80.150 59.025 80.175 ;
        RECT 57.925 80.120 58.995 80.150 ;
        RECT 57.925 80.090 58.975 80.120 ;
        RECT 57.925 80.060 58.955 80.090 ;
        RECT 57.925 80.050 58.885 80.060 ;
        RECT 57.925 80.040 58.860 80.050 ;
        RECT 57.925 80.025 58.840 80.040 ;
        RECT 57.925 80.010 58.820 80.025 ;
        RECT 58.030 80.000 58.815 80.010 ;
        RECT 58.030 79.965 58.800 80.000 ;
        RECT 57.585 79.135 57.860 79.835 ;
        RECT 58.030 79.715 58.785 79.965 ;
        RECT 58.955 79.645 59.285 79.890 ;
        RECT 59.455 79.790 59.715 80.240 ;
        RECT 59.885 80.225 60.405 80.765 ;
        RECT 61.305 80.695 61.535 81.515 ;
        RECT 61.705 80.715 62.035 81.345 ;
        RECT 60.575 80.055 61.095 80.595 ;
        RECT 61.285 80.275 61.615 80.525 ;
        RECT 61.785 80.115 62.035 80.715 ;
        RECT 62.205 80.695 62.415 81.515 ;
        RECT 62.650 80.675 62.910 81.515 ;
        RECT 63.085 80.770 63.340 81.345 ;
        RECT 63.510 81.135 63.840 81.515 ;
        RECT 64.055 80.965 64.225 81.345 ;
        RECT 64.505 81.005 64.745 81.515 ;
        RECT 64.915 81.005 65.205 81.345 ;
        RECT 65.435 81.005 65.750 81.515 ;
        RECT 63.510 80.795 64.225 80.965 ;
        RECT 59.100 79.620 59.285 79.645 ;
        RECT 59.100 79.520 59.715 79.620 ;
        RECT 58.030 78.965 58.285 79.510 ;
        RECT 58.455 79.135 58.935 79.475 ;
        RECT 59.110 78.965 59.715 79.520 ;
        RECT 59.885 78.965 61.095 80.055 ;
        RECT 61.305 78.965 61.535 80.105 ;
        RECT 61.705 79.135 62.035 80.115 ;
        RECT 62.205 78.965 62.415 80.105 ;
        RECT 62.650 78.965 62.910 80.115 ;
        RECT 63.085 80.040 63.255 80.770 ;
        RECT 63.510 80.605 63.680 80.795 ;
        RECT 63.425 80.275 63.680 80.605 ;
        RECT 63.510 80.065 63.680 80.275 ;
        RECT 63.960 80.245 64.315 80.615 ;
        RECT 64.550 80.495 64.745 80.835 ;
        RECT 64.545 80.325 64.745 80.495 ;
        RECT 64.550 80.275 64.745 80.325 ;
        RECT 64.915 80.105 65.095 81.005 ;
        RECT 65.920 80.945 66.090 81.215 ;
        RECT 66.260 81.115 66.590 81.515 ;
        RECT 65.265 80.275 65.675 80.835 ;
        RECT 65.920 80.775 66.615 80.945 ;
        RECT 65.845 80.105 66.015 80.605 ;
        RECT 63.085 79.135 63.340 80.040 ;
        RECT 63.510 79.895 64.225 80.065 ;
        RECT 63.510 78.965 63.840 79.725 ;
        RECT 64.055 79.135 64.225 79.895 ;
        RECT 64.555 79.935 66.015 80.105 ;
        RECT 64.555 79.760 64.915 79.935 ;
        RECT 66.185 79.765 66.615 80.775 ;
        RECT 66.790 80.695 67.065 81.515 ;
        RECT 67.235 80.875 67.565 81.345 ;
        RECT 67.735 81.045 67.905 81.515 ;
        RECT 68.075 80.875 68.405 81.345 ;
        RECT 68.575 81.045 68.865 81.515 ;
        RECT 67.235 80.865 68.405 80.875 ;
        RECT 67.235 80.695 68.835 80.865 ;
        RECT 66.790 80.325 67.510 80.525 ;
        RECT 67.680 80.325 68.450 80.525 ;
        RECT 68.620 80.155 68.835 80.695 ;
        RECT 65.500 78.965 65.670 79.765 ;
        RECT 65.840 79.595 66.615 79.765 ;
        RECT 66.790 79.935 67.905 80.145 ;
        RECT 65.840 79.135 66.170 79.595 ;
        RECT 66.340 78.965 66.510 79.425 ;
        RECT 66.790 79.135 67.065 79.935 ;
        RECT 67.235 78.965 67.565 79.765 ;
        RECT 67.735 79.305 67.905 79.935 ;
        RECT 68.075 79.935 68.835 80.155 ;
        RECT 70.040 80.775 70.655 81.345 ;
        RECT 70.825 81.005 71.040 81.515 ;
        RECT 71.270 81.005 71.550 81.335 ;
        RECT 71.730 81.005 71.970 81.515 ;
        RECT 72.305 81.055 72.865 81.345 ;
        RECT 73.035 81.055 73.285 81.515 ;
        RECT 68.075 79.475 68.405 79.935 ;
        RECT 68.575 79.305 68.875 79.765 ;
        RECT 67.735 79.135 68.875 79.305 ;
        RECT 70.040 79.755 70.355 80.775 ;
        RECT 70.525 80.105 70.695 80.605 ;
        RECT 70.945 80.275 71.210 80.835 ;
        RECT 71.380 80.105 71.550 81.005 ;
        RECT 71.720 80.275 72.075 80.835 ;
        RECT 70.525 79.935 71.950 80.105 ;
        RECT 70.040 79.135 70.575 79.755 ;
        RECT 70.745 78.965 71.075 79.765 ;
        RECT 71.560 79.760 71.950 79.935 ;
        RECT 72.305 79.685 72.555 81.055 ;
        RECT 73.905 80.885 74.235 81.245 ;
        RECT 72.845 80.695 74.235 80.885 ;
        RECT 74.695 80.965 74.865 81.255 ;
        RECT 75.035 81.135 75.365 81.515 ;
        RECT 74.695 80.795 75.360 80.965 ;
        RECT 72.845 80.605 73.015 80.695 ;
        RECT 72.725 80.275 73.015 80.605 ;
        RECT 73.185 80.275 73.525 80.525 ;
        RECT 73.745 80.275 74.420 80.525 ;
        RECT 72.845 80.025 73.015 80.275 ;
        RECT 72.845 79.855 73.785 80.025 ;
        RECT 74.155 79.915 74.420 80.275 ;
        RECT 74.610 79.975 74.960 80.625 ;
        RECT 72.305 79.135 72.765 79.685 ;
        RECT 72.955 78.965 73.285 79.685 ;
        RECT 73.485 79.305 73.785 79.855 ;
        RECT 75.130 79.805 75.360 80.795 ;
        RECT 74.695 79.635 75.360 79.805 ;
        RECT 73.955 78.965 74.235 79.635 ;
        RECT 74.695 79.135 74.865 79.635 ;
        RECT 75.035 78.965 75.365 79.465 ;
        RECT 75.535 79.135 75.720 81.255 ;
        RECT 75.975 81.055 76.225 81.515 ;
        RECT 76.395 81.065 76.730 81.235 ;
        RECT 76.925 81.065 77.600 81.235 ;
        RECT 76.395 80.925 76.565 81.065 ;
        RECT 75.890 79.935 76.170 80.885 ;
        RECT 76.340 80.795 76.565 80.925 ;
        RECT 76.340 79.690 76.510 80.795 ;
        RECT 76.735 80.645 77.260 80.865 ;
        RECT 76.680 79.880 76.920 80.475 ;
        RECT 77.090 79.945 77.260 80.645 ;
        RECT 77.430 80.285 77.600 81.065 ;
        RECT 77.920 81.015 78.290 81.515 ;
        RECT 78.470 81.065 78.875 81.235 ;
        RECT 79.045 81.065 79.830 81.235 ;
        RECT 78.470 80.835 78.640 81.065 ;
        RECT 77.810 80.535 78.640 80.835 ;
        RECT 79.025 80.565 79.490 80.895 ;
        RECT 77.810 80.505 78.010 80.535 ;
        RECT 78.130 80.285 78.300 80.355 ;
        RECT 77.430 80.115 78.300 80.285 ;
        RECT 77.790 80.025 78.300 80.115 ;
        RECT 76.340 79.560 76.645 79.690 ;
        RECT 77.090 79.580 77.620 79.945 ;
        RECT 75.960 78.965 76.225 79.425 ;
        RECT 76.395 79.135 76.645 79.560 ;
        RECT 77.790 79.410 77.960 80.025 ;
        RECT 76.855 79.240 77.960 79.410 ;
        RECT 78.130 78.965 78.300 79.765 ;
        RECT 78.470 79.465 78.640 80.535 ;
        RECT 78.810 79.635 79.000 80.355 ;
        RECT 79.170 79.605 79.490 80.565 ;
        RECT 79.660 80.605 79.830 81.065 ;
        RECT 80.105 80.985 80.315 81.515 ;
        RECT 80.575 80.775 80.905 81.300 ;
        RECT 81.075 80.905 81.245 81.515 ;
        RECT 81.415 80.860 81.745 81.295 ;
        RECT 81.415 80.775 81.795 80.860 ;
        RECT 80.705 80.605 80.905 80.775 ;
        RECT 81.570 80.735 81.795 80.775 ;
        RECT 81.965 80.765 83.175 81.515 ;
        RECT 79.660 80.275 80.535 80.605 ;
        RECT 80.705 80.275 81.455 80.605 ;
        RECT 78.470 79.135 78.720 79.465 ;
        RECT 79.660 79.435 79.830 80.275 ;
        RECT 80.705 80.070 80.895 80.275 ;
        RECT 81.625 80.155 81.795 80.735 ;
        RECT 81.580 80.105 81.795 80.155 ;
        RECT 80.000 79.695 80.895 80.070 ;
        RECT 81.405 80.025 81.795 80.105 ;
        RECT 81.965 80.055 82.485 80.595 ;
        RECT 82.655 80.225 83.175 80.765 ;
        RECT 78.945 79.265 79.830 79.435 ;
        RECT 80.010 78.965 80.325 79.465 ;
        RECT 80.555 79.135 80.895 79.695 ;
        RECT 81.065 78.965 81.235 79.975 ;
        RECT 81.405 79.180 81.735 80.025 ;
        RECT 81.965 78.965 83.175 80.055 ;
        RECT 5.520 78.795 83.260 78.965 ;
        RECT 5.605 77.705 6.815 78.795 ;
        RECT 5.605 76.995 6.125 77.535 ;
        RECT 6.295 77.165 6.815 77.705 ;
        RECT 7.905 77.925 8.180 78.625 ;
        RECT 8.390 78.250 8.605 78.795 ;
        RECT 8.775 78.285 9.250 78.625 ;
        RECT 9.420 78.290 10.035 78.795 ;
        RECT 9.420 78.115 9.615 78.290 ;
        RECT 5.605 76.245 6.815 76.995 ;
        RECT 7.905 76.895 8.075 77.925 ;
        RECT 8.350 77.755 9.065 78.050 ;
        RECT 9.285 77.925 9.615 78.115 ;
        RECT 9.785 77.755 10.035 78.120 ;
        RECT 8.245 77.585 10.035 77.755 ;
        RECT 8.245 77.155 8.475 77.585 ;
        RECT 7.905 76.415 8.165 76.895 ;
        RECT 8.645 76.885 9.055 77.405 ;
        RECT 8.335 76.245 8.665 76.705 ;
        RECT 8.855 76.465 9.055 76.885 ;
        RECT 9.225 76.730 9.480 77.585 ;
        RECT 10.275 77.405 10.445 78.625 ;
        RECT 10.695 78.285 10.955 78.795 ;
        RECT 9.650 77.155 10.445 77.405 ;
        RECT 10.615 77.235 10.955 78.115 ;
        RECT 12.045 77.655 12.305 78.795 ;
        RECT 12.545 78.285 14.160 78.615 ;
        RECT 12.555 77.485 12.725 78.045 ;
        RECT 12.985 77.945 14.160 78.115 ;
        RECT 14.330 77.995 14.610 78.795 ;
        RECT 12.985 77.655 13.315 77.945 ;
        RECT 13.990 77.825 14.160 77.945 ;
        RECT 13.485 77.485 13.730 77.775 ;
        RECT 13.990 77.655 14.650 77.825 ;
        RECT 14.820 77.655 15.095 78.625 ;
        RECT 15.265 78.285 15.525 78.795 ;
        RECT 14.480 77.485 14.650 77.655 ;
        RECT 12.050 77.235 12.385 77.485 ;
        RECT 10.195 77.065 10.445 77.155 ;
        RECT 12.555 77.155 13.270 77.485 ;
        RECT 13.485 77.155 14.310 77.485 ;
        RECT 14.480 77.155 14.755 77.485 ;
        RECT 12.555 77.065 12.805 77.155 ;
        RECT 9.225 76.465 10.015 76.730 ;
        RECT 10.195 76.645 10.525 77.065 ;
        RECT 10.695 76.245 10.955 77.065 ;
        RECT 12.045 76.245 12.305 77.065 ;
        RECT 12.475 76.645 12.805 77.065 ;
        RECT 14.480 76.985 14.650 77.155 ;
        RECT 12.985 76.815 14.650 76.985 ;
        RECT 14.925 76.920 15.095 77.655 ;
        RECT 15.265 77.235 15.605 78.115 ;
        RECT 15.775 77.405 15.945 78.625 ;
        RECT 16.185 78.290 16.800 78.795 ;
        RECT 16.185 77.755 16.435 78.120 ;
        RECT 16.605 78.115 16.800 78.290 ;
        RECT 16.970 78.285 17.445 78.625 ;
        RECT 17.615 78.250 17.830 78.795 ;
        RECT 16.605 77.925 16.935 78.115 ;
        RECT 17.155 77.755 17.870 78.050 ;
        RECT 18.040 77.925 18.315 78.625 ;
        RECT 16.185 77.585 17.975 77.755 ;
        RECT 15.775 77.155 16.570 77.405 ;
        RECT 15.775 77.065 16.025 77.155 ;
        RECT 12.985 76.415 13.245 76.815 ;
        RECT 13.415 76.245 13.745 76.645 ;
        RECT 13.915 76.465 14.085 76.815 ;
        RECT 14.255 76.245 14.630 76.645 ;
        RECT 14.820 76.575 15.095 76.920 ;
        RECT 15.265 76.245 15.525 77.065 ;
        RECT 15.695 76.645 16.025 77.065 ;
        RECT 16.740 76.730 16.995 77.585 ;
        RECT 16.205 76.465 16.995 76.730 ;
        RECT 17.165 76.885 17.575 77.405 ;
        RECT 17.745 77.155 17.975 77.585 ;
        RECT 18.145 76.895 18.315 77.925 ;
        RECT 18.485 77.630 18.775 78.795 ;
        RECT 19.150 77.825 19.480 78.625 ;
        RECT 19.650 77.995 19.980 78.795 ;
        RECT 20.280 77.825 20.610 78.625 ;
        RECT 21.255 77.995 21.505 78.795 ;
        RECT 19.150 77.655 21.585 77.825 ;
        RECT 21.775 77.655 21.945 78.795 ;
        RECT 22.115 77.655 22.455 78.625 ;
        RECT 22.675 78.335 22.885 78.795 ;
        RECT 23.375 78.205 23.875 78.625 ;
        RECT 18.945 77.235 19.295 77.485 ;
        RECT 19.480 77.025 19.650 77.655 ;
        RECT 19.820 77.235 20.150 77.435 ;
        RECT 20.320 77.235 20.650 77.435 ;
        RECT 20.820 77.235 21.240 77.435 ;
        RECT 21.415 77.405 21.585 77.655 ;
        RECT 21.415 77.235 22.110 77.405 ;
        RECT 17.165 76.465 17.365 76.885 ;
        RECT 17.555 76.245 17.885 76.705 ;
        RECT 18.055 76.415 18.315 76.895 ;
        RECT 18.485 76.245 18.775 76.970 ;
        RECT 19.150 76.415 19.650 77.025 ;
        RECT 20.280 76.895 21.505 77.065 ;
        RECT 22.280 77.045 22.455 77.655 ;
        RECT 20.280 76.415 20.610 76.895 ;
        RECT 20.780 76.245 21.005 76.705 ;
        RECT 21.175 76.415 21.505 76.895 ;
        RECT 21.695 76.245 21.945 77.045 ;
        RECT 22.115 76.415 22.455 77.045 ;
        RECT 22.625 76.825 22.865 78.150 ;
        RECT 23.035 77.995 23.875 78.205 ;
        RECT 23.035 76.985 23.205 77.995 ;
        RECT 23.375 77.575 23.775 77.825 ;
        RECT 24.065 77.775 24.265 78.565 ;
        RECT 23.945 77.605 24.265 77.775 ;
        RECT 24.435 77.615 24.755 78.795 ;
        RECT 24.925 77.655 25.205 78.795 ;
        RECT 25.375 77.645 25.705 78.625 ;
        RECT 25.875 77.655 26.135 78.795 ;
        RECT 27.260 78.005 27.795 78.625 ;
        RECT 23.375 77.155 23.545 77.575 ;
        RECT 23.945 77.405 24.125 77.605 ;
        RECT 23.760 77.235 24.125 77.405 ;
        RECT 24.295 77.235 24.755 77.435 ;
        RECT 24.935 77.215 25.270 77.485 ;
        RECT 25.440 77.045 25.610 77.645 ;
        RECT 25.780 77.235 26.115 77.485 ;
        RECT 23.725 76.985 24.755 77.025 ;
        RECT 23.035 76.805 23.385 76.985 ;
        RECT 23.555 76.855 24.755 76.985 ;
        RECT 23.555 76.635 23.885 76.855 ;
        RECT 22.625 76.455 23.885 76.635 ;
        RECT 24.075 76.245 24.245 76.685 ;
        RECT 24.415 76.440 24.755 76.855 ;
        RECT 24.925 76.245 25.235 77.045 ;
        RECT 25.440 76.415 26.135 77.045 ;
        RECT 27.260 76.985 27.575 78.005 ;
        RECT 27.965 77.995 28.295 78.795 ;
        RECT 28.780 77.825 29.170 78.000 ;
        RECT 27.745 77.655 29.170 77.825 ;
        RECT 29.615 77.785 29.785 78.625 ;
        RECT 29.955 78.455 31.125 78.625 ;
        RECT 29.955 77.955 30.285 78.455 ;
        RECT 30.795 78.415 31.125 78.455 ;
        RECT 31.315 78.375 31.670 78.795 ;
        RECT 30.455 78.195 30.685 78.285 ;
        RECT 31.840 78.195 32.090 78.625 ;
        RECT 30.455 77.955 32.090 78.195 ;
        RECT 32.260 78.035 32.590 78.795 ;
        RECT 32.760 77.955 33.015 78.625 ;
        RECT 27.745 77.155 27.915 77.655 ;
        RECT 27.260 76.415 27.875 76.985 ;
        RECT 28.165 76.925 28.430 77.485 ;
        RECT 28.600 76.755 28.770 77.655 ;
        RECT 29.615 77.615 32.675 77.785 ;
        RECT 28.940 76.925 29.295 77.485 ;
        RECT 29.530 77.235 29.880 77.445 ;
        RECT 30.050 77.235 30.495 77.435 ;
        RECT 30.665 77.235 31.140 77.435 ;
        RECT 29.615 76.895 30.680 77.065 ;
        RECT 28.045 76.245 28.260 76.755 ;
        RECT 28.490 76.425 28.770 76.755 ;
        RECT 28.950 76.245 29.190 76.755 ;
        RECT 29.615 76.415 29.785 76.895 ;
        RECT 29.955 76.245 30.285 76.725 ;
        RECT 30.510 76.665 30.680 76.895 ;
        RECT 30.860 76.835 31.140 77.235 ;
        RECT 31.410 77.235 31.740 77.435 ;
        RECT 31.910 77.235 32.275 77.435 ;
        RECT 31.410 76.835 31.695 77.235 ;
        RECT 32.505 77.065 32.675 77.615 ;
        RECT 31.875 76.895 32.675 77.065 ;
        RECT 31.875 76.665 32.045 76.895 ;
        RECT 32.845 76.825 33.015 77.955 ;
        RECT 33.265 77.735 33.595 78.580 ;
        RECT 33.765 77.785 33.935 78.795 ;
        RECT 34.105 78.065 34.445 78.625 ;
        RECT 34.675 78.295 34.990 78.795 ;
        RECT 35.170 78.325 36.055 78.495 ;
        RECT 33.205 77.655 33.595 77.735 ;
        RECT 34.105 77.690 35.000 78.065 ;
        RECT 33.205 77.605 33.420 77.655 ;
        RECT 33.205 77.025 33.375 77.605 ;
        RECT 34.105 77.485 34.295 77.690 ;
        RECT 35.170 77.485 35.340 78.325 ;
        RECT 36.280 78.295 36.530 78.625 ;
        RECT 33.545 77.155 34.295 77.485 ;
        RECT 34.465 77.155 35.340 77.485 ;
        RECT 33.205 76.985 33.430 77.025 ;
        RECT 34.095 76.985 34.295 77.155 ;
        RECT 33.205 76.900 33.585 76.985 ;
        RECT 32.830 76.755 33.015 76.825 ;
        RECT 32.805 76.745 33.015 76.755 ;
        RECT 30.510 76.415 32.045 76.665 ;
        RECT 32.215 76.245 32.545 76.725 ;
        RECT 32.760 76.415 33.015 76.745 ;
        RECT 33.255 76.465 33.585 76.900 ;
        RECT 33.755 76.245 33.925 76.855 ;
        RECT 34.095 76.460 34.425 76.985 ;
        RECT 34.685 76.245 34.895 76.775 ;
        RECT 35.170 76.695 35.340 77.155 ;
        RECT 35.510 77.195 35.830 78.155 ;
        RECT 36.000 77.405 36.190 78.125 ;
        RECT 36.360 77.225 36.530 78.295 ;
        RECT 36.700 77.995 36.870 78.795 ;
        RECT 37.040 78.350 38.145 78.520 ;
        RECT 37.040 77.735 37.210 78.350 ;
        RECT 38.355 78.200 38.605 78.625 ;
        RECT 38.775 78.335 39.040 78.795 ;
        RECT 37.380 77.815 37.910 78.180 ;
        RECT 38.355 78.070 38.660 78.200 ;
        RECT 36.700 77.645 37.210 77.735 ;
        RECT 36.700 77.475 37.570 77.645 ;
        RECT 36.700 77.405 36.870 77.475 ;
        RECT 36.990 77.225 37.190 77.255 ;
        RECT 35.510 76.865 35.975 77.195 ;
        RECT 36.360 76.925 37.190 77.225 ;
        RECT 36.360 76.695 36.530 76.925 ;
        RECT 35.170 76.525 35.955 76.695 ;
        RECT 36.125 76.525 36.530 76.695 ;
        RECT 36.710 76.245 37.080 76.745 ;
        RECT 37.400 76.695 37.570 77.475 ;
        RECT 37.740 77.115 37.910 77.815 ;
        RECT 38.080 77.285 38.320 77.880 ;
        RECT 37.740 76.895 38.265 77.115 ;
        RECT 38.490 76.965 38.660 78.070 ;
        RECT 38.435 76.835 38.660 76.965 ;
        RECT 38.830 76.875 39.110 77.825 ;
        RECT 38.435 76.695 38.605 76.835 ;
        RECT 37.400 76.525 38.075 76.695 ;
        RECT 38.270 76.525 38.605 76.695 ;
        RECT 38.775 76.245 39.025 76.705 ;
        RECT 39.280 76.505 39.465 78.625 ;
        RECT 39.635 78.295 39.965 78.795 ;
        RECT 40.135 78.125 40.305 78.625 ;
        RECT 39.640 77.955 40.305 78.125 ;
        RECT 39.640 76.965 39.870 77.955 ;
        RECT 40.565 77.925 40.840 78.625 ;
        RECT 41.050 78.250 41.265 78.795 ;
        RECT 41.435 78.285 41.910 78.625 ;
        RECT 42.080 78.290 42.695 78.795 ;
        RECT 42.080 78.115 42.275 78.290 ;
        RECT 40.040 77.135 40.390 77.785 ;
        RECT 39.640 76.795 40.305 76.965 ;
        RECT 39.635 76.245 39.965 76.625 ;
        RECT 40.135 76.505 40.305 76.795 ;
        RECT 40.565 76.895 40.735 77.925 ;
        RECT 41.010 77.755 41.725 78.050 ;
        RECT 41.945 77.925 42.275 78.115 ;
        RECT 42.445 77.755 42.695 78.120 ;
        RECT 40.905 77.585 42.695 77.755 ;
        RECT 40.905 77.155 41.135 77.585 ;
        RECT 40.565 76.415 40.825 76.895 ;
        RECT 41.305 76.885 41.715 77.405 ;
        RECT 40.995 76.245 41.325 76.705 ;
        RECT 41.515 76.465 41.715 76.885 ;
        RECT 41.885 76.730 42.140 77.585 ;
        RECT 42.935 77.405 43.105 78.625 ;
        RECT 43.355 78.285 43.615 78.795 ;
        RECT 42.310 77.155 43.105 77.405 ;
        RECT 43.275 77.235 43.615 78.115 ;
        RECT 44.245 77.630 44.535 78.795 ;
        RECT 44.710 77.655 45.030 78.795 ;
        RECT 45.210 77.485 45.405 78.535 ;
        RECT 45.585 77.945 45.915 78.625 ;
        RECT 46.115 77.995 46.370 78.795 ;
        RECT 45.585 77.665 45.935 77.945 ;
        RECT 44.770 77.435 45.030 77.485 ;
        RECT 44.765 77.265 45.030 77.435 ;
        RECT 44.770 77.155 45.030 77.265 ;
        RECT 45.210 77.155 45.595 77.485 ;
        RECT 45.765 77.285 45.935 77.665 ;
        RECT 46.125 77.455 46.370 77.815 ;
        RECT 42.855 77.065 43.105 77.155 ;
        RECT 45.765 77.115 46.285 77.285 ;
        RECT 41.885 76.465 42.675 76.730 ;
        RECT 42.855 76.645 43.185 77.065 ;
        RECT 43.355 76.245 43.615 77.065 ;
        RECT 44.245 76.245 44.535 76.970 ;
        RECT 44.710 76.775 45.925 76.945 ;
        RECT 44.710 76.425 45.000 76.775 ;
        RECT 45.195 76.245 45.525 76.605 ;
        RECT 45.695 76.470 45.925 76.775 ;
        RECT 46.115 76.550 46.285 77.115 ;
        RECT 46.545 76.525 46.825 78.625 ;
        RECT 47.015 78.035 47.800 78.795 ;
        RECT 48.195 77.965 48.580 78.625 ;
        RECT 48.195 77.865 48.605 77.965 ;
        RECT 46.995 77.655 48.605 77.865 ;
        RECT 48.905 77.775 49.105 78.565 ;
        RECT 46.995 77.055 47.270 77.655 ;
        RECT 48.775 77.605 49.105 77.775 ;
        RECT 49.275 77.615 49.595 78.795 ;
        RECT 49.805 77.655 50.035 78.795 ;
        RECT 50.205 77.645 50.535 78.625 ;
        RECT 50.705 77.655 50.915 78.795 ;
        RECT 51.350 77.825 51.680 78.625 ;
        RECT 51.850 77.995 52.180 78.795 ;
        RECT 52.480 77.825 52.810 78.625 ;
        RECT 53.455 77.995 53.705 78.795 ;
        RECT 51.350 77.655 53.785 77.825 ;
        RECT 53.975 77.655 54.145 78.795 ;
        RECT 54.315 77.655 54.655 78.625 ;
        RECT 48.775 77.485 48.955 77.605 ;
        RECT 47.440 77.235 47.795 77.485 ;
        RECT 47.990 77.235 48.455 77.485 ;
        RECT 48.625 77.235 48.955 77.485 ;
        RECT 49.130 77.235 49.595 77.435 ;
        RECT 49.785 77.235 50.115 77.485 ;
        RECT 46.995 76.875 48.245 77.055 ;
        RECT 47.880 76.805 48.245 76.875 ;
        RECT 48.415 76.855 49.595 77.025 ;
        RECT 47.055 76.245 47.225 76.705 ;
        RECT 48.415 76.635 48.745 76.855 ;
        RECT 47.495 76.455 48.745 76.635 ;
        RECT 48.915 76.245 49.085 76.685 ;
        RECT 49.255 76.440 49.595 76.855 ;
        RECT 49.805 76.245 50.035 77.065 ;
        RECT 50.285 77.045 50.535 77.645 ;
        RECT 51.145 77.235 51.495 77.485 ;
        RECT 50.205 76.415 50.535 77.045 ;
        RECT 50.705 76.245 50.915 77.065 ;
        RECT 51.680 77.025 51.850 77.655 ;
        RECT 52.020 77.235 52.350 77.435 ;
        RECT 52.520 77.235 52.850 77.435 ;
        RECT 53.020 77.235 53.440 77.435 ;
        RECT 53.615 77.405 53.785 77.655 ;
        RECT 53.615 77.235 54.310 77.405 ;
        RECT 51.350 76.415 51.850 77.025 ;
        RECT 52.480 76.895 53.705 77.065 ;
        RECT 54.480 77.045 54.655 77.655 ;
        RECT 55.900 77.785 56.200 78.625 ;
        RECT 56.395 77.955 56.645 78.795 ;
        RECT 57.235 78.205 58.040 78.625 ;
        RECT 56.815 78.035 58.380 78.205 ;
        RECT 56.815 77.785 56.985 78.035 ;
        RECT 55.900 77.615 56.985 77.785 ;
        RECT 55.745 77.155 56.075 77.445 ;
        RECT 52.480 76.415 52.810 76.895 ;
        RECT 52.980 76.245 53.205 76.705 ;
        RECT 53.375 76.415 53.705 76.895 ;
        RECT 53.895 76.245 54.145 77.045 ;
        RECT 54.315 76.415 54.655 77.045 ;
        RECT 56.245 76.985 56.415 77.615 ;
        RECT 57.155 77.485 57.475 77.865 ;
        RECT 57.665 77.775 58.040 77.865 ;
        RECT 57.645 77.605 58.040 77.775 ;
        RECT 58.210 77.785 58.380 78.035 ;
        RECT 58.550 77.955 58.880 78.795 ;
        RECT 59.050 78.035 59.715 78.625 ;
        RECT 58.210 77.615 59.130 77.785 ;
        RECT 56.585 77.235 56.915 77.445 ;
        RECT 57.095 77.235 57.475 77.485 ;
        RECT 57.665 77.445 58.040 77.605 ;
        RECT 58.960 77.445 59.130 77.615 ;
        RECT 57.665 77.235 58.150 77.445 ;
        RECT 58.340 77.235 58.790 77.445 ;
        RECT 58.960 77.235 59.295 77.445 ;
        RECT 59.465 77.065 59.715 78.035 ;
        RECT 59.890 78.405 60.225 78.625 ;
        RECT 61.230 78.415 61.585 78.795 ;
        RECT 59.890 77.785 60.145 78.405 ;
        RECT 60.395 78.245 60.625 78.285 ;
        RECT 61.755 78.245 62.005 78.625 ;
        RECT 60.395 78.045 62.005 78.245 ;
        RECT 60.395 77.955 60.580 78.045 ;
        RECT 61.170 78.035 62.005 78.045 ;
        RECT 62.255 78.015 62.505 78.795 ;
        RECT 62.675 77.945 62.935 78.625 ;
        RECT 60.735 77.845 61.065 77.875 ;
        RECT 60.735 77.785 62.535 77.845 ;
        RECT 59.890 77.675 62.595 77.785 ;
        RECT 59.890 77.615 61.065 77.675 ;
        RECT 62.395 77.640 62.595 77.675 ;
        RECT 59.885 77.235 60.375 77.435 ;
        RECT 60.565 77.235 61.040 77.445 ;
        RECT 55.905 76.805 56.415 76.985 ;
        RECT 56.820 76.895 58.520 77.065 ;
        RECT 56.820 76.805 57.205 76.895 ;
        RECT 55.905 76.415 56.235 76.805 ;
        RECT 56.405 76.465 57.590 76.635 ;
        RECT 57.850 76.245 58.020 76.715 ;
        RECT 58.190 76.430 58.520 76.895 ;
        RECT 58.690 76.245 58.860 77.065 ;
        RECT 59.030 76.425 59.715 77.065 ;
        RECT 59.890 76.245 60.345 77.010 ;
        RECT 60.820 76.835 61.040 77.235 ;
        RECT 61.285 77.235 61.615 77.445 ;
        RECT 61.285 76.835 61.495 77.235 ;
        RECT 61.785 77.200 62.195 77.505 ;
        RECT 62.425 77.065 62.595 77.640 ;
        RECT 62.325 76.945 62.595 77.065 ;
        RECT 61.750 76.900 62.595 76.945 ;
        RECT 61.750 76.775 62.505 76.900 ;
        RECT 61.750 76.625 61.920 76.775 ;
        RECT 62.765 76.755 62.935 77.945 ;
        RECT 63.290 77.825 63.680 78.000 ;
        RECT 64.165 77.995 64.495 78.795 ;
        RECT 64.665 78.005 65.200 78.625 ;
        RECT 66.325 78.290 66.955 78.795 ;
        RECT 63.290 77.655 64.715 77.825 ;
        RECT 63.165 76.925 63.520 77.485 ;
        RECT 63.690 76.755 63.860 77.655 ;
        RECT 64.030 76.925 64.295 77.485 ;
        RECT 64.545 77.155 64.715 77.655 ;
        RECT 64.885 76.985 65.200 78.005 ;
        RECT 66.340 77.755 66.595 78.120 ;
        RECT 66.765 78.115 66.955 78.290 ;
        RECT 67.135 78.285 67.610 78.625 ;
        RECT 66.765 77.925 67.095 78.115 ;
        RECT 67.320 77.755 67.570 78.050 ;
        RECT 67.795 77.950 68.010 78.795 ;
        RECT 68.210 77.955 68.485 78.625 ;
        RECT 66.340 77.585 68.130 77.755 ;
        RECT 68.315 77.605 68.485 77.955 ;
        RECT 68.655 77.785 68.915 78.795 ;
        RECT 70.005 77.630 70.295 78.795 ;
        RECT 70.465 78.290 71.095 78.795 ;
        RECT 70.480 77.755 70.735 78.120 ;
        RECT 70.905 78.115 71.095 78.290 ;
        RECT 71.275 78.285 71.750 78.625 ;
        RECT 70.905 77.925 71.235 78.115 ;
        RECT 71.460 77.755 71.710 78.050 ;
        RECT 71.935 77.950 72.150 78.795 ;
        RECT 72.350 77.955 72.625 78.625 ;
        RECT 62.705 76.745 62.935 76.755 ;
        RECT 60.620 76.415 61.920 76.625 ;
        RECT 62.175 76.245 62.505 76.605 ;
        RECT 62.675 76.415 62.935 76.745 ;
        RECT 63.270 76.245 63.510 76.755 ;
        RECT 63.690 76.425 63.970 76.755 ;
        RECT 64.200 76.245 64.415 76.755 ;
        RECT 64.585 76.415 65.200 76.985 ;
        RECT 66.325 76.925 66.710 77.405 ;
        RECT 66.880 76.730 67.135 77.585 ;
        RECT 66.345 76.465 67.135 76.730 ;
        RECT 67.305 76.910 67.715 77.405 ;
        RECT 67.900 77.155 68.130 77.585 ;
        RECT 68.300 77.085 68.915 77.605 ;
        RECT 70.480 77.585 72.270 77.755 ;
        RECT 72.455 77.605 72.625 77.955 ;
        RECT 72.795 77.785 73.055 78.795 ;
        RECT 73.225 77.655 73.485 78.795 ;
        RECT 73.655 77.825 73.985 78.625 ;
        RECT 74.155 77.995 74.325 78.795 ;
        RECT 74.495 77.825 74.825 78.625 ;
        RECT 74.995 77.995 75.250 78.795 ;
        RECT 75.530 77.845 75.795 78.615 ;
        RECT 75.965 78.075 76.295 78.795 ;
        RECT 76.485 78.255 76.745 78.615 ;
        RECT 76.915 78.425 77.245 78.795 ;
        RECT 77.415 78.255 77.675 78.615 ;
        RECT 76.485 78.025 77.675 78.255 ;
        RECT 78.245 77.845 78.535 78.615 ;
        RECT 73.655 77.655 75.355 77.825 ;
        RECT 67.305 76.465 67.535 76.910 ;
        RECT 68.300 76.875 68.470 77.085 ;
        RECT 67.715 76.245 68.045 76.740 ;
        RECT 68.220 76.415 68.470 76.875 ;
        RECT 68.640 76.245 68.915 76.905 ;
        RECT 70.005 76.245 70.295 76.970 ;
        RECT 70.465 76.925 70.850 77.405 ;
        RECT 71.020 76.730 71.275 77.585 ;
        RECT 70.485 76.465 71.275 76.730 ;
        RECT 71.445 76.910 71.855 77.405 ;
        RECT 72.040 77.155 72.270 77.585 ;
        RECT 72.440 77.085 73.055 77.605 ;
        RECT 73.225 77.235 73.985 77.485 ;
        RECT 74.155 77.235 74.905 77.485 ;
        RECT 71.445 76.465 71.675 76.910 ;
        RECT 72.440 76.875 72.610 77.085 ;
        RECT 75.075 77.065 75.355 77.655 ;
        RECT 71.855 76.245 72.185 76.740 ;
        RECT 72.360 76.415 72.610 76.875 ;
        RECT 72.780 76.245 73.055 76.905 ;
        RECT 73.225 76.875 74.325 77.045 ;
        RECT 73.225 76.415 73.565 76.875 ;
        RECT 73.735 76.245 73.905 76.705 ;
        RECT 74.075 76.625 74.325 76.875 ;
        RECT 74.495 76.815 75.355 77.065 ;
        RECT 74.915 76.625 75.245 76.645 ;
        RECT 74.075 76.415 75.245 76.625 ;
        RECT 75.530 76.425 75.865 77.845 ;
        RECT 76.040 77.665 78.535 77.845 ;
        RECT 78.745 77.945 79.005 78.625 ;
        RECT 79.175 78.015 79.425 78.795 ;
        RECT 79.675 78.245 79.925 78.625 ;
        RECT 80.095 78.415 80.450 78.795 ;
        RECT 81.455 78.405 81.790 78.625 ;
        RECT 81.055 78.245 81.285 78.285 ;
        RECT 79.675 78.045 81.285 78.245 ;
        RECT 79.675 78.035 80.510 78.045 ;
        RECT 81.100 77.955 81.285 78.045 ;
        RECT 76.040 76.975 76.265 77.665 ;
        RECT 76.465 77.155 76.745 77.485 ;
        RECT 76.925 77.155 77.500 77.485 ;
        RECT 77.680 77.155 78.115 77.485 ;
        RECT 78.295 77.155 78.565 77.485 ;
        RECT 76.040 76.785 78.525 76.975 ;
        RECT 76.045 76.245 76.790 76.615 ;
        RECT 77.355 76.425 77.610 76.785 ;
        RECT 77.790 76.245 78.120 76.615 ;
        RECT 78.300 76.425 78.525 76.785 ;
        RECT 78.745 76.745 78.915 77.945 ;
        RECT 80.615 77.845 80.945 77.875 ;
        RECT 79.145 77.785 80.945 77.845 ;
        RECT 81.535 77.785 81.790 78.405 ;
        RECT 79.085 77.675 81.790 77.785 ;
        RECT 79.085 77.640 79.285 77.675 ;
        RECT 79.085 77.065 79.255 77.640 ;
        RECT 80.615 77.615 81.790 77.675 ;
        RECT 81.965 77.705 83.175 78.795 ;
        RECT 79.485 77.200 79.895 77.505 ;
        RECT 80.065 77.235 80.395 77.445 ;
        RECT 79.085 76.945 79.355 77.065 ;
        RECT 79.085 76.900 79.930 76.945 ;
        RECT 79.175 76.775 79.930 76.900 ;
        RECT 80.185 76.835 80.395 77.235 ;
        RECT 80.640 77.235 81.115 77.445 ;
        RECT 81.305 77.235 81.795 77.435 ;
        RECT 80.640 76.835 80.860 77.235 ;
        RECT 81.965 77.165 82.485 77.705 ;
        RECT 78.745 76.415 79.005 76.745 ;
        RECT 79.760 76.625 79.930 76.775 ;
        RECT 79.175 76.245 79.505 76.605 ;
        RECT 79.760 76.415 81.060 76.625 ;
        RECT 81.335 76.245 81.790 77.010 ;
        RECT 82.655 76.995 83.175 77.535 ;
        RECT 81.965 76.245 83.175 76.995 ;
        RECT 5.520 76.075 83.260 76.245 ;
        RECT 5.605 75.325 6.815 76.075 ;
        RECT 5.605 74.785 6.125 75.325 ;
        RECT 6.985 75.305 9.575 76.075 ;
        RECT 6.295 74.615 6.815 75.155 ;
        RECT 6.985 74.785 8.195 75.305 ;
        RECT 9.755 75.265 10.025 76.075 ;
        RECT 10.195 75.265 10.525 75.905 ;
        RECT 10.695 75.265 10.935 76.075 ;
        RECT 11.125 75.325 12.335 76.075 ;
        RECT 8.365 74.615 9.575 75.135 ;
        RECT 9.745 74.835 10.095 75.085 ;
        RECT 10.265 74.665 10.435 75.265 ;
        RECT 10.605 74.835 10.955 75.085 ;
        RECT 11.125 74.785 11.645 75.325 ;
        RECT 12.515 75.265 12.785 76.075 ;
        RECT 12.955 75.265 13.285 75.905 ;
        RECT 13.455 75.265 13.695 76.075 ;
        RECT 13.885 75.530 19.230 76.075 ;
        RECT 5.605 73.525 6.815 74.615 ;
        RECT 6.985 73.525 9.575 74.615 ;
        RECT 9.755 73.525 10.085 74.665 ;
        RECT 10.265 74.495 10.945 74.665 ;
        RECT 11.815 74.615 12.335 75.155 ;
        RECT 12.505 74.835 12.855 75.085 ;
        RECT 13.025 74.665 13.195 75.265 ;
        RECT 13.365 74.835 13.715 75.085 ;
        RECT 15.470 74.700 15.810 75.530 ;
        RECT 19.405 75.305 22.915 76.075 ;
        RECT 23.085 75.325 24.295 76.075 ;
        RECT 24.500 75.335 25.115 75.905 ;
        RECT 25.285 75.565 25.500 76.075 ;
        RECT 25.730 75.565 26.010 75.895 ;
        RECT 26.190 75.565 26.430 76.075 ;
        RECT 10.615 73.710 10.945 74.495 ;
        RECT 11.125 73.525 12.335 74.615 ;
        RECT 12.515 73.525 12.845 74.665 ;
        RECT 13.025 74.495 13.705 74.665 ;
        RECT 13.375 73.710 13.705 74.495 ;
        RECT 17.290 73.960 17.640 75.210 ;
        RECT 19.405 74.785 21.055 75.305 ;
        RECT 21.225 74.615 22.915 75.135 ;
        RECT 23.085 74.785 23.605 75.325 ;
        RECT 23.775 74.615 24.295 75.155 ;
        RECT 13.885 73.525 19.230 73.960 ;
        RECT 19.405 73.525 22.915 74.615 ;
        RECT 23.085 73.525 24.295 74.615 ;
        RECT 24.500 74.315 24.815 75.335 ;
        RECT 24.985 74.665 25.155 75.165 ;
        RECT 25.405 74.835 25.670 75.395 ;
        RECT 25.840 74.665 26.010 75.565 ;
        RECT 26.965 75.445 27.295 75.805 ;
        RECT 27.915 75.615 28.165 76.075 ;
        RECT 28.335 75.615 28.895 75.905 ;
        RECT 26.180 74.835 26.535 75.395 ;
        RECT 26.965 75.255 28.355 75.445 ;
        RECT 28.185 75.165 28.355 75.255 ;
        RECT 26.780 74.835 27.455 75.085 ;
        RECT 27.675 74.835 28.015 75.085 ;
        RECT 28.185 74.835 28.475 75.165 ;
        RECT 24.985 74.495 26.410 74.665 ;
        RECT 24.500 73.695 25.035 74.315 ;
        RECT 25.205 73.525 25.535 74.325 ;
        RECT 26.020 74.320 26.410 74.495 ;
        RECT 26.780 74.475 27.045 74.835 ;
        RECT 28.185 74.585 28.355 74.835 ;
        RECT 27.415 74.415 28.355 74.585 ;
        RECT 26.965 73.525 27.245 74.195 ;
        RECT 27.415 73.865 27.715 74.415 ;
        RECT 28.645 74.245 28.895 75.615 ;
        RECT 29.230 75.565 29.470 76.075 ;
        RECT 29.650 75.565 29.930 75.895 ;
        RECT 30.160 75.565 30.375 76.075 ;
        RECT 29.125 74.835 29.480 75.395 ;
        RECT 29.650 74.665 29.820 75.565 ;
        RECT 29.990 74.835 30.255 75.395 ;
        RECT 30.545 75.335 31.160 75.905 ;
        RECT 31.365 75.350 31.655 76.075 ;
        RECT 32.375 75.525 32.545 75.815 ;
        RECT 32.715 75.695 33.045 76.075 ;
        RECT 32.375 75.355 33.040 75.525 ;
        RECT 30.505 74.665 30.675 75.165 ;
        RECT 29.250 74.495 30.675 74.665 ;
        RECT 29.250 74.320 29.640 74.495 ;
        RECT 27.915 73.525 28.245 74.245 ;
        RECT 28.435 73.695 28.895 74.245 ;
        RECT 30.125 73.525 30.455 74.325 ;
        RECT 30.845 74.315 31.160 75.335 ;
        RECT 30.625 73.695 31.160 74.315 ;
        RECT 31.365 73.525 31.655 74.690 ;
        RECT 32.290 74.535 32.640 75.185 ;
        RECT 32.810 74.365 33.040 75.355 ;
        RECT 32.375 74.195 33.040 74.365 ;
        RECT 32.375 73.695 32.545 74.195 ;
        RECT 32.715 73.525 33.045 74.025 ;
        RECT 33.215 73.695 33.400 75.815 ;
        RECT 33.655 75.615 33.905 76.075 ;
        RECT 34.075 75.625 34.410 75.795 ;
        RECT 34.605 75.625 35.280 75.795 ;
        RECT 34.075 75.485 34.245 75.625 ;
        RECT 33.570 74.495 33.850 75.445 ;
        RECT 34.020 75.355 34.245 75.485 ;
        RECT 34.020 74.250 34.190 75.355 ;
        RECT 34.415 75.205 34.940 75.425 ;
        RECT 34.360 74.440 34.600 75.035 ;
        RECT 34.770 74.505 34.940 75.205 ;
        RECT 35.110 74.845 35.280 75.625 ;
        RECT 35.600 75.575 35.970 76.075 ;
        RECT 36.150 75.625 36.555 75.795 ;
        RECT 36.725 75.625 37.510 75.795 ;
        RECT 36.150 75.395 36.320 75.625 ;
        RECT 35.490 75.095 36.320 75.395 ;
        RECT 36.705 75.125 37.170 75.455 ;
        RECT 35.490 75.065 35.690 75.095 ;
        RECT 35.810 74.845 35.980 74.915 ;
        RECT 35.110 74.675 35.980 74.845 ;
        RECT 35.470 74.585 35.980 74.675 ;
        RECT 34.020 74.120 34.325 74.250 ;
        RECT 34.770 74.140 35.300 74.505 ;
        RECT 33.640 73.525 33.905 73.985 ;
        RECT 34.075 73.695 34.325 74.120 ;
        RECT 35.470 73.970 35.640 74.585 ;
        RECT 34.535 73.800 35.640 73.970 ;
        RECT 35.810 73.525 35.980 74.325 ;
        RECT 36.150 74.025 36.320 75.095 ;
        RECT 36.490 74.195 36.680 74.915 ;
        RECT 36.850 74.165 37.170 75.125 ;
        RECT 37.340 75.165 37.510 75.625 ;
        RECT 37.785 75.545 37.995 76.075 ;
        RECT 38.255 75.335 38.585 75.860 ;
        RECT 38.755 75.465 38.925 76.075 ;
        RECT 39.095 75.420 39.425 75.855 ;
        RECT 39.095 75.335 39.475 75.420 ;
        RECT 38.385 75.165 38.585 75.335 ;
        RECT 39.250 75.295 39.475 75.335 ;
        RECT 37.340 74.835 38.215 75.165 ;
        RECT 38.385 74.835 39.135 75.165 ;
        RECT 36.150 73.695 36.400 74.025 ;
        RECT 37.340 73.995 37.510 74.835 ;
        RECT 38.385 74.630 38.575 74.835 ;
        RECT 39.305 74.715 39.475 75.295 ;
        RECT 39.645 75.325 40.855 76.075 ;
        RECT 41.115 75.525 41.285 75.815 ;
        RECT 41.455 75.695 41.785 76.075 ;
        RECT 41.115 75.355 41.780 75.525 ;
        RECT 39.645 74.785 40.165 75.325 ;
        RECT 39.260 74.665 39.475 74.715 ;
        RECT 37.680 74.255 38.575 74.630 ;
        RECT 39.085 74.585 39.475 74.665 ;
        RECT 40.335 74.615 40.855 75.155 ;
        RECT 36.625 73.825 37.510 73.995 ;
        RECT 37.690 73.525 38.005 74.025 ;
        RECT 38.235 73.695 38.575 74.255 ;
        RECT 38.745 73.525 38.915 74.535 ;
        RECT 39.085 73.740 39.415 74.585 ;
        RECT 39.645 73.525 40.855 74.615 ;
        RECT 41.030 74.535 41.380 75.185 ;
        RECT 41.550 74.365 41.780 75.355 ;
        RECT 41.115 74.195 41.780 74.365 ;
        RECT 41.115 73.695 41.285 74.195 ;
        RECT 41.455 73.525 41.785 74.025 ;
        RECT 41.955 73.695 42.140 75.815 ;
        RECT 42.395 75.615 42.645 76.075 ;
        RECT 42.815 75.625 43.150 75.795 ;
        RECT 43.345 75.625 44.020 75.795 ;
        RECT 42.815 75.485 42.985 75.625 ;
        RECT 42.310 74.495 42.590 75.445 ;
        RECT 42.760 75.355 42.985 75.485 ;
        RECT 42.760 74.250 42.930 75.355 ;
        RECT 43.155 75.205 43.680 75.425 ;
        RECT 43.100 74.440 43.340 75.035 ;
        RECT 43.510 74.505 43.680 75.205 ;
        RECT 43.850 74.845 44.020 75.625 ;
        RECT 44.340 75.575 44.710 76.075 ;
        RECT 44.890 75.625 45.295 75.795 ;
        RECT 45.465 75.625 46.250 75.795 ;
        RECT 44.890 75.395 45.060 75.625 ;
        RECT 44.230 75.095 45.060 75.395 ;
        RECT 45.445 75.125 45.910 75.455 ;
        RECT 44.230 75.065 44.430 75.095 ;
        RECT 44.550 74.845 44.720 74.915 ;
        RECT 43.850 74.675 44.720 74.845 ;
        RECT 44.210 74.585 44.720 74.675 ;
        RECT 42.760 74.120 43.065 74.250 ;
        RECT 43.510 74.140 44.040 74.505 ;
        RECT 42.380 73.525 42.645 73.985 ;
        RECT 42.815 73.695 43.065 74.120 ;
        RECT 44.210 73.970 44.380 74.585 ;
        RECT 43.275 73.800 44.380 73.970 ;
        RECT 44.550 73.525 44.720 74.325 ;
        RECT 44.890 74.025 45.060 75.095 ;
        RECT 45.230 74.195 45.420 74.915 ;
        RECT 45.590 74.165 45.910 75.125 ;
        RECT 46.080 75.165 46.250 75.625 ;
        RECT 46.525 75.545 46.735 76.075 ;
        RECT 46.995 75.335 47.325 75.860 ;
        RECT 47.495 75.465 47.665 76.075 ;
        RECT 47.835 75.420 48.165 75.855 ;
        RECT 48.390 75.600 48.725 75.860 ;
        RECT 48.895 75.675 49.225 76.075 ;
        RECT 49.395 75.675 51.010 75.845 ;
        RECT 47.835 75.335 48.215 75.420 ;
        RECT 47.125 75.165 47.325 75.335 ;
        RECT 47.990 75.295 48.215 75.335 ;
        RECT 46.080 74.835 46.955 75.165 ;
        RECT 47.125 74.835 47.875 75.165 ;
        RECT 44.890 73.695 45.140 74.025 ;
        RECT 46.080 73.995 46.250 74.835 ;
        RECT 47.125 74.630 47.315 74.835 ;
        RECT 48.045 74.715 48.215 75.295 ;
        RECT 48.000 74.665 48.215 74.715 ;
        RECT 46.420 74.255 47.315 74.630 ;
        RECT 47.825 74.585 48.215 74.665 ;
        RECT 45.365 73.825 46.250 73.995 ;
        RECT 46.430 73.525 46.745 74.025 ;
        RECT 46.975 73.695 47.315 74.255 ;
        RECT 47.485 73.525 47.655 74.535 ;
        RECT 47.825 73.740 48.155 74.585 ;
        RECT 48.390 74.245 48.645 75.600 ;
        RECT 49.395 75.505 49.565 75.675 ;
        RECT 49.005 75.335 49.565 75.505 ;
        RECT 49.830 75.395 50.100 75.495 ;
        RECT 50.290 75.395 50.580 75.495 ;
        RECT 49.005 75.165 49.175 75.335 ;
        RECT 49.825 75.225 50.100 75.395 ;
        RECT 50.285 75.225 50.580 75.395 ;
        RECT 48.870 74.835 49.175 75.165 ;
        RECT 49.370 75.055 49.620 75.165 ;
        RECT 49.365 74.885 49.620 75.055 ;
        RECT 49.370 74.835 49.620 74.885 ;
        RECT 49.830 74.835 50.100 75.225 ;
        RECT 50.290 74.835 50.580 75.225 ;
        RECT 50.750 74.835 51.170 75.500 ;
        RECT 51.555 75.355 51.885 76.075 ;
        RECT 52.065 75.275 52.375 76.075 ;
        RECT 52.580 75.275 53.275 75.905 ;
        RECT 53.650 75.295 54.150 75.905 ;
        RECT 51.480 74.835 51.830 75.165 ;
        RECT 52.075 74.835 52.410 75.105 ;
        RECT 49.005 74.665 49.175 74.835 ;
        RECT 51.625 74.715 51.830 74.835 ;
        RECT 49.005 74.495 51.375 74.665 ;
        RECT 51.625 74.545 51.835 74.715 ;
        RECT 52.580 74.675 52.750 75.275 ;
        RECT 52.920 74.835 53.255 75.085 ;
        RECT 53.445 74.835 53.795 75.085 ;
        RECT 48.390 73.735 48.725 74.245 ;
        RECT 48.975 73.525 49.305 74.325 ;
        RECT 49.550 74.115 50.975 74.285 ;
        RECT 49.550 73.695 49.835 74.115 ;
        RECT 50.090 73.525 50.420 73.945 ;
        RECT 50.645 73.865 50.975 74.115 ;
        RECT 51.205 74.035 51.375 74.495 ;
        RECT 51.635 73.865 51.805 74.365 ;
        RECT 50.645 73.695 51.805 73.865 ;
        RECT 52.065 73.525 52.345 74.665 ;
        RECT 52.515 73.695 52.845 74.675 ;
        RECT 53.980 74.665 54.150 75.295 ;
        RECT 54.780 75.425 55.110 75.905 ;
        RECT 55.280 75.615 55.505 76.075 ;
        RECT 55.675 75.425 56.005 75.905 ;
        RECT 54.780 75.255 56.005 75.425 ;
        RECT 56.195 75.275 56.445 76.075 ;
        RECT 56.615 75.275 56.955 75.905 ;
        RECT 57.125 75.350 57.415 76.075 ;
        RECT 57.590 75.310 58.045 76.075 ;
        RECT 58.320 75.695 59.620 75.905 ;
        RECT 59.875 75.715 60.205 76.075 ;
        RECT 59.450 75.545 59.620 75.695 ;
        RECT 60.375 75.575 60.635 75.905 ;
        RECT 60.405 75.565 60.635 75.575 ;
        RECT 54.320 74.885 54.650 75.085 ;
        RECT 54.820 74.885 55.150 75.085 ;
        RECT 55.320 74.885 55.740 75.085 ;
        RECT 55.915 74.915 56.610 75.085 ;
        RECT 55.915 74.665 56.085 74.915 ;
        RECT 56.780 74.665 56.955 75.275 ;
        RECT 58.520 75.085 58.740 75.485 ;
        RECT 57.585 74.885 58.075 75.085 ;
        RECT 58.265 74.875 58.740 75.085 ;
        RECT 58.985 75.085 59.195 75.485 ;
        RECT 59.450 75.420 60.205 75.545 ;
        RECT 59.450 75.375 60.295 75.420 ;
        RECT 60.025 75.255 60.295 75.375 ;
        RECT 58.985 74.875 59.315 75.085 ;
        RECT 59.485 74.815 59.895 75.120 ;
        RECT 53.015 73.525 53.275 74.665 ;
        RECT 53.650 74.495 56.085 74.665 ;
        RECT 53.650 73.695 53.980 74.495 ;
        RECT 54.150 73.525 54.480 74.325 ;
        RECT 54.780 73.695 55.110 74.495 ;
        RECT 55.755 73.525 56.005 74.325 ;
        RECT 56.275 73.525 56.445 74.665 ;
        RECT 56.615 73.695 56.955 74.665 ;
        RECT 57.125 73.525 57.415 74.690 ;
        RECT 57.590 74.645 58.765 74.705 ;
        RECT 60.125 74.680 60.295 75.255 ;
        RECT 60.095 74.645 60.295 74.680 ;
        RECT 57.590 74.535 60.295 74.645 ;
        RECT 57.590 73.915 57.845 74.535 ;
        RECT 58.435 74.475 60.235 74.535 ;
        RECT 58.435 74.445 58.765 74.475 ;
        RECT 60.465 74.375 60.635 75.565 ;
        RECT 58.095 74.275 58.280 74.365 ;
        RECT 58.870 74.275 59.705 74.285 ;
        RECT 58.095 74.075 59.705 74.275 ;
        RECT 58.095 74.035 58.325 74.075 ;
        RECT 57.590 73.695 57.925 73.915 ;
        RECT 58.930 73.525 59.285 73.905 ;
        RECT 59.455 73.695 59.705 74.075 ;
        RECT 59.955 73.525 60.205 74.305 ;
        RECT 60.375 73.695 60.635 74.375 ;
        RECT 60.810 75.335 61.065 75.905 ;
        RECT 61.235 75.675 61.565 76.075 ;
        RECT 61.990 75.540 62.520 75.905 ;
        RECT 61.990 75.505 62.165 75.540 ;
        RECT 61.235 75.335 62.165 75.505 ;
        RECT 60.810 74.665 60.980 75.335 ;
        RECT 61.235 75.165 61.405 75.335 ;
        RECT 61.150 74.835 61.405 75.165 ;
        RECT 61.630 74.835 61.825 75.165 ;
        RECT 60.810 73.695 61.145 74.665 ;
        RECT 61.315 73.525 61.485 74.665 ;
        RECT 61.655 73.865 61.825 74.835 ;
        RECT 61.995 74.205 62.165 75.335 ;
        RECT 62.335 74.545 62.505 75.345 ;
        RECT 62.710 75.055 62.985 75.905 ;
        RECT 62.705 74.885 62.985 75.055 ;
        RECT 62.710 74.745 62.985 74.885 ;
        RECT 63.155 74.545 63.345 75.905 ;
        RECT 63.525 75.540 64.035 76.075 ;
        RECT 64.255 75.265 64.500 75.870 ;
        RECT 64.945 75.335 65.330 75.905 ;
        RECT 65.500 75.615 65.825 76.075 ;
        RECT 66.345 75.445 66.625 75.905 ;
        RECT 63.545 75.095 64.775 75.265 ;
        RECT 62.335 74.375 63.345 74.545 ;
        RECT 63.515 74.530 64.265 74.720 ;
        RECT 61.995 74.035 63.120 74.205 ;
        RECT 63.515 73.865 63.685 74.530 ;
        RECT 64.435 74.285 64.775 75.095 ;
        RECT 61.655 73.695 63.685 73.865 ;
        RECT 63.855 73.525 64.025 74.285 ;
        RECT 64.260 73.875 64.775 74.285 ;
        RECT 64.945 74.665 65.225 75.335 ;
        RECT 65.500 75.275 66.625 75.445 ;
        RECT 65.500 75.165 65.950 75.275 ;
        RECT 65.395 74.835 65.950 75.165 ;
        RECT 66.815 75.105 67.215 75.905 ;
        RECT 67.615 75.615 67.885 76.075 ;
        RECT 68.055 75.445 68.340 75.905 ;
        RECT 64.945 73.695 65.330 74.665 ;
        RECT 65.500 74.375 65.950 74.835 ;
        RECT 66.120 74.545 67.215 75.105 ;
        RECT 65.500 74.155 66.625 74.375 ;
        RECT 65.500 73.525 65.825 73.985 ;
        RECT 66.345 73.695 66.625 74.155 ;
        RECT 66.815 73.695 67.215 74.545 ;
        RECT 67.385 75.275 68.340 75.445 ;
        RECT 69.285 75.445 69.615 75.805 ;
        RECT 70.245 75.615 70.495 76.075 ;
        RECT 70.665 75.615 71.215 75.905 ;
        RECT 67.385 74.375 67.595 75.275 ;
        RECT 69.285 75.255 70.675 75.445 ;
        RECT 70.505 75.165 70.675 75.255 ;
        RECT 67.765 74.545 68.455 75.105 ;
        RECT 69.085 74.835 69.775 75.085 ;
        RECT 70.005 74.835 70.335 75.085 ;
        RECT 70.505 74.835 70.795 75.165 ;
        RECT 69.085 74.395 69.400 74.835 ;
        RECT 70.505 74.585 70.675 74.835 ;
        RECT 69.735 74.415 70.675 74.585 ;
        RECT 67.385 74.155 68.340 74.375 ;
        RECT 67.615 73.525 67.885 73.985 ;
        RECT 68.055 73.695 68.340 74.155 ;
        RECT 69.285 73.525 69.565 74.195 ;
        RECT 69.735 73.865 70.035 74.415 ;
        RECT 70.965 74.245 71.215 75.615 ;
        RECT 71.385 75.275 71.675 76.075 ;
        RECT 71.845 75.275 72.185 75.905 ;
        RECT 72.355 75.275 72.605 76.075 ;
        RECT 72.795 75.425 73.125 75.905 ;
        RECT 73.295 75.615 73.520 76.075 ;
        RECT 73.690 75.425 74.020 75.905 ;
        RECT 71.845 74.665 72.020 75.275 ;
        RECT 72.795 75.255 74.020 75.425 ;
        RECT 74.650 75.295 75.150 75.905 ;
        RECT 72.190 74.915 72.885 75.085 ;
        RECT 72.715 74.665 72.885 74.915 ;
        RECT 73.060 74.885 73.480 75.085 ;
        RECT 73.650 74.885 73.980 75.085 ;
        RECT 74.150 74.885 74.480 75.085 ;
        RECT 74.650 74.665 74.820 75.295 ;
        RECT 75.525 75.275 75.865 75.905 ;
        RECT 76.035 75.275 76.285 76.075 ;
        RECT 76.475 75.425 76.805 75.905 ;
        RECT 76.975 75.615 77.200 76.075 ;
        RECT 77.370 75.425 77.700 75.905 ;
        RECT 75.005 74.835 75.355 75.085 ;
        RECT 75.525 74.665 75.700 75.275 ;
        RECT 76.475 75.255 77.700 75.425 ;
        RECT 78.330 75.295 78.830 75.905 ;
        RECT 79.240 75.335 79.855 75.905 ;
        RECT 80.025 75.565 80.240 76.075 ;
        RECT 80.470 75.565 80.750 75.895 ;
        RECT 80.930 75.565 81.170 76.075 ;
        RECT 75.870 74.915 76.565 75.085 ;
        RECT 76.395 74.665 76.565 74.915 ;
        RECT 76.740 74.885 77.160 75.085 ;
        RECT 77.330 74.885 77.660 75.085 ;
        RECT 77.830 74.885 78.160 75.085 ;
        RECT 78.330 74.665 78.500 75.295 ;
        RECT 78.685 74.835 79.035 75.085 ;
        RECT 70.245 73.525 70.575 74.245 ;
        RECT 70.765 73.695 71.215 74.245 ;
        RECT 71.385 73.525 71.675 74.665 ;
        RECT 71.845 73.695 72.185 74.665 ;
        RECT 72.355 73.525 72.525 74.665 ;
        RECT 72.715 74.495 75.150 74.665 ;
        RECT 72.795 73.525 73.045 74.325 ;
        RECT 73.690 73.695 74.020 74.495 ;
        RECT 74.320 73.525 74.650 74.325 ;
        RECT 74.820 73.695 75.150 74.495 ;
        RECT 75.525 73.695 75.865 74.665 ;
        RECT 76.035 73.525 76.205 74.665 ;
        RECT 76.395 74.495 78.830 74.665 ;
        RECT 76.475 73.525 76.725 74.325 ;
        RECT 77.370 73.695 77.700 74.495 ;
        RECT 78.000 73.525 78.330 74.325 ;
        RECT 78.500 73.695 78.830 74.495 ;
        RECT 79.240 74.315 79.555 75.335 ;
        RECT 79.725 74.665 79.895 75.165 ;
        RECT 80.145 74.835 80.410 75.395 ;
        RECT 80.580 74.665 80.750 75.565 ;
        RECT 80.920 74.835 81.275 75.395 ;
        RECT 81.965 75.325 83.175 76.075 ;
        RECT 79.725 74.495 81.150 74.665 ;
        RECT 79.240 73.695 79.775 74.315 ;
        RECT 79.945 73.525 80.275 74.325 ;
        RECT 80.760 74.320 81.150 74.495 ;
        RECT 81.965 74.615 82.485 75.155 ;
        RECT 82.655 74.785 83.175 75.325 ;
        RECT 81.965 73.525 83.175 74.615 ;
        RECT 5.520 73.355 83.260 73.525 ;
        RECT 5.605 72.265 6.815 73.355 ;
        RECT 6.985 72.920 12.330 73.355 ;
        RECT 5.605 71.555 6.125 72.095 ;
        RECT 6.295 71.725 6.815 72.265 ;
        RECT 5.605 70.805 6.815 71.555 ;
        RECT 8.570 71.350 8.910 72.180 ;
        RECT 10.390 71.670 10.740 72.920 ;
        RECT 12.505 72.265 16.015 73.355 ;
        RECT 12.505 71.575 14.155 72.095 ;
        RECT 14.325 71.745 16.015 72.265 ;
        RECT 16.685 72.215 16.915 73.355 ;
        RECT 17.085 72.205 17.415 73.185 ;
        RECT 17.585 72.215 17.795 73.355 ;
        RECT 16.665 71.795 16.995 72.045 ;
        RECT 6.985 70.805 12.330 71.350 ;
        RECT 12.505 70.805 16.015 71.575 ;
        RECT 16.685 70.805 16.915 71.625 ;
        RECT 17.165 71.605 17.415 72.205 ;
        RECT 18.485 72.190 18.775 73.355 ;
        RECT 18.945 72.265 20.615 73.355 ;
        RECT 21.250 72.555 21.565 73.355 ;
        RECT 21.830 73.000 22.910 73.170 ;
        RECT 21.830 72.385 22.000 73.000 ;
        RECT 17.085 70.975 17.415 71.605 ;
        RECT 17.585 70.805 17.795 71.625 ;
        RECT 18.945 71.575 19.695 72.095 ;
        RECT 19.865 71.745 20.615 72.265 ;
        RECT 18.485 70.805 18.775 71.530 ;
        RECT 18.945 70.805 20.615 71.575 ;
        RECT 21.245 71.375 21.515 72.385 ;
        RECT 21.685 72.215 22.000 72.385 ;
        RECT 21.685 71.545 21.855 72.215 ;
        RECT 22.170 72.045 22.405 72.725 ;
        RECT 22.575 72.215 22.910 73.000 ;
        RECT 23.130 72.215 23.425 73.355 ;
        RECT 23.685 72.385 24.015 73.185 ;
        RECT 24.185 72.555 24.355 73.355 ;
        RECT 24.525 72.385 24.855 73.185 ;
        RECT 25.025 72.555 25.195 73.355 ;
        RECT 25.365 72.405 25.695 73.185 ;
        RECT 25.865 72.895 26.035 73.355 ;
        RECT 25.365 72.385 26.135 72.405 ;
        RECT 23.685 72.215 26.135 72.385 ;
        RECT 22.025 71.715 22.405 72.045 ;
        RECT 22.575 71.715 22.910 72.045 ;
        RECT 23.105 71.795 25.615 72.045 ;
        RECT 25.785 71.625 26.135 72.215 ;
        RECT 21.685 71.375 22.910 71.545 ;
        RECT 21.315 70.805 21.645 71.205 ;
        RECT 21.815 71.105 21.985 71.375 ;
        RECT 22.155 70.805 22.485 71.205 ;
        RECT 22.655 71.105 22.910 71.375 ;
        RECT 23.765 71.445 26.135 71.625 ;
        RECT 26.305 71.750 26.585 73.185 ;
        RECT 26.755 72.580 27.465 73.355 ;
        RECT 27.635 72.410 27.965 73.185 ;
        RECT 26.815 72.195 27.965 72.410 ;
        RECT 23.130 70.805 23.395 71.265 ;
        RECT 23.765 70.975 23.935 71.445 ;
        RECT 24.185 70.805 24.355 71.265 ;
        RECT 24.605 70.975 24.775 71.445 ;
        RECT 25.025 70.805 25.195 71.265 ;
        RECT 25.445 70.975 25.615 71.445 ;
        RECT 25.785 70.805 26.035 71.270 ;
        RECT 26.305 70.975 26.645 71.750 ;
        RECT 26.815 71.625 27.100 72.195 ;
        RECT 27.285 71.795 27.755 72.025 ;
        RECT 28.160 71.995 28.375 73.110 ;
        RECT 28.555 72.635 28.885 73.355 ;
        RECT 28.665 71.995 28.895 72.335 ;
        RECT 27.925 71.815 28.375 71.995 ;
        RECT 27.925 71.795 28.255 71.815 ;
        RECT 28.565 71.795 28.895 71.995 ;
        RECT 29.065 71.750 29.345 73.185 ;
        RECT 29.515 72.580 30.225 73.355 ;
        RECT 30.395 72.410 30.725 73.185 ;
        RECT 29.575 72.195 30.725 72.410 ;
        RECT 26.815 71.435 27.525 71.625 ;
        RECT 27.225 71.295 27.525 71.435 ;
        RECT 27.715 71.435 28.895 71.625 ;
        RECT 27.715 71.355 28.045 71.435 ;
        RECT 27.225 71.285 27.540 71.295 ;
        RECT 27.225 71.275 27.550 71.285 ;
        RECT 27.225 71.270 27.560 71.275 ;
        RECT 26.815 70.805 26.985 71.265 ;
        RECT 27.225 71.260 27.565 71.270 ;
        RECT 27.225 71.255 27.570 71.260 ;
        RECT 27.225 71.245 27.575 71.255 ;
        RECT 27.225 71.240 27.580 71.245 ;
        RECT 27.225 70.975 27.585 71.240 ;
        RECT 28.215 70.805 28.385 71.265 ;
        RECT 28.555 70.975 28.895 71.435 ;
        RECT 29.065 70.975 29.405 71.750 ;
        RECT 29.575 71.625 29.860 72.195 ;
        RECT 30.045 71.795 30.515 72.025 ;
        RECT 30.920 71.995 31.135 73.110 ;
        RECT 31.315 72.635 31.645 73.355 ;
        RECT 32.305 72.465 32.565 73.175 ;
        RECT 32.735 72.645 33.065 73.355 ;
        RECT 33.235 72.465 33.465 73.175 ;
        RECT 31.425 71.995 31.655 72.335 ;
        RECT 32.305 72.225 33.465 72.465 ;
        RECT 33.645 72.445 33.915 73.175 ;
        RECT 34.095 72.625 34.435 73.355 ;
        RECT 33.645 72.225 34.415 72.445 ;
        RECT 30.685 71.815 31.135 71.995 ;
        RECT 30.685 71.795 31.015 71.815 ;
        RECT 31.325 71.795 31.655 71.995 ;
        RECT 32.295 71.715 32.595 72.045 ;
        RECT 32.775 71.735 33.300 72.045 ;
        RECT 33.480 71.735 33.945 72.045 ;
        RECT 29.575 71.435 30.285 71.625 ;
        RECT 29.985 71.295 30.285 71.435 ;
        RECT 30.475 71.435 31.655 71.625 ;
        RECT 30.475 71.355 30.805 71.435 ;
        RECT 29.985 71.285 30.300 71.295 ;
        RECT 29.985 71.275 30.310 71.285 ;
        RECT 29.985 71.270 30.320 71.275 ;
        RECT 29.575 70.805 29.745 71.265 ;
        RECT 29.985 71.260 30.325 71.270 ;
        RECT 29.985 71.255 30.330 71.260 ;
        RECT 29.985 71.245 30.335 71.255 ;
        RECT 29.985 71.240 30.340 71.245 ;
        RECT 29.985 70.975 30.345 71.240 ;
        RECT 30.975 70.805 31.145 71.265 ;
        RECT 31.315 70.975 31.655 71.435 ;
        RECT 32.305 70.805 32.595 71.535 ;
        RECT 32.775 71.095 33.005 71.735 ;
        RECT 34.125 71.555 34.415 72.225 ;
        RECT 33.185 71.355 34.415 71.555 ;
        RECT 33.185 70.985 33.495 71.355 ;
        RECT 33.675 70.805 34.345 71.175 ;
        RECT 34.605 70.985 34.865 73.175 ;
        RECT 35.045 72.265 36.715 73.355 ;
        RECT 36.885 72.520 37.230 73.355 ;
        RECT 37.405 72.350 37.660 73.155 ;
        RECT 37.830 72.520 38.090 73.355 ;
        RECT 38.265 72.350 38.520 73.155 ;
        RECT 38.690 72.520 38.950 73.355 ;
        RECT 39.120 72.350 39.380 73.155 ;
        RECT 39.550 72.520 39.935 73.355 ;
        RECT 40.110 72.785 40.430 73.185 ;
        RECT 35.045 71.575 35.795 72.095 ;
        RECT 35.965 71.745 36.715 72.265 ;
        RECT 36.905 72.180 39.935 72.350 ;
        RECT 36.905 71.615 37.075 72.180 ;
        RECT 37.245 71.785 39.460 72.010 ;
        RECT 39.635 71.615 39.935 72.180 ;
        RECT 35.045 70.805 36.715 71.575 ;
        RECT 36.905 71.445 39.935 71.615 ;
        RECT 40.110 72.335 40.280 72.785 ;
        RECT 40.600 72.555 40.910 73.355 ;
        RECT 41.080 72.725 41.410 73.185 ;
        RECT 41.580 72.895 41.750 73.355 ;
        RECT 41.920 72.725 42.250 73.185 ;
        RECT 42.420 72.895 42.670 73.355 ;
        RECT 42.860 72.895 43.110 73.355 ;
        RECT 41.080 72.675 42.250 72.725 ;
        RECT 43.280 72.725 43.530 73.185 ;
        RECT 43.780 72.895 44.070 73.355 ;
        RECT 43.280 72.675 44.070 72.725 ;
        RECT 41.080 72.505 44.070 72.675 ;
        RECT 40.110 72.165 43.670 72.335 ;
        RECT 37.365 70.805 37.660 71.275 ;
        RECT 37.830 71.000 38.090 71.445 ;
        RECT 38.260 70.805 38.520 71.275 ;
        RECT 38.690 71.000 38.945 71.445 ;
        RECT 40.110 71.375 40.280 72.165 ;
        RECT 40.450 71.795 40.800 71.995 ;
        RECT 41.080 71.795 41.760 71.995 ;
        RECT 41.970 71.795 43.160 71.995 ;
        RECT 43.340 71.795 43.670 72.165 ;
        RECT 43.870 71.625 44.070 72.505 ;
        RECT 44.245 72.190 44.535 73.355 ;
        RECT 44.710 72.215 45.045 73.185 ;
        RECT 45.215 72.215 45.385 73.355 ;
        RECT 45.555 73.015 47.585 73.185 ;
        RECT 39.115 70.805 39.415 71.275 ;
        RECT 40.110 70.975 40.430 71.375 ;
        RECT 40.600 70.805 40.910 71.625 ;
        RECT 41.080 71.435 42.770 71.625 ;
        RECT 41.080 70.975 41.410 71.435 ;
        RECT 42.020 71.355 42.770 71.435 ;
        RECT 41.580 70.805 41.830 71.265 ;
        RECT 42.940 71.185 43.110 71.625 ;
        RECT 43.280 71.355 44.070 71.625 ;
        RECT 44.710 71.545 44.880 72.215 ;
        RECT 45.555 72.045 45.725 73.015 ;
        RECT 45.050 71.715 45.305 72.045 ;
        RECT 45.530 71.715 45.725 72.045 ;
        RECT 45.895 72.675 47.020 72.845 ;
        RECT 45.135 71.545 45.305 71.715 ;
        RECT 45.895 71.545 46.065 72.675 ;
        RECT 42.020 70.975 44.070 71.185 ;
        RECT 44.245 70.805 44.535 71.530 ;
        RECT 44.710 70.975 44.965 71.545 ;
        RECT 45.135 71.375 46.065 71.545 ;
        RECT 46.235 72.335 47.245 72.505 ;
        RECT 46.235 71.535 46.405 72.335 ;
        RECT 46.610 71.995 46.885 72.135 ;
        RECT 46.605 71.825 46.885 71.995 ;
        RECT 45.890 71.340 46.065 71.375 ;
        RECT 45.135 70.805 45.465 71.205 ;
        RECT 45.890 70.975 46.420 71.340 ;
        RECT 46.610 70.975 46.885 71.825 ;
        RECT 47.055 70.975 47.245 72.335 ;
        RECT 47.415 72.350 47.585 73.015 ;
        RECT 47.755 72.595 47.925 73.355 ;
        RECT 48.160 72.595 48.675 73.005 ;
        RECT 47.415 72.160 48.165 72.350 ;
        RECT 48.335 71.785 48.675 72.595 ;
        RECT 48.845 72.265 50.055 73.355 ;
        RECT 50.225 72.845 50.485 73.355 ;
        RECT 47.445 71.615 48.675 71.785 ;
        RECT 47.425 70.805 47.935 71.340 ;
        RECT 48.155 71.010 48.400 71.615 ;
        RECT 48.845 71.555 49.365 72.095 ;
        RECT 49.535 71.725 50.055 72.265 ;
        RECT 50.225 71.795 50.565 72.675 ;
        RECT 50.735 71.965 50.905 73.185 ;
        RECT 51.145 72.850 51.760 73.355 ;
        RECT 51.145 72.315 51.395 72.680 ;
        RECT 51.565 72.675 51.760 72.850 ;
        RECT 51.930 72.845 52.405 73.185 ;
        RECT 52.575 72.810 52.790 73.355 ;
        RECT 51.565 72.485 51.895 72.675 ;
        RECT 52.115 72.315 52.830 72.610 ;
        RECT 53.000 72.485 53.275 73.185 ;
        RECT 53.445 72.845 54.635 73.135 ;
        RECT 51.145 72.145 52.935 72.315 ;
        RECT 50.735 71.715 51.530 71.965 ;
        RECT 50.735 71.625 50.985 71.715 ;
        RECT 48.845 70.805 50.055 71.555 ;
        RECT 50.225 70.805 50.485 71.625 ;
        RECT 50.655 71.205 50.985 71.625 ;
        RECT 51.700 71.290 51.955 72.145 ;
        RECT 51.165 71.025 51.955 71.290 ;
        RECT 52.125 71.445 52.535 71.965 ;
        RECT 52.705 71.715 52.935 72.145 ;
        RECT 53.105 71.455 53.275 72.485 ;
        RECT 53.465 72.505 54.635 72.675 ;
        RECT 54.805 72.555 55.085 73.355 ;
        RECT 53.465 72.215 53.790 72.505 ;
        RECT 54.465 72.385 54.635 72.505 ;
        RECT 53.960 72.045 54.155 72.335 ;
        RECT 54.465 72.215 55.125 72.385 ;
        RECT 55.295 72.215 55.570 73.185 ;
        RECT 54.955 72.045 55.125 72.215 ;
        RECT 53.445 71.715 53.790 72.045 ;
        RECT 53.960 71.715 54.785 72.045 ;
        RECT 54.955 71.715 55.230 72.045 ;
        RECT 54.955 71.545 55.125 71.715 ;
        RECT 52.125 71.025 52.325 71.445 ;
        RECT 52.515 70.805 52.845 71.265 ;
        RECT 53.015 70.975 53.275 71.455 ;
        RECT 53.460 71.375 55.125 71.545 ;
        RECT 55.400 71.480 55.570 72.215 ;
        RECT 55.750 72.965 56.085 73.185 ;
        RECT 57.090 72.975 57.445 73.355 ;
        RECT 55.750 72.345 56.005 72.965 ;
        RECT 56.255 72.805 56.485 72.845 ;
        RECT 57.615 72.805 57.865 73.185 ;
        RECT 56.255 72.605 57.865 72.805 ;
        RECT 56.255 72.515 56.440 72.605 ;
        RECT 57.030 72.595 57.865 72.605 ;
        RECT 58.115 72.575 58.365 73.355 ;
        RECT 58.535 72.505 58.795 73.185 ;
        RECT 59.055 72.685 59.225 73.185 ;
        RECT 59.395 72.855 59.725 73.355 ;
        RECT 59.055 72.515 59.720 72.685 ;
        RECT 56.595 72.405 56.925 72.435 ;
        RECT 56.595 72.345 58.395 72.405 ;
        RECT 55.750 72.235 58.455 72.345 ;
        RECT 55.750 72.175 56.925 72.235 ;
        RECT 58.255 72.200 58.455 72.235 ;
        RECT 55.745 71.795 56.235 71.995 ;
        RECT 56.425 71.795 56.900 72.005 ;
        RECT 53.460 71.025 53.715 71.375 ;
        RECT 53.885 70.805 54.215 71.205 ;
        RECT 54.385 71.025 54.555 71.375 ;
        RECT 54.725 70.805 55.105 71.205 ;
        RECT 55.295 71.135 55.570 71.480 ;
        RECT 55.750 70.805 56.205 71.570 ;
        RECT 56.680 71.395 56.900 71.795 ;
        RECT 57.145 71.795 57.475 72.005 ;
        RECT 57.145 71.395 57.355 71.795 ;
        RECT 57.645 71.760 58.055 72.065 ;
        RECT 58.285 71.625 58.455 72.200 ;
        RECT 58.185 71.505 58.455 71.625 ;
        RECT 57.610 71.460 58.455 71.505 ;
        RECT 57.610 71.335 58.365 71.460 ;
        RECT 57.610 71.185 57.780 71.335 ;
        RECT 58.625 71.315 58.795 72.505 ;
        RECT 58.970 71.695 59.320 72.345 ;
        RECT 59.490 71.525 59.720 72.515 ;
        RECT 58.565 71.305 58.795 71.315 ;
        RECT 56.480 70.975 57.780 71.185 ;
        RECT 58.035 70.805 58.365 71.165 ;
        RECT 58.535 70.975 58.795 71.305 ;
        RECT 59.055 71.355 59.720 71.525 ;
        RECT 59.055 71.065 59.225 71.355 ;
        RECT 59.395 70.805 59.725 71.185 ;
        RECT 59.895 71.065 60.080 73.185 ;
        RECT 60.320 72.895 60.585 73.355 ;
        RECT 60.755 72.760 61.005 73.185 ;
        RECT 61.215 72.910 62.320 73.080 ;
        RECT 60.700 72.630 61.005 72.760 ;
        RECT 60.250 71.435 60.530 72.385 ;
        RECT 60.700 71.525 60.870 72.630 ;
        RECT 61.040 71.845 61.280 72.440 ;
        RECT 61.450 72.375 61.980 72.740 ;
        RECT 61.450 71.675 61.620 72.375 ;
        RECT 62.150 72.295 62.320 72.910 ;
        RECT 62.490 72.555 62.660 73.355 ;
        RECT 62.830 72.855 63.080 73.185 ;
        RECT 63.305 72.885 64.190 73.055 ;
        RECT 62.150 72.205 62.660 72.295 ;
        RECT 60.700 71.395 60.925 71.525 ;
        RECT 61.095 71.455 61.620 71.675 ;
        RECT 61.790 72.035 62.660 72.205 ;
        RECT 60.335 70.805 60.585 71.265 ;
        RECT 60.755 71.255 60.925 71.395 ;
        RECT 61.790 71.255 61.960 72.035 ;
        RECT 62.490 71.965 62.660 72.035 ;
        RECT 62.170 71.785 62.370 71.815 ;
        RECT 62.830 71.785 63.000 72.855 ;
        RECT 63.170 71.965 63.360 72.685 ;
        RECT 62.170 71.485 63.000 71.785 ;
        RECT 63.530 71.755 63.850 72.715 ;
        RECT 60.755 71.085 61.090 71.255 ;
        RECT 61.285 71.085 61.960 71.255 ;
        RECT 62.280 70.805 62.650 71.305 ;
        RECT 62.830 71.255 63.000 71.485 ;
        RECT 63.385 71.425 63.850 71.755 ;
        RECT 64.020 72.045 64.190 72.885 ;
        RECT 64.370 72.855 64.685 73.355 ;
        RECT 64.915 72.625 65.255 73.185 ;
        RECT 64.360 72.250 65.255 72.625 ;
        RECT 65.425 72.345 65.595 73.355 ;
        RECT 65.065 72.045 65.255 72.250 ;
        RECT 65.765 72.295 66.095 73.140 ;
        RECT 66.510 72.385 66.900 72.560 ;
        RECT 67.385 72.555 67.715 73.355 ;
        RECT 67.885 72.565 68.420 73.185 ;
        RECT 65.765 72.215 66.155 72.295 ;
        RECT 66.510 72.215 67.935 72.385 ;
        RECT 65.940 72.165 66.155 72.215 ;
        RECT 64.020 71.715 64.895 72.045 ;
        RECT 65.065 71.715 65.815 72.045 ;
        RECT 64.020 71.255 64.190 71.715 ;
        RECT 65.065 71.545 65.265 71.715 ;
        RECT 65.985 71.585 66.155 72.165 ;
        RECT 65.930 71.545 66.155 71.585 ;
        RECT 62.830 71.085 63.235 71.255 ;
        RECT 63.405 71.085 64.190 71.255 ;
        RECT 64.465 70.805 64.675 71.335 ;
        RECT 64.935 71.020 65.265 71.545 ;
        RECT 65.775 71.460 66.155 71.545 ;
        RECT 66.385 71.485 66.740 72.045 ;
        RECT 65.435 70.805 65.605 71.415 ;
        RECT 65.775 71.025 66.105 71.460 ;
        RECT 66.910 71.315 67.080 72.215 ;
        RECT 67.250 71.485 67.515 72.045 ;
        RECT 67.765 71.715 67.935 72.215 ;
        RECT 68.105 71.545 68.420 72.565 ;
        RECT 68.665 72.215 68.895 73.355 ;
        RECT 69.065 72.205 69.395 73.185 ;
        RECT 69.565 72.215 69.775 73.355 ;
        RECT 68.645 71.795 68.975 72.045 ;
        RECT 66.490 70.805 66.730 71.315 ;
        RECT 66.910 70.985 67.190 71.315 ;
        RECT 67.420 70.805 67.635 71.315 ;
        RECT 67.805 70.975 68.420 71.545 ;
        RECT 68.665 70.805 68.895 71.625 ;
        RECT 69.145 71.605 69.395 72.205 ;
        RECT 70.005 72.190 70.295 73.355 ;
        RECT 70.470 73.015 71.550 73.170 ;
        RECT 70.470 73.000 71.615 73.015 ;
        RECT 70.470 72.215 70.805 73.000 ;
        RECT 71.380 72.845 71.615 73.000 ;
        RECT 70.975 72.045 71.210 72.725 ;
        RECT 71.380 72.385 71.550 72.845 ;
        RECT 71.815 72.555 72.130 73.355 ;
        RECT 72.395 72.685 72.565 73.185 ;
        RECT 72.735 72.855 73.065 73.355 ;
        RECT 72.395 72.515 73.060 72.685 ;
        RECT 71.380 72.215 71.695 72.385 ;
        RECT 70.470 71.715 70.805 72.045 ;
        RECT 70.975 71.715 71.355 72.045 ;
        RECT 69.065 70.975 69.395 71.605 ;
        RECT 69.565 70.805 69.775 71.625 ;
        RECT 71.525 71.545 71.695 72.215 ;
        RECT 70.005 70.805 70.295 71.530 ;
        RECT 70.470 71.375 71.695 71.545 ;
        RECT 71.865 71.375 72.135 72.385 ;
        RECT 72.310 71.695 72.660 72.345 ;
        RECT 72.830 71.525 73.060 72.515 ;
        RECT 70.470 71.105 70.725 71.375 ;
        RECT 70.895 70.805 71.225 71.205 ;
        RECT 71.395 71.105 71.565 71.375 ;
        RECT 72.395 71.355 73.060 71.525 ;
        RECT 71.735 70.805 72.065 71.205 ;
        RECT 72.395 71.065 72.565 71.355 ;
        RECT 72.735 70.805 73.065 71.185 ;
        RECT 73.235 71.065 73.420 73.185 ;
        RECT 73.660 72.895 73.925 73.355 ;
        RECT 74.095 72.760 74.345 73.185 ;
        RECT 74.555 72.910 75.660 73.080 ;
        RECT 74.040 72.630 74.345 72.760 ;
        RECT 73.590 71.435 73.870 72.385 ;
        RECT 74.040 71.525 74.210 72.630 ;
        RECT 74.380 71.845 74.620 72.440 ;
        RECT 74.790 72.375 75.320 72.740 ;
        RECT 74.790 71.675 74.960 72.375 ;
        RECT 75.490 72.295 75.660 72.910 ;
        RECT 75.830 72.555 76.000 73.355 ;
        RECT 76.170 72.855 76.420 73.185 ;
        RECT 76.645 72.885 77.530 73.055 ;
        RECT 75.490 72.205 76.000 72.295 ;
        RECT 74.040 71.395 74.265 71.525 ;
        RECT 74.435 71.455 74.960 71.675 ;
        RECT 75.130 72.035 76.000 72.205 ;
        RECT 73.675 70.805 73.925 71.265 ;
        RECT 74.095 71.255 74.265 71.395 ;
        RECT 75.130 71.255 75.300 72.035 ;
        RECT 75.830 71.965 76.000 72.035 ;
        RECT 75.510 71.785 75.710 71.815 ;
        RECT 76.170 71.785 76.340 72.855 ;
        RECT 76.510 71.965 76.700 72.685 ;
        RECT 75.510 71.485 76.340 71.785 ;
        RECT 76.870 71.755 77.190 72.715 ;
        RECT 74.095 71.085 74.430 71.255 ;
        RECT 74.625 71.085 75.300 71.255 ;
        RECT 75.620 70.805 75.990 71.305 ;
        RECT 76.170 71.255 76.340 71.485 ;
        RECT 76.725 71.425 77.190 71.755 ;
        RECT 77.360 72.045 77.530 72.885 ;
        RECT 77.710 72.855 78.025 73.355 ;
        RECT 78.255 72.625 78.595 73.185 ;
        RECT 77.700 72.250 78.595 72.625 ;
        RECT 78.765 72.345 78.935 73.355 ;
        RECT 78.405 72.045 78.595 72.250 ;
        RECT 79.105 72.295 79.435 73.140 ;
        RECT 79.850 72.385 80.240 72.560 ;
        RECT 80.725 72.555 81.055 73.355 ;
        RECT 81.225 72.565 81.760 73.185 ;
        RECT 79.105 72.215 79.495 72.295 ;
        RECT 79.850 72.215 81.275 72.385 ;
        RECT 79.280 72.165 79.495 72.215 ;
        RECT 77.360 71.715 78.235 72.045 ;
        RECT 78.405 71.715 79.155 72.045 ;
        RECT 77.360 71.255 77.530 71.715 ;
        RECT 78.405 71.545 78.605 71.715 ;
        RECT 79.325 71.585 79.495 72.165 ;
        RECT 79.270 71.545 79.495 71.585 ;
        RECT 76.170 71.085 76.575 71.255 ;
        RECT 76.745 71.085 77.530 71.255 ;
        RECT 77.805 70.805 78.015 71.335 ;
        RECT 78.275 71.020 78.605 71.545 ;
        RECT 79.115 71.460 79.495 71.545 ;
        RECT 79.725 71.485 80.080 72.045 ;
        RECT 78.775 70.805 78.945 71.415 ;
        RECT 79.115 71.025 79.445 71.460 ;
        RECT 80.250 71.315 80.420 72.215 ;
        RECT 80.590 71.485 80.855 72.045 ;
        RECT 81.105 71.715 81.275 72.215 ;
        RECT 81.445 71.545 81.760 72.565 ;
        RECT 81.965 72.265 83.175 73.355 ;
        RECT 81.965 71.725 82.485 72.265 ;
        RECT 82.655 71.555 83.175 72.095 ;
        RECT 79.830 70.805 80.070 71.315 ;
        RECT 80.250 70.985 80.530 71.315 ;
        RECT 80.760 70.805 80.975 71.315 ;
        RECT 81.145 70.975 81.760 71.545 ;
        RECT 81.965 70.805 83.175 71.555 ;
        RECT 5.520 70.635 83.260 70.805 ;
        RECT 5.605 69.885 6.815 70.635 ;
        RECT 5.605 69.345 6.125 69.885 ;
        RECT 6.985 69.865 8.655 70.635 ;
        RECT 6.295 69.175 6.815 69.715 ;
        RECT 6.985 69.345 7.735 69.865 ;
        RECT 9.285 69.835 9.980 70.465 ;
        RECT 10.185 69.835 10.495 70.635 ;
        RECT 10.665 70.090 16.010 70.635 ;
        RECT 7.905 69.175 8.655 69.695 ;
        RECT 9.305 69.395 9.640 69.645 ;
        RECT 9.810 69.235 9.980 69.835 ;
        RECT 10.150 69.395 10.485 69.665 ;
        RECT 12.250 69.260 12.590 70.090 ;
        RECT 17.105 69.835 17.415 70.635 ;
        RECT 17.620 69.835 18.315 70.465 ;
        RECT 18.485 70.255 19.375 70.425 ;
        RECT 5.605 68.085 6.815 69.175 ;
        RECT 6.985 68.085 8.655 69.175 ;
        RECT 9.285 68.085 9.545 69.225 ;
        RECT 9.715 68.255 10.045 69.235 ;
        RECT 10.215 68.085 10.495 69.225 ;
        RECT 14.070 68.520 14.420 69.770 ;
        RECT 17.115 69.395 17.450 69.665 ;
        RECT 17.620 69.235 17.790 69.835 ;
        RECT 18.485 69.700 19.035 70.085 ;
        RECT 17.960 69.395 18.295 69.645 ;
        RECT 19.205 69.530 19.375 70.255 ;
        RECT 18.485 69.460 19.375 69.530 ;
        RECT 19.545 69.930 19.765 70.415 ;
        RECT 19.935 70.095 20.185 70.635 ;
        RECT 20.355 69.985 20.615 70.465 ;
        RECT 19.545 69.505 19.875 69.930 ;
        RECT 18.485 69.435 19.380 69.460 ;
        RECT 18.485 69.420 19.390 69.435 ;
        RECT 18.485 69.405 19.395 69.420 ;
        RECT 18.485 69.400 19.405 69.405 ;
        RECT 18.485 69.390 19.410 69.400 ;
        RECT 18.485 69.380 19.415 69.390 ;
        RECT 18.485 69.375 19.425 69.380 ;
        RECT 18.485 69.365 19.435 69.375 ;
        RECT 18.485 69.360 19.445 69.365 ;
        RECT 10.665 68.085 16.010 68.520 ;
        RECT 17.105 68.085 17.385 69.225 ;
        RECT 17.555 68.255 17.885 69.235 ;
        RECT 18.055 68.085 18.315 69.225 ;
        RECT 18.485 68.910 18.745 69.360 ;
        RECT 19.110 69.355 19.445 69.360 ;
        RECT 19.110 69.350 19.460 69.355 ;
        RECT 19.110 69.340 19.475 69.350 ;
        RECT 19.110 69.335 19.500 69.340 ;
        RECT 20.045 69.335 20.275 69.730 ;
        RECT 19.110 69.330 20.275 69.335 ;
        RECT 19.140 69.295 20.275 69.330 ;
        RECT 19.175 69.270 20.275 69.295 ;
        RECT 19.205 69.240 20.275 69.270 ;
        RECT 19.225 69.210 20.275 69.240 ;
        RECT 19.245 69.180 20.275 69.210 ;
        RECT 19.315 69.170 20.275 69.180 ;
        RECT 19.340 69.160 20.275 69.170 ;
        RECT 19.360 69.145 20.275 69.160 ;
        RECT 19.380 69.130 20.275 69.145 ;
        RECT 19.385 69.120 20.170 69.130 ;
        RECT 19.400 69.085 20.170 69.120 ;
        RECT 18.915 68.765 19.245 69.010 ;
        RECT 19.415 68.835 20.170 69.085 ;
        RECT 20.445 68.955 20.615 69.985 ;
        RECT 20.985 70.005 21.315 70.365 ;
        RECT 21.935 70.175 22.185 70.635 ;
        RECT 22.355 70.175 22.915 70.465 ;
        RECT 20.985 69.815 22.375 70.005 ;
        RECT 22.205 69.725 22.375 69.815 ;
        RECT 20.800 69.395 21.475 69.645 ;
        RECT 21.695 69.395 22.035 69.645 ;
        RECT 22.205 69.395 22.495 69.725 ;
        RECT 20.800 69.035 21.065 69.395 ;
        RECT 22.205 69.145 22.375 69.395 ;
        RECT 18.915 68.740 19.100 68.765 ;
        RECT 18.485 68.640 19.100 68.740 ;
        RECT 18.485 68.085 19.090 68.640 ;
        RECT 19.265 68.255 19.745 68.595 ;
        RECT 19.915 68.085 20.170 68.630 ;
        RECT 20.340 68.255 20.615 68.955 ;
        RECT 21.435 68.975 22.375 69.145 ;
        RECT 20.985 68.085 21.265 68.755 ;
        RECT 21.435 68.425 21.735 68.975 ;
        RECT 22.665 68.805 22.915 70.175 ;
        RECT 23.135 69.980 23.465 70.415 ;
        RECT 23.635 70.025 23.805 70.635 ;
        RECT 23.085 69.895 23.465 69.980 ;
        RECT 23.975 69.895 24.305 70.420 ;
        RECT 24.565 70.105 24.775 70.635 ;
        RECT 25.050 70.185 25.835 70.355 ;
        RECT 26.005 70.185 26.410 70.355 ;
        RECT 23.085 69.855 23.310 69.895 ;
        RECT 23.085 69.275 23.255 69.855 ;
        RECT 23.975 69.725 24.175 69.895 ;
        RECT 25.050 69.725 25.220 70.185 ;
        RECT 23.425 69.395 24.175 69.725 ;
        RECT 24.345 69.395 25.220 69.725 ;
        RECT 23.085 69.225 23.300 69.275 ;
        RECT 23.085 69.145 23.475 69.225 ;
        RECT 21.935 68.085 22.265 68.805 ;
        RECT 22.455 68.255 22.915 68.805 ;
        RECT 23.145 68.300 23.475 69.145 ;
        RECT 23.985 69.190 24.175 69.395 ;
        RECT 23.645 68.085 23.815 69.095 ;
        RECT 23.985 68.815 24.880 69.190 ;
        RECT 23.985 68.255 24.325 68.815 ;
        RECT 24.555 68.085 24.870 68.585 ;
        RECT 25.050 68.555 25.220 69.395 ;
        RECT 25.390 69.685 25.855 70.015 ;
        RECT 26.240 69.955 26.410 70.185 ;
        RECT 26.590 70.135 26.960 70.635 ;
        RECT 27.280 70.185 27.955 70.355 ;
        RECT 28.150 70.185 28.485 70.355 ;
        RECT 25.390 68.725 25.710 69.685 ;
        RECT 26.240 69.655 27.070 69.955 ;
        RECT 25.880 68.755 26.070 69.475 ;
        RECT 26.240 68.585 26.410 69.655 ;
        RECT 26.870 69.625 27.070 69.655 ;
        RECT 26.580 69.405 26.750 69.475 ;
        RECT 27.280 69.405 27.450 70.185 ;
        RECT 28.315 70.045 28.485 70.185 ;
        RECT 28.655 70.175 28.905 70.635 ;
        RECT 26.580 69.235 27.450 69.405 ;
        RECT 27.620 69.765 28.145 69.985 ;
        RECT 28.315 69.915 28.540 70.045 ;
        RECT 26.580 69.145 27.090 69.235 ;
        RECT 25.050 68.385 25.935 68.555 ;
        RECT 26.160 68.255 26.410 68.585 ;
        RECT 26.580 68.085 26.750 68.885 ;
        RECT 26.920 68.530 27.090 69.145 ;
        RECT 27.620 69.065 27.790 69.765 ;
        RECT 27.260 68.700 27.790 69.065 ;
        RECT 27.960 69.000 28.200 69.595 ;
        RECT 28.370 68.810 28.540 69.915 ;
        RECT 28.710 69.055 28.990 70.005 ;
        RECT 28.235 68.680 28.540 68.810 ;
        RECT 26.920 68.360 28.025 68.530 ;
        RECT 28.235 68.255 28.485 68.680 ;
        RECT 28.655 68.085 28.920 68.545 ;
        RECT 29.160 68.255 29.345 70.375 ;
        RECT 29.515 70.255 29.845 70.635 ;
        RECT 30.015 70.085 30.185 70.375 ;
        RECT 29.520 69.915 30.185 70.085 ;
        RECT 29.520 68.925 29.750 69.915 ;
        RECT 31.365 69.910 31.655 70.635 ;
        RECT 32.000 69.985 32.330 70.465 ;
        RECT 32.500 70.155 32.750 70.635 ;
        RECT 32.920 69.985 33.250 70.465 ;
        RECT 33.420 70.155 33.670 70.635 ;
        RECT 33.840 70.155 34.170 70.465 ;
        RECT 33.840 69.985 34.010 70.155 ;
        RECT 34.535 69.985 34.875 70.465 ;
        RECT 35.105 70.175 35.350 70.635 ;
        RECT 32.000 69.815 34.010 69.985 ;
        RECT 34.180 69.815 34.875 69.985 ;
        RECT 29.920 69.095 30.270 69.745 ;
        RECT 31.880 69.395 32.460 69.645 ;
        RECT 32.630 69.305 32.960 69.645 ;
        RECT 33.130 69.475 33.460 69.645 ;
        RECT 29.520 68.755 30.185 68.925 ;
        RECT 29.515 68.085 29.845 68.585 ;
        RECT 30.015 68.255 30.185 68.755 ;
        RECT 31.365 68.085 31.655 69.250 ;
        RECT 32.000 68.085 32.330 69.225 ;
        RECT 32.630 68.595 32.970 69.305 ;
        RECT 32.575 68.425 32.970 68.595 ;
        RECT 32.630 68.365 32.970 68.425 ;
        RECT 33.140 68.365 33.460 69.475 ;
        RECT 33.640 69.475 33.970 69.645 ;
        RECT 33.640 68.365 33.945 69.475 ;
        RECT 34.180 69.235 34.350 69.815 ;
        RECT 34.520 69.445 34.855 69.645 ;
        RECT 35.045 69.395 35.360 70.005 ;
        RECT 35.530 69.645 35.780 70.455 ;
        RECT 35.950 70.110 36.210 70.635 ;
        RECT 36.380 69.985 36.640 70.440 ;
        RECT 36.810 70.155 37.070 70.635 ;
        RECT 37.240 69.985 37.500 70.440 ;
        RECT 37.670 70.155 37.930 70.635 ;
        RECT 38.100 69.985 38.360 70.440 ;
        RECT 38.530 70.155 38.790 70.635 ;
        RECT 38.960 69.985 39.220 70.440 ;
        RECT 39.390 70.155 39.690 70.635 ;
        RECT 40.195 70.085 40.365 70.375 ;
        RECT 40.535 70.255 40.865 70.635 ;
        RECT 36.380 69.815 39.690 69.985 ;
        RECT 40.195 69.915 40.860 70.085 ;
        RECT 35.530 69.395 38.550 69.645 ;
        RECT 34.115 68.255 34.445 69.235 ;
        RECT 34.615 68.085 34.875 69.275 ;
        RECT 35.055 68.085 35.350 69.195 ;
        RECT 35.530 68.260 35.780 69.395 ;
        RECT 38.720 69.225 39.690 69.815 ;
        RECT 35.950 68.085 36.210 69.195 ;
        RECT 36.380 68.985 39.690 69.225 ;
        RECT 40.110 69.095 40.460 69.745 ;
        RECT 36.380 68.260 36.640 68.985 ;
        RECT 36.810 68.085 37.070 68.815 ;
        RECT 37.240 68.260 37.500 68.985 ;
        RECT 37.670 68.085 37.930 68.815 ;
        RECT 38.100 68.260 38.360 68.985 ;
        RECT 38.530 68.085 38.790 68.815 ;
        RECT 38.960 68.260 39.220 68.985 ;
        RECT 40.630 68.925 40.860 69.915 ;
        RECT 39.390 68.085 39.685 68.815 ;
        RECT 40.195 68.755 40.860 68.925 ;
        RECT 40.195 68.255 40.365 68.755 ;
        RECT 40.535 68.085 40.865 68.585 ;
        RECT 41.035 68.255 41.220 70.375 ;
        RECT 41.475 70.175 41.725 70.635 ;
        RECT 41.895 70.185 42.230 70.355 ;
        RECT 42.425 70.185 43.100 70.355 ;
        RECT 41.895 70.045 42.065 70.185 ;
        RECT 41.390 69.055 41.670 70.005 ;
        RECT 41.840 69.915 42.065 70.045 ;
        RECT 41.840 68.810 42.010 69.915 ;
        RECT 42.235 69.765 42.760 69.985 ;
        RECT 42.180 69.000 42.420 69.595 ;
        RECT 42.590 69.065 42.760 69.765 ;
        RECT 42.930 69.405 43.100 70.185 ;
        RECT 43.420 70.135 43.790 70.635 ;
        RECT 43.970 70.185 44.375 70.355 ;
        RECT 44.545 70.185 45.330 70.355 ;
        RECT 43.970 69.955 44.140 70.185 ;
        RECT 43.310 69.655 44.140 69.955 ;
        RECT 44.525 69.685 44.990 70.015 ;
        RECT 43.310 69.625 43.510 69.655 ;
        RECT 43.630 69.405 43.800 69.475 ;
        RECT 42.930 69.235 43.800 69.405 ;
        RECT 43.290 69.145 43.800 69.235 ;
        RECT 41.840 68.680 42.145 68.810 ;
        RECT 42.590 68.700 43.120 69.065 ;
        RECT 41.460 68.085 41.725 68.545 ;
        RECT 41.895 68.255 42.145 68.680 ;
        RECT 43.290 68.530 43.460 69.145 ;
        RECT 42.355 68.360 43.460 68.530 ;
        RECT 43.630 68.085 43.800 68.885 ;
        RECT 43.970 68.585 44.140 69.655 ;
        RECT 44.310 68.755 44.500 69.475 ;
        RECT 44.670 68.725 44.990 69.685 ;
        RECT 45.160 69.725 45.330 70.185 ;
        RECT 45.605 70.105 45.815 70.635 ;
        RECT 46.075 69.895 46.405 70.420 ;
        RECT 46.575 70.025 46.745 70.635 ;
        RECT 46.915 69.980 47.245 70.415 ;
        RECT 46.915 69.895 47.295 69.980 ;
        RECT 46.205 69.725 46.405 69.895 ;
        RECT 47.070 69.855 47.295 69.895 ;
        RECT 45.160 69.395 46.035 69.725 ;
        RECT 46.205 69.395 46.955 69.725 ;
        RECT 43.970 68.255 44.220 68.585 ;
        RECT 45.160 68.555 45.330 69.395 ;
        RECT 46.205 69.190 46.395 69.395 ;
        RECT 47.125 69.275 47.295 69.855 ;
        RECT 47.465 69.885 48.675 70.635 ;
        RECT 48.880 69.895 49.495 70.465 ;
        RECT 49.665 70.125 49.880 70.635 ;
        RECT 50.110 70.125 50.390 70.455 ;
        RECT 50.570 70.125 50.810 70.635 ;
        RECT 47.465 69.345 47.985 69.885 ;
        RECT 47.080 69.225 47.295 69.275 ;
        RECT 45.500 68.815 46.395 69.190 ;
        RECT 46.905 69.145 47.295 69.225 ;
        RECT 48.155 69.175 48.675 69.715 ;
        RECT 44.445 68.385 45.330 68.555 ;
        RECT 45.510 68.085 45.825 68.585 ;
        RECT 46.055 68.255 46.395 68.815 ;
        RECT 46.565 68.085 46.735 69.095 ;
        RECT 46.905 68.300 47.235 69.145 ;
        RECT 47.465 68.085 48.675 69.175 ;
        RECT 48.880 68.875 49.195 69.895 ;
        RECT 49.365 69.225 49.535 69.725 ;
        RECT 49.785 69.395 50.050 69.955 ;
        RECT 50.220 69.225 50.390 70.125 ;
        RECT 52.265 70.005 52.595 70.365 ;
        RECT 53.215 70.175 53.465 70.635 ;
        RECT 53.635 70.175 54.195 70.465 ;
        RECT 50.560 69.395 50.915 69.955 ;
        RECT 52.265 69.815 53.655 70.005 ;
        RECT 53.485 69.725 53.655 69.815 ;
        RECT 52.080 69.395 52.755 69.645 ;
        RECT 52.975 69.395 53.315 69.645 ;
        RECT 53.485 69.395 53.775 69.725 ;
        RECT 49.365 69.055 50.790 69.225 ;
        RECT 48.880 68.255 49.415 68.875 ;
        RECT 49.585 68.085 49.915 68.885 ;
        RECT 50.400 68.880 50.790 69.055 ;
        RECT 52.080 69.035 52.345 69.395 ;
        RECT 53.485 69.145 53.655 69.395 ;
        RECT 52.715 68.975 53.655 69.145 ;
        RECT 52.265 68.085 52.545 68.755 ;
        RECT 52.715 68.425 53.015 68.975 ;
        RECT 53.945 68.805 54.195 70.175 ;
        RECT 53.215 68.085 53.545 68.805 ;
        RECT 53.735 68.255 54.195 68.805 ;
        RECT 54.365 70.135 54.665 70.465 ;
        RECT 54.835 70.155 55.110 70.635 ;
        RECT 54.365 69.225 54.535 70.135 ;
        RECT 55.290 69.985 55.585 70.375 ;
        RECT 55.755 70.155 56.010 70.635 ;
        RECT 56.185 69.985 56.445 70.375 ;
        RECT 56.615 70.155 56.895 70.635 ;
        RECT 54.705 69.395 55.055 69.965 ;
        RECT 55.290 69.815 56.940 69.985 ;
        RECT 57.125 69.910 57.415 70.635 ;
        RECT 57.700 70.005 57.985 70.465 ;
        RECT 58.155 70.175 58.425 70.635 ;
        RECT 57.700 69.835 58.655 70.005 ;
        RECT 55.225 69.475 56.365 69.645 ;
        RECT 55.225 69.225 55.395 69.475 ;
        RECT 56.535 69.305 56.940 69.815 ;
        RECT 54.365 69.055 55.395 69.225 ;
        RECT 56.185 69.135 56.940 69.305 ;
        RECT 54.365 68.255 54.675 69.055 ;
        RECT 56.185 68.885 56.445 69.135 ;
        RECT 54.845 68.085 55.155 68.885 ;
        RECT 55.325 68.715 56.445 68.885 ;
        RECT 55.325 68.255 55.585 68.715 ;
        RECT 55.755 68.085 56.010 68.545 ;
        RECT 56.185 68.255 56.445 68.715 ;
        RECT 56.615 68.085 56.900 68.955 ;
        RECT 57.125 68.085 57.415 69.250 ;
        RECT 57.585 69.105 58.275 69.665 ;
        RECT 58.445 68.935 58.655 69.835 ;
        RECT 57.700 68.715 58.655 68.935 ;
        RECT 58.825 69.665 59.225 70.465 ;
        RECT 59.415 70.005 59.695 70.465 ;
        RECT 60.215 70.175 60.540 70.635 ;
        RECT 59.415 69.835 60.540 70.005 ;
        RECT 60.710 69.895 61.095 70.465 ;
        RECT 60.090 69.725 60.540 69.835 ;
        RECT 58.825 69.105 59.920 69.665 ;
        RECT 60.090 69.395 60.645 69.725 ;
        RECT 57.700 68.255 57.985 68.715 ;
        RECT 58.155 68.085 58.425 68.545 ;
        RECT 58.825 68.255 59.225 69.105 ;
        RECT 60.090 68.935 60.540 69.395 ;
        RECT 60.815 69.225 61.095 69.895 ;
        RECT 59.415 68.715 60.540 68.935 ;
        RECT 59.415 68.255 59.695 68.715 ;
        RECT 60.215 68.085 60.540 68.545 ;
        RECT 60.710 68.255 61.095 69.225 ;
        RECT 61.730 69.895 61.985 70.465 ;
        RECT 62.155 70.235 62.485 70.635 ;
        RECT 62.910 70.100 63.440 70.465 ;
        RECT 62.910 70.065 63.085 70.100 ;
        RECT 62.155 69.895 63.085 70.065 ;
        RECT 61.730 69.225 61.900 69.895 ;
        RECT 62.155 69.725 62.325 69.895 ;
        RECT 62.070 69.395 62.325 69.725 ;
        RECT 62.550 69.395 62.745 69.725 ;
        RECT 61.730 68.255 62.065 69.225 ;
        RECT 62.235 68.085 62.405 69.225 ;
        RECT 62.575 68.425 62.745 69.395 ;
        RECT 62.915 68.765 63.085 69.895 ;
        RECT 63.255 69.105 63.425 69.905 ;
        RECT 63.630 69.615 63.905 70.465 ;
        RECT 63.625 69.445 63.905 69.615 ;
        RECT 63.630 69.305 63.905 69.445 ;
        RECT 64.075 69.105 64.265 70.465 ;
        RECT 64.445 70.100 64.955 70.635 ;
        RECT 65.175 69.825 65.420 70.430 ;
        RECT 65.865 69.895 66.250 70.465 ;
        RECT 66.420 70.175 66.745 70.635 ;
        RECT 67.265 70.005 67.545 70.465 ;
        RECT 64.465 69.655 65.695 69.825 ;
        RECT 63.255 68.935 64.265 69.105 ;
        RECT 64.435 69.090 65.185 69.280 ;
        RECT 62.915 68.595 64.040 68.765 ;
        RECT 64.435 68.425 64.605 69.090 ;
        RECT 65.355 68.845 65.695 69.655 ;
        RECT 62.575 68.255 64.605 68.425 ;
        RECT 64.775 68.085 64.945 68.845 ;
        RECT 65.180 68.435 65.695 68.845 ;
        RECT 65.865 69.225 66.145 69.895 ;
        RECT 66.420 69.835 67.545 70.005 ;
        RECT 66.420 69.725 66.870 69.835 ;
        RECT 66.315 69.395 66.870 69.725 ;
        RECT 67.735 69.665 68.135 70.465 ;
        RECT 68.535 70.175 68.805 70.635 ;
        RECT 68.975 70.005 69.260 70.465 ;
        RECT 69.615 70.235 69.945 70.635 ;
        RECT 70.115 70.065 70.285 70.335 ;
        RECT 70.455 70.235 70.785 70.635 ;
        RECT 70.955 70.065 71.210 70.335 ;
        RECT 65.865 68.255 66.250 69.225 ;
        RECT 66.420 68.935 66.870 69.395 ;
        RECT 67.040 69.105 68.135 69.665 ;
        RECT 66.420 68.715 67.545 68.935 ;
        RECT 66.420 68.085 66.745 68.545 ;
        RECT 67.265 68.255 67.545 68.715 ;
        RECT 67.735 68.255 68.135 69.105 ;
        RECT 68.305 69.835 69.260 70.005 ;
        RECT 68.305 68.935 68.515 69.835 ;
        RECT 68.685 69.105 69.375 69.665 ;
        RECT 69.545 69.055 69.815 70.065 ;
        RECT 69.985 69.895 71.210 70.065 ;
        RECT 71.475 70.085 71.645 70.465 ;
        RECT 71.825 70.255 72.155 70.635 ;
        RECT 71.475 69.915 72.140 70.085 ;
        RECT 72.335 69.960 72.595 70.465 ;
        RECT 69.985 69.225 70.155 69.895 ;
        RECT 70.325 69.395 70.705 69.725 ;
        RECT 70.875 69.395 71.210 69.725 ;
        RECT 69.985 69.055 70.300 69.225 ;
        RECT 68.305 68.715 69.260 68.935 ;
        RECT 68.535 68.085 68.805 68.545 ;
        RECT 68.975 68.255 69.260 68.715 ;
        RECT 69.550 68.085 69.865 68.885 ;
        RECT 70.130 68.440 70.300 69.055 ;
        RECT 70.470 68.715 70.705 69.395 ;
        RECT 71.405 69.365 71.735 69.735 ;
        RECT 71.970 69.660 72.140 69.915 ;
        RECT 71.970 69.330 72.255 69.660 ;
        RECT 70.875 68.440 71.210 69.225 ;
        RECT 71.970 69.185 72.140 69.330 ;
        RECT 70.130 68.270 71.210 68.440 ;
        RECT 71.475 69.015 72.140 69.185 ;
        RECT 72.425 69.160 72.595 69.960 ;
        RECT 72.855 70.085 73.025 70.375 ;
        RECT 73.195 70.255 73.525 70.635 ;
        RECT 72.855 69.915 73.520 70.085 ;
        RECT 71.475 68.255 71.645 69.015 ;
        RECT 71.825 68.085 72.155 68.845 ;
        RECT 72.325 68.255 72.595 69.160 ;
        RECT 72.770 69.095 73.120 69.745 ;
        RECT 73.290 68.925 73.520 69.915 ;
        RECT 72.855 68.755 73.520 68.925 ;
        RECT 72.855 68.255 73.025 68.755 ;
        RECT 73.195 68.085 73.525 68.585 ;
        RECT 73.695 68.255 73.880 70.375 ;
        RECT 74.135 70.175 74.385 70.635 ;
        RECT 74.555 70.185 74.890 70.355 ;
        RECT 75.085 70.185 75.760 70.355 ;
        RECT 74.555 70.045 74.725 70.185 ;
        RECT 74.050 69.055 74.330 70.005 ;
        RECT 74.500 69.915 74.725 70.045 ;
        RECT 74.500 68.810 74.670 69.915 ;
        RECT 74.895 69.765 75.420 69.985 ;
        RECT 74.840 69.000 75.080 69.595 ;
        RECT 75.250 69.065 75.420 69.765 ;
        RECT 75.590 69.405 75.760 70.185 ;
        RECT 76.080 70.135 76.450 70.635 ;
        RECT 76.630 70.185 77.035 70.355 ;
        RECT 77.205 70.185 77.990 70.355 ;
        RECT 76.630 69.955 76.800 70.185 ;
        RECT 75.970 69.655 76.800 69.955 ;
        RECT 77.185 69.685 77.650 70.015 ;
        RECT 75.970 69.625 76.170 69.655 ;
        RECT 76.290 69.405 76.460 69.475 ;
        RECT 75.590 69.235 76.460 69.405 ;
        RECT 75.950 69.145 76.460 69.235 ;
        RECT 74.500 68.680 74.805 68.810 ;
        RECT 75.250 68.700 75.780 69.065 ;
        RECT 74.120 68.085 74.385 68.545 ;
        RECT 74.555 68.255 74.805 68.680 ;
        RECT 75.950 68.530 76.120 69.145 ;
        RECT 75.015 68.360 76.120 68.530 ;
        RECT 76.290 68.085 76.460 68.885 ;
        RECT 76.630 68.585 76.800 69.655 ;
        RECT 76.970 68.755 77.160 69.475 ;
        RECT 77.330 68.725 77.650 69.685 ;
        RECT 77.820 69.725 77.990 70.185 ;
        RECT 78.265 70.105 78.475 70.635 ;
        RECT 78.735 69.895 79.065 70.420 ;
        RECT 79.235 70.025 79.405 70.635 ;
        RECT 79.575 69.980 79.905 70.415 ;
        RECT 80.215 70.085 80.385 70.465 ;
        RECT 80.600 70.255 80.930 70.635 ;
        RECT 79.575 69.895 79.955 69.980 ;
        RECT 80.215 69.915 80.930 70.085 ;
        RECT 78.865 69.725 79.065 69.895 ;
        RECT 79.730 69.855 79.955 69.895 ;
        RECT 77.820 69.395 78.695 69.725 ;
        RECT 78.865 69.395 79.615 69.725 ;
        RECT 76.630 68.255 76.880 68.585 ;
        RECT 77.820 68.555 77.990 69.395 ;
        RECT 78.865 69.190 79.055 69.395 ;
        RECT 79.785 69.275 79.955 69.855 ;
        RECT 80.125 69.365 80.480 69.735 ;
        RECT 80.760 69.725 80.930 69.915 ;
        RECT 81.100 69.890 81.355 70.465 ;
        RECT 80.760 69.395 81.015 69.725 ;
        RECT 79.740 69.225 79.955 69.275 ;
        RECT 78.160 68.815 79.055 69.190 ;
        RECT 79.565 69.145 79.955 69.225 ;
        RECT 80.760 69.185 80.930 69.395 ;
        RECT 77.105 68.385 77.990 68.555 ;
        RECT 78.170 68.085 78.485 68.585 ;
        RECT 78.715 68.255 79.055 68.815 ;
        RECT 79.225 68.085 79.395 69.095 ;
        RECT 79.565 68.300 79.895 69.145 ;
        RECT 80.215 69.015 80.930 69.185 ;
        RECT 81.185 69.160 81.355 69.890 ;
        RECT 81.530 69.795 81.790 70.635 ;
        RECT 81.965 69.885 83.175 70.635 ;
        RECT 80.215 68.255 80.385 69.015 ;
        RECT 80.600 68.085 80.930 68.845 ;
        RECT 81.100 68.255 81.355 69.160 ;
        RECT 81.530 68.085 81.790 69.235 ;
        RECT 81.965 69.175 82.485 69.715 ;
        RECT 82.655 69.345 83.175 69.885 ;
        RECT 81.965 68.085 83.175 69.175 ;
        RECT 5.520 67.915 83.260 68.085 ;
        RECT 5.605 66.825 6.815 67.915 ;
        RECT 7.075 67.245 7.245 67.745 ;
        RECT 7.415 67.415 7.745 67.915 ;
        RECT 7.075 67.075 7.740 67.245 ;
        RECT 5.605 66.115 6.125 66.655 ;
        RECT 6.295 66.285 6.815 66.825 ;
        RECT 6.990 66.255 7.340 66.905 ;
        RECT 5.605 65.365 6.815 66.115 ;
        RECT 7.510 66.085 7.740 67.075 ;
        RECT 7.075 65.915 7.740 66.085 ;
        RECT 7.075 65.625 7.245 65.915 ;
        RECT 7.415 65.365 7.745 65.745 ;
        RECT 7.915 65.625 8.100 67.745 ;
        RECT 8.340 67.455 8.605 67.915 ;
        RECT 8.775 67.320 9.025 67.745 ;
        RECT 9.235 67.470 10.340 67.640 ;
        RECT 8.720 67.190 9.025 67.320 ;
        RECT 8.270 65.995 8.550 66.945 ;
        RECT 8.720 66.085 8.890 67.190 ;
        RECT 9.060 66.405 9.300 67.000 ;
        RECT 9.470 66.935 10.000 67.300 ;
        RECT 9.470 66.235 9.640 66.935 ;
        RECT 10.170 66.855 10.340 67.470 ;
        RECT 10.510 67.115 10.680 67.915 ;
        RECT 10.850 67.415 11.100 67.745 ;
        RECT 11.325 67.445 12.210 67.615 ;
        RECT 10.170 66.765 10.680 66.855 ;
        RECT 8.720 65.955 8.945 66.085 ;
        RECT 9.115 66.015 9.640 66.235 ;
        RECT 9.810 66.595 10.680 66.765 ;
        RECT 8.355 65.365 8.605 65.825 ;
        RECT 8.775 65.815 8.945 65.955 ;
        RECT 9.810 65.815 9.980 66.595 ;
        RECT 10.510 66.525 10.680 66.595 ;
        RECT 10.190 66.345 10.390 66.375 ;
        RECT 10.850 66.345 11.020 67.415 ;
        RECT 11.190 66.525 11.380 67.245 ;
        RECT 10.190 66.045 11.020 66.345 ;
        RECT 11.550 66.315 11.870 67.275 ;
        RECT 8.775 65.645 9.110 65.815 ;
        RECT 9.305 65.645 9.980 65.815 ;
        RECT 10.300 65.365 10.670 65.865 ;
        RECT 10.850 65.815 11.020 66.045 ;
        RECT 11.405 65.985 11.870 66.315 ;
        RECT 12.040 66.605 12.210 67.445 ;
        RECT 12.390 67.415 12.705 67.915 ;
        RECT 12.935 67.185 13.275 67.745 ;
        RECT 12.380 66.810 13.275 67.185 ;
        RECT 13.445 66.905 13.615 67.915 ;
        RECT 13.085 66.605 13.275 66.810 ;
        RECT 13.785 66.855 14.115 67.700 ;
        RECT 14.815 67.305 15.145 67.735 ;
        RECT 15.325 67.475 15.520 67.915 ;
        RECT 15.690 67.305 16.020 67.735 ;
        RECT 14.815 67.135 16.020 67.305 ;
        RECT 13.785 66.775 14.175 66.855 ;
        RECT 14.815 66.805 15.710 67.135 ;
        RECT 16.190 66.965 16.465 67.735 ;
        RECT 16.650 67.115 16.905 67.915 ;
        RECT 17.105 67.065 17.435 67.745 ;
        RECT 13.960 66.725 14.175 66.775 ;
        RECT 12.040 66.275 12.915 66.605 ;
        RECT 13.085 66.275 13.835 66.605 ;
        RECT 12.040 65.815 12.210 66.275 ;
        RECT 13.085 66.105 13.285 66.275 ;
        RECT 14.005 66.145 14.175 66.725 ;
        RECT 15.880 66.775 16.465 66.965 ;
        RECT 14.820 66.275 15.115 66.605 ;
        RECT 15.295 66.275 15.710 66.605 ;
        RECT 13.950 66.105 14.175 66.145 ;
        RECT 10.850 65.645 11.255 65.815 ;
        RECT 11.425 65.645 12.210 65.815 ;
        RECT 12.485 65.365 12.695 65.895 ;
        RECT 12.955 65.580 13.285 66.105 ;
        RECT 13.795 66.020 14.175 66.105 ;
        RECT 13.455 65.365 13.625 65.975 ;
        RECT 13.795 65.585 14.125 66.020 ;
        RECT 14.815 65.365 15.115 66.095 ;
        RECT 15.295 65.655 15.525 66.275 ;
        RECT 15.880 66.105 16.055 66.775 ;
        RECT 15.725 65.925 16.055 66.105 ;
        RECT 16.225 65.955 16.465 66.605 ;
        RECT 16.650 66.575 16.895 66.935 ;
        RECT 17.085 66.785 17.435 67.065 ;
        RECT 17.085 66.405 17.255 66.785 ;
        RECT 17.615 66.605 17.810 67.655 ;
        RECT 17.990 66.775 18.310 67.915 ;
        RECT 18.485 66.750 18.775 67.915 ;
        RECT 18.945 66.945 19.235 67.745 ;
        RECT 19.405 67.115 19.640 67.915 ;
        RECT 19.825 67.575 21.360 67.745 ;
        RECT 19.825 66.945 20.155 67.575 ;
        RECT 18.945 66.775 20.155 66.945 ;
        RECT 16.735 66.235 17.255 66.405 ;
        RECT 17.425 66.275 17.810 66.605 ;
        RECT 17.990 66.555 18.250 66.605 ;
        RECT 17.990 66.385 18.255 66.555 ;
        RECT 17.990 66.275 18.250 66.385 ;
        RECT 18.945 66.275 19.190 66.605 ;
        RECT 16.735 66.215 16.905 66.235 ;
        RECT 16.705 66.045 16.905 66.215 ;
        RECT 19.360 66.105 19.530 66.775 ;
        RECT 20.325 66.605 20.560 67.350 ;
        RECT 19.700 66.275 20.100 66.605 ;
        RECT 20.270 66.275 20.560 66.605 ;
        RECT 20.750 66.605 21.020 67.350 ;
        RECT 21.190 66.945 21.360 67.575 ;
        RECT 21.530 67.115 21.935 67.915 ;
        RECT 21.190 66.775 21.935 66.945 ;
        RECT 20.750 66.275 21.090 66.605 ;
        RECT 21.260 66.275 21.595 66.605 ;
        RECT 21.765 66.275 21.935 66.775 ;
        RECT 22.105 66.350 22.455 67.745 ;
        RECT 23.095 66.805 23.390 67.915 ;
        RECT 23.570 66.605 23.820 67.740 ;
        RECT 23.990 66.805 24.250 67.915 ;
        RECT 24.420 67.015 24.680 67.740 ;
        RECT 24.850 67.185 25.110 67.915 ;
        RECT 25.280 67.015 25.540 67.740 ;
        RECT 25.710 67.185 25.970 67.915 ;
        RECT 26.140 67.015 26.400 67.740 ;
        RECT 26.570 67.185 26.830 67.915 ;
        RECT 27.000 67.015 27.260 67.740 ;
        RECT 27.430 67.185 27.725 67.915 ;
        RECT 24.420 66.775 27.730 67.015 ;
        RECT 28.145 66.825 29.815 67.915 ;
        RECT 30.560 67.285 30.845 67.745 ;
        RECT 31.015 67.455 31.285 67.915 ;
        RECT 30.560 67.065 31.515 67.285 ;
        RECT 15.725 65.545 15.950 65.925 ;
        RECT 16.120 65.365 16.450 65.755 ;
        RECT 16.735 65.670 16.905 66.045 ;
        RECT 17.095 65.895 18.310 66.065 ;
        RECT 17.095 65.590 17.325 65.895 ;
        RECT 17.495 65.365 17.825 65.725 ;
        RECT 18.020 65.545 18.310 65.895 ;
        RECT 18.485 65.365 18.775 66.090 ;
        RECT 18.945 65.535 19.530 66.105 ;
        RECT 19.780 65.935 21.175 66.105 ;
        RECT 19.780 65.590 20.110 65.935 ;
        RECT 20.325 65.365 20.700 65.765 ;
        RECT 20.880 65.590 21.175 65.935 ;
        RECT 21.345 65.365 22.015 66.105 ;
        RECT 22.185 65.535 22.455 66.350 ;
        RECT 23.085 65.995 23.400 66.605 ;
        RECT 23.570 66.355 26.590 66.605 ;
        RECT 23.145 65.365 23.390 65.825 ;
        RECT 23.570 65.545 23.820 66.355 ;
        RECT 26.760 66.185 27.730 66.775 ;
        RECT 24.420 66.015 27.730 66.185 ;
        RECT 28.145 66.135 28.895 66.655 ;
        RECT 29.065 66.305 29.815 66.825 ;
        RECT 30.445 66.335 31.135 66.895 ;
        RECT 31.305 66.165 31.515 67.065 ;
        RECT 23.990 65.365 24.250 65.890 ;
        RECT 24.420 65.560 24.680 66.015 ;
        RECT 24.850 65.365 25.110 65.845 ;
        RECT 25.280 65.560 25.540 66.015 ;
        RECT 25.710 65.365 25.970 65.845 ;
        RECT 26.140 65.560 26.400 66.015 ;
        RECT 26.570 65.365 26.830 65.845 ;
        RECT 27.000 65.560 27.260 66.015 ;
        RECT 27.430 65.365 27.730 65.845 ;
        RECT 28.145 65.365 29.815 66.135 ;
        RECT 30.560 65.995 31.515 66.165 ;
        RECT 31.685 66.895 32.085 67.745 ;
        RECT 32.275 67.285 32.555 67.745 ;
        RECT 33.075 67.455 33.400 67.915 ;
        RECT 32.275 67.065 33.400 67.285 ;
        RECT 31.685 66.335 32.780 66.895 ;
        RECT 32.950 66.605 33.400 67.065 ;
        RECT 33.570 66.775 33.955 67.745 ;
        RECT 34.125 66.840 34.465 67.915 ;
        RECT 34.650 67.405 36.700 67.695 ;
        RECT 30.560 65.535 30.845 65.995 ;
        RECT 31.015 65.365 31.285 65.825 ;
        RECT 31.685 65.535 32.085 66.335 ;
        RECT 32.950 66.275 33.505 66.605 ;
        RECT 32.950 66.165 33.400 66.275 ;
        RECT 32.275 65.995 33.400 66.165 ;
        RECT 33.675 66.105 33.955 66.775 ;
        RECT 34.635 66.605 34.875 67.200 ;
        RECT 35.070 67.065 36.700 67.235 ;
        RECT 36.870 67.115 37.150 67.915 ;
        RECT 35.070 66.775 35.390 67.065 ;
        RECT 36.530 66.945 36.700 67.065 ;
        RECT 32.275 65.535 32.555 65.995 ;
        RECT 33.075 65.365 33.400 65.825 ;
        RECT 33.570 65.535 33.955 66.105 ;
        RECT 34.125 66.035 34.465 66.605 ;
        RECT 34.635 66.275 35.290 66.605 ;
        RECT 35.560 66.275 36.300 66.895 ;
        RECT 36.530 66.775 37.190 66.945 ;
        RECT 37.360 66.775 37.635 67.745 ;
        RECT 37.805 66.825 39.015 67.915 ;
        RECT 37.020 66.605 37.190 66.775 ;
        RECT 36.470 66.275 36.850 66.605 ;
        RECT 37.020 66.275 37.295 66.605 ;
        RECT 34.125 65.365 34.465 65.865 ;
        RECT 34.635 65.585 34.880 66.275 ;
        RECT 37.020 66.105 37.190 66.275 ;
        RECT 35.605 65.935 37.190 66.105 ;
        RECT 37.465 66.040 37.635 66.775 ;
        RECT 35.075 65.365 35.405 65.865 ;
        RECT 35.605 65.585 35.775 65.935 ;
        RECT 35.950 65.365 36.280 65.765 ;
        RECT 36.450 65.585 36.620 65.935 ;
        RECT 36.790 65.365 37.170 65.765 ;
        RECT 37.360 65.695 37.635 66.040 ;
        RECT 37.805 66.115 38.325 66.655 ;
        RECT 38.495 66.285 39.015 66.825 ;
        RECT 39.185 66.775 39.570 67.745 ;
        RECT 39.740 67.455 40.065 67.915 ;
        RECT 40.585 67.285 40.865 67.745 ;
        RECT 39.740 67.065 40.865 67.285 ;
        RECT 37.805 65.365 39.015 66.115 ;
        RECT 39.185 66.105 39.465 66.775 ;
        RECT 39.740 66.605 40.190 67.065 ;
        RECT 41.055 66.895 41.455 67.745 ;
        RECT 41.855 67.455 42.125 67.915 ;
        RECT 42.295 67.285 42.580 67.745 ;
        RECT 39.635 66.275 40.190 66.605 ;
        RECT 40.360 66.335 41.455 66.895 ;
        RECT 39.740 66.165 40.190 66.275 ;
        RECT 39.185 65.535 39.570 66.105 ;
        RECT 39.740 65.995 40.865 66.165 ;
        RECT 39.740 65.365 40.065 65.825 ;
        RECT 40.585 65.535 40.865 65.995 ;
        RECT 41.055 65.535 41.455 66.335 ;
        RECT 41.625 67.065 42.580 67.285 ;
        RECT 41.625 66.165 41.835 67.065 ;
        RECT 42.005 66.335 42.695 66.895 ;
        RECT 42.865 66.825 44.075 67.915 ;
        RECT 41.625 65.995 42.580 66.165 ;
        RECT 41.855 65.365 42.125 65.825 ;
        RECT 42.295 65.535 42.580 65.995 ;
        RECT 42.865 66.115 43.385 66.655 ;
        RECT 43.555 66.285 44.075 66.825 ;
        RECT 44.245 66.750 44.535 67.915 ;
        RECT 44.705 66.825 48.215 67.915 ;
        RECT 44.705 66.135 46.355 66.655 ;
        RECT 46.525 66.305 48.215 66.825 ;
        RECT 49.395 66.985 49.565 67.745 ;
        RECT 49.780 67.155 50.110 67.915 ;
        RECT 49.395 66.815 50.110 66.985 ;
        RECT 50.280 66.840 50.535 67.745 ;
        RECT 49.305 66.265 49.660 66.635 ;
        RECT 49.940 66.605 50.110 66.815 ;
        RECT 49.940 66.275 50.195 66.605 ;
        RECT 42.865 65.365 44.075 66.115 ;
        RECT 44.245 65.365 44.535 66.090 ;
        RECT 44.705 65.365 48.215 66.135 ;
        RECT 49.940 66.085 50.110 66.275 ;
        RECT 50.365 66.110 50.535 66.840 ;
        RECT 50.710 66.765 50.970 67.915 ;
        RECT 51.155 66.945 51.485 67.745 ;
        RECT 51.655 67.115 51.885 67.915 ;
        RECT 52.055 66.945 52.385 67.745 ;
        RECT 51.155 66.775 52.385 66.945 ;
        RECT 52.555 66.775 52.810 67.915 ;
        RECT 53.100 67.285 53.385 67.745 ;
        RECT 53.555 67.455 53.825 67.915 ;
        RECT 53.100 67.065 54.055 67.285 ;
        RECT 51.145 66.275 51.455 66.605 ;
        RECT 49.395 65.915 50.110 66.085 ;
        RECT 49.395 65.535 49.565 65.915 ;
        RECT 49.780 65.365 50.110 65.745 ;
        RECT 50.280 65.535 50.535 66.110 ;
        RECT 50.710 65.365 50.970 66.205 ;
        RECT 51.155 65.875 51.485 66.105 ;
        RECT 51.660 66.045 52.035 66.605 ;
        RECT 52.205 65.875 52.385 66.775 ;
        RECT 52.570 66.025 52.790 66.605 ;
        RECT 52.985 66.335 53.675 66.895 ;
        RECT 53.845 66.165 54.055 67.065 ;
        RECT 51.155 65.535 52.385 65.875 ;
        RECT 53.100 65.995 54.055 66.165 ;
        RECT 54.225 66.895 54.625 67.745 ;
        RECT 54.815 67.285 55.095 67.745 ;
        RECT 55.615 67.455 55.940 67.915 ;
        RECT 54.815 67.065 55.940 67.285 ;
        RECT 54.225 66.335 55.320 66.895 ;
        RECT 55.490 66.605 55.940 67.065 ;
        RECT 56.110 66.775 56.495 67.745 ;
        RECT 52.555 65.365 52.810 65.855 ;
        RECT 53.100 65.535 53.385 65.995 ;
        RECT 53.555 65.365 53.825 65.825 ;
        RECT 54.225 65.535 54.625 66.335 ;
        RECT 55.490 66.275 56.045 66.605 ;
        RECT 55.490 66.165 55.940 66.275 ;
        RECT 54.815 65.995 55.940 66.165 ;
        RECT 56.215 66.105 56.495 66.775 ;
        RECT 56.670 67.525 57.005 67.745 ;
        RECT 58.010 67.535 58.365 67.915 ;
        RECT 56.670 66.905 56.925 67.525 ;
        RECT 57.175 67.365 57.405 67.405 ;
        RECT 58.535 67.365 58.785 67.745 ;
        RECT 57.175 67.165 58.785 67.365 ;
        RECT 57.175 67.075 57.360 67.165 ;
        RECT 57.950 67.155 58.785 67.165 ;
        RECT 59.035 67.135 59.285 67.915 ;
        RECT 59.455 67.065 59.715 67.745 ;
        RECT 59.975 67.245 60.145 67.745 ;
        RECT 60.315 67.415 60.645 67.915 ;
        RECT 59.975 67.075 60.640 67.245 ;
        RECT 57.515 66.965 57.845 66.995 ;
        RECT 57.515 66.905 59.315 66.965 ;
        RECT 56.670 66.795 59.375 66.905 ;
        RECT 56.670 66.735 57.845 66.795 ;
        RECT 59.175 66.760 59.375 66.795 ;
        RECT 56.665 66.355 57.155 66.555 ;
        RECT 57.345 66.355 57.820 66.565 ;
        RECT 54.815 65.535 55.095 65.995 ;
        RECT 55.615 65.365 55.940 65.825 ;
        RECT 56.110 65.535 56.495 66.105 ;
        RECT 56.670 65.365 57.125 66.130 ;
        RECT 57.600 65.955 57.820 66.355 ;
        RECT 58.065 66.355 58.395 66.565 ;
        RECT 58.065 65.955 58.275 66.355 ;
        RECT 58.565 66.320 58.975 66.625 ;
        RECT 59.205 66.185 59.375 66.760 ;
        RECT 59.105 66.065 59.375 66.185 ;
        RECT 58.530 66.020 59.375 66.065 ;
        RECT 58.530 65.895 59.285 66.020 ;
        RECT 58.530 65.745 58.700 65.895 ;
        RECT 59.545 65.875 59.715 67.065 ;
        RECT 59.890 66.255 60.240 66.905 ;
        RECT 60.410 66.085 60.640 67.075 ;
        RECT 59.485 65.865 59.715 65.875 ;
        RECT 57.400 65.535 58.700 65.745 ;
        RECT 58.955 65.365 59.285 65.725 ;
        RECT 59.455 65.535 59.715 65.865 ;
        RECT 59.975 65.915 60.640 66.085 ;
        RECT 59.975 65.625 60.145 65.915 ;
        RECT 60.315 65.365 60.645 65.745 ;
        RECT 60.815 65.625 61.000 67.745 ;
        RECT 61.240 67.455 61.505 67.915 ;
        RECT 61.675 67.320 61.925 67.745 ;
        RECT 62.135 67.470 63.240 67.640 ;
        RECT 61.620 67.190 61.925 67.320 ;
        RECT 61.170 65.995 61.450 66.945 ;
        RECT 61.620 66.085 61.790 67.190 ;
        RECT 61.960 66.405 62.200 67.000 ;
        RECT 62.370 66.935 62.900 67.300 ;
        RECT 62.370 66.235 62.540 66.935 ;
        RECT 63.070 66.855 63.240 67.470 ;
        RECT 63.410 67.115 63.580 67.915 ;
        RECT 63.750 67.415 64.000 67.745 ;
        RECT 64.225 67.445 65.110 67.615 ;
        RECT 63.070 66.765 63.580 66.855 ;
        RECT 61.620 65.955 61.845 66.085 ;
        RECT 62.015 66.015 62.540 66.235 ;
        RECT 62.710 66.595 63.580 66.765 ;
        RECT 61.255 65.365 61.505 65.825 ;
        RECT 61.675 65.815 61.845 65.955 ;
        RECT 62.710 65.815 62.880 66.595 ;
        RECT 63.410 66.525 63.580 66.595 ;
        RECT 63.090 66.345 63.290 66.375 ;
        RECT 63.750 66.345 63.920 67.415 ;
        RECT 64.090 66.525 64.280 67.245 ;
        RECT 63.090 66.045 63.920 66.345 ;
        RECT 64.450 66.315 64.770 67.275 ;
        RECT 61.675 65.645 62.010 65.815 ;
        RECT 62.205 65.645 62.880 65.815 ;
        RECT 63.200 65.365 63.570 65.865 ;
        RECT 63.750 65.815 63.920 66.045 ;
        RECT 64.305 65.985 64.770 66.315 ;
        RECT 64.940 66.605 65.110 67.445 ;
        RECT 65.290 67.415 65.605 67.915 ;
        RECT 65.835 67.185 66.175 67.745 ;
        RECT 65.280 66.810 66.175 67.185 ;
        RECT 66.345 66.905 66.515 67.915 ;
        RECT 65.985 66.605 66.175 66.810 ;
        RECT 66.685 66.855 67.015 67.700 ;
        RECT 66.685 66.775 67.075 66.855 ;
        RECT 66.860 66.725 67.075 66.775 ;
        RECT 68.170 66.765 68.430 67.915 ;
        RECT 68.605 66.840 68.860 67.745 ;
        RECT 69.030 67.155 69.360 67.915 ;
        RECT 69.575 66.985 69.745 67.745 ;
        RECT 64.940 66.275 65.815 66.605 ;
        RECT 65.985 66.275 66.735 66.605 ;
        RECT 64.940 65.815 65.110 66.275 ;
        RECT 65.985 66.105 66.185 66.275 ;
        RECT 66.905 66.145 67.075 66.725 ;
        RECT 66.850 66.105 67.075 66.145 ;
        RECT 63.750 65.645 64.155 65.815 ;
        RECT 64.325 65.645 65.110 65.815 ;
        RECT 65.385 65.365 65.595 65.895 ;
        RECT 65.855 65.580 66.185 66.105 ;
        RECT 66.695 66.020 67.075 66.105 ;
        RECT 66.355 65.365 66.525 65.975 ;
        RECT 66.695 65.585 67.025 66.020 ;
        RECT 68.170 65.365 68.430 66.205 ;
        RECT 68.605 66.110 68.775 66.840 ;
        RECT 69.030 66.815 69.745 66.985 ;
        RECT 69.030 66.605 69.200 66.815 ;
        RECT 70.005 66.750 70.295 67.915 ;
        RECT 70.465 66.775 70.850 67.745 ;
        RECT 71.020 67.455 71.345 67.915 ;
        RECT 71.865 67.285 72.145 67.745 ;
        RECT 71.020 67.065 72.145 67.285 ;
        RECT 68.945 66.275 69.200 66.605 ;
        RECT 68.605 65.535 68.860 66.110 ;
        RECT 69.030 66.085 69.200 66.275 ;
        RECT 69.480 66.265 69.835 66.635 ;
        RECT 70.465 66.105 70.745 66.775 ;
        RECT 71.020 66.605 71.470 67.065 ;
        RECT 72.335 66.895 72.735 67.745 ;
        RECT 73.135 67.455 73.405 67.915 ;
        RECT 73.575 67.285 73.860 67.745 ;
        RECT 74.150 67.490 74.485 67.915 ;
        RECT 74.655 67.310 74.840 67.715 ;
        RECT 70.915 66.275 71.470 66.605 ;
        RECT 71.640 66.335 72.735 66.895 ;
        RECT 71.020 66.165 71.470 66.275 ;
        RECT 69.030 65.915 69.745 66.085 ;
        RECT 69.030 65.365 69.360 65.745 ;
        RECT 69.575 65.535 69.745 65.915 ;
        RECT 70.005 65.365 70.295 66.090 ;
        RECT 70.465 65.535 70.850 66.105 ;
        RECT 71.020 65.995 72.145 66.165 ;
        RECT 71.020 65.365 71.345 65.825 ;
        RECT 71.865 65.535 72.145 65.995 ;
        RECT 72.335 65.535 72.735 66.335 ;
        RECT 72.905 67.065 73.860 67.285 ;
        RECT 74.175 67.135 74.840 67.310 ;
        RECT 75.045 67.135 75.375 67.915 ;
        RECT 72.905 66.165 73.115 67.065 ;
        RECT 73.285 66.335 73.975 66.895 ;
        RECT 72.905 65.995 73.860 66.165 ;
        RECT 73.135 65.365 73.405 65.825 ;
        RECT 73.575 65.535 73.860 65.995 ;
        RECT 74.175 66.105 74.515 67.135 ;
        RECT 75.545 66.945 75.815 67.715 ;
        RECT 74.685 66.775 75.815 66.945 ;
        RECT 76.075 66.985 76.245 67.745 ;
        RECT 76.460 67.155 76.790 67.915 ;
        RECT 76.075 66.815 76.790 66.985 ;
        RECT 76.960 66.840 77.215 67.745 ;
        RECT 74.685 66.275 74.935 66.775 ;
        RECT 74.175 65.935 74.860 66.105 ;
        RECT 75.115 66.025 75.475 66.605 ;
        RECT 74.150 65.365 74.485 65.765 ;
        RECT 74.655 65.535 74.860 65.935 ;
        RECT 75.645 65.865 75.815 66.775 ;
        RECT 75.985 66.265 76.340 66.635 ;
        RECT 76.620 66.605 76.790 66.815 ;
        RECT 76.620 66.275 76.875 66.605 ;
        RECT 76.620 66.085 76.790 66.275 ;
        RECT 77.045 66.110 77.215 66.840 ;
        RECT 77.390 66.765 77.650 67.915 ;
        RECT 77.825 67.065 78.085 67.745 ;
        RECT 78.255 67.135 78.505 67.915 ;
        RECT 78.755 67.365 79.005 67.745 ;
        RECT 79.175 67.535 79.530 67.915 ;
        RECT 80.535 67.525 80.870 67.745 ;
        RECT 80.135 67.365 80.365 67.405 ;
        RECT 78.755 67.165 80.365 67.365 ;
        RECT 78.755 67.155 79.590 67.165 ;
        RECT 80.180 67.075 80.365 67.165 ;
        RECT 75.070 65.365 75.345 65.845 ;
        RECT 75.555 65.535 75.815 65.865 ;
        RECT 76.075 65.915 76.790 66.085 ;
        RECT 76.075 65.535 76.245 65.915 ;
        RECT 76.460 65.365 76.790 65.745 ;
        RECT 76.960 65.535 77.215 66.110 ;
        RECT 77.390 65.365 77.650 66.205 ;
        RECT 77.825 65.865 77.995 67.065 ;
        RECT 79.695 66.965 80.025 66.995 ;
        RECT 78.225 66.905 80.025 66.965 ;
        RECT 80.615 66.905 80.870 67.525 ;
        RECT 78.165 66.795 80.870 66.905 ;
        RECT 78.165 66.760 78.365 66.795 ;
        RECT 78.165 66.185 78.335 66.760 ;
        RECT 79.695 66.735 80.870 66.795 ;
        RECT 81.965 66.825 83.175 67.915 ;
        RECT 78.565 66.320 78.975 66.625 ;
        RECT 79.145 66.355 79.475 66.565 ;
        RECT 78.165 66.065 78.435 66.185 ;
        RECT 78.165 66.020 79.010 66.065 ;
        RECT 78.255 65.895 79.010 66.020 ;
        RECT 79.265 65.955 79.475 66.355 ;
        RECT 79.720 66.355 80.195 66.565 ;
        RECT 80.385 66.355 80.875 66.555 ;
        RECT 79.720 65.955 79.940 66.355 ;
        RECT 81.965 66.285 82.485 66.825 ;
        RECT 77.825 65.535 78.085 65.865 ;
        RECT 78.840 65.745 79.010 65.895 ;
        RECT 78.255 65.365 78.585 65.725 ;
        RECT 78.840 65.535 80.140 65.745 ;
        RECT 80.415 65.365 80.870 66.130 ;
        RECT 82.655 66.115 83.175 66.655 ;
        RECT 81.965 65.365 83.175 66.115 ;
        RECT 5.520 65.195 83.260 65.365 ;
        RECT 5.605 64.445 6.815 65.195 ;
        RECT 7.905 64.475 8.245 64.985 ;
        RECT 5.605 63.905 6.125 64.445 ;
        RECT 6.295 63.735 6.815 64.275 ;
        RECT 5.605 62.645 6.815 63.735 ;
        RECT 7.905 63.075 8.165 64.475 ;
        RECT 8.415 64.395 8.685 65.195 ;
        RECT 8.340 63.955 8.670 64.205 ;
        RECT 8.865 63.955 9.145 64.925 ;
        RECT 9.325 63.955 9.625 64.925 ;
        RECT 9.805 63.955 10.155 64.920 ;
        RECT 10.375 64.695 10.870 65.025 ;
        RECT 8.355 63.785 8.670 63.955 ;
        RECT 10.375 63.785 10.545 64.695 ;
        RECT 8.355 63.615 10.545 63.785 ;
        RECT 7.905 62.815 8.245 63.075 ;
        RECT 8.415 62.645 8.745 63.445 ;
        RECT 9.210 62.815 9.460 63.615 ;
        RECT 9.645 62.645 9.975 63.365 ;
        RECT 10.195 62.815 10.445 63.615 ;
        RECT 10.715 63.205 10.955 64.515 ;
        RECT 11.160 64.455 11.775 65.025 ;
        RECT 11.945 64.685 12.160 65.195 ;
        RECT 12.390 64.685 12.670 65.015 ;
        RECT 12.850 64.685 13.090 65.195 ;
        RECT 11.160 63.435 11.475 64.455 ;
        RECT 11.645 63.785 11.815 64.285 ;
        RECT 12.065 63.955 12.330 64.515 ;
        RECT 12.500 63.785 12.670 64.685 ;
        RECT 12.840 63.955 13.195 64.515 ;
        RECT 13.435 64.465 13.735 65.195 ;
        RECT 13.915 64.285 14.145 64.905 ;
        RECT 14.345 64.635 14.570 65.015 ;
        RECT 14.740 64.805 15.070 65.195 ;
        RECT 14.345 64.455 14.675 64.635 ;
        RECT 13.440 63.955 13.735 64.285 ;
        RECT 13.915 63.955 14.330 64.285 ;
        RECT 14.500 63.785 14.675 64.455 ;
        RECT 14.845 63.955 15.085 64.605 ;
        RECT 15.465 64.565 15.795 64.925 ;
        RECT 16.415 64.735 16.665 65.195 ;
        RECT 16.835 64.735 17.395 65.025 ;
        RECT 15.465 64.375 16.855 64.565 ;
        RECT 16.685 64.285 16.855 64.375 ;
        RECT 15.280 63.955 15.955 64.205 ;
        RECT 16.175 63.955 16.515 64.205 ;
        RECT 16.685 63.955 16.975 64.285 ;
        RECT 11.645 63.615 13.070 63.785 ;
        RECT 10.615 62.645 10.950 63.025 ;
        RECT 11.160 62.815 11.695 63.435 ;
        RECT 11.865 62.645 12.195 63.445 ;
        RECT 12.680 63.440 13.070 63.615 ;
        RECT 13.435 63.425 14.330 63.755 ;
        RECT 14.500 63.595 15.085 63.785 ;
        RECT 15.280 63.595 15.545 63.955 ;
        RECT 16.685 63.705 16.855 63.955 ;
        RECT 13.435 63.255 14.640 63.425 ;
        RECT 13.435 62.825 13.765 63.255 ;
        RECT 13.945 62.645 14.140 63.085 ;
        RECT 14.310 62.825 14.640 63.255 ;
        RECT 14.810 62.825 15.085 63.595 ;
        RECT 15.915 63.535 16.855 63.705 ;
        RECT 15.465 62.645 15.745 63.315 ;
        RECT 15.915 62.985 16.215 63.535 ;
        RECT 17.145 63.365 17.395 64.735 ;
        RECT 16.415 62.645 16.745 63.365 ;
        RECT 16.935 62.815 17.395 63.365 ;
        RECT 17.565 64.610 17.875 65.025 ;
        RECT 18.070 64.815 18.400 65.195 ;
        RECT 18.570 64.855 19.975 65.025 ;
        RECT 18.570 64.625 18.740 64.855 ;
        RECT 17.565 63.495 17.735 64.610 ;
        RECT 18.045 64.455 18.740 64.625 ;
        RECT 19.805 64.625 19.975 64.855 ;
        RECT 20.245 64.795 20.575 65.195 ;
        RECT 20.815 64.625 20.985 65.025 ;
        RECT 18.045 64.285 18.215 64.455 ;
        RECT 17.905 63.955 18.215 64.285 ;
        RECT 18.385 63.955 18.720 64.285 ;
        RECT 18.990 63.955 19.185 64.530 ;
        RECT 19.445 64.285 19.635 64.515 ;
        RECT 19.805 64.455 20.985 64.625 ;
        RECT 22.165 64.375 22.425 65.195 ;
        RECT 22.595 64.375 22.925 64.795 ;
        RECT 23.105 64.710 23.895 64.975 ;
        RECT 22.675 64.285 22.925 64.375 ;
        RECT 19.445 63.955 19.790 64.285 ;
        RECT 20.100 63.955 20.575 64.285 ;
        RECT 20.830 63.955 21.015 64.285 ;
        RECT 18.045 63.785 18.215 63.955 ;
        RECT 18.045 63.615 20.985 63.785 ;
        RECT 17.565 62.855 17.905 63.495 ;
        RECT 18.495 63.275 20.055 63.445 ;
        RECT 18.075 62.645 18.320 63.105 ;
        RECT 18.495 62.815 18.745 63.275 ;
        RECT 18.935 62.645 19.605 63.025 ;
        RECT 19.805 62.815 20.055 63.275 ;
        RECT 20.815 62.815 20.985 63.615 ;
        RECT 22.165 63.325 22.505 64.205 ;
        RECT 22.675 64.035 23.470 64.285 ;
        RECT 22.165 62.645 22.425 63.155 ;
        RECT 22.675 62.815 22.845 64.035 ;
        RECT 23.640 63.855 23.895 64.710 ;
        RECT 24.065 64.555 24.265 64.975 ;
        RECT 24.455 64.735 24.785 65.195 ;
        RECT 24.065 64.035 24.475 64.555 ;
        RECT 24.955 64.545 25.215 65.025 ;
        RECT 24.645 63.855 24.875 64.285 ;
        RECT 23.085 63.685 24.875 63.855 ;
        RECT 23.085 63.320 23.335 63.685 ;
        RECT 23.505 63.325 23.835 63.515 ;
        RECT 24.055 63.390 24.770 63.685 ;
        RECT 25.045 63.515 25.215 64.545 ;
        RECT 25.545 64.635 25.875 65.025 ;
        RECT 26.045 64.805 27.230 64.975 ;
        RECT 27.490 64.725 27.660 65.195 ;
        RECT 25.545 64.455 26.055 64.635 ;
        RECT 25.385 63.995 25.715 64.285 ;
        RECT 25.885 63.825 26.055 64.455 ;
        RECT 26.460 64.545 26.845 64.635 ;
        RECT 27.830 64.545 28.160 65.010 ;
        RECT 26.460 64.375 28.160 64.545 ;
        RECT 28.330 64.375 28.500 65.195 ;
        RECT 28.670 64.375 29.355 65.015 ;
        RECT 29.985 64.395 30.295 65.195 ;
        RECT 30.500 64.395 31.195 65.025 ;
        RECT 31.365 64.470 31.655 65.195 ;
        RECT 26.225 63.995 26.555 64.205 ;
        RECT 26.735 63.955 27.115 64.205 ;
        RECT 23.505 63.150 23.700 63.325 ;
        RECT 23.085 62.645 23.700 63.150 ;
        RECT 23.870 62.815 24.345 63.155 ;
        RECT 24.515 62.645 24.730 63.190 ;
        RECT 24.940 62.815 25.215 63.515 ;
        RECT 25.540 63.655 26.625 63.825 ;
        RECT 25.540 62.815 25.840 63.655 ;
        RECT 26.035 62.645 26.285 63.485 ;
        RECT 26.455 63.405 26.625 63.655 ;
        RECT 26.795 63.575 27.115 63.955 ;
        RECT 27.305 63.995 27.790 64.205 ;
        RECT 27.980 63.995 28.430 64.205 ;
        RECT 28.600 63.995 28.935 64.205 ;
        RECT 27.305 63.835 27.680 63.995 ;
        RECT 27.285 63.665 27.680 63.835 ;
        RECT 28.600 63.825 28.770 63.995 ;
        RECT 27.305 63.575 27.680 63.665 ;
        RECT 27.850 63.655 28.770 63.825 ;
        RECT 27.850 63.405 28.020 63.655 ;
        RECT 26.455 63.235 28.020 63.405 ;
        RECT 26.875 62.815 27.680 63.235 ;
        RECT 28.190 62.645 28.520 63.485 ;
        RECT 29.105 63.405 29.355 64.375 ;
        RECT 29.995 63.955 30.330 64.225 ;
        RECT 30.500 63.835 30.670 64.395 ;
        RECT 31.885 64.375 32.095 65.195 ;
        RECT 32.265 64.395 32.595 65.025 ;
        RECT 30.840 63.955 31.175 64.205 ;
        RECT 30.500 63.795 30.675 63.835 ;
        RECT 28.690 62.815 29.355 63.405 ;
        RECT 29.985 62.645 30.265 63.785 ;
        RECT 30.435 62.815 30.765 63.795 ;
        RECT 30.935 62.645 31.195 63.785 ;
        RECT 31.365 62.645 31.655 63.810 ;
        RECT 32.265 63.795 32.515 64.395 ;
        RECT 32.765 64.375 32.995 65.195 ;
        RECT 33.255 64.540 33.585 64.975 ;
        RECT 33.755 64.585 33.925 65.195 ;
        RECT 33.205 64.455 33.585 64.540 ;
        RECT 34.095 64.455 34.425 64.980 ;
        RECT 34.685 64.665 34.895 65.195 ;
        RECT 35.170 64.745 35.955 64.915 ;
        RECT 36.125 64.745 36.530 64.915 ;
        RECT 33.205 64.415 33.430 64.455 ;
        RECT 32.685 63.955 33.015 64.205 ;
        RECT 33.205 63.835 33.375 64.415 ;
        RECT 34.095 64.285 34.295 64.455 ;
        RECT 35.170 64.285 35.340 64.745 ;
        RECT 33.545 63.955 34.295 64.285 ;
        RECT 34.465 63.955 35.340 64.285 ;
        RECT 31.885 62.645 32.095 63.785 ;
        RECT 32.265 62.815 32.595 63.795 ;
        RECT 33.205 63.785 33.420 63.835 ;
        RECT 32.765 62.645 32.995 63.785 ;
        RECT 33.205 63.705 33.595 63.785 ;
        RECT 33.265 62.860 33.595 63.705 ;
        RECT 34.105 63.750 34.295 63.955 ;
        RECT 33.765 62.645 33.935 63.655 ;
        RECT 34.105 63.375 35.000 63.750 ;
        RECT 34.105 62.815 34.445 63.375 ;
        RECT 34.675 62.645 34.990 63.145 ;
        RECT 35.170 63.115 35.340 63.955 ;
        RECT 35.510 64.245 35.975 64.575 ;
        RECT 36.360 64.515 36.530 64.745 ;
        RECT 36.710 64.695 37.080 65.195 ;
        RECT 37.400 64.745 38.075 64.915 ;
        RECT 38.270 64.745 38.605 64.915 ;
        RECT 35.510 63.285 35.830 64.245 ;
        RECT 36.360 64.215 37.190 64.515 ;
        RECT 36.000 63.315 36.190 64.035 ;
        RECT 36.360 63.145 36.530 64.215 ;
        RECT 36.990 64.185 37.190 64.215 ;
        RECT 36.700 63.965 36.870 64.035 ;
        RECT 37.400 63.965 37.570 64.745 ;
        RECT 38.435 64.605 38.605 64.745 ;
        RECT 38.775 64.735 39.025 65.195 ;
        RECT 36.700 63.795 37.570 63.965 ;
        RECT 37.740 64.325 38.265 64.545 ;
        RECT 38.435 64.475 38.660 64.605 ;
        RECT 36.700 63.705 37.210 63.795 ;
        RECT 35.170 62.945 36.055 63.115 ;
        RECT 36.280 62.815 36.530 63.145 ;
        RECT 36.700 62.645 36.870 63.445 ;
        RECT 37.040 63.090 37.210 63.705 ;
        RECT 37.740 63.625 37.910 64.325 ;
        RECT 37.380 63.260 37.910 63.625 ;
        RECT 38.080 63.560 38.320 64.155 ;
        RECT 38.490 63.370 38.660 64.475 ;
        RECT 38.830 63.615 39.110 64.565 ;
        RECT 38.355 63.240 38.660 63.370 ;
        RECT 37.040 62.920 38.145 63.090 ;
        RECT 38.355 62.815 38.605 63.240 ;
        RECT 38.775 62.645 39.040 63.105 ;
        RECT 39.280 62.815 39.465 64.935 ;
        RECT 39.635 64.815 39.965 65.195 ;
        RECT 40.135 64.645 40.305 64.935 ;
        RECT 39.640 64.475 40.305 64.645 ;
        RECT 39.640 63.485 39.870 64.475 ;
        RECT 40.585 64.465 40.915 65.195 ;
        RECT 40.040 63.655 40.390 64.305 ;
        RECT 41.085 64.285 41.295 64.905 ;
        RECT 41.475 64.485 41.905 65.015 ;
        RECT 40.600 63.935 40.890 64.285 ;
        RECT 41.085 63.935 41.480 64.285 ;
        RECT 41.660 64.235 41.905 64.485 ;
        RECT 42.085 64.415 42.315 65.195 ;
        RECT 42.495 64.565 42.875 65.015 ;
        RECT 41.660 63.935 42.195 64.235 ;
        RECT 42.495 64.115 42.725 64.565 ;
        RECT 43.330 64.455 43.585 65.025 ;
        RECT 43.755 64.795 44.085 65.195 ;
        RECT 44.510 64.660 45.040 65.025 ;
        RECT 44.510 64.625 44.685 64.660 ;
        RECT 43.755 64.455 44.685 64.625 ;
        RECT 40.655 63.555 41.695 63.755 ;
        RECT 39.640 63.315 40.305 63.485 ;
        RECT 39.635 62.645 39.965 63.145 ;
        RECT 40.135 62.815 40.305 63.315 ;
        RECT 40.655 62.825 40.825 63.555 ;
        RECT 41.005 62.645 41.335 63.375 ;
        RECT 41.505 62.825 41.695 63.555 ;
        RECT 41.865 62.825 42.195 63.935 ;
        RECT 42.385 63.435 42.725 64.115 ;
        RECT 42.905 63.615 43.135 64.305 ;
        RECT 43.330 63.785 43.500 64.455 ;
        RECT 43.755 64.285 43.925 64.455 ;
        RECT 43.670 63.955 43.925 64.285 ;
        RECT 44.150 63.955 44.345 64.285 ;
        RECT 42.385 63.235 43.145 63.435 ;
        RECT 42.385 62.645 42.715 63.055 ;
        RECT 42.885 62.845 43.145 63.235 ;
        RECT 43.330 62.815 43.665 63.785 ;
        RECT 43.835 62.645 44.005 63.785 ;
        RECT 44.175 62.985 44.345 63.955 ;
        RECT 44.515 63.325 44.685 64.455 ;
        RECT 44.855 63.665 45.025 64.465 ;
        RECT 45.230 64.175 45.505 65.025 ;
        RECT 45.225 64.005 45.505 64.175 ;
        RECT 45.230 63.865 45.505 64.005 ;
        RECT 45.675 63.665 45.865 65.025 ;
        RECT 46.045 64.660 46.555 65.195 ;
        RECT 46.775 64.385 47.020 64.990 ;
        RECT 47.465 64.455 47.850 65.025 ;
        RECT 48.020 64.735 48.345 65.195 ;
        RECT 48.865 64.565 49.145 65.025 ;
        RECT 46.065 64.215 47.295 64.385 ;
        RECT 44.855 63.495 45.865 63.665 ;
        RECT 46.035 63.650 46.785 63.840 ;
        RECT 44.515 63.155 45.640 63.325 ;
        RECT 46.035 62.985 46.205 63.650 ;
        RECT 46.955 63.405 47.295 64.215 ;
        RECT 44.175 62.815 46.205 62.985 ;
        RECT 46.375 62.645 46.545 63.405 ;
        RECT 46.780 62.995 47.295 63.405 ;
        RECT 47.465 63.785 47.745 64.455 ;
        RECT 48.020 64.395 49.145 64.565 ;
        RECT 48.020 64.285 48.470 64.395 ;
        RECT 47.915 63.955 48.470 64.285 ;
        RECT 49.335 64.225 49.735 65.025 ;
        RECT 50.135 64.735 50.405 65.195 ;
        RECT 50.575 64.565 50.860 65.025 ;
        RECT 47.465 62.815 47.850 63.785 ;
        RECT 48.020 63.495 48.470 63.955 ;
        RECT 48.640 63.665 49.735 64.225 ;
        RECT 48.020 63.275 49.145 63.495 ;
        RECT 48.020 62.645 48.345 63.105 ;
        RECT 48.865 62.815 49.145 63.275 ;
        RECT 49.335 62.815 49.735 63.665 ;
        RECT 49.905 64.395 50.860 64.565 ;
        RECT 52.070 64.455 52.325 65.025 ;
        RECT 52.495 64.795 52.825 65.195 ;
        RECT 53.250 64.660 53.780 65.025 ;
        RECT 53.250 64.625 53.425 64.660 ;
        RECT 52.495 64.455 53.425 64.625 ;
        RECT 53.970 64.515 54.245 65.025 ;
        RECT 49.905 63.495 50.115 64.395 ;
        RECT 50.285 63.665 50.975 64.225 ;
        RECT 52.070 63.785 52.240 64.455 ;
        RECT 52.495 64.285 52.665 64.455 ;
        RECT 52.410 63.955 52.665 64.285 ;
        RECT 52.890 63.955 53.085 64.285 ;
        RECT 49.905 63.275 50.860 63.495 ;
        RECT 50.135 62.645 50.405 63.105 ;
        RECT 50.575 62.815 50.860 63.275 ;
        RECT 52.070 62.815 52.405 63.785 ;
        RECT 52.575 62.645 52.745 63.785 ;
        RECT 52.915 62.985 53.085 63.955 ;
        RECT 53.255 63.325 53.425 64.455 ;
        RECT 53.595 63.665 53.765 64.465 ;
        RECT 53.965 64.345 54.245 64.515 ;
        RECT 53.970 63.865 54.245 64.345 ;
        RECT 54.415 63.665 54.605 65.025 ;
        RECT 54.785 64.660 55.295 65.195 ;
        RECT 55.515 64.385 55.760 64.990 ;
        RECT 57.125 64.470 57.415 65.195 ;
        RECT 57.590 64.455 57.845 65.025 ;
        RECT 58.015 64.795 58.345 65.195 ;
        RECT 58.770 64.660 59.300 65.025 ;
        RECT 59.490 64.855 59.765 65.025 ;
        RECT 59.485 64.685 59.765 64.855 ;
        RECT 58.770 64.625 58.945 64.660 ;
        RECT 58.015 64.455 58.945 64.625 ;
        RECT 54.805 64.215 56.035 64.385 ;
        RECT 53.595 63.495 54.605 63.665 ;
        RECT 54.775 63.650 55.525 63.840 ;
        RECT 53.255 63.155 54.380 63.325 ;
        RECT 54.775 62.985 54.945 63.650 ;
        RECT 55.695 63.405 56.035 64.215 ;
        RECT 52.915 62.815 54.945 62.985 ;
        RECT 55.115 62.645 55.285 63.405 ;
        RECT 55.520 62.995 56.035 63.405 ;
        RECT 57.125 62.645 57.415 63.810 ;
        RECT 57.590 63.785 57.760 64.455 ;
        RECT 58.015 64.285 58.185 64.455 ;
        RECT 57.930 63.955 58.185 64.285 ;
        RECT 58.410 63.955 58.605 64.285 ;
        RECT 57.590 62.815 57.925 63.785 ;
        RECT 58.095 62.645 58.265 63.785 ;
        RECT 58.435 62.985 58.605 63.955 ;
        RECT 58.775 63.325 58.945 64.455 ;
        RECT 59.115 63.665 59.285 64.465 ;
        RECT 59.490 63.865 59.765 64.685 ;
        RECT 59.935 63.665 60.125 65.025 ;
        RECT 60.305 64.660 60.815 65.195 ;
        RECT 61.035 64.385 61.280 64.990 ;
        RECT 62.190 64.455 62.445 65.025 ;
        RECT 62.615 64.795 62.945 65.195 ;
        RECT 63.370 64.660 63.900 65.025 ;
        RECT 64.090 64.855 64.365 65.025 ;
        RECT 64.085 64.685 64.365 64.855 ;
        RECT 63.370 64.625 63.545 64.660 ;
        RECT 62.615 64.455 63.545 64.625 ;
        RECT 60.325 64.215 61.555 64.385 ;
        RECT 59.115 63.495 60.125 63.665 ;
        RECT 60.295 63.650 61.045 63.840 ;
        RECT 58.775 63.155 59.900 63.325 ;
        RECT 60.295 62.985 60.465 63.650 ;
        RECT 61.215 63.405 61.555 64.215 ;
        RECT 58.435 62.815 60.465 62.985 ;
        RECT 60.635 62.645 60.805 63.405 ;
        RECT 61.040 62.995 61.555 63.405 ;
        RECT 62.190 63.785 62.360 64.455 ;
        RECT 62.615 64.285 62.785 64.455 ;
        RECT 62.530 63.955 62.785 64.285 ;
        RECT 63.010 63.955 63.205 64.285 ;
        RECT 62.190 62.815 62.525 63.785 ;
        RECT 62.695 62.645 62.865 63.785 ;
        RECT 63.035 62.985 63.205 63.955 ;
        RECT 63.375 63.325 63.545 64.455 ;
        RECT 63.715 63.665 63.885 64.465 ;
        RECT 64.090 63.865 64.365 64.685 ;
        RECT 64.535 63.665 64.725 65.025 ;
        RECT 64.905 64.660 65.415 65.195 ;
        RECT 65.635 64.385 65.880 64.990 ;
        RECT 66.330 64.455 66.585 65.025 ;
        RECT 66.755 64.795 67.085 65.195 ;
        RECT 67.510 64.660 68.040 65.025 ;
        RECT 68.230 64.855 68.505 65.025 ;
        RECT 68.225 64.685 68.505 64.855 ;
        RECT 67.510 64.625 67.685 64.660 ;
        RECT 66.755 64.455 67.685 64.625 ;
        RECT 64.925 64.215 66.155 64.385 ;
        RECT 63.715 63.495 64.725 63.665 ;
        RECT 64.895 63.650 65.645 63.840 ;
        RECT 63.375 63.155 64.500 63.325 ;
        RECT 64.895 62.985 65.065 63.650 ;
        RECT 65.815 63.405 66.155 64.215 ;
        RECT 63.035 62.815 65.065 62.985 ;
        RECT 65.235 62.645 65.405 63.405 ;
        RECT 65.640 62.995 66.155 63.405 ;
        RECT 66.330 63.785 66.500 64.455 ;
        RECT 66.755 64.285 66.925 64.455 ;
        RECT 66.670 63.955 66.925 64.285 ;
        RECT 67.150 63.955 67.345 64.285 ;
        RECT 66.330 62.815 66.665 63.785 ;
        RECT 66.835 62.645 67.005 63.785 ;
        RECT 67.175 62.985 67.345 63.955 ;
        RECT 67.515 63.325 67.685 64.455 ;
        RECT 67.855 63.665 68.025 64.465 ;
        RECT 68.230 63.865 68.505 64.685 ;
        RECT 68.675 63.665 68.865 65.025 ;
        RECT 69.045 64.660 69.555 65.195 ;
        RECT 69.775 64.385 70.020 64.990 ;
        RECT 70.465 64.455 70.850 65.025 ;
        RECT 71.020 64.735 71.345 65.195 ;
        RECT 71.865 64.565 72.145 65.025 ;
        RECT 69.065 64.215 70.295 64.385 ;
        RECT 67.855 63.495 68.865 63.665 ;
        RECT 69.035 63.650 69.785 63.840 ;
        RECT 67.515 63.155 68.640 63.325 ;
        RECT 69.035 62.985 69.205 63.650 ;
        RECT 69.955 63.405 70.295 64.215 ;
        RECT 67.175 62.815 69.205 62.985 ;
        RECT 69.375 62.645 69.545 63.405 ;
        RECT 69.780 62.995 70.295 63.405 ;
        RECT 70.465 63.785 70.745 64.455 ;
        RECT 71.020 64.395 72.145 64.565 ;
        RECT 71.020 64.285 71.470 64.395 ;
        RECT 70.915 63.955 71.470 64.285 ;
        RECT 72.335 64.225 72.735 65.025 ;
        RECT 73.135 64.735 73.405 65.195 ;
        RECT 73.575 64.565 73.860 65.025 ;
        RECT 74.255 64.815 75.425 65.025 ;
        RECT 74.255 64.795 74.585 64.815 ;
        RECT 70.465 62.815 70.850 63.785 ;
        RECT 71.020 63.495 71.470 63.955 ;
        RECT 71.640 63.665 72.735 64.225 ;
        RECT 71.020 63.275 72.145 63.495 ;
        RECT 71.020 62.645 71.345 63.105 ;
        RECT 71.865 62.815 72.145 63.275 ;
        RECT 72.335 62.815 72.735 63.665 ;
        RECT 72.905 64.395 73.860 64.565 ;
        RECT 72.905 63.495 73.115 64.395 ;
        RECT 74.145 64.375 75.005 64.625 ;
        RECT 75.175 64.565 75.425 64.815 ;
        RECT 75.595 64.735 75.765 65.195 ;
        RECT 75.935 64.565 76.275 65.025 ;
        RECT 75.175 64.395 76.275 64.565 ;
        RECT 76.535 64.645 76.705 65.025 ;
        RECT 76.885 64.815 77.215 65.195 ;
        RECT 76.535 64.475 77.200 64.645 ;
        RECT 77.395 64.520 77.655 65.025 ;
        RECT 73.285 63.665 73.975 64.225 ;
        RECT 74.145 63.785 74.425 64.375 ;
        RECT 74.595 63.955 75.345 64.205 ;
        RECT 75.515 63.955 76.275 64.205 ;
        RECT 76.465 63.925 76.795 64.295 ;
        RECT 77.030 64.220 77.200 64.475 ;
        RECT 77.030 63.890 77.315 64.220 ;
        RECT 74.145 63.615 75.845 63.785 ;
        RECT 72.905 63.275 73.860 63.495 ;
        RECT 73.135 62.645 73.405 63.105 ;
        RECT 73.575 62.815 73.860 63.275 ;
        RECT 74.250 62.645 74.505 63.445 ;
        RECT 74.675 62.815 75.005 63.615 ;
        RECT 75.175 62.645 75.345 63.445 ;
        RECT 75.515 62.815 75.845 63.615 ;
        RECT 76.015 62.645 76.275 63.785 ;
        RECT 77.030 63.745 77.200 63.890 ;
        RECT 76.535 63.575 77.200 63.745 ;
        RECT 77.485 63.720 77.655 64.520 ;
        RECT 77.830 64.430 78.285 65.195 ;
        RECT 78.560 64.815 79.860 65.025 ;
        RECT 80.115 64.835 80.445 65.195 ;
        RECT 79.690 64.665 79.860 64.815 ;
        RECT 80.615 64.695 80.875 65.025 ;
        RECT 78.760 64.205 78.980 64.605 ;
        RECT 77.825 64.005 78.315 64.205 ;
        RECT 78.505 63.995 78.980 64.205 ;
        RECT 79.225 64.205 79.435 64.605 ;
        RECT 79.690 64.540 80.445 64.665 ;
        RECT 79.690 64.495 80.535 64.540 ;
        RECT 80.265 64.375 80.535 64.495 ;
        RECT 79.225 63.995 79.555 64.205 ;
        RECT 79.725 63.935 80.135 64.240 ;
        RECT 76.535 62.815 76.705 63.575 ;
        RECT 76.885 62.645 77.215 63.405 ;
        RECT 77.385 62.815 77.655 63.720 ;
        RECT 77.830 63.765 79.005 63.825 ;
        RECT 80.365 63.800 80.535 64.375 ;
        RECT 80.335 63.765 80.535 63.800 ;
        RECT 77.830 63.655 80.535 63.765 ;
        RECT 77.830 63.035 78.085 63.655 ;
        RECT 78.675 63.595 80.475 63.655 ;
        RECT 78.675 63.565 79.005 63.595 ;
        RECT 80.705 63.495 80.875 64.695 ;
        RECT 81.965 64.445 83.175 65.195 ;
        RECT 78.335 63.395 78.520 63.485 ;
        RECT 79.110 63.395 79.945 63.405 ;
        RECT 78.335 63.195 79.945 63.395 ;
        RECT 78.335 63.155 78.565 63.195 ;
        RECT 77.830 62.815 78.165 63.035 ;
        RECT 79.170 62.645 79.525 63.025 ;
        RECT 79.695 62.815 79.945 63.195 ;
        RECT 80.195 62.645 80.445 63.425 ;
        RECT 80.615 62.815 80.875 63.495 ;
        RECT 81.965 63.735 82.485 64.275 ;
        RECT 82.655 63.905 83.175 64.445 ;
        RECT 81.965 62.645 83.175 63.735 ;
        RECT 5.520 62.475 83.260 62.645 ;
        RECT 5.605 61.385 6.815 62.475 ;
        RECT 5.605 60.675 6.125 61.215 ;
        RECT 6.295 60.845 6.815 61.385 ;
        RECT 7.455 61.525 7.730 62.295 ;
        RECT 7.900 61.865 8.230 62.295 ;
        RECT 8.400 62.035 8.595 62.475 ;
        RECT 8.775 61.865 9.105 62.295 ;
        RECT 7.900 61.695 9.105 61.865 ;
        RECT 9.285 61.920 9.890 62.475 ;
        RECT 10.065 61.965 10.545 62.305 ;
        RECT 10.715 61.930 10.970 62.475 ;
        RECT 9.285 61.820 9.900 61.920 ;
        RECT 7.455 61.335 8.040 61.525 ;
        RECT 8.210 61.365 9.105 61.695 ;
        RECT 9.715 61.795 9.900 61.820 ;
        RECT 5.605 59.925 6.815 60.675 ;
        RECT 7.455 60.515 7.695 61.165 ;
        RECT 7.865 60.665 8.040 61.335 ;
        RECT 9.285 61.200 9.545 61.650 ;
        RECT 9.715 61.550 10.045 61.795 ;
        RECT 10.215 61.475 10.970 61.725 ;
        RECT 11.140 61.605 11.415 62.305 ;
        RECT 10.200 61.440 10.970 61.475 ;
        RECT 10.185 61.430 10.970 61.440 ;
        RECT 10.180 61.415 11.075 61.430 ;
        RECT 10.160 61.400 11.075 61.415 ;
        RECT 10.140 61.390 11.075 61.400 ;
        RECT 10.115 61.380 11.075 61.390 ;
        RECT 10.045 61.350 11.075 61.380 ;
        RECT 10.025 61.320 11.075 61.350 ;
        RECT 10.005 61.290 11.075 61.320 ;
        RECT 9.975 61.265 11.075 61.290 ;
        RECT 9.940 61.230 11.075 61.265 ;
        RECT 9.910 61.225 11.075 61.230 ;
        RECT 9.910 61.220 10.300 61.225 ;
        RECT 9.910 61.210 10.275 61.220 ;
        RECT 9.910 61.205 10.260 61.210 ;
        RECT 9.910 61.200 10.245 61.205 ;
        RECT 9.285 61.195 10.245 61.200 ;
        RECT 9.285 61.185 10.235 61.195 ;
        RECT 9.285 61.180 10.225 61.185 ;
        RECT 9.285 61.170 10.215 61.180 ;
        RECT 8.210 60.835 8.625 61.165 ;
        RECT 8.805 60.835 9.100 61.165 ;
        RECT 9.285 61.160 10.210 61.170 ;
        RECT 9.285 61.155 10.205 61.160 ;
        RECT 9.285 61.140 10.195 61.155 ;
        RECT 9.285 61.125 10.190 61.140 ;
        RECT 9.285 61.100 10.180 61.125 ;
        RECT 9.285 61.030 10.175 61.100 ;
        RECT 7.865 60.485 8.195 60.665 ;
        RECT 7.470 59.925 7.800 60.315 ;
        RECT 7.970 60.105 8.195 60.485 ;
        RECT 8.395 60.215 8.625 60.835 ;
        RECT 8.805 59.925 9.105 60.655 ;
        RECT 9.285 60.475 9.835 60.860 ;
        RECT 10.005 60.305 10.175 61.030 ;
        RECT 9.285 60.135 10.175 60.305 ;
        RECT 10.345 60.630 10.675 61.055 ;
        RECT 10.845 60.830 11.075 61.225 ;
        RECT 10.345 60.145 10.565 60.630 ;
        RECT 11.245 60.575 11.415 61.605 ;
        RECT 10.735 59.925 10.985 60.465 ;
        RECT 11.155 60.095 11.415 60.575 ;
        RECT 11.585 62.045 11.925 62.305 ;
        RECT 11.585 60.645 11.845 62.045 ;
        RECT 12.095 61.675 12.425 62.475 ;
        RECT 12.890 61.505 13.140 62.305 ;
        RECT 13.325 61.755 13.655 62.475 ;
        RECT 13.875 61.505 14.125 62.305 ;
        RECT 14.295 62.095 14.630 62.475 ;
        RECT 12.035 61.335 14.225 61.505 ;
        RECT 12.035 61.165 12.350 61.335 ;
        RECT 12.020 60.915 12.350 61.165 ;
        RECT 11.585 60.135 11.925 60.645 ;
        RECT 12.095 59.925 12.365 60.725 ;
        RECT 12.545 60.195 12.825 61.165 ;
        RECT 13.005 60.195 13.305 61.165 ;
        RECT 13.485 60.200 13.835 61.165 ;
        RECT 14.055 60.425 14.225 61.335 ;
        RECT 14.395 60.605 14.635 61.915 ;
        RECT 15.725 60.870 16.005 62.305 ;
        RECT 16.175 61.700 16.885 62.475 ;
        RECT 17.055 61.530 17.385 62.305 ;
        RECT 16.235 61.315 17.385 61.530 ;
        RECT 14.055 60.095 14.550 60.425 ;
        RECT 15.725 60.095 16.065 60.870 ;
        RECT 16.235 60.745 16.520 61.315 ;
        RECT 16.705 60.915 17.175 61.145 ;
        RECT 17.580 61.115 17.795 62.230 ;
        RECT 17.975 61.755 18.305 62.475 ;
        RECT 18.085 61.115 18.315 61.455 ;
        RECT 18.485 61.310 18.775 62.475 ;
        RECT 18.945 61.385 20.615 62.475 ;
        RECT 20.790 62.095 21.125 62.475 ;
        RECT 17.345 60.935 17.795 61.115 ;
        RECT 17.345 60.915 17.675 60.935 ;
        RECT 17.985 60.915 18.315 61.115 ;
        RECT 16.235 60.555 16.945 60.745 ;
        RECT 16.645 60.415 16.945 60.555 ;
        RECT 17.135 60.555 18.315 60.745 ;
        RECT 18.945 60.695 19.695 61.215 ;
        RECT 19.865 60.865 20.615 61.385 ;
        RECT 17.135 60.475 17.465 60.555 ;
        RECT 16.645 60.405 16.960 60.415 ;
        RECT 16.645 60.395 16.970 60.405 ;
        RECT 16.645 60.390 16.980 60.395 ;
        RECT 16.235 59.925 16.405 60.385 ;
        RECT 16.645 60.380 16.985 60.390 ;
        RECT 16.645 60.375 16.990 60.380 ;
        RECT 16.645 60.365 16.995 60.375 ;
        RECT 16.645 60.360 17.000 60.365 ;
        RECT 16.645 60.095 17.005 60.360 ;
        RECT 17.635 59.925 17.805 60.385 ;
        RECT 17.975 60.095 18.315 60.555 ;
        RECT 18.485 59.925 18.775 60.650 ;
        RECT 18.945 59.925 20.615 60.695 ;
        RECT 20.785 60.605 21.025 61.915 ;
        RECT 21.295 61.505 21.545 62.305 ;
        RECT 21.765 61.755 22.095 62.475 ;
        RECT 22.280 61.505 22.530 62.305 ;
        RECT 22.995 61.675 23.325 62.475 ;
        RECT 23.495 62.045 23.835 62.305 ;
        RECT 21.195 61.335 23.385 61.505 ;
        RECT 21.195 60.425 21.365 61.335 ;
        RECT 23.070 61.165 23.385 61.335 ;
        RECT 20.870 60.095 21.365 60.425 ;
        RECT 21.585 60.200 21.935 61.165 ;
        RECT 22.115 60.195 22.415 61.165 ;
        RECT 22.595 60.195 22.875 61.165 ;
        RECT 23.070 60.915 23.400 61.165 ;
        RECT 23.055 59.925 23.325 60.725 ;
        RECT 23.575 60.645 23.835 62.045 ;
        RECT 24.095 61.805 24.265 62.305 ;
        RECT 24.435 61.975 24.765 62.475 ;
        RECT 24.095 61.635 24.760 61.805 ;
        RECT 24.010 60.815 24.360 61.465 ;
        RECT 24.530 60.645 24.760 61.635 ;
        RECT 23.495 60.135 23.835 60.645 ;
        RECT 24.095 60.475 24.760 60.645 ;
        RECT 24.095 60.185 24.265 60.475 ;
        RECT 24.435 59.925 24.765 60.305 ;
        RECT 24.935 60.185 25.120 62.305 ;
        RECT 25.360 62.015 25.625 62.475 ;
        RECT 25.795 61.880 26.045 62.305 ;
        RECT 26.255 62.030 27.360 62.200 ;
        RECT 25.740 61.750 26.045 61.880 ;
        RECT 25.290 60.555 25.570 61.505 ;
        RECT 25.740 60.645 25.910 61.750 ;
        RECT 26.080 60.965 26.320 61.560 ;
        RECT 26.490 61.495 27.020 61.860 ;
        RECT 26.490 60.795 26.660 61.495 ;
        RECT 27.190 61.415 27.360 62.030 ;
        RECT 27.530 61.675 27.700 62.475 ;
        RECT 27.870 61.975 28.120 62.305 ;
        RECT 28.345 62.005 29.230 62.175 ;
        RECT 27.190 61.325 27.700 61.415 ;
        RECT 25.740 60.515 25.965 60.645 ;
        RECT 26.135 60.575 26.660 60.795 ;
        RECT 26.830 61.155 27.700 61.325 ;
        RECT 25.375 59.925 25.625 60.385 ;
        RECT 25.795 60.375 25.965 60.515 ;
        RECT 26.830 60.375 27.000 61.155 ;
        RECT 27.530 61.085 27.700 61.155 ;
        RECT 27.210 60.905 27.410 60.935 ;
        RECT 27.870 60.905 28.040 61.975 ;
        RECT 28.210 61.085 28.400 61.805 ;
        RECT 27.210 60.605 28.040 60.905 ;
        RECT 28.570 60.875 28.890 61.835 ;
        RECT 25.795 60.205 26.130 60.375 ;
        RECT 26.325 60.205 27.000 60.375 ;
        RECT 27.320 59.925 27.690 60.425 ;
        RECT 27.870 60.375 28.040 60.605 ;
        RECT 28.425 60.545 28.890 60.875 ;
        RECT 29.060 61.165 29.230 62.005 ;
        RECT 29.410 61.975 29.725 62.475 ;
        RECT 29.955 61.745 30.295 62.305 ;
        RECT 29.400 61.370 30.295 61.745 ;
        RECT 30.465 61.465 30.635 62.475 ;
        RECT 30.105 61.165 30.295 61.370 ;
        RECT 30.805 61.415 31.135 62.260 ;
        RECT 30.805 61.335 31.195 61.415 ;
        RECT 30.980 61.285 31.195 61.335 ;
        RECT 29.060 60.835 29.935 61.165 ;
        RECT 30.105 60.835 30.855 61.165 ;
        RECT 29.060 60.375 29.230 60.835 ;
        RECT 30.105 60.665 30.305 60.835 ;
        RECT 31.025 60.705 31.195 61.285 ;
        RECT 30.970 60.665 31.195 60.705 ;
        RECT 27.870 60.205 28.275 60.375 ;
        RECT 28.445 60.205 29.230 60.375 ;
        RECT 29.505 59.925 29.715 60.455 ;
        RECT 29.975 60.140 30.305 60.665 ;
        RECT 30.815 60.580 31.195 60.665 ;
        RECT 30.475 59.925 30.645 60.535 ;
        RECT 30.815 60.145 31.145 60.580 ;
        RECT 31.375 60.105 31.635 62.295 ;
        RECT 31.805 61.745 32.145 62.475 ;
        RECT 32.325 61.565 32.595 62.295 ;
        RECT 31.825 61.345 32.595 61.565 ;
        RECT 32.775 61.585 33.005 62.295 ;
        RECT 33.175 61.765 33.505 62.475 ;
        RECT 33.675 61.585 33.935 62.295 ;
        RECT 34.215 61.805 34.385 62.305 ;
        RECT 34.555 61.975 34.885 62.475 ;
        RECT 34.215 61.635 34.880 61.805 ;
        RECT 32.775 61.345 33.935 61.585 ;
        RECT 31.825 60.675 32.115 61.345 ;
        RECT 32.295 60.855 32.760 61.165 ;
        RECT 32.940 60.855 33.465 61.165 ;
        RECT 31.825 60.475 33.055 60.675 ;
        RECT 31.895 59.925 32.565 60.295 ;
        RECT 32.745 60.105 33.055 60.475 ;
        RECT 33.235 60.215 33.465 60.855 ;
        RECT 33.645 60.835 33.945 61.165 ;
        RECT 34.130 60.815 34.480 61.465 ;
        RECT 33.645 59.925 33.935 60.655 ;
        RECT 34.650 60.645 34.880 61.635 ;
        RECT 34.215 60.475 34.880 60.645 ;
        RECT 34.215 60.185 34.385 60.475 ;
        RECT 34.555 59.925 34.885 60.305 ;
        RECT 35.055 60.185 35.240 62.305 ;
        RECT 35.480 62.015 35.745 62.475 ;
        RECT 35.915 61.880 36.165 62.305 ;
        RECT 36.375 62.030 37.480 62.200 ;
        RECT 35.860 61.750 36.165 61.880 ;
        RECT 35.410 60.555 35.690 61.505 ;
        RECT 35.860 60.645 36.030 61.750 ;
        RECT 36.200 60.965 36.440 61.560 ;
        RECT 36.610 61.495 37.140 61.860 ;
        RECT 36.610 60.795 36.780 61.495 ;
        RECT 37.310 61.415 37.480 62.030 ;
        RECT 37.650 61.675 37.820 62.475 ;
        RECT 37.990 61.975 38.240 62.305 ;
        RECT 38.465 62.005 39.350 62.175 ;
        RECT 37.310 61.325 37.820 61.415 ;
        RECT 35.860 60.515 36.085 60.645 ;
        RECT 36.255 60.575 36.780 60.795 ;
        RECT 36.950 61.155 37.820 61.325 ;
        RECT 35.495 59.925 35.745 60.385 ;
        RECT 35.915 60.375 36.085 60.515 ;
        RECT 36.950 60.375 37.120 61.155 ;
        RECT 37.650 61.085 37.820 61.155 ;
        RECT 37.330 60.905 37.530 60.935 ;
        RECT 37.990 60.905 38.160 61.975 ;
        RECT 38.330 61.085 38.520 61.805 ;
        RECT 37.330 60.605 38.160 60.905 ;
        RECT 38.690 60.875 39.010 61.835 ;
        RECT 35.915 60.205 36.250 60.375 ;
        RECT 36.445 60.205 37.120 60.375 ;
        RECT 37.440 59.925 37.810 60.425 ;
        RECT 37.990 60.375 38.160 60.605 ;
        RECT 38.545 60.545 39.010 60.875 ;
        RECT 39.180 61.165 39.350 62.005 ;
        RECT 39.530 61.975 39.845 62.475 ;
        RECT 40.075 61.745 40.415 62.305 ;
        RECT 39.520 61.370 40.415 61.745 ;
        RECT 40.585 61.465 40.755 62.475 ;
        RECT 40.225 61.165 40.415 61.370 ;
        RECT 40.925 61.415 41.255 62.260 ;
        RECT 41.670 61.505 42.060 61.680 ;
        RECT 42.545 61.675 42.875 62.475 ;
        RECT 43.045 61.685 43.580 62.305 ;
        RECT 40.925 61.335 41.315 61.415 ;
        RECT 41.670 61.335 43.095 61.505 ;
        RECT 41.100 61.285 41.315 61.335 ;
        RECT 39.180 60.835 40.055 61.165 ;
        RECT 40.225 60.835 40.975 61.165 ;
        RECT 39.180 60.375 39.350 60.835 ;
        RECT 40.225 60.665 40.425 60.835 ;
        RECT 41.145 60.705 41.315 61.285 ;
        RECT 41.090 60.665 41.315 60.705 ;
        RECT 37.990 60.205 38.395 60.375 ;
        RECT 38.565 60.205 39.350 60.375 ;
        RECT 39.625 59.925 39.835 60.455 ;
        RECT 40.095 60.140 40.425 60.665 ;
        RECT 40.935 60.580 41.315 60.665 ;
        RECT 41.545 60.605 41.900 61.165 ;
        RECT 40.595 59.925 40.765 60.535 ;
        RECT 40.935 60.145 41.265 60.580 ;
        RECT 42.070 60.435 42.240 61.335 ;
        RECT 42.410 60.605 42.675 61.165 ;
        RECT 42.925 60.835 43.095 61.335 ;
        RECT 43.265 60.665 43.580 61.685 ;
        RECT 44.245 61.310 44.535 62.475 ;
        RECT 44.765 61.335 44.975 62.475 ;
        RECT 45.145 61.325 45.475 62.305 ;
        RECT 45.645 61.335 45.875 62.475 ;
        RECT 46.090 61.335 46.425 62.305 ;
        RECT 46.595 61.335 46.765 62.475 ;
        RECT 46.935 62.135 48.965 62.305 ;
        RECT 41.650 59.925 41.890 60.435 ;
        RECT 42.070 60.105 42.350 60.435 ;
        RECT 42.580 59.925 42.795 60.435 ;
        RECT 42.965 60.095 43.580 60.665 ;
        RECT 44.245 59.925 44.535 60.650 ;
        RECT 44.765 59.925 44.975 60.745 ;
        RECT 45.145 60.725 45.395 61.325 ;
        RECT 45.565 60.915 45.895 61.165 ;
        RECT 45.145 60.095 45.475 60.725 ;
        RECT 45.645 59.925 45.875 60.745 ;
        RECT 46.090 60.665 46.260 61.335 ;
        RECT 46.935 61.165 47.105 62.135 ;
        RECT 46.430 60.835 46.685 61.165 ;
        RECT 46.910 60.835 47.105 61.165 ;
        RECT 47.275 61.795 48.400 61.965 ;
        RECT 46.515 60.665 46.685 60.835 ;
        RECT 47.275 60.665 47.445 61.795 ;
        RECT 46.090 60.095 46.345 60.665 ;
        RECT 46.515 60.495 47.445 60.665 ;
        RECT 47.615 61.455 48.625 61.625 ;
        RECT 47.615 60.655 47.785 61.455 ;
        RECT 47.990 61.115 48.265 61.255 ;
        RECT 47.985 60.945 48.265 61.115 ;
        RECT 47.270 60.460 47.445 60.495 ;
        RECT 46.515 59.925 46.845 60.325 ;
        RECT 47.270 60.095 47.800 60.460 ;
        RECT 47.990 60.095 48.265 60.945 ;
        RECT 48.435 60.095 48.625 61.455 ;
        RECT 48.795 61.470 48.965 62.135 ;
        RECT 49.135 61.715 49.305 62.475 ;
        RECT 49.540 61.715 50.055 62.125 ;
        RECT 48.795 61.280 49.545 61.470 ;
        RECT 49.715 60.905 50.055 61.715 ;
        RECT 50.285 61.415 50.615 62.260 ;
        RECT 50.785 61.465 50.955 62.475 ;
        RECT 51.125 61.745 51.465 62.305 ;
        RECT 51.695 61.975 52.010 62.475 ;
        RECT 52.190 62.005 53.075 62.175 ;
        RECT 48.825 60.735 50.055 60.905 ;
        RECT 50.225 61.335 50.615 61.415 ;
        RECT 51.125 61.370 52.020 61.745 ;
        RECT 50.225 61.285 50.440 61.335 ;
        RECT 48.805 59.925 49.315 60.460 ;
        RECT 49.535 60.130 49.780 60.735 ;
        RECT 50.225 60.705 50.395 61.285 ;
        RECT 51.125 61.165 51.315 61.370 ;
        RECT 52.190 61.165 52.360 62.005 ;
        RECT 53.300 61.975 53.550 62.305 ;
        RECT 50.565 60.835 51.315 61.165 ;
        RECT 51.485 60.835 52.360 61.165 ;
        RECT 50.225 60.665 50.450 60.705 ;
        RECT 51.115 60.665 51.315 60.835 ;
        RECT 50.225 60.580 50.605 60.665 ;
        RECT 50.275 60.145 50.605 60.580 ;
        RECT 50.775 59.925 50.945 60.535 ;
        RECT 51.115 60.140 51.445 60.665 ;
        RECT 51.705 59.925 51.915 60.455 ;
        RECT 52.190 60.375 52.360 60.835 ;
        RECT 52.530 60.875 52.850 61.835 ;
        RECT 53.020 61.085 53.210 61.805 ;
        RECT 53.380 60.905 53.550 61.975 ;
        RECT 53.720 61.675 53.890 62.475 ;
        RECT 54.060 62.030 55.165 62.200 ;
        RECT 54.060 61.415 54.230 62.030 ;
        RECT 55.375 61.880 55.625 62.305 ;
        RECT 55.795 62.015 56.060 62.475 ;
        RECT 54.400 61.495 54.930 61.860 ;
        RECT 55.375 61.750 55.680 61.880 ;
        RECT 53.720 61.325 54.230 61.415 ;
        RECT 53.720 61.155 54.590 61.325 ;
        RECT 53.720 61.085 53.890 61.155 ;
        RECT 54.010 60.905 54.210 60.935 ;
        RECT 52.530 60.545 52.995 60.875 ;
        RECT 53.380 60.605 54.210 60.905 ;
        RECT 53.380 60.375 53.550 60.605 ;
        RECT 52.190 60.205 52.975 60.375 ;
        RECT 53.145 60.205 53.550 60.375 ;
        RECT 53.730 59.925 54.100 60.425 ;
        RECT 54.420 60.375 54.590 61.155 ;
        RECT 54.760 60.795 54.930 61.495 ;
        RECT 55.100 60.965 55.340 61.560 ;
        RECT 54.760 60.575 55.285 60.795 ;
        RECT 55.510 60.645 55.680 61.750 ;
        RECT 55.455 60.515 55.680 60.645 ;
        RECT 55.850 60.555 56.130 61.505 ;
        RECT 55.455 60.375 55.625 60.515 ;
        RECT 54.420 60.205 55.095 60.375 ;
        RECT 55.290 60.205 55.625 60.375 ;
        RECT 55.795 59.925 56.045 60.385 ;
        RECT 56.300 60.185 56.485 62.305 ;
        RECT 56.655 61.975 56.985 62.475 ;
        RECT 57.155 61.805 57.325 62.305 ;
        RECT 56.660 61.635 57.325 61.805 ;
        RECT 56.660 60.645 56.890 61.635 ;
        RECT 57.060 60.815 57.410 61.465 ;
        RECT 58.050 61.325 58.310 62.475 ;
        RECT 58.485 61.400 58.740 62.305 ;
        RECT 58.910 61.715 59.240 62.475 ;
        RECT 59.455 61.545 59.625 62.305 ;
        RECT 59.975 61.805 60.145 62.305 ;
        RECT 60.315 61.975 60.645 62.475 ;
        RECT 59.975 61.635 60.640 61.805 ;
        RECT 56.660 60.475 57.325 60.645 ;
        RECT 56.655 59.925 56.985 60.305 ;
        RECT 57.155 60.185 57.325 60.475 ;
        RECT 58.050 59.925 58.310 60.765 ;
        RECT 58.485 60.670 58.655 61.400 ;
        RECT 58.910 61.375 59.625 61.545 ;
        RECT 58.910 61.165 59.080 61.375 ;
        RECT 58.825 60.835 59.080 61.165 ;
        RECT 58.485 60.095 58.740 60.670 ;
        RECT 58.910 60.645 59.080 60.835 ;
        RECT 59.360 60.825 59.715 61.195 ;
        RECT 59.890 60.815 60.240 61.465 ;
        RECT 60.410 60.645 60.640 61.635 ;
        RECT 58.910 60.475 59.625 60.645 ;
        RECT 58.910 59.925 59.240 60.305 ;
        RECT 59.455 60.095 59.625 60.475 ;
        RECT 59.975 60.475 60.640 60.645 ;
        RECT 59.975 60.185 60.145 60.475 ;
        RECT 60.315 59.925 60.645 60.305 ;
        RECT 60.815 60.185 61.000 62.305 ;
        RECT 61.240 62.015 61.505 62.475 ;
        RECT 61.675 61.880 61.925 62.305 ;
        RECT 62.135 62.030 63.240 62.200 ;
        RECT 61.620 61.750 61.925 61.880 ;
        RECT 61.170 60.555 61.450 61.505 ;
        RECT 61.620 60.645 61.790 61.750 ;
        RECT 61.960 60.965 62.200 61.560 ;
        RECT 62.370 61.495 62.900 61.860 ;
        RECT 62.370 60.795 62.540 61.495 ;
        RECT 63.070 61.415 63.240 62.030 ;
        RECT 63.410 61.675 63.580 62.475 ;
        RECT 63.750 61.975 64.000 62.305 ;
        RECT 64.225 62.005 65.110 62.175 ;
        RECT 63.070 61.325 63.580 61.415 ;
        RECT 61.620 60.515 61.845 60.645 ;
        RECT 62.015 60.575 62.540 60.795 ;
        RECT 62.710 61.155 63.580 61.325 ;
        RECT 61.255 59.925 61.505 60.385 ;
        RECT 61.675 60.375 61.845 60.515 ;
        RECT 62.710 60.375 62.880 61.155 ;
        RECT 63.410 61.085 63.580 61.155 ;
        RECT 63.090 60.905 63.290 60.935 ;
        RECT 63.750 60.905 63.920 61.975 ;
        RECT 64.090 61.085 64.280 61.805 ;
        RECT 63.090 60.605 63.920 60.905 ;
        RECT 64.450 60.875 64.770 61.835 ;
        RECT 61.675 60.205 62.010 60.375 ;
        RECT 62.205 60.205 62.880 60.375 ;
        RECT 63.200 59.925 63.570 60.425 ;
        RECT 63.750 60.375 63.920 60.605 ;
        RECT 64.305 60.545 64.770 60.875 ;
        RECT 64.940 61.165 65.110 62.005 ;
        RECT 65.290 61.975 65.605 62.475 ;
        RECT 65.835 61.745 66.175 62.305 ;
        RECT 65.280 61.370 66.175 61.745 ;
        RECT 66.345 61.465 66.515 62.475 ;
        RECT 65.985 61.165 66.175 61.370 ;
        RECT 66.685 61.415 67.015 62.260 ;
        RECT 66.685 61.335 67.075 61.415 ;
        RECT 67.255 61.335 67.585 62.475 ;
        RECT 66.860 61.285 67.075 61.335 ;
        RECT 64.940 60.835 65.815 61.165 ;
        RECT 65.985 60.835 66.735 61.165 ;
        RECT 64.940 60.375 65.110 60.835 ;
        RECT 65.985 60.665 66.185 60.835 ;
        RECT 66.905 60.705 67.075 61.285 ;
        RECT 66.850 60.665 67.075 60.705 ;
        RECT 63.750 60.205 64.155 60.375 ;
        RECT 64.325 60.205 65.110 60.375 ;
        RECT 65.385 59.925 65.595 60.455 ;
        RECT 65.855 60.140 66.185 60.665 ;
        RECT 66.695 60.580 67.075 60.665 ;
        RECT 67.245 60.585 67.585 61.165 ;
        RECT 67.755 61.135 68.115 62.305 ;
        RECT 68.315 61.305 68.645 62.475 ;
        RECT 68.845 61.135 69.175 62.305 ;
        RECT 69.375 61.305 69.705 62.475 ;
        RECT 70.005 61.310 70.295 62.475 ;
        RECT 70.475 61.365 70.770 62.475 ;
        RECT 70.950 61.165 71.200 62.300 ;
        RECT 71.370 61.365 71.630 62.475 ;
        RECT 71.800 61.575 72.060 62.300 ;
        RECT 72.230 61.745 72.490 62.475 ;
        RECT 72.660 61.575 72.920 62.300 ;
        RECT 73.090 61.745 73.350 62.475 ;
        RECT 73.520 61.575 73.780 62.300 ;
        RECT 73.950 61.745 74.210 62.475 ;
        RECT 74.380 61.575 74.640 62.300 ;
        RECT 74.810 61.745 75.105 62.475 ;
        RECT 71.800 61.335 75.110 61.575 ;
        RECT 67.755 60.855 69.175 61.135 ;
        RECT 66.355 59.925 66.525 60.535 ;
        RECT 66.695 60.145 67.025 60.580 ;
        RECT 67.755 60.520 68.115 60.855 ;
        RECT 67.255 59.925 67.585 60.415 ;
        RECT 67.755 60.095 68.375 60.520 ;
        RECT 68.835 59.925 69.165 60.615 ;
        RECT 70.005 59.925 70.295 60.650 ;
        RECT 70.465 60.555 70.780 61.165 ;
        RECT 70.950 60.915 73.970 61.165 ;
        RECT 70.525 59.925 70.770 60.385 ;
        RECT 70.950 60.105 71.200 60.915 ;
        RECT 74.140 60.745 75.110 61.335 ;
        RECT 71.800 60.575 75.110 60.745 ;
        RECT 75.525 61.335 75.865 62.305 ;
        RECT 76.035 61.335 76.205 62.475 ;
        RECT 76.475 61.675 76.725 62.475 ;
        RECT 77.370 61.505 77.700 62.305 ;
        RECT 78.000 61.675 78.330 62.475 ;
        RECT 78.500 61.505 78.830 62.305 ;
        RECT 76.395 61.335 78.830 61.505 ;
        RECT 79.390 61.505 79.780 61.680 ;
        RECT 80.265 61.675 80.595 62.475 ;
        RECT 80.765 61.685 81.300 62.305 ;
        RECT 79.390 61.335 80.815 61.505 ;
        RECT 75.525 60.725 75.700 61.335 ;
        RECT 76.395 61.085 76.565 61.335 ;
        RECT 75.870 60.915 76.565 61.085 ;
        RECT 76.740 60.915 77.160 61.115 ;
        RECT 77.330 60.915 77.660 61.115 ;
        RECT 77.830 60.915 78.160 61.115 ;
        RECT 71.370 59.925 71.630 60.450 ;
        RECT 71.800 60.120 72.060 60.575 ;
        RECT 72.230 59.925 72.490 60.405 ;
        RECT 72.660 60.120 72.920 60.575 ;
        RECT 73.090 59.925 73.350 60.405 ;
        RECT 73.520 60.120 73.780 60.575 ;
        RECT 73.950 59.925 74.210 60.405 ;
        RECT 74.380 60.120 74.640 60.575 ;
        RECT 74.810 59.925 75.110 60.405 ;
        RECT 75.525 60.095 75.865 60.725 ;
        RECT 76.035 59.925 76.285 60.725 ;
        RECT 76.475 60.575 77.700 60.745 ;
        RECT 76.475 60.095 76.805 60.575 ;
        RECT 76.975 59.925 77.200 60.385 ;
        RECT 77.370 60.095 77.700 60.575 ;
        RECT 78.330 60.705 78.500 61.335 ;
        RECT 78.685 60.915 79.035 61.165 ;
        RECT 78.330 60.095 78.830 60.705 ;
        RECT 79.265 60.605 79.620 61.165 ;
        RECT 79.790 60.435 79.960 61.335 ;
        RECT 80.130 60.605 80.395 61.165 ;
        RECT 80.645 60.835 80.815 61.335 ;
        RECT 80.985 60.665 81.300 61.685 ;
        RECT 81.965 61.385 83.175 62.475 ;
        RECT 81.965 60.845 82.485 61.385 ;
        RECT 82.655 60.675 83.175 61.215 ;
        RECT 79.370 59.925 79.610 60.435 ;
        RECT 79.790 60.105 80.070 60.435 ;
        RECT 80.300 59.925 80.515 60.435 ;
        RECT 80.685 60.095 81.300 60.665 ;
        RECT 81.965 59.925 83.175 60.675 ;
        RECT 5.520 59.755 83.260 59.925 ;
        RECT 5.605 59.005 6.815 59.755 ;
        RECT 7.035 59.100 7.365 59.535 ;
        RECT 7.535 59.145 7.705 59.755 ;
        RECT 6.985 59.015 7.365 59.100 ;
        RECT 7.875 59.015 8.205 59.540 ;
        RECT 8.465 59.225 8.675 59.755 ;
        RECT 8.950 59.305 9.735 59.475 ;
        RECT 9.905 59.305 10.310 59.475 ;
        RECT 5.605 58.465 6.125 59.005 ;
        RECT 6.985 58.975 7.210 59.015 ;
        RECT 6.295 58.295 6.815 58.835 ;
        RECT 5.605 57.205 6.815 58.295 ;
        RECT 6.985 58.395 7.155 58.975 ;
        RECT 7.875 58.845 8.075 59.015 ;
        RECT 8.950 58.845 9.120 59.305 ;
        RECT 7.325 58.515 8.075 58.845 ;
        RECT 8.245 58.515 9.120 58.845 ;
        RECT 6.985 58.345 7.200 58.395 ;
        RECT 6.985 58.265 7.375 58.345 ;
        RECT 7.045 57.420 7.375 58.265 ;
        RECT 7.885 58.310 8.075 58.515 ;
        RECT 7.545 57.205 7.715 58.215 ;
        RECT 7.885 57.935 8.780 58.310 ;
        RECT 7.885 57.375 8.225 57.935 ;
        RECT 8.455 57.205 8.770 57.705 ;
        RECT 8.950 57.675 9.120 58.515 ;
        RECT 9.290 58.805 9.755 59.135 ;
        RECT 10.140 59.075 10.310 59.305 ;
        RECT 10.490 59.255 10.860 59.755 ;
        RECT 11.180 59.305 11.855 59.475 ;
        RECT 12.050 59.305 12.385 59.475 ;
        RECT 9.290 57.845 9.610 58.805 ;
        RECT 10.140 58.775 10.970 59.075 ;
        RECT 9.780 57.875 9.970 58.595 ;
        RECT 10.140 57.705 10.310 58.775 ;
        RECT 10.770 58.745 10.970 58.775 ;
        RECT 10.480 58.525 10.650 58.595 ;
        RECT 11.180 58.525 11.350 59.305 ;
        RECT 12.215 59.165 12.385 59.305 ;
        RECT 12.555 59.295 12.805 59.755 ;
        RECT 10.480 58.355 11.350 58.525 ;
        RECT 11.520 58.885 12.045 59.105 ;
        RECT 12.215 59.035 12.440 59.165 ;
        RECT 10.480 58.265 10.990 58.355 ;
        RECT 8.950 57.505 9.835 57.675 ;
        RECT 10.060 57.375 10.310 57.705 ;
        RECT 10.480 57.205 10.650 58.005 ;
        RECT 10.820 57.650 10.990 58.265 ;
        RECT 11.520 58.185 11.690 58.885 ;
        RECT 11.160 57.820 11.690 58.185 ;
        RECT 11.860 58.120 12.100 58.715 ;
        RECT 12.270 57.930 12.440 59.035 ;
        RECT 12.610 58.175 12.890 59.125 ;
        RECT 12.135 57.800 12.440 57.930 ;
        RECT 10.820 57.480 11.925 57.650 ;
        RECT 12.135 57.375 12.385 57.800 ;
        RECT 12.555 57.205 12.820 57.665 ;
        RECT 13.060 57.375 13.245 59.495 ;
        RECT 13.415 59.375 13.745 59.755 ;
        RECT 13.915 59.205 14.085 59.495 ;
        RECT 13.420 59.035 14.085 59.205 ;
        RECT 14.345 59.105 14.605 59.585 ;
        RECT 14.775 59.215 15.025 59.755 ;
        RECT 13.420 58.045 13.650 59.035 ;
        RECT 13.820 58.215 14.170 58.865 ;
        RECT 14.345 58.075 14.515 59.105 ;
        RECT 15.195 59.050 15.415 59.535 ;
        RECT 14.685 58.455 14.915 58.850 ;
        RECT 15.085 58.625 15.415 59.050 ;
        RECT 15.585 59.375 16.475 59.545 ;
        RECT 15.585 58.650 15.755 59.375 ;
        RECT 16.645 59.255 16.905 59.585 ;
        RECT 17.115 59.275 17.390 59.755 ;
        RECT 15.925 58.820 16.475 59.205 ;
        RECT 15.585 58.580 16.475 58.650 ;
        RECT 15.580 58.555 16.475 58.580 ;
        RECT 15.570 58.540 16.475 58.555 ;
        RECT 15.565 58.525 16.475 58.540 ;
        RECT 15.555 58.520 16.475 58.525 ;
        RECT 15.550 58.510 16.475 58.520 ;
        RECT 15.545 58.500 16.475 58.510 ;
        RECT 15.535 58.495 16.475 58.500 ;
        RECT 15.525 58.485 16.475 58.495 ;
        RECT 15.515 58.480 16.475 58.485 ;
        RECT 15.515 58.475 15.850 58.480 ;
        RECT 15.500 58.470 15.850 58.475 ;
        RECT 15.485 58.460 15.850 58.470 ;
        RECT 15.460 58.455 15.850 58.460 ;
        RECT 14.685 58.450 15.850 58.455 ;
        RECT 14.685 58.415 15.820 58.450 ;
        RECT 14.685 58.390 15.785 58.415 ;
        RECT 14.685 58.360 15.755 58.390 ;
        RECT 14.685 58.330 15.735 58.360 ;
        RECT 14.685 58.300 15.715 58.330 ;
        RECT 14.685 58.290 15.645 58.300 ;
        RECT 14.685 58.280 15.620 58.290 ;
        RECT 14.685 58.265 15.600 58.280 ;
        RECT 14.685 58.250 15.580 58.265 ;
        RECT 14.790 58.240 15.575 58.250 ;
        RECT 14.790 58.205 15.560 58.240 ;
        RECT 13.420 57.875 14.085 58.045 ;
        RECT 13.415 57.205 13.745 57.705 ;
        RECT 13.915 57.375 14.085 57.875 ;
        RECT 14.345 57.375 14.620 58.075 ;
        RECT 14.790 57.955 15.545 58.205 ;
        RECT 15.715 57.885 16.045 58.130 ;
        RECT 16.215 58.030 16.475 58.480 ;
        RECT 16.645 58.345 16.815 59.255 ;
        RECT 17.600 59.185 17.805 59.585 ;
        RECT 17.975 59.355 18.310 59.755 ;
        RECT 16.985 58.515 17.345 59.095 ;
        RECT 17.600 59.015 18.285 59.185 ;
        RECT 17.525 58.345 17.775 58.845 ;
        RECT 16.645 58.175 17.775 58.345 ;
        RECT 15.860 57.860 16.045 57.885 ;
        RECT 15.860 57.760 16.475 57.860 ;
        RECT 14.790 57.205 15.045 57.750 ;
        RECT 15.215 57.375 15.695 57.715 ;
        RECT 15.870 57.205 16.475 57.760 ;
        RECT 16.645 57.405 16.915 58.175 ;
        RECT 17.945 57.985 18.285 59.015 ;
        RECT 18.945 59.145 19.285 59.560 ;
        RECT 19.455 59.315 19.625 59.755 ;
        RECT 19.795 59.365 21.045 59.545 ;
        RECT 19.795 59.145 20.125 59.365 ;
        RECT 21.315 59.295 21.485 59.755 ;
        RECT 18.945 58.975 20.125 59.145 ;
        RECT 20.295 59.125 20.660 59.195 ;
        RECT 20.295 58.945 21.545 59.125 ;
        RECT 18.945 58.565 19.410 58.765 ;
        RECT 19.585 58.515 19.915 58.765 ;
        RECT 20.085 58.735 20.550 58.765 ;
        RECT 20.085 58.565 20.555 58.735 ;
        RECT 20.085 58.515 20.550 58.565 ;
        RECT 20.745 58.515 21.100 58.765 ;
        RECT 19.585 58.395 19.765 58.515 ;
        RECT 17.085 57.205 17.415 57.985 ;
        RECT 17.620 57.810 18.285 57.985 ;
        RECT 17.620 57.405 17.805 57.810 ;
        RECT 17.975 57.205 18.310 57.630 ;
        RECT 18.945 57.205 19.265 58.385 ;
        RECT 19.435 58.225 19.765 58.395 ;
        RECT 21.270 58.345 21.545 58.945 ;
        RECT 19.435 57.435 19.635 58.225 ;
        RECT 19.935 58.135 21.545 58.345 ;
        RECT 19.935 58.035 20.345 58.135 ;
        RECT 19.960 57.375 20.345 58.035 ;
        RECT 20.740 57.205 21.525 57.965 ;
        RECT 21.715 57.375 21.995 59.475 ;
        RECT 22.185 58.945 22.425 59.755 ;
        RECT 22.595 58.945 22.925 59.585 ;
        RECT 23.095 58.945 23.365 59.755 ;
        RECT 23.545 59.005 24.755 59.755 ;
        RECT 24.925 59.105 25.185 59.585 ;
        RECT 25.355 59.295 25.685 59.755 ;
        RECT 25.875 59.115 26.075 59.535 ;
        RECT 22.165 58.515 22.515 58.765 ;
        RECT 22.685 58.345 22.855 58.945 ;
        RECT 23.025 58.515 23.375 58.765 ;
        RECT 23.545 58.465 24.065 59.005 ;
        RECT 22.175 58.175 22.855 58.345 ;
        RECT 22.175 57.390 22.505 58.175 ;
        RECT 23.035 57.205 23.365 58.345 ;
        RECT 24.235 58.295 24.755 58.835 ;
        RECT 23.545 57.205 24.755 58.295 ;
        RECT 24.925 58.075 25.095 59.105 ;
        RECT 25.265 58.415 25.495 58.845 ;
        RECT 25.665 58.595 26.075 59.115 ;
        RECT 26.245 59.270 27.035 59.535 ;
        RECT 26.245 58.415 26.500 59.270 ;
        RECT 27.215 58.935 27.545 59.355 ;
        RECT 27.715 58.935 27.975 59.755 ;
        RECT 27.215 58.845 27.465 58.935 ;
        RECT 26.670 58.595 27.465 58.845 ;
        RECT 25.265 58.245 27.055 58.415 ;
        RECT 24.925 57.375 25.200 58.075 ;
        RECT 25.370 57.950 26.085 58.245 ;
        RECT 26.305 57.885 26.635 58.075 ;
        RECT 25.410 57.205 25.625 57.750 ;
        RECT 25.795 57.375 26.270 57.715 ;
        RECT 26.440 57.710 26.635 57.885 ;
        RECT 26.805 57.880 27.055 58.245 ;
        RECT 26.440 57.205 27.055 57.710 ;
        RECT 27.295 57.375 27.465 58.595 ;
        RECT 27.635 57.885 27.975 58.765 ;
        RECT 27.715 57.205 27.975 57.715 ;
        RECT 28.155 57.385 28.415 59.575 ;
        RECT 28.675 59.385 29.345 59.755 ;
        RECT 29.525 59.205 29.835 59.575 ;
        RECT 28.605 59.005 29.835 59.205 ;
        RECT 28.605 58.335 28.895 59.005 ;
        RECT 30.015 58.825 30.245 59.465 ;
        RECT 30.425 59.025 30.715 59.755 ;
        RECT 31.365 59.030 31.655 59.755 ;
        RECT 31.825 59.005 33.035 59.755 ;
        RECT 33.295 59.205 33.465 59.585 ;
        RECT 33.645 59.375 33.975 59.755 ;
        RECT 33.295 59.035 33.960 59.205 ;
        RECT 34.155 59.080 34.415 59.585 ;
        RECT 34.585 59.375 35.475 59.545 ;
        RECT 29.075 58.515 29.540 58.825 ;
        RECT 29.720 58.515 30.245 58.825 ;
        RECT 30.425 58.515 30.725 58.845 ;
        RECT 31.825 58.465 32.345 59.005 ;
        RECT 28.605 58.115 29.375 58.335 ;
        RECT 28.585 57.205 28.925 57.935 ;
        RECT 29.105 57.385 29.375 58.115 ;
        RECT 29.555 58.095 30.715 58.335 ;
        RECT 29.555 57.385 29.785 58.095 ;
        RECT 29.955 57.205 30.285 57.915 ;
        RECT 30.455 57.385 30.715 58.095 ;
        RECT 31.365 57.205 31.655 58.370 ;
        RECT 32.515 58.295 33.035 58.835 ;
        RECT 33.225 58.485 33.555 58.855 ;
        RECT 33.790 58.780 33.960 59.035 ;
        RECT 33.790 58.450 34.075 58.780 ;
        RECT 33.790 58.305 33.960 58.450 ;
        RECT 31.825 57.205 33.035 58.295 ;
        RECT 33.295 58.135 33.960 58.305 ;
        RECT 34.245 58.280 34.415 59.080 ;
        RECT 34.585 58.820 35.135 59.205 ;
        RECT 35.305 58.650 35.475 59.375 ;
        RECT 33.295 57.375 33.465 58.135 ;
        RECT 33.645 57.205 33.975 57.965 ;
        RECT 34.145 57.375 34.415 58.280 ;
        RECT 34.585 58.580 35.475 58.650 ;
        RECT 35.645 59.050 35.865 59.535 ;
        RECT 36.035 59.215 36.285 59.755 ;
        RECT 36.455 59.105 36.715 59.585 ;
        RECT 35.645 58.625 35.975 59.050 ;
        RECT 34.585 58.555 35.480 58.580 ;
        RECT 34.585 58.540 35.490 58.555 ;
        RECT 34.585 58.525 35.495 58.540 ;
        RECT 34.585 58.520 35.505 58.525 ;
        RECT 34.585 58.510 35.510 58.520 ;
        RECT 34.585 58.500 35.515 58.510 ;
        RECT 34.585 58.495 35.525 58.500 ;
        RECT 34.585 58.485 35.535 58.495 ;
        RECT 34.585 58.480 35.545 58.485 ;
        RECT 34.585 58.030 34.845 58.480 ;
        RECT 35.210 58.475 35.545 58.480 ;
        RECT 35.210 58.470 35.560 58.475 ;
        RECT 35.210 58.460 35.575 58.470 ;
        RECT 35.210 58.455 35.600 58.460 ;
        RECT 36.145 58.455 36.375 58.850 ;
        RECT 35.210 58.450 36.375 58.455 ;
        RECT 35.240 58.415 36.375 58.450 ;
        RECT 35.275 58.390 36.375 58.415 ;
        RECT 35.305 58.360 36.375 58.390 ;
        RECT 35.325 58.330 36.375 58.360 ;
        RECT 35.345 58.300 36.375 58.330 ;
        RECT 35.415 58.290 36.375 58.300 ;
        RECT 35.440 58.280 36.375 58.290 ;
        RECT 35.460 58.265 36.375 58.280 ;
        RECT 35.480 58.250 36.375 58.265 ;
        RECT 35.485 58.240 36.270 58.250 ;
        RECT 35.500 58.205 36.270 58.240 ;
        RECT 35.015 57.885 35.345 58.130 ;
        RECT 35.515 57.955 36.270 58.205 ;
        RECT 36.545 58.075 36.715 59.105 ;
        RECT 36.885 58.985 38.555 59.755 ;
        RECT 39.275 59.205 39.445 59.495 ;
        RECT 39.615 59.375 39.945 59.755 ;
        RECT 39.275 59.035 39.940 59.205 ;
        RECT 36.885 58.465 37.635 58.985 ;
        RECT 37.805 58.295 38.555 58.815 ;
        RECT 35.015 57.860 35.200 57.885 ;
        RECT 34.585 57.760 35.200 57.860 ;
        RECT 34.585 57.205 35.190 57.760 ;
        RECT 35.365 57.375 35.845 57.715 ;
        RECT 36.015 57.205 36.270 57.750 ;
        RECT 36.440 57.375 36.715 58.075 ;
        RECT 36.885 57.205 38.555 58.295 ;
        RECT 39.190 58.215 39.540 58.865 ;
        RECT 39.710 58.045 39.940 59.035 ;
        RECT 39.275 57.875 39.940 58.045 ;
        RECT 39.275 57.375 39.445 57.875 ;
        RECT 39.615 57.205 39.945 57.705 ;
        RECT 40.115 57.375 40.300 59.495 ;
        RECT 40.555 59.295 40.805 59.755 ;
        RECT 40.975 59.305 41.310 59.475 ;
        RECT 41.505 59.305 42.180 59.475 ;
        RECT 40.975 59.165 41.145 59.305 ;
        RECT 40.470 58.175 40.750 59.125 ;
        RECT 40.920 59.035 41.145 59.165 ;
        RECT 40.920 57.930 41.090 59.035 ;
        RECT 41.315 58.885 41.840 59.105 ;
        RECT 41.260 58.120 41.500 58.715 ;
        RECT 41.670 58.185 41.840 58.885 ;
        RECT 42.010 58.525 42.180 59.305 ;
        RECT 42.500 59.255 42.870 59.755 ;
        RECT 43.050 59.305 43.455 59.475 ;
        RECT 43.625 59.305 44.410 59.475 ;
        RECT 43.050 59.075 43.220 59.305 ;
        RECT 42.390 58.775 43.220 59.075 ;
        RECT 43.605 58.805 44.070 59.135 ;
        RECT 42.390 58.745 42.590 58.775 ;
        RECT 42.710 58.525 42.880 58.595 ;
        RECT 42.010 58.355 42.880 58.525 ;
        RECT 42.370 58.265 42.880 58.355 ;
        RECT 40.920 57.800 41.225 57.930 ;
        RECT 41.670 57.820 42.200 58.185 ;
        RECT 40.540 57.205 40.805 57.665 ;
        RECT 40.975 57.375 41.225 57.800 ;
        RECT 42.370 57.650 42.540 58.265 ;
        RECT 41.435 57.480 42.540 57.650 ;
        RECT 42.710 57.205 42.880 58.005 ;
        RECT 43.050 57.705 43.220 58.775 ;
        RECT 43.390 57.875 43.580 58.595 ;
        RECT 43.750 57.845 44.070 58.805 ;
        RECT 44.240 58.845 44.410 59.305 ;
        RECT 44.685 59.225 44.895 59.755 ;
        RECT 45.155 59.015 45.485 59.540 ;
        RECT 45.655 59.145 45.825 59.755 ;
        RECT 45.995 59.100 46.325 59.535 ;
        RECT 46.565 59.245 46.805 59.755 ;
        RECT 45.995 59.015 46.375 59.100 ;
        RECT 45.285 58.845 45.485 59.015 ;
        RECT 46.150 58.975 46.375 59.015 ;
        RECT 44.240 58.515 45.115 58.845 ;
        RECT 45.285 58.515 46.035 58.845 ;
        RECT 43.050 57.375 43.300 57.705 ;
        RECT 44.240 57.675 44.410 58.515 ;
        RECT 45.285 58.310 45.475 58.515 ;
        RECT 46.205 58.395 46.375 58.975 ;
        RECT 46.550 58.515 46.805 59.075 ;
        RECT 46.975 59.015 47.305 59.550 ;
        RECT 47.520 59.015 47.690 59.755 ;
        RECT 47.900 59.105 48.230 59.575 ;
        RECT 48.400 59.275 48.570 59.755 ;
        RECT 48.740 59.105 49.070 59.575 ;
        RECT 49.240 59.275 49.410 59.755 ;
        RECT 46.160 58.345 46.375 58.395 ;
        RECT 46.975 58.345 47.155 59.015 ;
        RECT 47.900 58.935 49.595 59.105 ;
        RECT 49.815 59.100 50.145 59.535 ;
        RECT 50.315 59.145 50.485 59.755 ;
        RECT 47.325 58.515 47.700 58.845 ;
        RECT 47.870 58.595 49.080 58.765 ;
        RECT 47.870 58.345 48.075 58.595 ;
        RECT 49.250 58.345 49.595 58.935 ;
        RECT 44.580 57.935 45.475 58.310 ;
        RECT 45.985 58.265 46.375 58.345 ;
        RECT 43.525 57.505 44.410 57.675 ;
        RECT 44.590 57.205 44.905 57.705 ;
        RECT 45.135 57.375 45.475 57.935 ;
        RECT 45.645 57.205 45.815 58.215 ;
        RECT 45.985 57.420 46.315 58.265 ;
        RECT 46.615 58.175 48.075 58.345 ;
        RECT 48.740 58.175 49.595 58.345 ;
        RECT 49.765 59.015 50.145 59.100 ;
        RECT 50.655 59.015 50.985 59.540 ;
        RECT 51.245 59.225 51.455 59.755 ;
        RECT 51.730 59.305 52.515 59.475 ;
        RECT 52.685 59.305 53.090 59.475 ;
        RECT 49.765 58.975 49.990 59.015 ;
        RECT 49.765 58.395 49.935 58.975 ;
        RECT 50.655 58.845 50.855 59.015 ;
        RECT 51.730 58.845 51.900 59.305 ;
        RECT 50.105 58.515 50.855 58.845 ;
        RECT 51.025 58.515 51.900 58.845 ;
        RECT 49.765 58.345 49.980 58.395 ;
        RECT 49.765 58.265 50.155 58.345 ;
        RECT 46.615 57.375 46.975 58.175 ;
        RECT 48.740 58.005 49.070 58.175 ;
        RECT 47.520 57.205 47.690 58.005 ;
        RECT 47.900 57.835 49.070 58.005 ;
        RECT 47.900 57.375 48.230 57.835 ;
        RECT 48.400 57.205 48.570 57.665 ;
        RECT 48.740 57.375 49.070 57.835 ;
        RECT 49.240 57.205 49.410 58.005 ;
        RECT 49.825 57.420 50.155 58.265 ;
        RECT 50.665 58.310 50.855 58.515 ;
        RECT 50.325 57.205 50.495 58.215 ;
        RECT 50.665 57.935 51.560 58.310 ;
        RECT 50.665 57.375 51.005 57.935 ;
        RECT 51.235 57.205 51.550 57.705 ;
        RECT 51.730 57.675 51.900 58.515 ;
        RECT 52.070 58.805 52.535 59.135 ;
        RECT 52.920 59.075 53.090 59.305 ;
        RECT 53.270 59.255 53.640 59.755 ;
        RECT 53.960 59.305 54.635 59.475 ;
        RECT 54.830 59.305 55.165 59.475 ;
        RECT 52.070 57.845 52.390 58.805 ;
        RECT 52.920 58.775 53.750 59.075 ;
        RECT 52.560 57.875 52.750 58.595 ;
        RECT 52.920 57.705 53.090 58.775 ;
        RECT 53.550 58.745 53.750 58.775 ;
        RECT 53.260 58.525 53.430 58.595 ;
        RECT 53.960 58.525 54.130 59.305 ;
        RECT 54.995 59.165 55.165 59.305 ;
        RECT 55.335 59.295 55.585 59.755 ;
        RECT 53.260 58.355 54.130 58.525 ;
        RECT 54.300 58.885 54.825 59.105 ;
        RECT 54.995 59.035 55.220 59.165 ;
        RECT 53.260 58.265 53.770 58.355 ;
        RECT 51.730 57.505 52.615 57.675 ;
        RECT 52.840 57.375 53.090 57.705 ;
        RECT 53.260 57.205 53.430 58.005 ;
        RECT 53.600 57.650 53.770 58.265 ;
        RECT 54.300 58.185 54.470 58.885 ;
        RECT 53.940 57.820 54.470 58.185 ;
        RECT 54.640 58.120 54.880 58.715 ;
        RECT 55.050 57.930 55.220 59.035 ;
        RECT 55.390 58.175 55.670 59.125 ;
        RECT 54.915 57.800 55.220 57.930 ;
        RECT 53.600 57.480 54.705 57.650 ;
        RECT 54.915 57.375 55.165 57.800 ;
        RECT 55.335 57.205 55.600 57.665 ;
        RECT 55.840 57.375 56.025 59.495 ;
        RECT 56.195 59.375 56.525 59.755 ;
        RECT 56.695 59.205 56.865 59.495 ;
        RECT 56.200 59.035 56.865 59.205 ;
        RECT 56.200 58.045 56.430 59.035 ;
        RECT 57.125 59.030 57.415 59.755 ;
        RECT 57.585 58.985 60.175 59.755 ;
        RECT 60.435 59.205 60.605 59.495 ;
        RECT 60.775 59.375 61.105 59.755 ;
        RECT 60.435 59.035 61.100 59.205 ;
        RECT 56.600 58.215 56.950 58.865 ;
        RECT 57.585 58.465 58.795 58.985 ;
        RECT 56.200 57.875 56.865 58.045 ;
        RECT 56.195 57.205 56.525 57.705 ;
        RECT 56.695 57.375 56.865 57.875 ;
        RECT 57.125 57.205 57.415 58.370 ;
        RECT 58.965 58.295 60.175 58.815 ;
        RECT 57.585 57.205 60.175 58.295 ;
        RECT 60.350 58.215 60.700 58.865 ;
        RECT 60.870 58.045 61.100 59.035 ;
        RECT 60.435 57.875 61.100 58.045 ;
        RECT 60.435 57.375 60.605 57.875 ;
        RECT 60.775 57.205 61.105 57.705 ;
        RECT 61.275 57.375 61.460 59.495 ;
        RECT 61.715 59.295 61.965 59.755 ;
        RECT 62.135 59.305 62.470 59.475 ;
        RECT 62.665 59.305 63.340 59.475 ;
        RECT 62.135 59.165 62.305 59.305 ;
        RECT 61.630 58.175 61.910 59.125 ;
        RECT 62.080 59.035 62.305 59.165 ;
        RECT 62.080 57.930 62.250 59.035 ;
        RECT 62.475 58.885 63.000 59.105 ;
        RECT 62.420 58.120 62.660 58.715 ;
        RECT 62.830 58.185 63.000 58.885 ;
        RECT 63.170 58.525 63.340 59.305 ;
        RECT 63.660 59.255 64.030 59.755 ;
        RECT 64.210 59.305 64.615 59.475 ;
        RECT 64.785 59.305 65.570 59.475 ;
        RECT 64.210 59.075 64.380 59.305 ;
        RECT 63.550 58.775 64.380 59.075 ;
        RECT 64.765 58.805 65.230 59.135 ;
        RECT 63.550 58.745 63.750 58.775 ;
        RECT 63.870 58.525 64.040 58.595 ;
        RECT 63.170 58.355 64.040 58.525 ;
        RECT 63.530 58.265 64.040 58.355 ;
        RECT 62.080 57.800 62.385 57.930 ;
        RECT 62.830 57.820 63.360 58.185 ;
        RECT 61.700 57.205 61.965 57.665 ;
        RECT 62.135 57.375 62.385 57.800 ;
        RECT 63.530 57.650 63.700 58.265 ;
        RECT 62.595 57.480 63.700 57.650 ;
        RECT 63.870 57.205 64.040 58.005 ;
        RECT 64.210 57.705 64.380 58.775 ;
        RECT 64.550 57.875 64.740 58.595 ;
        RECT 64.910 57.845 65.230 58.805 ;
        RECT 65.400 58.845 65.570 59.305 ;
        RECT 65.845 59.225 66.055 59.755 ;
        RECT 66.315 59.015 66.645 59.540 ;
        RECT 66.815 59.145 66.985 59.755 ;
        RECT 67.155 59.100 67.485 59.535 ;
        RECT 67.155 59.015 67.535 59.100 ;
        RECT 66.445 58.845 66.645 59.015 ;
        RECT 67.310 58.975 67.535 59.015 ;
        RECT 65.400 58.515 66.275 58.845 ;
        RECT 66.445 58.515 67.195 58.845 ;
        RECT 64.210 57.375 64.460 57.705 ;
        RECT 65.400 57.675 65.570 58.515 ;
        RECT 66.445 58.310 66.635 58.515 ;
        RECT 67.365 58.395 67.535 58.975 ;
        RECT 67.710 58.915 67.970 59.755 ;
        RECT 68.145 59.010 68.400 59.585 ;
        RECT 68.570 59.375 68.900 59.755 ;
        RECT 69.115 59.205 69.285 59.585 ;
        RECT 68.570 59.035 69.285 59.205 ;
        RECT 69.745 59.125 70.075 59.485 ;
        RECT 70.695 59.295 70.945 59.755 ;
        RECT 71.115 59.295 71.675 59.585 ;
        RECT 67.320 58.345 67.535 58.395 ;
        RECT 65.740 57.935 66.635 58.310 ;
        RECT 67.145 58.265 67.535 58.345 ;
        RECT 64.685 57.505 65.570 57.675 ;
        RECT 65.750 57.205 66.065 57.705 ;
        RECT 66.295 57.375 66.635 57.935 ;
        RECT 66.805 57.205 66.975 58.215 ;
        RECT 67.145 57.420 67.475 58.265 ;
        RECT 67.710 57.205 67.970 58.355 ;
        RECT 68.145 58.280 68.315 59.010 ;
        RECT 68.570 58.845 68.740 59.035 ;
        RECT 69.745 58.935 71.135 59.125 ;
        RECT 68.485 58.515 68.740 58.845 ;
        RECT 68.570 58.305 68.740 58.515 ;
        RECT 69.020 58.485 69.375 58.855 ;
        RECT 70.965 58.845 71.135 58.935 ;
        RECT 69.560 58.515 70.235 58.765 ;
        RECT 70.455 58.515 70.795 58.765 ;
        RECT 70.965 58.515 71.255 58.845 ;
        RECT 68.145 57.375 68.400 58.280 ;
        RECT 68.570 58.135 69.285 58.305 ;
        RECT 69.560 58.155 69.825 58.515 ;
        RECT 70.965 58.265 71.135 58.515 ;
        RECT 68.570 57.205 68.900 57.965 ;
        RECT 69.115 57.375 69.285 58.135 ;
        RECT 70.195 58.095 71.135 58.265 ;
        RECT 69.745 57.205 70.025 57.875 ;
        RECT 70.195 57.545 70.495 58.095 ;
        RECT 71.425 57.925 71.675 59.295 ;
        RECT 72.010 59.245 72.250 59.755 ;
        RECT 72.430 59.245 72.710 59.575 ;
        RECT 72.940 59.245 73.155 59.755 ;
        RECT 71.905 58.515 72.260 59.075 ;
        RECT 72.430 58.345 72.600 59.245 ;
        RECT 72.770 58.515 73.035 59.075 ;
        RECT 73.325 59.015 73.940 59.585 ;
        RECT 74.695 59.205 74.865 59.495 ;
        RECT 75.035 59.375 75.365 59.755 ;
        RECT 74.695 59.035 75.360 59.205 ;
        RECT 73.285 58.345 73.455 58.845 ;
        RECT 72.030 58.175 73.455 58.345 ;
        RECT 72.030 58.000 72.420 58.175 ;
        RECT 70.695 57.205 71.025 57.925 ;
        RECT 71.215 57.375 71.675 57.925 ;
        RECT 72.905 57.205 73.235 58.005 ;
        RECT 73.625 57.995 73.940 59.015 ;
        RECT 74.610 58.215 74.960 58.865 ;
        RECT 75.130 58.045 75.360 59.035 ;
        RECT 73.405 57.375 73.940 57.995 ;
        RECT 74.695 57.875 75.360 58.045 ;
        RECT 74.695 57.375 74.865 57.875 ;
        RECT 75.035 57.205 75.365 57.705 ;
        RECT 75.535 57.375 75.720 59.495 ;
        RECT 75.975 59.295 76.225 59.755 ;
        RECT 76.395 59.305 76.730 59.475 ;
        RECT 76.925 59.305 77.600 59.475 ;
        RECT 76.395 59.165 76.565 59.305 ;
        RECT 75.890 58.175 76.170 59.125 ;
        RECT 76.340 59.035 76.565 59.165 ;
        RECT 76.340 57.930 76.510 59.035 ;
        RECT 76.735 58.885 77.260 59.105 ;
        RECT 76.680 58.120 76.920 58.715 ;
        RECT 77.090 58.185 77.260 58.885 ;
        RECT 77.430 58.525 77.600 59.305 ;
        RECT 77.920 59.255 78.290 59.755 ;
        RECT 78.470 59.305 78.875 59.475 ;
        RECT 79.045 59.305 79.830 59.475 ;
        RECT 78.470 59.075 78.640 59.305 ;
        RECT 77.810 58.775 78.640 59.075 ;
        RECT 79.025 58.805 79.490 59.135 ;
        RECT 77.810 58.745 78.010 58.775 ;
        RECT 78.130 58.525 78.300 58.595 ;
        RECT 77.430 58.355 78.300 58.525 ;
        RECT 77.790 58.265 78.300 58.355 ;
        RECT 76.340 57.800 76.645 57.930 ;
        RECT 77.090 57.820 77.620 58.185 ;
        RECT 75.960 57.205 76.225 57.665 ;
        RECT 76.395 57.375 76.645 57.800 ;
        RECT 77.790 57.650 77.960 58.265 ;
        RECT 76.855 57.480 77.960 57.650 ;
        RECT 78.130 57.205 78.300 58.005 ;
        RECT 78.470 57.705 78.640 58.775 ;
        RECT 78.810 57.875 79.000 58.595 ;
        RECT 79.170 57.845 79.490 58.805 ;
        RECT 79.660 58.845 79.830 59.305 ;
        RECT 80.105 59.225 80.315 59.755 ;
        RECT 80.575 59.015 80.905 59.540 ;
        RECT 81.075 59.145 81.245 59.755 ;
        RECT 81.415 59.100 81.745 59.535 ;
        RECT 81.415 59.015 81.795 59.100 ;
        RECT 80.705 58.845 80.905 59.015 ;
        RECT 81.570 58.975 81.795 59.015 ;
        RECT 81.965 59.005 83.175 59.755 ;
        RECT 79.660 58.515 80.535 58.845 ;
        RECT 80.705 58.515 81.455 58.845 ;
        RECT 78.470 57.375 78.720 57.705 ;
        RECT 79.660 57.675 79.830 58.515 ;
        RECT 80.705 58.310 80.895 58.515 ;
        RECT 81.625 58.395 81.795 58.975 ;
        RECT 81.580 58.345 81.795 58.395 ;
        RECT 80.000 57.935 80.895 58.310 ;
        RECT 81.405 58.265 81.795 58.345 ;
        RECT 81.965 58.295 82.485 58.835 ;
        RECT 82.655 58.465 83.175 59.005 ;
        RECT 78.945 57.505 79.830 57.675 ;
        RECT 80.010 57.205 80.325 57.705 ;
        RECT 80.555 57.375 80.895 57.935 ;
        RECT 81.065 57.205 81.235 58.215 ;
        RECT 81.405 57.420 81.735 58.265 ;
        RECT 81.965 57.205 83.175 58.295 ;
        RECT 5.520 57.035 83.260 57.205 ;
        RECT 5.605 55.945 6.815 57.035 ;
        RECT 7.075 56.365 7.245 56.865 ;
        RECT 7.415 56.535 7.745 57.035 ;
        RECT 7.075 56.195 7.740 56.365 ;
        RECT 5.605 55.235 6.125 55.775 ;
        RECT 6.295 55.405 6.815 55.945 ;
        RECT 6.990 55.375 7.340 56.025 ;
        RECT 5.605 54.485 6.815 55.235 ;
        RECT 7.510 55.205 7.740 56.195 ;
        RECT 7.075 55.035 7.740 55.205 ;
        RECT 7.075 54.745 7.245 55.035 ;
        RECT 7.415 54.485 7.745 54.865 ;
        RECT 7.915 54.745 8.100 56.865 ;
        RECT 8.340 56.575 8.605 57.035 ;
        RECT 8.775 56.440 9.025 56.865 ;
        RECT 9.235 56.590 10.340 56.760 ;
        RECT 8.720 56.310 9.025 56.440 ;
        RECT 8.270 55.115 8.550 56.065 ;
        RECT 8.720 55.205 8.890 56.310 ;
        RECT 9.060 55.525 9.300 56.120 ;
        RECT 9.470 56.055 10.000 56.420 ;
        RECT 9.470 55.355 9.640 56.055 ;
        RECT 10.170 55.975 10.340 56.590 ;
        RECT 10.510 56.235 10.680 57.035 ;
        RECT 10.850 56.535 11.100 56.865 ;
        RECT 11.325 56.565 12.210 56.735 ;
        RECT 10.170 55.885 10.680 55.975 ;
        RECT 8.720 55.075 8.945 55.205 ;
        RECT 9.115 55.135 9.640 55.355 ;
        RECT 9.810 55.715 10.680 55.885 ;
        RECT 8.355 54.485 8.605 54.945 ;
        RECT 8.775 54.935 8.945 55.075 ;
        RECT 9.810 54.935 9.980 55.715 ;
        RECT 10.510 55.645 10.680 55.715 ;
        RECT 10.190 55.465 10.390 55.495 ;
        RECT 10.850 55.465 11.020 56.535 ;
        RECT 11.190 55.645 11.380 56.365 ;
        RECT 10.190 55.165 11.020 55.465 ;
        RECT 11.550 55.435 11.870 56.395 ;
        RECT 8.775 54.765 9.110 54.935 ;
        RECT 9.305 54.765 9.980 54.935 ;
        RECT 10.300 54.485 10.670 54.985 ;
        RECT 10.850 54.935 11.020 55.165 ;
        RECT 11.405 55.105 11.870 55.435 ;
        RECT 12.040 55.725 12.210 56.565 ;
        RECT 12.390 56.535 12.705 57.035 ;
        RECT 12.935 56.305 13.275 56.865 ;
        RECT 12.380 55.930 13.275 56.305 ;
        RECT 13.445 56.025 13.615 57.035 ;
        RECT 13.085 55.725 13.275 55.930 ;
        RECT 13.785 55.975 14.115 56.820 ;
        RECT 14.355 56.065 14.685 56.850 ;
        RECT 13.785 55.895 14.175 55.975 ;
        RECT 14.355 55.895 15.035 56.065 ;
        RECT 15.215 55.895 15.545 57.035 ;
        RECT 15.725 55.945 18.315 57.035 ;
        RECT 13.960 55.845 14.175 55.895 ;
        RECT 12.040 55.395 12.915 55.725 ;
        RECT 13.085 55.395 13.835 55.725 ;
        RECT 12.040 54.935 12.210 55.395 ;
        RECT 13.085 55.225 13.285 55.395 ;
        RECT 14.005 55.265 14.175 55.845 ;
        RECT 14.345 55.475 14.695 55.725 ;
        RECT 14.865 55.295 15.035 55.895 ;
        RECT 15.205 55.475 15.555 55.725 ;
        RECT 13.950 55.225 14.175 55.265 ;
        RECT 10.850 54.765 11.255 54.935 ;
        RECT 11.425 54.765 12.210 54.935 ;
        RECT 12.485 54.485 12.695 55.015 ;
        RECT 12.955 54.700 13.285 55.225 ;
        RECT 13.795 55.140 14.175 55.225 ;
        RECT 13.455 54.485 13.625 55.095 ;
        RECT 13.795 54.705 14.125 55.140 ;
        RECT 14.365 54.485 14.605 55.295 ;
        RECT 14.775 54.655 15.105 55.295 ;
        RECT 15.275 54.485 15.545 55.295 ;
        RECT 15.725 55.255 16.935 55.775 ;
        RECT 17.105 55.425 18.315 55.945 ;
        RECT 18.485 55.870 18.775 57.035 ;
        RECT 18.945 55.945 21.535 57.035 ;
        RECT 18.945 55.255 20.155 55.775 ;
        RECT 20.325 55.425 21.535 55.945 ;
        RECT 21.705 55.895 21.965 57.035 ;
        RECT 22.135 55.885 22.465 56.865 ;
        RECT 22.635 55.895 22.915 57.035 ;
        RECT 23.085 55.895 23.365 57.035 ;
        RECT 23.535 55.885 23.865 56.865 ;
        RECT 24.035 55.895 24.295 57.035 ;
        RECT 24.465 55.945 26.135 57.035 ;
        RECT 21.725 55.475 22.060 55.725 ;
        RECT 22.230 55.285 22.400 55.885 ;
        RECT 23.600 55.845 23.775 55.885 ;
        RECT 22.570 55.455 22.905 55.725 ;
        RECT 23.095 55.455 23.430 55.725 ;
        RECT 23.600 55.285 23.770 55.845 ;
        RECT 23.940 55.475 24.275 55.725 ;
        RECT 15.725 54.485 18.315 55.255 ;
        RECT 18.485 54.485 18.775 55.210 ;
        RECT 18.945 54.485 21.535 55.255 ;
        RECT 21.705 54.655 22.400 55.285 ;
        RECT 22.605 54.485 22.915 55.285 ;
        RECT 23.085 54.485 23.395 55.285 ;
        RECT 23.600 54.655 24.295 55.285 ;
        RECT 24.465 55.255 25.215 55.775 ;
        RECT 25.385 55.425 26.135 55.945 ;
        RECT 26.305 56.165 26.580 56.865 ;
        RECT 26.750 56.490 27.005 57.035 ;
        RECT 27.175 56.525 27.655 56.865 ;
        RECT 27.830 56.480 28.435 57.035 ;
        RECT 28.605 56.600 33.950 57.035 ;
        RECT 34.125 56.600 39.470 57.035 ;
        RECT 27.820 56.380 28.435 56.480 ;
        RECT 27.820 56.355 28.005 56.380 ;
        RECT 24.465 54.485 26.135 55.255 ;
        RECT 26.305 55.135 26.475 56.165 ;
        RECT 26.750 56.035 27.505 56.285 ;
        RECT 27.675 56.110 28.005 56.355 ;
        RECT 26.750 56.000 27.520 56.035 ;
        RECT 26.750 55.990 27.535 56.000 ;
        RECT 26.645 55.975 27.540 55.990 ;
        RECT 26.645 55.960 27.560 55.975 ;
        RECT 26.645 55.950 27.580 55.960 ;
        RECT 26.645 55.940 27.605 55.950 ;
        RECT 26.645 55.910 27.675 55.940 ;
        RECT 26.645 55.880 27.695 55.910 ;
        RECT 26.645 55.850 27.715 55.880 ;
        RECT 26.645 55.825 27.745 55.850 ;
        RECT 26.645 55.790 27.780 55.825 ;
        RECT 26.645 55.785 27.810 55.790 ;
        RECT 26.645 55.390 26.875 55.785 ;
        RECT 27.420 55.780 27.810 55.785 ;
        RECT 27.445 55.770 27.810 55.780 ;
        RECT 27.460 55.765 27.810 55.770 ;
        RECT 27.475 55.760 27.810 55.765 ;
        RECT 28.175 55.760 28.435 56.210 ;
        RECT 27.475 55.755 28.435 55.760 ;
        RECT 27.485 55.745 28.435 55.755 ;
        RECT 27.495 55.740 28.435 55.745 ;
        RECT 27.505 55.730 28.435 55.740 ;
        RECT 27.510 55.720 28.435 55.730 ;
        RECT 27.515 55.715 28.435 55.720 ;
        RECT 27.525 55.700 28.435 55.715 ;
        RECT 27.530 55.685 28.435 55.700 ;
        RECT 27.540 55.660 28.435 55.685 ;
        RECT 27.045 55.190 27.375 55.615 ;
        RECT 26.305 54.655 26.565 55.135 ;
        RECT 26.735 54.485 26.985 55.025 ;
        RECT 27.155 54.705 27.375 55.190 ;
        RECT 27.545 55.590 28.435 55.660 ;
        RECT 27.545 54.865 27.715 55.590 ;
        RECT 27.885 55.035 28.435 55.420 ;
        RECT 30.190 55.030 30.530 55.860 ;
        RECT 32.010 55.350 32.360 56.600 ;
        RECT 35.710 55.030 36.050 55.860 ;
        RECT 37.530 55.350 37.880 56.600 ;
        RECT 39.645 55.945 41.315 57.035 ;
        RECT 41.945 56.480 42.550 57.035 ;
        RECT 42.725 56.525 43.205 56.865 ;
        RECT 43.375 56.490 43.630 57.035 ;
        RECT 41.945 56.380 42.560 56.480 ;
        RECT 42.375 56.355 42.560 56.380 ;
        RECT 39.645 55.255 40.395 55.775 ;
        RECT 40.565 55.425 41.315 55.945 ;
        RECT 41.945 55.760 42.205 56.210 ;
        RECT 42.375 56.110 42.705 56.355 ;
        RECT 42.875 56.035 43.630 56.285 ;
        RECT 43.800 56.165 44.075 56.865 ;
        RECT 42.860 56.000 43.630 56.035 ;
        RECT 42.845 55.990 43.630 56.000 ;
        RECT 42.840 55.975 43.735 55.990 ;
        RECT 42.820 55.960 43.735 55.975 ;
        RECT 42.800 55.950 43.735 55.960 ;
        RECT 42.775 55.940 43.735 55.950 ;
        RECT 42.705 55.910 43.735 55.940 ;
        RECT 42.685 55.880 43.735 55.910 ;
        RECT 42.665 55.850 43.735 55.880 ;
        RECT 42.635 55.825 43.735 55.850 ;
        RECT 42.600 55.790 43.735 55.825 ;
        RECT 42.570 55.785 43.735 55.790 ;
        RECT 42.570 55.780 42.960 55.785 ;
        RECT 42.570 55.770 42.935 55.780 ;
        RECT 42.570 55.765 42.920 55.770 ;
        RECT 42.570 55.760 42.905 55.765 ;
        RECT 41.945 55.755 42.905 55.760 ;
        RECT 41.945 55.745 42.895 55.755 ;
        RECT 41.945 55.740 42.885 55.745 ;
        RECT 41.945 55.730 42.875 55.740 ;
        RECT 41.945 55.720 42.870 55.730 ;
        RECT 41.945 55.715 42.865 55.720 ;
        RECT 41.945 55.700 42.855 55.715 ;
        RECT 41.945 55.685 42.850 55.700 ;
        RECT 41.945 55.660 42.840 55.685 ;
        RECT 41.945 55.590 42.835 55.660 ;
        RECT 27.545 54.695 28.435 54.865 ;
        RECT 28.605 54.485 33.950 55.030 ;
        RECT 34.125 54.485 39.470 55.030 ;
        RECT 39.645 54.485 41.315 55.255 ;
        RECT 41.945 55.035 42.495 55.420 ;
        RECT 42.665 54.865 42.835 55.590 ;
        RECT 41.945 54.695 42.835 54.865 ;
        RECT 43.005 55.190 43.335 55.615 ;
        RECT 43.505 55.390 43.735 55.785 ;
        RECT 43.005 54.705 43.225 55.190 ;
        RECT 43.905 55.135 44.075 56.165 ;
        RECT 44.245 55.870 44.535 57.035 ;
        RECT 44.705 56.525 45.905 56.765 ;
        RECT 46.085 56.610 46.415 57.035 ;
        RECT 46.930 56.610 47.290 57.035 ;
        RECT 47.495 56.440 47.755 56.620 ;
        RECT 46.120 56.355 47.755 56.440 ;
        RECT 47.925 56.480 48.530 57.035 ;
        RECT 48.705 56.525 49.185 56.865 ;
        RECT 49.355 56.490 49.610 57.035 ;
        RECT 47.925 56.380 48.540 56.480 ;
        RECT 44.705 55.895 45.010 56.325 ;
        RECT 45.180 56.270 47.755 56.355 ;
        RECT 45.180 56.185 46.290 56.270 ;
        RECT 47.075 56.210 47.755 56.270 ;
        RECT 48.355 56.355 48.540 56.380 ;
        RECT 44.705 55.225 44.875 55.895 ;
        RECT 45.180 55.725 45.350 56.185 ;
        RECT 45.050 55.395 45.350 55.725 ;
        RECT 45.610 55.475 46.145 56.015 ;
        RECT 46.510 55.895 46.905 56.100 ;
        RECT 46.395 55.335 46.565 55.725 ;
        RECT 46.245 55.305 46.565 55.335 ;
        RECT 45.680 55.225 46.565 55.305 ;
        RECT 43.395 54.485 43.645 55.025 ;
        RECT 43.815 54.655 44.075 55.135 ;
        RECT 44.245 54.485 44.535 55.210 ;
        RECT 44.705 55.165 46.565 55.225 ;
        RECT 44.705 55.135 46.415 55.165 ;
        RECT 44.705 55.055 45.850 55.135 ;
        RECT 44.705 55.005 45.010 55.055 ;
        RECT 44.755 54.705 45.010 55.005 ;
        RECT 45.180 54.485 45.510 54.885 ;
        RECT 45.680 54.705 45.850 55.055 ;
        RECT 46.735 54.995 46.905 55.895 ;
        RECT 47.075 55.305 47.245 56.210 ;
        RECT 47.415 55.475 47.755 56.040 ;
        RECT 47.925 55.760 48.185 56.210 ;
        RECT 48.355 56.110 48.685 56.355 ;
        RECT 48.855 56.035 49.610 56.285 ;
        RECT 49.780 56.165 50.055 56.865 ;
        RECT 50.225 56.600 55.570 57.035 ;
        RECT 48.840 56.000 49.610 56.035 ;
        RECT 48.825 55.990 49.610 56.000 ;
        RECT 48.820 55.975 49.715 55.990 ;
        RECT 48.800 55.960 49.715 55.975 ;
        RECT 48.780 55.950 49.715 55.960 ;
        RECT 48.755 55.940 49.715 55.950 ;
        RECT 48.685 55.910 49.715 55.940 ;
        RECT 48.665 55.880 49.715 55.910 ;
        RECT 48.645 55.850 49.715 55.880 ;
        RECT 48.615 55.825 49.715 55.850 ;
        RECT 48.580 55.790 49.715 55.825 ;
        RECT 48.550 55.785 49.715 55.790 ;
        RECT 48.550 55.780 48.940 55.785 ;
        RECT 48.550 55.770 48.915 55.780 ;
        RECT 48.550 55.765 48.900 55.770 ;
        RECT 48.550 55.760 48.885 55.765 ;
        RECT 47.925 55.755 48.885 55.760 ;
        RECT 47.925 55.745 48.875 55.755 ;
        RECT 47.925 55.740 48.865 55.745 ;
        RECT 47.925 55.730 48.855 55.740 ;
        RECT 47.925 55.720 48.850 55.730 ;
        RECT 47.925 55.715 48.845 55.720 ;
        RECT 47.925 55.700 48.835 55.715 ;
        RECT 47.925 55.685 48.830 55.700 ;
        RECT 47.925 55.660 48.820 55.685 ;
        RECT 47.925 55.590 48.815 55.660 ;
        RECT 47.075 55.135 47.755 55.305 ;
        RECT 46.150 54.485 46.320 54.965 ;
        RECT 46.555 54.665 46.905 54.995 ;
        RECT 47.075 54.485 47.245 54.965 ;
        RECT 47.495 54.690 47.755 55.135 ;
        RECT 47.925 55.035 48.475 55.420 ;
        RECT 48.645 54.865 48.815 55.590 ;
        RECT 47.925 54.695 48.815 54.865 ;
        RECT 48.985 55.190 49.315 55.615 ;
        RECT 49.485 55.390 49.715 55.785 ;
        RECT 48.985 54.705 49.205 55.190 ;
        RECT 49.885 55.135 50.055 56.165 ;
        RECT 49.375 54.485 49.625 55.025 ;
        RECT 49.795 54.655 50.055 55.135 ;
        RECT 51.810 55.030 52.150 55.860 ;
        RECT 53.630 55.350 53.980 56.600 ;
        RECT 55.745 55.945 58.335 57.035 ;
        RECT 55.745 55.255 56.955 55.775 ;
        RECT 57.125 55.425 58.335 55.945 ;
        RECT 58.515 55.925 58.810 57.035 ;
        RECT 58.990 55.725 59.240 56.860 ;
        RECT 59.410 55.925 59.670 57.035 ;
        RECT 59.840 56.135 60.100 56.860 ;
        RECT 60.270 56.305 60.530 57.035 ;
        RECT 60.700 56.135 60.960 56.860 ;
        RECT 61.130 56.305 61.390 57.035 ;
        RECT 61.560 56.135 61.820 56.860 ;
        RECT 61.990 56.305 62.250 57.035 ;
        RECT 62.420 56.135 62.680 56.860 ;
        RECT 62.850 56.305 63.145 57.035 ;
        RECT 59.840 55.895 63.150 56.135 ;
        RECT 63.565 55.945 65.235 57.035 ;
        RECT 65.510 56.235 65.765 57.035 ;
        RECT 65.935 56.065 66.265 56.865 ;
        RECT 66.435 56.235 66.605 57.035 ;
        RECT 66.775 56.065 67.105 56.865 ;
        RECT 50.225 54.485 55.570 55.030 ;
        RECT 55.745 54.485 58.335 55.255 ;
        RECT 58.505 55.115 58.820 55.725 ;
        RECT 58.990 55.475 62.010 55.725 ;
        RECT 58.565 54.485 58.810 54.945 ;
        RECT 58.990 54.665 59.240 55.475 ;
        RECT 62.180 55.305 63.150 55.895 ;
        RECT 59.840 55.135 63.150 55.305 ;
        RECT 63.565 55.255 64.315 55.775 ;
        RECT 64.485 55.425 65.235 55.945 ;
        RECT 65.405 55.895 67.105 56.065 ;
        RECT 67.275 55.895 67.535 57.035 ;
        RECT 67.705 56.315 68.165 56.865 ;
        RECT 68.355 56.315 68.685 57.035 ;
        RECT 65.405 55.305 65.685 55.895 ;
        RECT 65.855 55.475 66.605 55.725 ;
        RECT 66.775 55.475 67.535 55.725 ;
        RECT 59.410 54.485 59.670 55.010 ;
        RECT 59.840 54.680 60.100 55.135 ;
        RECT 60.270 54.485 60.530 54.965 ;
        RECT 60.700 54.680 60.960 55.135 ;
        RECT 61.130 54.485 61.390 54.965 ;
        RECT 61.560 54.680 61.820 55.135 ;
        RECT 61.990 54.485 62.250 54.965 ;
        RECT 62.420 54.680 62.680 55.135 ;
        RECT 62.850 54.485 63.150 54.965 ;
        RECT 63.565 54.485 65.235 55.255 ;
        RECT 65.405 55.055 66.265 55.305 ;
        RECT 66.435 55.115 67.535 55.285 ;
        RECT 65.515 54.865 65.845 54.885 ;
        RECT 66.435 54.865 66.685 55.115 ;
        RECT 65.515 54.655 66.685 54.865 ;
        RECT 66.855 54.485 67.025 54.945 ;
        RECT 67.195 54.655 67.535 55.115 ;
        RECT 67.705 54.945 67.955 56.315 ;
        RECT 68.885 56.145 69.185 56.695 ;
        RECT 69.355 56.365 69.635 57.035 ;
        RECT 68.245 55.975 69.185 56.145 ;
        RECT 68.245 55.725 68.415 55.975 ;
        RECT 69.555 55.725 69.820 56.085 ;
        RECT 70.005 55.870 70.295 57.035 ;
        RECT 71.130 56.065 71.460 56.865 ;
        RECT 71.630 56.235 71.960 57.035 ;
        RECT 72.260 56.065 72.590 56.865 ;
        RECT 73.235 56.235 73.485 57.035 ;
        RECT 71.130 55.895 73.565 56.065 ;
        RECT 73.755 55.895 73.925 57.035 ;
        RECT 74.095 55.895 74.435 56.865 ;
        RECT 74.695 56.365 74.865 56.865 ;
        RECT 75.035 56.535 75.365 57.035 ;
        RECT 74.695 56.195 75.360 56.365 ;
        RECT 68.125 55.395 68.415 55.725 ;
        RECT 68.585 55.475 68.925 55.725 ;
        RECT 69.145 55.475 69.820 55.725 ;
        RECT 70.925 55.475 71.275 55.725 ;
        RECT 68.245 55.305 68.415 55.395 ;
        RECT 68.245 55.115 69.635 55.305 ;
        RECT 71.460 55.265 71.630 55.895 ;
        RECT 71.800 55.475 72.130 55.675 ;
        RECT 72.300 55.475 72.630 55.675 ;
        RECT 72.800 55.475 73.220 55.675 ;
        RECT 73.395 55.645 73.565 55.895 ;
        RECT 73.395 55.475 74.090 55.645 ;
        RECT 67.705 54.655 68.265 54.945 ;
        RECT 68.435 54.485 68.685 54.945 ;
        RECT 69.305 54.755 69.635 55.115 ;
        RECT 70.005 54.485 70.295 55.210 ;
        RECT 71.130 54.655 71.630 55.265 ;
        RECT 72.260 55.135 73.485 55.305 ;
        RECT 74.260 55.285 74.435 55.895 ;
        RECT 74.610 55.375 74.960 56.025 ;
        RECT 72.260 54.655 72.590 55.135 ;
        RECT 72.760 54.485 72.985 54.945 ;
        RECT 73.155 54.655 73.485 55.135 ;
        RECT 73.675 54.485 73.925 55.285 ;
        RECT 74.095 54.655 74.435 55.285 ;
        RECT 75.130 55.205 75.360 56.195 ;
        RECT 74.695 55.035 75.360 55.205 ;
        RECT 74.695 54.745 74.865 55.035 ;
        RECT 75.035 54.485 75.365 54.865 ;
        RECT 75.535 54.745 75.720 56.865 ;
        RECT 75.960 56.575 76.225 57.035 ;
        RECT 76.395 56.440 76.645 56.865 ;
        RECT 76.855 56.590 77.960 56.760 ;
        RECT 76.340 56.310 76.645 56.440 ;
        RECT 75.890 55.115 76.170 56.065 ;
        RECT 76.340 55.205 76.510 56.310 ;
        RECT 76.680 55.525 76.920 56.120 ;
        RECT 77.090 56.055 77.620 56.420 ;
        RECT 77.090 55.355 77.260 56.055 ;
        RECT 77.790 55.975 77.960 56.590 ;
        RECT 78.130 56.235 78.300 57.035 ;
        RECT 78.470 56.535 78.720 56.865 ;
        RECT 78.945 56.565 79.830 56.735 ;
        RECT 77.790 55.885 78.300 55.975 ;
        RECT 76.340 55.075 76.565 55.205 ;
        RECT 76.735 55.135 77.260 55.355 ;
        RECT 77.430 55.715 78.300 55.885 ;
        RECT 75.975 54.485 76.225 54.945 ;
        RECT 76.395 54.935 76.565 55.075 ;
        RECT 77.430 54.935 77.600 55.715 ;
        RECT 78.130 55.645 78.300 55.715 ;
        RECT 77.810 55.465 78.010 55.495 ;
        RECT 78.470 55.465 78.640 56.535 ;
        RECT 78.810 55.645 79.000 56.365 ;
        RECT 77.810 55.165 78.640 55.465 ;
        RECT 79.170 55.435 79.490 56.395 ;
        RECT 76.395 54.765 76.730 54.935 ;
        RECT 76.925 54.765 77.600 54.935 ;
        RECT 77.920 54.485 78.290 54.985 ;
        RECT 78.470 54.935 78.640 55.165 ;
        RECT 79.025 55.105 79.490 55.435 ;
        RECT 79.660 55.725 79.830 56.565 ;
        RECT 80.010 56.535 80.325 57.035 ;
        RECT 80.555 56.305 80.895 56.865 ;
        RECT 80.000 55.930 80.895 56.305 ;
        RECT 81.065 56.025 81.235 57.035 ;
        RECT 80.705 55.725 80.895 55.930 ;
        RECT 81.405 55.975 81.735 56.820 ;
        RECT 81.405 55.895 81.795 55.975 ;
        RECT 81.580 55.845 81.795 55.895 ;
        RECT 79.660 55.395 80.535 55.725 ;
        RECT 80.705 55.395 81.455 55.725 ;
        RECT 79.660 54.935 79.830 55.395 ;
        RECT 80.705 55.225 80.905 55.395 ;
        RECT 81.625 55.265 81.795 55.845 ;
        RECT 81.965 55.945 83.175 57.035 ;
        RECT 81.965 55.405 82.485 55.945 ;
        RECT 81.570 55.225 81.795 55.265 ;
        RECT 82.655 55.235 83.175 55.775 ;
        RECT 78.470 54.765 78.875 54.935 ;
        RECT 79.045 54.765 79.830 54.935 ;
        RECT 80.105 54.485 80.315 55.015 ;
        RECT 80.575 54.700 80.905 55.225 ;
        RECT 81.415 55.140 81.795 55.225 ;
        RECT 81.075 54.485 81.245 55.095 ;
        RECT 81.415 54.705 81.745 55.140 ;
        RECT 81.965 54.485 83.175 55.235 ;
        RECT 5.520 54.315 83.260 54.485 ;
        RECT 5.605 53.565 6.815 54.315 ;
        RECT 6.985 53.565 8.195 54.315 ;
        RECT 8.365 53.665 8.625 54.145 ;
        RECT 8.795 53.775 9.045 54.315 ;
        RECT 5.605 53.025 6.125 53.565 ;
        RECT 6.295 52.855 6.815 53.395 ;
        RECT 6.985 53.025 7.505 53.565 ;
        RECT 7.675 52.855 8.195 53.395 ;
        RECT 5.605 51.765 6.815 52.855 ;
        RECT 6.985 51.765 8.195 52.855 ;
        RECT 8.365 52.635 8.535 53.665 ;
        RECT 9.215 53.610 9.435 54.095 ;
        RECT 8.705 53.015 8.935 53.410 ;
        RECT 9.105 53.185 9.435 53.610 ;
        RECT 9.605 53.935 10.495 54.105 ;
        RECT 9.605 53.210 9.775 53.935 ;
        RECT 10.665 53.815 10.925 54.145 ;
        RECT 11.135 53.835 11.410 54.315 ;
        RECT 9.945 53.380 10.495 53.765 ;
        RECT 9.605 53.140 10.495 53.210 ;
        RECT 9.600 53.115 10.495 53.140 ;
        RECT 9.590 53.100 10.495 53.115 ;
        RECT 9.585 53.085 10.495 53.100 ;
        RECT 9.575 53.080 10.495 53.085 ;
        RECT 9.570 53.070 10.495 53.080 ;
        RECT 9.565 53.060 10.495 53.070 ;
        RECT 9.555 53.055 10.495 53.060 ;
        RECT 9.545 53.045 10.495 53.055 ;
        RECT 9.535 53.040 10.495 53.045 ;
        RECT 9.535 53.035 9.870 53.040 ;
        RECT 9.520 53.030 9.870 53.035 ;
        RECT 9.505 53.020 9.870 53.030 ;
        RECT 9.480 53.015 9.870 53.020 ;
        RECT 8.705 53.010 9.870 53.015 ;
        RECT 8.705 52.975 9.840 53.010 ;
        RECT 8.705 52.950 9.805 52.975 ;
        RECT 8.705 52.920 9.775 52.950 ;
        RECT 8.705 52.890 9.755 52.920 ;
        RECT 8.705 52.860 9.735 52.890 ;
        RECT 8.705 52.850 9.665 52.860 ;
        RECT 8.705 52.840 9.640 52.850 ;
        RECT 8.705 52.825 9.620 52.840 ;
        RECT 8.705 52.810 9.600 52.825 ;
        RECT 8.810 52.800 9.595 52.810 ;
        RECT 8.810 52.765 9.580 52.800 ;
        RECT 8.365 51.935 8.640 52.635 ;
        RECT 8.810 52.515 9.565 52.765 ;
        RECT 9.735 52.445 10.065 52.690 ;
        RECT 10.235 52.590 10.495 53.040 ;
        RECT 10.665 52.905 10.835 53.815 ;
        RECT 11.620 53.745 11.825 54.145 ;
        RECT 11.995 53.915 12.330 54.315 ;
        RECT 11.005 53.075 11.365 53.655 ;
        RECT 11.620 53.575 12.305 53.745 ;
        RECT 11.545 52.905 11.795 53.405 ;
        RECT 10.665 52.735 11.795 52.905 ;
        RECT 9.880 52.420 10.065 52.445 ;
        RECT 9.880 52.320 10.495 52.420 ;
        RECT 8.810 51.765 9.065 52.310 ;
        RECT 9.235 51.935 9.715 52.275 ;
        RECT 9.890 51.765 10.495 52.320 ;
        RECT 10.665 51.965 10.935 52.735 ;
        RECT 11.965 52.545 12.305 53.575 ;
        RECT 12.515 53.505 12.785 54.315 ;
        RECT 12.955 53.505 13.285 54.145 ;
        RECT 13.455 53.505 13.695 54.315 ;
        RECT 13.885 53.770 19.230 54.315 ;
        RECT 12.505 53.075 12.855 53.325 ;
        RECT 13.025 52.905 13.195 53.505 ;
        RECT 13.365 53.075 13.715 53.325 ;
        RECT 15.470 52.940 15.810 53.770 ;
        RECT 19.875 53.675 20.205 54.145 ;
        RECT 20.375 53.845 20.545 54.315 ;
        RECT 20.715 53.675 21.045 54.145 ;
        RECT 21.215 53.845 21.385 54.315 ;
        RECT 21.555 53.925 23.565 54.145 ;
        RECT 23.755 53.925 25.765 54.145 ;
        RECT 21.555 53.675 21.805 53.925 ;
        RECT 19.875 53.495 21.805 53.675 ;
        RECT 21.975 53.515 25.345 53.755 ;
        RECT 25.515 53.675 25.765 53.925 ;
        RECT 25.935 53.845 26.105 54.315 ;
        RECT 26.275 53.675 26.605 54.145 ;
        RECT 26.775 53.845 26.945 54.315 ;
        RECT 27.115 53.675 27.445 54.145 ;
        RECT 27.850 53.805 28.090 54.315 ;
        RECT 28.270 53.805 28.550 54.135 ;
        RECT 28.780 53.805 28.995 54.315 ;
        RECT 11.105 51.765 11.435 52.545 ;
        RECT 11.640 52.370 12.305 52.545 ;
        RECT 11.640 51.965 11.825 52.370 ;
        RECT 11.995 51.765 12.330 52.190 ;
        RECT 12.515 51.765 12.845 52.905 ;
        RECT 13.025 52.735 13.705 52.905 ;
        RECT 13.375 51.950 13.705 52.735 ;
        RECT 17.290 52.200 17.640 53.450 ;
        RECT 19.870 53.125 21.675 53.325 ;
        RECT 21.975 52.955 22.225 53.515 ;
        RECT 25.515 53.495 27.445 53.675 ;
        RECT 22.395 53.125 23.820 53.325 ;
        RECT 24.055 53.115 25.465 53.325 ;
        RECT 25.690 53.115 27.515 53.325 ;
        RECT 27.745 53.075 28.100 53.635 ;
        RECT 13.885 51.765 19.230 52.200 ;
        RECT 19.870 52.105 20.205 52.945 ;
        RECT 20.375 52.775 23.105 52.955 ;
        RECT 20.375 52.275 20.585 52.775 ;
        RECT 20.755 52.105 21.005 52.605 ;
        RECT 21.175 52.275 21.425 52.775 ;
        RECT 21.595 52.105 21.845 52.605 ;
        RECT 22.015 52.275 22.265 52.775 ;
        RECT 22.435 52.105 22.685 52.605 ;
        RECT 22.855 52.275 23.105 52.775 ;
        RECT 23.275 52.775 27.405 52.945 ;
        RECT 28.270 52.905 28.440 53.805 ;
        RECT 28.610 53.075 28.875 53.635 ;
        RECT 29.165 53.575 29.780 54.145 ;
        RECT 29.125 52.905 29.295 53.405 ;
        RECT 23.275 52.105 24.045 52.775 ;
        RECT 19.870 51.935 24.045 52.105 ;
        RECT 24.215 51.765 24.465 52.605 ;
        RECT 24.635 51.935 24.885 52.775 ;
        RECT 25.055 51.765 25.305 52.605 ;
        RECT 25.475 51.935 25.725 52.775 ;
        RECT 25.895 51.765 26.145 52.605 ;
        RECT 26.315 51.935 26.565 52.775 ;
        RECT 26.735 51.765 26.985 52.605 ;
        RECT 27.155 51.935 27.405 52.775 ;
        RECT 27.870 52.735 29.295 52.905 ;
        RECT 27.870 52.560 28.260 52.735 ;
        RECT 28.745 51.765 29.075 52.565 ;
        RECT 29.465 52.555 29.780 53.575 ;
        RECT 29.985 53.565 31.195 54.315 ;
        RECT 31.365 53.590 31.655 54.315 ;
        RECT 29.985 53.025 30.505 53.565 ;
        RECT 31.825 53.545 35.335 54.315 ;
        RECT 35.505 53.565 36.715 54.315 ;
        RECT 36.895 53.585 37.195 54.315 ;
        RECT 30.675 52.855 31.195 53.395 ;
        RECT 31.825 53.025 33.475 53.545 ;
        RECT 29.245 51.935 29.780 52.555 ;
        RECT 29.985 51.765 31.195 52.855 ;
        RECT 31.365 51.765 31.655 52.930 ;
        RECT 33.645 52.855 35.335 53.375 ;
        RECT 35.505 53.025 36.025 53.565 ;
        RECT 37.375 53.405 37.605 54.025 ;
        RECT 37.805 53.755 38.030 54.135 ;
        RECT 38.200 53.925 38.530 54.315 ;
        RECT 37.805 53.575 38.135 53.755 ;
        RECT 36.195 52.855 36.715 53.395 ;
        RECT 36.900 53.075 37.195 53.405 ;
        RECT 37.375 53.075 37.790 53.405 ;
        RECT 37.960 52.905 38.135 53.575 ;
        RECT 38.305 53.075 38.545 53.725 ;
        RECT 38.725 53.545 41.315 54.315 ;
        RECT 38.725 53.025 39.935 53.545 ;
        RECT 41.495 53.505 41.765 54.315 ;
        RECT 41.935 53.505 42.265 54.145 ;
        RECT 42.435 53.505 42.675 54.315 ;
        RECT 42.865 53.545 44.535 54.315 ;
        RECT 44.740 53.575 45.355 54.145 ;
        RECT 45.525 53.805 45.740 54.315 ;
        RECT 45.970 53.805 46.250 54.135 ;
        RECT 46.430 53.805 46.670 54.315 ;
        RECT 31.825 51.765 35.335 52.855 ;
        RECT 35.505 51.765 36.715 52.855 ;
        RECT 36.895 52.545 37.790 52.875 ;
        RECT 37.960 52.715 38.545 52.905 ;
        RECT 40.105 52.855 41.315 53.375 ;
        RECT 41.485 53.075 41.835 53.325 ;
        RECT 42.005 52.905 42.175 53.505 ;
        RECT 42.345 53.075 42.695 53.325 ;
        RECT 42.865 53.025 43.615 53.545 ;
        RECT 36.895 52.375 38.100 52.545 ;
        RECT 36.895 51.945 37.225 52.375 ;
        RECT 37.405 51.765 37.600 52.205 ;
        RECT 37.770 51.945 38.100 52.375 ;
        RECT 38.270 51.945 38.545 52.715 ;
        RECT 38.725 51.765 41.315 52.855 ;
        RECT 41.495 51.765 41.825 52.905 ;
        RECT 42.005 52.735 42.685 52.905 ;
        RECT 43.785 52.855 44.535 53.375 ;
        RECT 42.355 51.950 42.685 52.735 ;
        RECT 42.865 51.765 44.535 52.855 ;
        RECT 44.740 52.555 45.055 53.575 ;
        RECT 45.225 52.905 45.395 53.405 ;
        RECT 45.645 53.075 45.910 53.635 ;
        RECT 46.080 52.905 46.250 53.805 ;
        RECT 46.420 53.075 46.775 53.635 ;
        RECT 47.095 53.445 47.265 54.010 ;
        RECT 47.455 53.785 47.685 54.090 ;
        RECT 47.855 53.955 48.185 54.315 ;
        RECT 48.380 53.785 48.670 54.135 ;
        RECT 47.455 53.615 48.670 53.785 ;
        RECT 48.845 53.770 54.190 54.315 ;
        RECT 47.095 53.275 47.615 53.445 ;
        RECT 45.225 52.735 46.650 52.905 ;
        RECT 47.010 52.745 47.255 53.105 ;
        RECT 47.445 52.895 47.615 53.275 ;
        RECT 47.785 53.075 48.170 53.405 ;
        RECT 48.350 53.295 48.610 53.405 ;
        RECT 48.350 53.125 48.615 53.295 ;
        RECT 48.350 53.075 48.610 53.125 ;
        RECT 44.740 51.935 45.275 52.555 ;
        RECT 45.445 51.765 45.775 52.565 ;
        RECT 46.260 52.560 46.650 52.735 ;
        RECT 47.445 52.615 47.795 52.895 ;
        RECT 47.010 51.765 47.265 52.565 ;
        RECT 47.465 51.935 47.795 52.615 ;
        RECT 47.975 52.025 48.170 53.075 ;
        RECT 50.430 52.940 50.770 53.770 ;
        RECT 54.365 53.545 56.955 54.315 ;
        RECT 57.125 53.590 57.415 54.315 ;
        RECT 58.550 53.855 58.815 54.315 ;
        RECT 59.185 53.675 59.355 54.145 ;
        RECT 59.605 53.855 59.775 54.315 ;
        RECT 60.025 53.675 60.195 54.145 ;
        RECT 60.445 53.855 60.615 54.315 ;
        RECT 60.865 53.675 61.035 54.145 ;
        RECT 61.205 53.850 61.455 54.315 ;
        RECT 48.350 51.765 48.670 52.905 ;
        RECT 52.250 52.200 52.600 53.450 ;
        RECT 54.365 53.025 55.575 53.545 ;
        RECT 59.185 53.495 61.555 53.675 ;
        RECT 55.745 52.855 56.955 53.375 ;
        RECT 58.525 53.075 61.035 53.325 ;
        RECT 48.845 51.765 54.190 52.200 ;
        RECT 54.365 51.765 56.955 52.855 ;
        RECT 57.125 51.765 57.415 52.930 ;
        RECT 61.205 52.905 61.555 53.495 ;
        RECT 61.725 53.545 65.235 54.315 ;
        RECT 61.725 53.025 63.375 53.545 ;
        RECT 65.870 53.475 66.130 54.315 ;
        RECT 66.305 53.570 66.560 54.145 ;
        RECT 66.730 53.935 67.060 54.315 ;
        RECT 67.275 53.765 67.445 54.145 ;
        RECT 66.730 53.595 67.445 53.765 ;
        RECT 58.550 51.765 58.845 52.905 ;
        RECT 59.105 52.735 61.555 52.905 ;
        RECT 63.545 52.855 65.235 53.375 ;
        RECT 59.105 51.935 59.435 52.735 ;
        RECT 59.605 51.765 59.775 52.565 ;
        RECT 59.945 51.935 60.275 52.735 ;
        RECT 60.785 52.715 61.555 52.735 ;
        RECT 60.445 51.765 60.615 52.565 ;
        RECT 60.785 51.935 61.115 52.715 ;
        RECT 61.285 51.765 61.455 52.225 ;
        RECT 61.725 51.765 65.235 52.855 ;
        RECT 65.870 51.765 66.130 52.915 ;
        RECT 66.305 52.840 66.475 53.570 ;
        RECT 66.730 53.405 66.900 53.595 ;
        RECT 67.710 53.475 67.970 54.315 ;
        RECT 68.145 53.570 68.400 54.145 ;
        RECT 68.570 53.935 68.900 54.315 ;
        RECT 69.115 53.765 69.285 54.145 ;
        RECT 68.570 53.595 69.285 53.765 ;
        RECT 69.545 53.640 69.805 54.145 ;
        RECT 69.985 53.935 70.315 54.315 ;
        RECT 70.495 53.765 70.665 54.145 ;
        RECT 66.645 53.075 66.900 53.405 ;
        RECT 66.730 52.865 66.900 53.075 ;
        RECT 67.180 53.045 67.535 53.415 ;
        RECT 66.305 51.935 66.560 52.840 ;
        RECT 66.730 52.695 67.445 52.865 ;
        RECT 66.730 51.765 67.060 52.525 ;
        RECT 67.275 51.935 67.445 52.695 ;
        RECT 67.710 51.765 67.970 52.915 ;
        RECT 68.145 52.840 68.315 53.570 ;
        RECT 68.570 53.405 68.740 53.595 ;
        RECT 68.485 53.075 68.740 53.405 ;
        RECT 68.570 52.865 68.740 53.075 ;
        RECT 69.020 53.045 69.375 53.415 ;
        RECT 68.145 51.935 68.400 52.840 ;
        RECT 68.570 52.695 69.285 52.865 ;
        RECT 68.570 51.765 68.900 52.525 ;
        RECT 69.115 51.935 69.285 52.695 ;
        RECT 69.545 52.840 69.725 53.640 ;
        RECT 70.000 53.595 70.665 53.765 ;
        RECT 70.000 53.340 70.170 53.595 ;
        RECT 71.130 53.535 71.630 54.145 ;
        RECT 69.895 53.010 70.170 53.340 ;
        RECT 70.395 53.045 70.735 53.415 ;
        RECT 70.925 53.075 71.275 53.325 ;
        RECT 70.000 52.865 70.170 53.010 ;
        RECT 71.460 52.905 71.630 53.535 ;
        RECT 72.260 53.665 72.590 54.145 ;
        RECT 72.760 53.855 72.985 54.315 ;
        RECT 73.155 53.665 73.485 54.145 ;
        RECT 72.260 53.495 73.485 53.665 ;
        RECT 73.675 53.515 73.925 54.315 ;
        RECT 74.095 53.515 74.435 54.145 ;
        RECT 74.695 53.765 74.865 54.055 ;
        RECT 75.035 53.935 75.365 54.315 ;
        RECT 74.695 53.595 75.360 53.765 ;
        RECT 74.205 53.465 74.435 53.515 ;
        RECT 71.800 53.125 72.130 53.325 ;
        RECT 72.300 53.125 72.630 53.325 ;
        RECT 72.800 53.125 73.220 53.325 ;
        RECT 73.395 53.155 74.090 53.325 ;
        RECT 73.395 52.905 73.565 53.155 ;
        RECT 74.260 52.905 74.435 53.465 ;
        RECT 69.545 51.935 69.815 52.840 ;
        RECT 70.000 52.695 70.675 52.865 ;
        RECT 69.985 51.765 70.315 52.525 ;
        RECT 70.495 51.935 70.675 52.695 ;
        RECT 71.130 52.735 73.565 52.905 ;
        RECT 71.130 51.935 71.460 52.735 ;
        RECT 71.630 51.765 71.960 52.565 ;
        RECT 72.260 51.935 72.590 52.735 ;
        RECT 73.235 51.765 73.485 52.565 ;
        RECT 73.755 51.765 73.925 52.905 ;
        RECT 74.095 51.935 74.435 52.905 ;
        RECT 74.610 52.775 74.960 53.425 ;
        RECT 75.130 52.605 75.360 53.595 ;
        RECT 74.695 52.435 75.360 52.605 ;
        RECT 74.695 51.935 74.865 52.435 ;
        RECT 75.035 51.765 75.365 52.265 ;
        RECT 75.535 51.935 75.720 54.055 ;
        RECT 75.975 53.855 76.225 54.315 ;
        RECT 76.395 53.865 76.730 54.035 ;
        RECT 76.925 53.865 77.600 54.035 ;
        RECT 76.395 53.725 76.565 53.865 ;
        RECT 75.890 52.735 76.170 53.685 ;
        RECT 76.340 53.595 76.565 53.725 ;
        RECT 76.340 52.490 76.510 53.595 ;
        RECT 76.735 53.445 77.260 53.665 ;
        RECT 76.680 52.680 76.920 53.275 ;
        RECT 77.090 52.745 77.260 53.445 ;
        RECT 77.430 53.085 77.600 53.865 ;
        RECT 77.920 53.815 78.290 54.315 ;
        RECT 78.470 53.865 78.875 54.035 ;
        RECT 79.045 53.865 79.830 54.035 ;
        RECT 78.470 53.635 78.640 53.865 ;
        RECT 77.810 53.335 78.640 53.635 ;
        RECT 79.025 53.365 79.490 53.695 ;
        RECT 77.810 53.305 78.010 53.335 ;
        RECT 78.130 53.085 78.300 53.155 ;
        RECT 77.430 52.915 78.300 53.085 ;
        RECT 77.790 52.825 78.300 52.915 ;
        RECT 76.340 52.360 76.645 52.490 ;
        RECT 77.090 52.380 77.620 52.745 ;
        RECT 75.960 51.765 76.225 52.225 ;
        RECT 76.395 51.935 76.645 52.360 ;
        RECT 77.790 52.210 77.960 52.825 ;
        RECT 76.855 52.040 77.960 52.210 ;
        RECT 78.130 51.765 78.300 52.565 ;
        RECT 78.470 52.265 78.640 53.335 ;
        RECT 78.810 52.435 79.000 53.155 ;
        RECT 79.170 52.405 79.490 53.365 ;
        RECT 79.660 53.405 79.830 53.865 ;
        RECT 80.105 53.785 80.315 54.315 ;
        RECT 80.575 53.575 80.905 54.100 ;
        RECT 81.075 53.705 81.245 54.315 ;
        RECT 81.415 53.660 81.745 54.095 ;
        RECT 81.415 53.575 81.795 53.660 ;
        RECT 80.705 53.405 80.905 53.575 ;
        RECT 81.570 53.535 81.795 53.575 ;
        RECT 81.965 53.565 83.175 54.315 ;
        RECT 79.660 53.075 80.535 53.405 ;
        RECT 80.705 53.075 81.455 53.405 ;
        RECT 78.470 51.935 78.720 52.265 ;
        RECT 79.660 52.235 79.830 53.075 ;
        RECT 80.705 52.870 80.895 53.075 ;
        RECT 81.625 52.955 81.795 53.535 ;
        RECT 81.580 52.905 81.795 52.955 ;
        RECT 80.000 52.495 80.895 52.870 ;
        RECT 81.405 52.825 81.795 52.905 ;
        RECT 81.965 52.855 82.485 53.395 ;
        RECT 82.655 53.025 83.175 53.565 ;
        RECT 78.945 52.065 79.830 52.235 ;
        RECT 80.010 51.765 80.325 52.265 ;
        RECT 80.555 51.935 80.895 52.495 ;
        RECT 81.065 51.765 81.235 52.775 ;
        RECT 81.405 51.980 81.735 52.825 ;
        RECT 81.965 51.765 83.175 52.855 ;
        RECT 5.520 51.595 83.260 51.765 ;
        RECT 5.605 50.505 6.815 51.595 ;
        RECT 6.985 51.160 12.330 51.595 ;
        RECT 5.605 49.795 6.125 50.335 ;
        RECT 6.295 49.965 6.815 50.505 ;
        RECT 5.605 49.045 6.815 49.795 ;
        RECT 8.570 49.590 8.910 50.420 ;
        RECT 10.390 49.910 10.740 51.160 ;
        RECT 12.505 50.505 15.095 51.595 ;
        RECT 12.505 49.815 13.715 50.335 ;
        RECT 13.885 49.985 15.095 50.505 ;
        RECT 6.985 49.045 12.330 49.590 ;
        RECT 12.505 49.045 15.095 49.815 ;
        RECT 15.735 49.225 15.995 51.415 ;
        RECT 16.165 50.865 16.505 51.595 ;
        RECT 16.685 50.685 16.955 51.415 ;
        RECT 16.185 50.465 16.955 50.685 ;
        RECT 17.135 50.705 17.365 51.415 ;
        RECT 17.535 50.885 17.865 51.595 ;
        RECT 18.035 50.705 18.295 51.415 ;
        RECT 17.135 50.465 18.295 50.705 ;
        RECT 16.185 49.795 16.475 50.465 ;
        RECT 18.485 50.430 18.775 51.595 ;
        RECT 19.405 50.625 19.675 51.395 ;
        RECT 19.845 50.815 20.175 51.595 ;
        RECT 20.380 50.990 20.565 51.395 ;
        RECT 20.735 51.170 21.070 51.595 ;
        RECT 20.380 50.815 21.045 50.990 ;
        RECT 21.495 50.865 21.790 51.595 ;
        RECT 19.405 50.455 20.535 50.625 ;
        RECT 16.655 49.975 17.120 50.285 ;
        RECT 17.300 49.975 17.825 50.285 ;
        RECT 16.185 49.595 17.415 49.795 ;
        RECT 16.255 49.045 16.925 49.415 ;
        RECT 17.105 49.225 17.415 49.595 ;
        RECT 17.595 49.335 17.825 49.975 ;
        RECT 18.005 49.955 18.305 50.285 ;
        RECT 18.005 49.045 18.295 49.775 ;
        RECT 18.485 49.045 18.775 49.770 ;
        RECT 19.405 49.545 19.575 50.455 ;
        RECT 19.745 49.705 20.105 50.285 ;
        RECT 20.285 49.955 20.535 50.455 ;
        RECT 20.705 49.785 21.045 50.815 ;
        RECT 21.960 50.695 22.220 51.420 ;
        RECT 22.390 50.865 22.650 51.595 ;
        RECT 22.820 50.695 23.080 51.420 ;
        RECT 23.250 50.865 23.510 51.595 ;
        RECT 23.680 50.695 23.940 51.420 ;
        RECT 24.110 50.865 24.370 51.595 ;
        RECT 24.540 50.695 24.800 51.420 ;
        RECT 20.360 49.615 21.045 49.785 ;
        RECT 21.490 50.455 24.800 50.695 ;
        RECT 24.970 50.485 25.230 51.595 ;
        RECT 21.490 49.865 22.460 50.455 ;
        RECT 25.400 50.285 25.650 51.420 ;
        RECT 25.830 50.485 26.125 51.595 ;
        RECT 26.365 50.535 26.695 51.380 ;
        RECT 26.865 50.585 27.035 51.595 ;
        RECT 27.205 50.865 27.545 51.425 ;
        RECT 27.775 51.095 28.090 51.595 ;
        RECT 28.270 51.125 29.155 51.295 ;
        RECT 26.305 50.455 26.695 50.535 ;
        RECT 27.205 50.490 28.100 50.865 ;
        RECT 26.305 50.405 26.520 50.455 ;
        RECT 22.630 50.035 25.650 50.285 ;
        RECT 21.490 49.695 24.800 49.865 ;
        RECT 19.405 49.215 19.665 49.545 ;
        RECT 19.875 49.045 20.150 49.525 ;
        RECT 20.360 49.215 20.565 49.615 ;
        RECT 20.735 49.045 21.070 49.445 ;
        RECT 21.490 49.045 21.790 49.525 ;
        RECT 21.960 49.240 22.220 49.695 ;
        RECT 22.390 49.045 22.650 49.525 ;
        RECT 22.820 49.240 23.080 49.695 ;
        RECT 23.250 49.045 23.510 49.525 ;
        RECT 23.680 49.240 23.940 49.695 ;
        RECT 24.110 49.045 24.370 49.525 ;
        RECT 24.540 49.240 24.800 49.695 ;
        RECT 24.970 49.045 25.230 49.570 ;
        RECT 25.400 49.225 25.650 50.035 ;
        RECT 25.820 49.675 26.135 50.285 ;
        RECT 26.305 49.825 26.475 50.405 ;
        RECT 27.205 50.285 27.395 50.490 ;
        RECT 28.270 50.285 28.440 51.125 ;
        RECT 29.380 51.095 29.630 51.425 ;
        RECT 26.645 49.955 27.395 50.285 ;
        RECT 27.565 49.955 28.440 50.285 ;
        RECT 26.305 49.785 26.530 49.825 ;
        RECT 27.195 49.785 27.395 49.955 ;
        RECT 26.305 49.700 26.685 49.785 ;
        RECT 25.830 49.045 26.075 49.505 ;
        RECT 26.355 49.265 26.685 49.700 ;
        RECT 26.855 49.045 27.025 49.655 ;
        RECT 27.195 49.260 27.525 49.785 ;
        RECT 27.785 49.045 27.995 49.575 ;
        RECT 28.270 49.495 28.440 49.955 ;
        RECT 28.610 49.995 28.930 50.955 ;
        RECT 29.100 50.205 29.290 50.925 ;
        RECT 29.460 50.025 29.630 51.095 ;
        RECT 29.800 50.795 29.970 51.595 ;
        RECT 30.140 51.150 31.245 51.320 ;
        RECT 30.140 50.535 30.310 51.150 ;
        RECT 31.455 51.000 31.705 51.425 ;
        RECT 31.875 51.135 32.140 51.595 ;
        RECT 30.480 50.615 31.010 50.980 ;
        RECT 31.455 50.870 31.760 51.000 ;
        RECT 29.800 50.445 30.310 50.535 ;
        RECT 29.800 50.275 30.670 50.445 ;
        RECT 29.800 50.205 29.970 50.275 ;
        RECT 30.090 50.025 30.290 50.055 ;
        RECT 28.610 49.665 29.075 49.995 ;
        RECT 29.460 49.725 30.290 50.025 ;
        RECT 29.460 49.495 29.630 49.725 ;
        RECT 28.270 49.325 29.055 49.495 ;
        RECT 29.225 49.325 29.630 49.495 ;
        RECT 29.810 49.045 30.180 49.545 ;
        RECT 30.500 49.495 30.670 50.275 ;
        RECT 30.840 49.915 31.010 50.615 ;
        RECT 31.180 50.085 31.420 50.680 ;
        RECT 30.840 49.695 31.365 49.915 ;
        RECT 31.590 49.765 31.760 50.870 ;
        RECT 31.535 49.635 31.760 49.765 ;
        RECT 31.930 49.675 32.210 50.625 ;
        RECT 31.535 49.495 31.705 49.635 ;
        RECT 30.500 49.325 31.175 49.495 ;
        RECT 31.370 49.325 31.705 49.495 ;
        RECT 31.875 49.045 32.125 49.505 ;
        RECT 32.380 49.305 32.565 51.425 ;
        RECT 32.735 51.095 33.065 51.595 ;
        RECT 33.235 50.925 33.405 51.425 ;
        RECT 33.665 51.085 33.925 51.595 ;
        RECT 32.740 50.755 33.405 50.925 ;
        RECT 32.740 49.765 32.970 50.755 ;
        RECT 33.140 49.935 33.490 50.585 ;
        RECT 33.665 50.035 34.005 50.915 ;
        RECT 34.175 50.205 34.345 51.425 ;
        RECT 34.585 51.090 35.200 51.595 ;
        RECT 34.585 50.555 34.835 50.920 ;
        RECT 35.005 50.915 35.200 51.090 ;
        RECT 35.370 51.085 35.845 51.425 ;
        RECT 36.015 51.050 36.230 51.595 ;
        RECT 35.005 50.725 35.335 50.915 ;
        RECT 35.555 50.555 36.270 50.850 ;
        RECT 36.440 50.725 36.715 51.425 ;
        RECT 37.000 50.965 37.285 51.425 ;
        RECT 37.455 51.135 37.725 51.595 ;
        RECT 37.000 50.745 37.955 50.965 ;
        RECT 34.585 50.385 36.375 50.555 ;
        RECT 34.175 49.955 34.970 50.205 ;
        RECT 34.175 49.865 34.425 49.955 ;
        RECT 32.740 49.595 33.405 49.765 ;
        RECT 32.735 49.045 33.065 49.425 ;
        RECT 33.235 49.305 33.405 49.595 ;
        RECT 33.665 49.045 33.925 49.865 ;
        RECT 34.095 49.445 34.425 49.865 ;
        RECT 35.140 49.530 35.395 50.385 ;
        RECT 34.605 49.265 35.395 49.530 ;
        RECT 35.565 49.685 35.975 50.205 ;
        RECT 36.145 49.955 36.375 50.385 ;
        RECT 36.545 49.695 36.715 50.725 ;
        RECT 36.885 50.015 37.575 50.575 ;
        RECT 37.745 49.845 37.955 50.745 ;
        RECT 35.565 49.265 35.765 49.685 ;
        RECT 35.955 49.045 36.285 49.505 ;
        RECT 36.455 49.215 36.715 49.695 ;
        RECT 37.000 49.675 37.955 49.845 ;
        RECT 38.125 50.575 38.525 51.425 ;
        RECT 38.715 50.965 38.995 51.425 ;
        RECT 39.515 51.135 39.840 51.595 ;
        RECT 38.715 50.745 39.840 50.965 ;
        RECT 38.125 50.015 39.220 50.575 ;
        RECT 39.390 50.285 39.840 50.745 ;
        RECT 40.010 50.455 40.395 51.425 ;
        RECT 40.575 50.645 40.850 51.415 ;
        RECT 41.020 50.985 41.350 51.415 ;
        RECT 41.520 51.155 41.715 51.595 ;
        RECT 41.895 50.985 42.225 51.415 ;
        RECT 41.020 50.815 42.225 50.985 ;
        RECT 40.575 50.455 41.160 50.645 ;
        RECT 41.330 50.485 42.225 50.815 ;
        RECT 42.875 50.455 43.205 51.595 ;
        RECT 43.735 50.625 44.065 51.410 ;
        RECT 43.385 50.455 44.065 50.625 ;
        RECT 37.000 49.215 37.285 49.675 ;
        RECT 37.455 49.045 37.725 49.505 ;
        RECT 38.125 49.215 38.525 50.015 ;
        RECT 39.390 49.955 39.945 50.285 ;
        RECT 39.390 49.845 39.840 49.955 ;
        RECT 38.715 49.675 39.840 49.845 ;
        RECT 40.115 49.785 40.395 50.455 ;
        RECT 38.715 49.215 38.995 49.675 ;
        RECT 39.515 49.045 39.840 49.505 ;
        RECT 40.010 49.215 40.395 49.785 ;
        RECT 40.575 49.635 40.815 50.285 ;
        RECT 40.985 49.785 41.160 50.455 ;
        RECT 41.330 49.955 41.745 50.285 ;
        RECT 41.925 49.955 42.220 50.285 ;
        RECT 42.865 50.035 43.215 50.285 ;
        RECT 40.985 49.605 41.315 49.785 ;
        RECT 40.590 49.045 40.920 49.435 ;
        RECT 41.090 49.225 41.315 49.605 ;
        RECT 41.515 49.335 41.745 49.955 ;
        RECT 43.385 49.855 43.555 50.455 ;
        RECT 44.245 50.430 44.535 51.595 ;
        RECT 44.705 50.455 45.090 51.425 ;
        RECT 45.260 51.135 45.585 51.595 ;
        RECT 46.105 50.965 46.385 51.425 ;
        RECT 45.260 50.745 46.385 50.965 ;
        RECT 43.725 50.035 44.075 50.285 ;
        RECT 41.925 49.045 42.225 49.775 ;
        RECT 42.875 49.045 43.145 49.855 ;
        RECT 43.315 49.215 43.645 49.855 ;
        RECT 43.815 49.045 44.055 49.855 ;
        RECT 44.705 49.785 44.985 50.455 ;
        RECT 45.260 50.285 45.710 50.745 ;
        RECT 46.575 50.575 46.975 51.425 ;
        RECT 47.375 51.135 47.645 51.595 ;
        RECT 47.815 50.965 48.100 51.425 ;
        RECT 45.155 49.955 45.710 50.285 ;
        RECT 45.880 50.015 46.975 50.575 ;
        RECT 45.260 49.845 45.710 49.955 ;
        RECT 44.245 49.045 44.535 49.770 ;
        RECT 44.705 49.215 45.090 49.785 ;
        RECT 45.260 49.675 46.385 49.845 ;
        RECT 45.260 49.045 45.585 49.505 ;
        RECT 46.105 49.215 46.385 49.675 ;
        RECT 46.575 49.215 46.975 50.015 ;
        RECT 47.145 50.745 48.100 50.965 ;
        RECT 47.145 49.845 47.355 50.745 ;
        RECT 47.525 50.015 48.215 50.575 ;
        RECT 49.305 50.455 49.690 51.425 ;
        RECT 49.860 51.135 50.185 51.595 ;
        RECT 50.705 50.965 50.985 51.425 ;
        RECT 49.860 50.745 50.985 50.965 ;
        RECT 47.145 49.675 48.100 49.845 ;
        RECT 47.375 49.045 47.645 49.505 ;
        RECT 47.815 49.215 48.100 49.675 ;
        RECT 49.305 49.785 49.585 50.455 ;
        RECT 49.860 50.285 50.310 50.745 ;
        RECT 51.175 50.575 51.575 51.425 ;
        RECT 51.975 51.135 52.245 51.595 ;
        RECT 52.415 50.965 52.700 51.425 ;
        RECT 49.755 49.955 50.310 50.285 ;
        RECT 50.480 50.015 51.575 50.575 ;
        RECT 49.860 49.845 50.310 49.955 ;
        RECT 49.305 49.215 49.690 49.785 ;
        RECT 49.860 49.675 50.985 49.845 ;
        RECT 49.860 49.045 50.185 49.505 ;
        RECT 50.705 49.215 50.985 49.675 ;
        RECT 51.175 49.215 51.575 50.015 ;
        RECT 51.745 50.745 52.700 50.965 ;
        RECT 51.745 49.845 51.955 50.745 ;
        RECT 52.125 50.015 52.815 50.575 ;
        RECT 52.985 50.505 55.575 51.595 ;
        RECT 55.835 50.925 56.005 51.425 ;
        RECT 56.175 51.095 56.505 51.595 ;
        RECT 55.835 50.755 56.500 50.925 ;
        RECT 51.745 49.675 52.700 49.845 ;
        RECT 51.975 49.045 52.245 49.505 ;
        RECT 52.415 49.215 52.700 49.675 ;
        RECT 52.985 49.815 54.195 50.335 ;
        RECT 54.365 49.985 55.575 50.505 ;
        RECT 55.750 49.935 56.100 50.585 ;
        RECT 52.985 49.045 55.575 49.815 ;
        RECT 56.270 49.765 56.500 50.755 ;
        RECT 55.835 49.595 56.500 49.765 ;
        RECT 55.835 49.305 56.005 49.595 ;
        RECT 56.175 49.045 56.505 49.425 ;
        RECT 56.675 49.305 56.860 51.425 ;
        RECT 57.100 51.135 57.365 51.595 ;
        RECT 57.535 51.000 57.785 51.425 ;
        RECT 57.995 51.150 59.100 51.320 ;
        RECT 57.480 50.870 57.785 51.000 ;
        RECT 57.030 49.675 57.310 50.625 ;
        RECT 57.480 49.765 57.650 50.870 ;
        RECT 57.820 50.085 58.060 50.680 ;
        RECT 58.230 50.615 58.760 50.980 ;
        RECT 58.230 49.915 58.400 50.615 ;
        RECT 58.930 50.535 59.100 51.150 ;
        RECT 59.270 50.795 59.440 51.595 ;
        RECT 59.610 51.095 59.860 51.425 ;
        RECT 60.085 51.125 60.970 51.295 ;
        RECT 58.930 50.445 59.440 50.535 ;
        RECT 57.480 49.635 57.705 49.765 ;
        RECT 57.875 49.695 58.400 49.915 ;
        RECT 58.570 50.275 59.440 50.445 ;
        RECT 57.115 49.045 57.365 49.505 ;
        RECT 57.535 49.495 57.705 49.635 ;
        RECT 58.570 49.495 58.740 50.275 ;
        RECT 59.270 50.205 59.440 50.275 ;
        RECT 58.950 50.025 59.150 50.055 ;
        RECT 59.610 50.025 59.780 51.095 ;
        RECT 59.950 50.205 60.140 50.925 ;
        RECT 58.950 49.725 59.780 50.025 ;
        RECT 60.310 49.995 60.630 50.955 ;
        RECT 57.535 49.325 57.870 49.495 ;
        RECT 58.065 49.325 58.740 49.495 ;
        RECT 59.060 49.045 59.430 49.545 ;
        RECT 59.610 49.495 59.780 49.725 ;
        RECT 60.165 49.665 60.630 49.995 ;
        RECT 60.800 50.285 60.970 51.125 ;
        RECT 61.150 51.095 61.465 51.595 ;
        RECT 61.695 50.865 62.035 51.425 ;
        RECT 61.140 50.490 62.035 50.865 ;
        RECT 62.205 50.585 62.375 51.595 ;
        RECT 61.845 50.285 62.035 50.490 ;
        RECT 62.545 50.535 62.875 51.380 ;
        RECT 62.545 50.455 62.935 50.535 ;
        RECT 63.105 50.505 64.315 51.595 ;
        RECT 62.720 50.405 62.935 50.455 ;
        RECT 60.800 49.955 61.675 50.285 ;
        RECT 61.845 49.955 62.595 50.285 ;
        RECT 60.800 49.495 60.970 49.955 ;
        RECT 61.845 49.785 62.045 49.955 ;
        RECT 62.765 49.825 62.935 50.405 ;
        RECT 62.710 49.785 62.935 49.825 ;
        RECT 59.610 49.325 60.015 49.495 ;
        RECT 60.185 49.325 60.970 49.495 ;
        RECT 61.245 49.045 61.455 49.575 ;
        RECT 61.715 49.260 62.045 49.785 ;
        RECT 62.555 49.700 62.935 49.785 ;
        RECT 63.105 49.795 63.625 50.335 ;
        RECT 63.795 49.965 64.315 50.505 ;
        RECT 64.490 50.445 64.750 51.595 ;
        RECT 64.925 50.520 65.180 51.425 ;
        RECT 65.350 50.835 65.680 51.595 ;
        RECT 65.895 50.665 66.065 51.425 ;
        RECT 62.215 49.045 62.385 49.655 ;
        RECT 62.555 49.265 62.885 49.700 ;
        RECT 63.105 49.045 64.315 49.795 ;
        RECT 64.490 49.045 64.750 49.885 ;
        RECT 64.925 49.790 65.095 50.520 ;
        RECT 65.350 50.495 66.065 50.665 ;
        RECT 65.350 50.285 65.520 50.495 ;
        RECT 66.325 50.455 66.665 51.425 ;
        RECT 66.835 50.455 67.005 51.595 ;
        RECT 67.275 50.795 67.525 51.595 ;
        RECT 68.170 50.625 68.500 51.425 ;
        RECT 68.800 50.795 69.130 51.595 ;
        RECT 69.300 50.625 69.630 51.425 ;
        RECT 67.195 50.455 69.630 50.625 ;
        RECT 65.265 49.955 65.520 50.285 ;
        RECT 64.925 49.215 65.180 49.790 ;
        RECT 65.350 49.765 65.520 49.955 ;
        RECT 65.800 49.945 66.155 50.315 ;
        RECT 66.325 49.845 66.500 50.455 ;
        RECT 67.195 50.205 67.365 50.455 ;
        RECT 66.670 50.035 67.365 50.205 ;
        RECT 67.540 50.035 67.960 50.235 ;
        RECT 68.130 50.035 68.460 50.235 ;
        RECT 68.630 50.035 68.960 50.235 ;
        RECT 65.350 49.595 66.065 49.765 ;
        RECT 65.350 49.045 65.680 49.425 ;
        RECT 65.895 49.215 66.065 49.595 ;
        RECT 66.325 49.215 66.665 49.845 ;
        RECT 66.835 49.045 67.085 49.845 ;
        RECT 67.275 49.695 68.500 49.865 ;
        RECT 67.275 49.215 67.605 49.695 ;
        RECT 67.775 49.045 68.000 49.505 ;
        RECT 68.170 49.215 68.500 49.695 ;
        RECT 69.130 49.825 69.300 50.455 ;
        RECT 70.005 50.430 70.295 51.595 ;
        RECT 70.555 50.925 70.725 51.425 ;
        RECT 70.895 51.095 71.225 51.595 ;
        RECT 70.555 50.755 71.220 50.925 ;
        RECT 69.485 50.035 69.835 50.285 ;
        RECT 70.470 49.935 70.820 50.585 ;
        RECT 69.130 49.215 69.630 49.825 ;
        RECT 70.005 49.045 70.295 49.770 ;
        RECT 70.990 49.765 71.220 50.755 ;
        RECT 70.555 49.595 71.220 49.765 ;
        RECT 70.555 49.305 70.725 49.595 ;
        RECT 70.895 49.045 71.225 49.425 ;
        RECT 71.395 49.305 71.580 51.425 ;
        RECT 71.820 51.135 72.085 51.595 ;
        RECT 72.255 51.000 72.505 51.425 ;
        RECT 72.715 51.150 73.820 51.320 ;
        RECT 72.200 50.870 72.505 51.000 ;
        RECT 71.750 49.675 72.030 50.625 ;
        RECT 72.200 49.765 72.370 50.870 ;
        RECT 72.540 50.085 72.780 50.680 ;
        RECT 72.950 50.615 73.480 50.980 ;
        RECT 72.950 49.915 73.120 50.615 ;
        RECT 73.650 50.535 73.820 51.150 ;
        RECT 73.990 50.795 74.160 51.595 ;
        RECT 74.330 51.095 74.580 51.425 ;
        RECT 74.805 51.125 75.690 51.295 ;
        RECT 73.650 50.445 74.160 50.535 ;
        RECT 72.200 49.635 72.425 49.765 ;
        RECT 72.595 49.695 73.120 49.915 ;
        RECT 73.290 50.275 74.160 50.445 ;
        RECT 71.835 49.045 72.085 49.505 ;
        RECT 72.255 49.495 72.425 49.635 ;
        RECT 73.290 49.495 73.460 50.275 ;
        RECT 73.990 50.205 74.160 50.275 ;
        RECT 73.670 50.025 73.870 50.055 ;
        RECT 74.330 50.025 74.500 51.095 ;
        RECT 74.670 50.205 74.860 50.925 ;
        RECT 73.670 49.725 74.500 50.025 ;
        RECT 75.030 49.995 75.350 50.955 ;
        RECT 72.255 49.325 72.590 49.495 ;
        RECT 72.785 49.325 73.460 49.495 ;
        RECT 73.780 49.045 74.150 49.545 ;
        RECT 74.330 49.495 74.500 49.725 ;
        RECT 74.885 49.665 75.350 49.995 ;
        RECT 75.520 50.285 75.690 51.125 ;
        RECT 75.870 51.095 76.185 51.595 ;
        RECT 76.415 50.865 76.755 51.425 ;
        RECT 75.860 50.490 76.755 50.865 ;
        RECT 76.925 50.585 77.095 51.595 ;
        RECT 76.565 50.285 76.755 50.490 ;
        RECT 77.265 50.535 77.595 51.380 ;
        RECT 77.860 50.805 78.395 51.425 ;
        RECT 77.265 50.455 77.655 50.535 ;
        RECT 77.440 50.405 77.655 50.455 ;
        RECT 75.520 49.955 76.395 50.285 ;
        RECT 76.565 49.955 77.315 50.285 ;
        RECT 75.520 49.495 75.690 49.955 ;
        RECT 76.565 49.785 76.765 49.955 ;
        RECT 77.485 49.825 77.655 50.405 ;
        RECT 77.430 49.785 77.655 49.825 ;
        RECT 74.330 49.325 74.735 49.495 ;
        RECT 74.905 49.325 75.690 49.495 ;
        RECT 75.965 49.045 76.175 49.575 ;
        RECT 76.435 49.260 76.765 49.785 ;
        RECT 77.275 49.700 77.655 49.785 ;
        RECT 77.860 49.785 78.175 50.805 ;
        RECT 78.565 50.795 78.895 51.595 ;
        RECT 79.380 50.625 79.770 50.800 ;
        RECT 78.345 50.455 79.770 50.625 ;
        RECT 80.215 50.665 80.385 51.425 ;
        RECT 80.600 50.835 80.930 51.595 ;
        RECT 80.215 50.495 80.930 50.665 ;
        RECT 81.100 50.520 81.355 51.425 ;
        RECT 78.345 49.955 78.515 50.455 ;
        RECT 76.935 49.045 77.105 49.655 ;
        RECT 77.275 49.265 77.605 49.700 ;
        RECT 77.860 49.215 78.475 49.785 ;
        RECT 78.765 49.725 79.030 50.285 ;
        RECT 79.200 49.555 79.370 50.455 ;
        RECT 79.540 49.725 79.895 50.285 ;
        RECT 80.125 49.945 80.480 50.315 ;
        RECT 80.760 50.285 80.930 50.495 ;
        RECT 80.760 49.955 81.015 50.285 ;
        RECT 80.760 49.765 80.930 49.955 ;
        RECT 81.185 49.790 81.355 50.520 ;
        RECT 81.530 50.445 81.790 51.595 ;
        RECT 81.965 50.505 83.175 51.595 ;
        RECT 81.965 49.965 82.485 50.505 ;
        RECT 80.215 49.595 80.930 49.765 ;
        RECT 78.645 49.045 78.860 49.555 ;
        RECT 79.090 49.225 79.370 49.555 ;
        RECT 79.550 49.045 79.790 49.555 ;
        RECT 80.215 49.215 80.385 49.595 ;
        RECT 80.600 49.045 80.930 49.425 ;
        RECT 81.100 49.215 81.355 49.790 ;
        RECT 81.530 49.045 81.790 49.885 ;
        RECT 82.655 49.795 83.175 50.335 ;
        RECT 81.965 49.045 83.175 49.795 ;
        RECT 5.520 48.875 83.260 49.045 ;
        RECT 5.605 48.125 6.815 48.875 ;
        RECT 6.985 48.330 12.330 48.875 ;
        RECT 5.605 47.585 6.125 48.125 ;
        RECT 6.295 47.415 6.815 47.955 ;
        RECT 8.570 47.500 8.910 48.330 ;
        RECT 12.505 48.125 13.715 48.875 ;
        RECT 13.890 48.345 14.180 48.695 ;
        RECT 14.375 48.515 14.705 48.875 ;
        RECT 14.875 48.345 15.105 48.650 ;
        RECT 13.890 48.175 15.105 48.345 ;
        RECT 15.295 48.535 15.465 48.570 ;
        RECT 15.295 48.365 15.495 48.535 ;
        RECT 5.605 46.325 6.815 47.415 ;
        RECT 10.390 46.760 10.740 48.010 ;
        RECT 12.505 47.585 13.025 48.125 ;
        RECT 15.295 48.005 15.465 48.365 ;
        RECT 13.195 47.415 13.715 47.955 ;
        RECT 13.950 47.855 14.210 47.965 ;
        RECT 13.945 47.685 14.210 47.855 ;
        RECT 13.950 47.635 14.210 47.685 ;
        RECT 14.390 47.635 14.775 47.965 ;
        RECT 14.945 47.835 15.465 48.005 ;
        RECT 15.725 48.135 16.190 48.680 ;
        RECT 6.985 46.325 12.330 46.760 ;
        RECT 12.505 46.325 13.715 47.415 ;
        RECT 13.890 46.325 14.210 47.465 ;
        RECT 14.390 46.585 14.585 47.635 ;
        RECT 14.945 47.455 15.115 47.835 ;
        RECT 14.765 47.175 15.115 47.455 ;
        RECT 15.305 47.305 15.550 47.665 ;
        RECT 15.725 47.175 15.895 48.135 ;
        RECT 16.695 48.055 16.865 48.875 ;
        RECT 17.035 48.225 17.365 48.705 ;
        RECT 17.535 48.485 17.885 48.875 ;
        RECT 18.055 48.305 18.285 48.705 ;
        RECT 17.775 48.225 18.285 48.305 ;
        RECT 17.035 48.135 18.285 48.225 ;
        RECT 18.455 48.135 18.775 48.615 ;
        RECT 19.030 48.305 19.205 48.705 ;
        RECT 19.375 48.495 19.705 48.875 ;
        RECT 19.950 48.375 20.180 48.705 ;
        RECT 19.030 48.135 19.660 48.305 ;
        RECT 17.035 48.055 17.945 48.135 ;
        RECT 16.065 47.515 16.310 47.965 ;
        RECT 16.570 47.685 17.265 47.885 ;
        RECT 17.435 47.715 18.035 47.885 ;
        RECT 17.435 47.515 17.605 47.715 ;
        RECT 18.265 47.545 18.435 47.965 ;
        RECT 16.065 47.345 17.605 47.515 ;
        RECT 17.775 47.375 18.435 47.545 ;
        RECT 17.775 47.175 17.945 47.375 ;
        RECT 18.605 47.205 18.775 48.135 ;
        RECT 19.490 47.965 19.660 48.135 ;
        RECT 18.945 47.285 19.310 47.965 ;
        RECT 19.490 47.635 19.840 47.965 ;
        RECT 14.765 46.495 15.095 47.175 ;
        RECT 15.295 46.325 15.550 47.125 ;
        RECT 15.725 47.005 17.945 47.175 ;
        RECT 18.115 47.005 18.775 47.205 ;
        RECT 19.490 47.115 19.660 47.635 ;
        RECT 15.725 46.325 16.025 46.835 ;
        RECT 16.195 46.495 16.525 47.005 ;
        RECT 18.115 46.835 18.285 47.005 ;
        RECT 19.030 46.945 19.660 47.115 ;
        RECT 20.010 47.085 20.180 48.375 ;
        RECT 20.380 47.265 20.660 48.540 ;
        RECT 20.885 48.535 21.155 48.540 ;
        RECT 20.845 48.365 21.155 48.535 ;
        RECT 21.615 48.495 21.945 48.875 ;
        RECT 22.115 48.620 22.450 48.665 ;
        RECT 20.885 47.265 21.155 48.365 ;
        RECT 21.345 47.265 21.685 48.295 ;
        RECT 22.115 48.155 22.455 48.620 ;
        RECT 23.595 48.415 23.900 48.875 ;
        RECT 24.070 48.245 24.400 48.705 ;
        RECT 24.570 48.415 24.740 48.875 ;
        RECT 24.910 48.245 25.240 48.705 ;
        RECT 25.410 48.415 25.580 48.875 ;
        RECT 25.750 48.245 26.080 48.705 ;
        RECT 26.250 48.415 26.420 48.875 ;
        RECT 26.590 48.245 26.920 48.705 ;
        RECT 27.090 48.415 27.345 48.875 ;
        RECT 21.855 47.635 22.115 47.965 ;
        RECT 21.855 47.085 22.025 47.635 ;
        RECT 22.285 47.465 22.455 48.155 ;
        RECT 16.695 46.325 17.325 46.835 ;
        RECT 17.905 46.665 18.285 46.835 ;
        RECT 18.455 46.325 18.755 46.835 ;
        RECT 19.030 46.495 19.205 46.945 ;
        RECT 20.010 46.915 22.025 47.085 ;
        RECT 19.375 46.325 19.705 46.765 ;
        RECT 20.010 46.495 20.180 46.915 ;
        RECT 20.415 46.325 21.085 46.735 ;
        RECT 21.300 46.495 21.470 46.915 ;
        RECT 21.670 46.325 22.000 46.735 ;
        RECT 22.195 46.495 22.455 47.465 ;
        RECT 23.545 48.055 27.515 48.245 ;
        RECT 23.545 47.465 23.865 48.055 ;
        RECT 24.065 47.635 26.920 47.885 ;
        RECT 27.170 47.465 27.515 48.055 ;
        RECT 23.545 47.295 27.515 47.465 ;
        RECT 27.705 48.185 27.945 48.705 ;
        RECT 28.115 48.380 28.510 48.875 ;
        RECT 29.075 48.545 29.245 48.690 ;
        RECT 28.870 48.350 29.245 48.545 ;
        RECT 27.705 47.515 27.880 48.185 ;
        RECT 28.870 48.015 29.040 48.350 ;
        RECT 29.525 48.305 29.765 48.680 ;
        RECT 29.935 48.370 30.270 48.875 ;
        RECT 29.525 48.155 29.745 48.305 ;
        RECT 28.055 47.655 29.040 48.015 ;
        RECT 29.210 47.825 29.745 48.155 ;
        RECT 28.055 47.635 29.340 47.655 ;
        RECT 27.705 47.380 27.915 47.515 ;
        RECT 28.480 47.485 29.340 47.635 ;
        RECT 23.600 46.325 23.900 47.125 ;
        RECT 24.070 46.495 24.400 47.295 ;
        RECT 24.570 46.325 24.740 47.125 ;
        RECT 24.910 46.495 25.240 47.295 ;
        RECT 25.410 46.325 25.580 47.125 ;
        RECT 25.750 46.495 26.080 47.295 ;
        RECT 26.250 46.325 26.420 47.125 ;
        RECT 26.590 46.495 26.920 47.295 ;
        RECT 27.090 46.325 27.345 47.125 ;
        RECT 27.705 46.595 28.010 47.380 ;
        RECT 28.185 47.005 28.880 47.315 ;
        RECT 28.190 46.325 28.875 46.795 ;
        RECT 29.055 46.540 29.340 47.485 ;
        RECT 29.510 47.175 29.745 47.825 ;
        RECT 29.915 47.345 30.215 48.195 ;
        RECT 31.365 48.150 31.655 48.875 ;
        RECT 31.825 48.225 32.085 48.705 ;
        RECT 32.255 48.335 32.505 48.875 ;
        RECT 29.510 46.945 30.185 47.175 ;
        RECT 29.515 46.325 29.845 46.775 ;
        RECT 30.015 46.515 30.185 46.945 ;
        RECT 31.365 46.325 31.655 47.490 ;
        RECT 31.825 47.195 31.995 48.225 ;
        RECT 32.675 48.195 32.895 48.655 ;
        RECT 32.645 48.170 32.895 48.195 ;
        RECT 32.165 47.575 32.395 47.970 ;
        RECT 32.565 47.745 32.895 48.170 ;
        RECT 33.065 48.495 33.955 48.665 ;
        RECT 33.065 47.770 33.235 48.495 ;
        RECT 33.405 47.940 33.955 48.325 ;
        RECT 34.635 48.220 34.965 48.655 ;
        RECT 35.135 48.265 35.305 48.875 ;
        RECT 34.585 48.135 34.965 48.220 ;
        RECT 35.475 48.135 35.805 48.660 ;
        RECT 36.065 48.345 36.275 48.875 ;
        RECT 36.550 48.425 37.335 48.595 ;
        RECT 37.505 48.425 37.910 48.595 ;
        RECT 34.585 48.095 34.810 48.135 ;
        RECT 33.065 47.700 33.955 47.770 ;
        RECT 33.060 47.675 33.955 47.700 ;
        RECT 33.050 47.660 33.955 47.675 ;
        RECT 33.045 47.645 33.955 47.660 ;
        RECT 33.035 47.640 33.955 47.645 ;
        RECT 33.030 47.630 33.955 47.640 ;
        RECT 33.025 47.620 33.955 47.630 ;
        RECT 33.015 47.615 33.955 47.620 ;
        RECT 33.005 47.605 33.955 47.615 ;
        RECT 32.995 47.600 33.955 47.605 ;
        RECT 32.995 47.595 33.330 47.600 ;
        RECT 32.980 47.590 33.330 47.595 ;
        RECT 32.965 47.580 33.330 47.590 ;
        RECT 32.940 47.575 33.330 47.580 ;
        RECT 32.165 47.570 33.330 47.575 ;
        RECT 32.165 47.535 33.300 47.570 ;
        RECT 32.165 47.510 33.265 47.535 ;
        RECT 32.165 47.480 33.235 47.510 ;
        RECT 32.165 47.450 33.215 47.480 ;
        RECT 32.165 47.420 33.195 47.450 ;
        RECT 32.165 47.410 33.125 47.420 ;
        RECT 32.165 47.400 33.100 47.410 ;
        RECT 32.165 47.385 33.080 47.400 ;
        RECT 32.165 47.370 33.060 47.385 ;
        RECT 32.270 47.360 33.055 47.370 ;
        RECT 32.270 47.325 33.040 47.360 ;
        RECT 31.825 46.495 32.100 47.195 ;
        RECT 32.270 47.075 33.025 47.325 ;
        RECT 33.195 47.005 33.525 47.250 ;
        RECT 33.695 47.150 33.955 47.600 ;
        RECT 34.585 47.515 34.755 48.095 ;
        RECT 35.475 47.965 35.675 48.135 ;
        RECT 36.550 47.965 36.720 48.425 ;
        RECT 34.925 47.635 35.675 47.965 ;
        RECT 35.845 47.635 36.720 47.965 ;
        RECT 34.585 47.465 34.800 47.515 ;
        RECT 34.585 47.385 34.975 47.465 ;
        RECT 33.340 46.980 33.525 47.005 ;
        RECT 33.340 46.880 33.955 46.980 ;
        RECT 32.270 46.325 32.525 46.870 ;
        RECT 32.695 46.495 33.175 46.835 ;
        RECT 33.350 46.325 33.955 46.880 ;
        RECT 34.645 46.540 34.975 47.385 ;
        RECT 35.485 47.430 35.675 47.635 ;
        RECT 35.145 46.325 35.315 47.335 ;
        RECT 35.485 47.055 36.380 47.430 ;
        RECT 35.485 46.495 35.825 47.055 ;
        RECT 36.055 46.325 36.370 46.825 ;
        RECT 36.550 46.795 36.720 47.635 ;
        RECT 36.890 47.925 37.355 48.255 ;
        RECT 37.740 48.195 37.910 48.425 ;
        RECT 38.090 48.375 38.460 48.875 ;
        RECT 38.780 48.425 39.455 48.595 ;
        RECT 39.650 48.425 39.985 48.595 ;
        RECT 36.890 46.965 37.210 47.925 ;
        RECT 37.740 47.895 38.570 48.195 ;
        RECT 37.380 46.995 37.570 47.715 ;
        RECT 37.740 46.825 37.910 47.895 ;
        RECT 38.370 47.865 38.570 47.895 ;
        RECT 38.080 47.645 38.250 47.715 ;
        RECT 38.780 47.645 38.950 48.425 ;
        RECT 39.815 48.285 39.985 48.425 ;
        RECT 40.155 48.415 40.405 48.875 ;
        RECT 38.080 47.475 38.950 47.645 ;
        RECT 39.120 48.005 39.645 48.225 ;
        RECT 39.815 48.155 40.040 48.285 ;
        RECT 38.080 47.385 38.590 47.475 ;
        RECT 36.550 46.625 37.435 46.795 ;
        RECT 37.660 46.495 37.910 46.825 ;
        RECT 38.080 46.325 38.250 47.125 ;
        RECT 38.420 46.770 38.590 47.385 ;
        RECT 39.120 47.305 39.290 48.005 ;
        RECT 38.760 46.940 39.290 47.305 ;
        RECT 39.460 47.240 39.700 47.835 ;
        RECT 39.870 47.050 40.040 48.155 ;
        RECT 40.210 47.295 40.490 48.245 ;
        RECT 39.735 46.920 40.040 47.050 ;
        RECT 38.420 46.600 39.525 46.770 ;
        RECT 39.735 46.495 39.985 46.920 ;
        RECT 40.155 46.325 40.420 46.785 ;
        RECT 40.660 46.495 40.845 48.615 ;
        RECT 41.015 48.495 41.345 48.875 ;
        RECT 41.515 48.325 41.685 48.615 ;
        RECT 41.020 48.155 41.685 48.325 ;
        RECT 42.060 48.245 42.345 48.705 ;
        RECT 42.515 48.415 42.785 48.875 ;
        RECT 41.020 47.165 41.250 48.155 ;
        RECT 42.060 48.075 43.015 48.245 ;
        RECT 41.420 47.335 41.770 47.985 ;
        RECT 41.945 47.345 42.635 47.905 ;
        RECT 42.805 47.175 43.015 48.075 ;
        RECT 41.020 46.995 41.685 47.165 ;
        RECT 41.015 46.325 41.345 46.825 ;
        RECT 41.515 46.495 41.685 46.995 ;
        RECT 42.060 46.955 43.015 47.175 ;
        RECT 43.185 47.905 43.585 48.705 ;
        RECT 43.775 48.245 44.055 48.705 ;
        RECT 44.575 48.415 44.900 48.875 ;
        RECT 43.775 48.075 44.900 48.245 ;
        RECT 45.070 48.135 45.455 48.705 ;
        RECT 44.450 47.965 44.900 48.075 ;
        RECT 43.185 47.345 44.280 47.905 ;
        RECT 44.450 47.635 45.005 47.965 ;
        RECT 42.060 46.495 42.345 46.955 ;
        RECT 42.515 46.325 42.785 46.785 ;
        RECT 43.185 46.495 43.585 47.345 ;
        RECT 44.450 47.175 44.900 47.635 ;
        RECT 45.175 47.465 45.455 48.135 ;
        RECT 43.775 46.955 44.900 47.175 ;
        RECT 43.775 46.495 44.055 46.955 ;
        RECT 44.575 46.325 44.900 46.785 ;
        RECT 45.070 46.495 45.455 47.465 ;
        RECT 45.625 47.930 45.965 48.705 ;
        RECT 46.135 48.415 46.305 48.875 ;
        RECT 46.545 48.440 46.905 48.705 ;
        RECT 46.545 48.435 46.900 48.440 ;
        RECT 46.545 48.425 46.895 48.435 ;
        RECT 46.545 48.420 46.890 48.425 ;
        RECT 46.545 48.410 46.885 48.420 ;
        RECT 47.535 48.415 47.705 48.875 ;
        RECT 46.545 48.405 46.880 48.410 ;
        RECT 46.545 48.395 46.870 48.405 ;
        RECT 46.545 48.385 46.860 48.395 ;
        RECT 46.545 48.245 46.845 48.385 ;
        RECT 46.135 48.055 46.845 48.245 ;
        RECT 47.035 48.245 47.365 48.325 ;
        RECT 47.875 48.245 48.215 48.705 ;
        RECT 47.035 48.055 48.215 48.245 ;
        RECT 48.935 48.325 49.105 48.615 ;
        RECT 49.275 48.495 49.605 48.875 ;
        RECT 48.935 48.155 49.600 48.325 ;
        RECT 45.625 46.495 45.905 47.930 ;
        RECT 46.135 47.485 46.420 48.055 ;
        RECT 46.605 47.655 47.075 47.885 ;
        RECT 47.245 47.865 47.575 47.885 ;
        RECT 47.245 47.685 47.695 47.865 ;
        RECT 47.885 47.685 48.215 47.885 ;
        RECT 46.135 47.270 47.285 47.485 ;
        RECT 46.075 46.325 46.785 47.100 ;
        RECT 46.955 46.495 47.285 47.270 ;
        RECT 47.480 46.570 47.695 47.685 ;
        RECT 47.985 47.345 48.215 47.685 ;
        RECT 48.850 47.335 49.200 47.985 ;
        RECT 49.370 47.165 49.600 48.155 ;
        RECT 47.875 46.325 48.205 47.045 ;
        RECT 48.935 46.995 49.600 47.165 ;
        RECT 48.935 46.495 49.105 46.995 ;
        RECT 49.275 46.325 49.605 46.825 ;
        RECT 49.775 46.495 49.960 48.615 ;
        RECT 50.215 48.415 50.465 48.875 ;
        RECT 50.635 48.425 50.970 48.595 ;
        RECT 51.165 48.425 51.840 48.595 ;
        RECT 50.635 48.285 50.805 48.425 ;
        RECT 50.130 47.295 50.410 48.245 ;
        RECT 50.580 48.155 50.805 48.285 ;
        RECT 50.580 47.050 50.750 48.155 ;
        RECT 50.975 48.005 51.500 48.225 ;
        RECT 50.920 47.240 51.160 47.835 ;
        RECT 51.330 47.305 51.500 48.005 ;
        RECT 51.670 47.645 51.840 48.425 ;
        RECT 52.160 48.375 52.530 48.875 ;
        RECT 52.710 48.425 53.115 48.595 ;
        RECT 53.285 48.425 54.070 48.595 ;
        RECT 52.710 48.195 52.880 48.425 ;
        RECT 52.050 47.895 52.880 48.195 ;
        RECT 53.265 47.925 53.730 48.255 ;
        RECT 52.050 47.865 52.250 47.895 ;
        RECT 52.370 47.645 52.540 47.715 ;
        RECT 51.670 47.475 52.540 47.645 ;
        RECT 52.030 47.385 52.540 47.475 ;
        RECT 50.580 46.920 50.885 47.050 ;
        RECT 51.330 46.940 51.860 47.305 ;
        RECT 50.200 46.325 50.465 46.785 ;
        RECT 50.635 46.495 50.885 46.920 ;
        RECT 52.030 46.770 52.200 47.385 ;
        RECT 51.095 46.600 52.200 46.770 ;
        RECT 52.370 46.325 52.540 47.125 ;
        RECT 52.710 46.825 52.880 47.895 ;
        RECT 53.050 46.995 53.240 47.715 ;
        RECT 53.410 46.965 53.730 47.925 ;
        RECT 53.900 47.965 54.070 48.425 ;
        RECT 54.345 48.345 54.555 48.875 ;
        RECT 54.815 48.135 55.145 48.660 ;
        RECT 55.315 48.265 55.485 48.875 ;
        RECT 55.655 48.220 55.985 48.655 ;
        RECT 56.155 48.360 56.325 48.875 ;
        RECT 55.655 48.135 56.035 48.220 ;
        RECT 57.125 48.150 57.415 48.875 ;
        RECT 57.675 48.325 57.845 48.615 ;
        RECT 58.015 48.495 58.345 48.875 ;
        RECT 57.675 48.155 58.340 48.325 ;
        RECT 54.945 47.965 55.145 48.135 ;
        RECT 55.810 48.095 56.035 48.135 ;
        RECT 53.900 47.635 54.775 47.965 ;
        RECT 54.945 47.635 55.695 47.965 ;
        RECT 52.710 46.495 52.960 46.825 ;
        RECT 53.900 46.795 54.070 47.635 ;
        RECT 54.945 47.430 55.135 47.635 ;
        RECT 55.865 47.515 56.035 48.095 ;
        RECT 55.820 47.465 56.035 47.515 ;
        RECT 54.240 47.055 55.135 47.430 ;
        RECT 55.645 47.385 56.035 47.465 ;
        RECT 53.185 46.625 54.070 46.795 ;
        RECT 54.250 46.325 54.565 46.825 ;
        RECT 54.795 46.495 55.135 47.055 ;
        RECT 55.305 46.325 55.475 47.335 ;
        RECT 55.645 46.540 55.975 47.385 ;
        RECT 56.145 46.325 56.315 47.240 ;
        RECT 57.125 46.325 57.415 47.490 ;
        RECT 57.590 47.335 57.940 47.985 ;
        RECT 58.110 47.165 58.340 48.155 ;
        RECT 57.675 46.995 58.340 47.165 ;
        RECT 57.675 46.495 57.845 46.995 ;
        RECT 58.015 46.325 58.345 46.825 ;
        RECT 58.515 46.495 58.700 48.615 ;
        RECT 58.955 48.415 59.205 48.875 ;
        RECT 59.375 48.425 59.710 48.595 ;
        RECT 59.905 48.425 60.580 48.595 ;
        RECT 59.375 48.285 59.545 48.425 ;
        RECT 58.870 47.295 59.150 48.245 ;
        RECT 59.320 48.155 59.545 48.285 ;
        RECT 59.320 47.050 59.490 48.155 ;
        RECT 59.715 48.005 60.240 48.225 ;
        RECT 59.660 47.240 59.900 47.835 ;
        RECT 60.070 47.305 60.240 48.005 ;
        RECT 60.410 47.645 60.580 48.425 ;
        RECT 60.900 48.375 61.270 48.875 ;
        RECT 61.450 48.425 61.855 48.595 ;
        RECT 62.025 48.425 62.810 48.595 ;
        RECT 61.450 48.195 61.620 48.425 ;
        RECT 60.790 47.895 61.620 48.195 ;
        RECT 62.005 47.925 62.470 48.255 ;
        RECT 60.790 47.865 60.990 47.895 ;
        RECT 61.110 47.645 61.280 47.715 ;
        RECT 60.410 47.475 61.280 47.645 ;
        RECT 60.770 47.385 61.280 47.475 ;
        RECT 59.320 46.920 59.625 47.050 ;
        RECT 60.070 46.940 60.600 47.305 ;
        RECT 58.940 46.325 59.205 46.785 ;
        RECT 59.375 46.495 59.625 46.920 ;
        RECT 60.770 46.770 60.940 47.385 ;
        RECT 59.835 46.600 60.940 46.770 ;
        RECT 61.110 46.325 61.280 47.125 ;
        RECT 61.450 46.825 61.620 47.895 ;
        RECT 61.790 46.995 61.980 47.715 ;
        RECT 62.150 46.965 62.470 47.925 ;
        RECT 62.640 47.965 62.810 48.425 ;
        RECT 63.085 48.345 63.295 48.875 ;
        RECT 63.555 48.135 63.885 48.660 ;
        RECT 64.055 48.265 64.225 48.875 ;
        RECT 64.395 48.220 64.725 48.655 ;
        RECT 64.895 48.360 65.065 48.875 ;
        RECT 65.495 48.325 65.665 48.615 ;
        RECT 65.835 48.495 66.165 48.875 ;
        RECT 64.395 48.135 64.775 48.220 ;
        RECT 65.495 48.155 66.160 48.325 ;
        RECT 63.685 47.965 63.885 48.135 ;
        RECT 64.550 48.095 64.775 48.135 ;
        RECT 62.640 47.635 63.515 47.965 ;
        RECT 63.685 47.635 64.435 47.965 ;
        RECT 61.450 46.495 61.700 46.825 ;
        RECT 62.640 46.795 62.810 47.635 ;
        RECT 63.685 47.430 63.875 47.635 ;
        RECT 64.605 47.515 64.775 48.095 ;
        RECT 64.560 47.465 64.775 47.515 ;
        RECT 62.980 47.055 63.875 47.430 ;
        RECT 64.385 47.385 64.775 47.465 ;
        RECT 61.925 46.625 62.810 46.795 ;
        RECT 62.990 46.325 63.305 46.825 ;
        RECT 63.535 46.495 63.875 47.055 ;
        RECT 64.045 46.325 64.215 47.335 ;
        RECT 64.385 46.540 64.715 47.385 ;
        RECT 65.410 47.335 65.760 47.985 ;
        RECT 64.885 46.325 65.055 47.240 ;
        RECT 65.930 47.165 66.160 48.155 ;
        RECT 65.495 46.995 66.160 47.165 ;
        RECT 65.495 46.495 65.665 46.995 ;
        RECT 65.835 46.325 66.165 46.825 ;
        RECT 66.335 46.495 66.520 48.615 ;
        RECT 66.775 48.415 67.025 48.875 ;
        RECT 67.195 48.425 67.530 48.595 ;
        RECT 67.725 48.425 68.400 48.595 ;
        RECT 67.195 48.285 67.365 48.425 ;
        RECT 66.690 47.295 66.970 48.245 ;
        RECT 67.140 48.155 67.365 48.285 ;
        RECT 67.140 47.050 67.310 48.155 ;
        RECT 67.535 48.005 68.060 48.225 ;
        RECT 67.480 47.240 67.720 47.835 ;
        RECT 67.890 47.305 68.060 48.005 ;
        RECT 68.230 47.645 68.400 48.425 ;
        RECT 68.720 48.375 69.090 48.875 ;
        RECT 69.270 48.425 69.675 48.595 ;
        RECT 69.845 48.425 70.630 48.595 ;
        RECT 69.270 48.195 69.440 48.425 ;
        RECT 68.610 47.895 69.440 48.195 ;
        RECT 69.825 47.925 70.290 48.255 ;
        RECT 68.610 47.865 68.810 47.895 ;
        RECT 68.930 47.645 69.100 47.715 ;
        RECT 68.230 47.475 69.100 47.645 ;
        RECT 68.590 47.385 69.100 47.475 ;
        RECT 67.140 46.920 67.445 47.050 ;
        RECT 67.890 46.940 68.420 47.305 ;
        RECT 66.760 46.325 67.025 46.785 ;
        RECT 67.195 46.495 67.445 46.920 ;
        RECT 68.590 46.770 68.760 47.385 ;
        RECT 67.655 46.600 68.760 46.770 ;
        RECT 68.930 46.325 69.100 47.125 ;
        RECT 69.270 46.825 69.440 47.895 ;
        RECT 69.610 46.995 69.800 47.715 ;
        RECT 69.970 46.965 70.290 47.925 ;
        RECT 70.460 47.965 70.630 48.425 ;
        RECT 70.905 48.345 71.115 48.875 ;
        RECT 71.375 48.135 71.705 48.660 ;
        RECT 71.875 48.265 72.045 48.875 ;
        RECT 72.215 48.220 72.545 48.655 ;
        RECT 72.765 48.375 73.025 48.705 ;
        RECT 73.195 48.515 73.525 48.875 ;
        RECT 73.780 48.495 75.080 48.705 ;
        RECT 72.215 48.135 72.595 48.220 ;
        RECT 71.505 47.965 71.705 48.135 ;
        RECT 72.370 48.095 72.595 48.135 ;
        RECT 70.460 47.635 71.335 47.965 ;
        RECT 71.505 47.635 72.255 47.965 ;
        RECT 69.270 46.495 69.520 46.825 ;
        RECT 70.460 46.795 70.630 47.635 ;
        RECT 71.505 47.430 71.695 47.635 ;
        RECT 72.425 47.515 72.595 48.095 ;
        RECT 72.380 47.465 72.595 47.515 ;
        RECT 70.800 47.055 71.695 47.430 ;
        RECT 72.205 47.385 72.595 47.465 ;
        RECT 69.745 46.625 70.630 46.795 ;
        RECT 70.810 46.325 71.125 46.825 ;
        RECT 71.355 46.495 71.695 47.055 ;
        RECT 71.865 46.325 72.035 47.335 ;
        RECT 72.205 46.540 72.535 47.385 ;
        RECT 72.765 47.175 72.935 48.375 ;
        RECT 73.780 48.345 73.950 48.495 ;
        RECT 73.195 48.220 73.950 48.345 ;
        RECT 73.105 48.175 73.950 48.220 ;
        RECT 73.105 48.055 73.375 48.175 ;
        RECT 73.105 47.480 73.275 48.055 ;
        RECT 73.505 47.615 73.915 47.920 ;
        RECT 74.205 47.885 74.415 48.285 ;
        RECT 74.085 47.675 74.415 47.885 ;
        RECT 74.660 47.885 74.880 48.285 ;
        RECT 75.355 48.110 75.810 48.875 ;
        RECT 77.070 48.365 77.310 48.875 ;
        RECT 77.490 48.365 77.770 48.695 ;
        RECT 78.000 48.365 78.215 48.875 ;
        RECT 74.660 47.675 75.135 47.885 ;
        RECT 75.325 47.685 75.815 47.885 ;
        RECT 76.965 47.635 77.320 48.195 ;
        RECT 73.105 47.445 73.305 47.480 ;
        RECT 74.635 47.445 75.810 47.505 ;
        RECT 77.490 47.465 77.660 48.365 ;
        RECT 77.830 47.635 78.095 48.195 ;
        RECT 78.385 48.135 79.000 48.705 ;
        RECT 79.370 48.365 79.610 48.875 ;
        RECT 79.790 48.365 80.070 48.695 ;
        RECT 80.300 48.365 80.515 48.875 ;
        RECT 78.345 47.465 78.515 47.965 ;
        RECT 73.105 47.335 75.810 47.445 ;
        RECT 73.165 47.275 74.965 47.335 ;
        RECT 74.635 47.245 74.965 47.275 ;
        RECT 72.765 46.495 73.025 47.175 ;
        RECT 73.195 46.325 73.445 47.105 ;
        RECT 73.695 47.075 74.530 47.085 ;
        RECT 75.120 47.075 75.305 47.165 ;
        RECT 73.695 46.875 75.305 47.075 ;
        RECT 73.695 46.495 73.945 46.875 ;
        RECT 75.075 46.835 75.305 46.875 ;
        RECT 75.555 46.715 75.810 47.335 ;
        RECT 77.090 47.295 78.515 47.465 ;
        RECT 77.090 47.120 77.480 47.295 ;
        RECT 74.115 46.325 74.470 46.705 ;
        RECT 75.475 46.495 75.810 46.715 ;
        RECT 77.965 46.325 78.295 47.125 ;
        RECT 78.685 47.115 79.000 48.135 ;
        RECT 79.265 47.635 79.620 48.195 ;
        RECT 79.790 47.465 79.960 48.365 ;
        RECT 80.130 47.635 80.395 48.195 ;
        RECT 80.685 48.135 81.300 48.705 ;
        RECT 80.645 47.465 80.815 47.965 ;
        RECT 79.390 47.295 80.815 47.465 ;
        RECT 79.390 47.120 79.780 47.295 ;
        RECT 78.465 46.495 79.000 47.115 ;
        RECT 80.265 46.325 80.595 47.125 ;
        RECT 80.985 47.115 81.300 48.135 ;
        RECT 81.965 48.125 83.175 48.875 ;
        RECT 80.765 46.495 81.300 47.115 ;
        RECT 81.965 47.415 82.485 47.955 ;
        RECT 82.655 47.585 83.175 48.125 ;
        RECT 81.965 46.325 83.175 47.415 ;
        RECT 5.520 46.155 83.260 46.325 ;
        RECT 5.605 45.065 6.815 46.155 ;
        RECT 6.985 45.065 8.655 46.155 ;
        RECT 5.605 44.355 6.125 44.895 ;
        RECT 6.295 44.525 6.815 45.065 ;
        RECT 6.985 44.375 7.735 44.895 ;
        RECT 7.905 44.545 8.655 45.065 ;
        RECT 8.825 45.285 9.100 45.985 ;
        RECT 9.270 45.610 9.525 46.155 ;
        RECT 9.695 45.645 10.175 45.985 ;
        RECT 10.350 45.600 10.955 46.155 ;
        RECT 10.340 45.500 10.955 45.600 ;
        RECT 11.135 45.545 11.465 45.975 ;
        RECT 11.645 45.715 11.840 46.155 ;
        RECT 12.010 45.545 12.340 45.975 ;
        RECT 10.340 45.475 10.525 45.500 ;
        RECT 5.605 43.605 6.815 44.355 ;
        RECT 6.985 43.605 8.655 44.375 ;
        RECT 8.825 44.255 8.995 45.285 ;
        RECT 9.270 45.155 10.025 45.405 ;
        RECT 10.195 45.230 10.525 45.475 ;
        RECT 11.135 45.375 12.340 45.545 ;
        RECT 9.270 45.120 10.040 45.155 ;
        RECT 9.270 45.110 10.055 45.120 ;
        RECT 9.165 45.095 10.060 45.110 ;
        RECT 9.165 45.080 10.080 45.095 ;
        RECT 9.165 45.070 10.100 45.080 ;
        RECT 9.165 45.060 10.125 45.070 ;
        RECT 9.165 45.030 10.195 45.060 ;
        RECT 9.165 45.000 10.215 45.030 ;
        RECT 9.165 44.970 10.235 45.000 ;
        RECT 9.165 44.945 10.265 44.970 ;
        RECT 9.165 44.910 10.300 44.945 ;
        RECT 9.165 44.905 10.330 44.910 ;
        RECT 9.165 44.510 9.395 44.905 ;
        RECT 9.940 44.900 10.330 44.905 ;
        RECT 9.965 44.890 10.330 44.900 ;
        RECT 9.980 44.885 10.330 44.890 ;
        RECT 9.995 44.880 10.330 44.885 ;
        RECT 10.695 44.880 10.955 45.330 ;
        RECT 11.135 45.045 12.030 45.375 ;
        RECT 12.510 45.205 12.785 45.975 ;
        RECT 9.995 44.875 10.955 44.880 ;
        RECT 10.005 44.865 10.955 44.875 ;
        RECT 10.015 44.860 10.955 44.865 ;
        RECT 10.025 44.850 10.955 44.860 ;
        RECT 10.030 44.840 10.955 44.850 ;
        RECT 12.200 45.015 12.785 45.205 ;
        RECT 12.965 45.065 15.555 46.155 ;
        RECT 10.035 44.835 10.955 44.840 ;
        RECT 10.045 44.820 10.955 44.835 ;
        RECT 10.050 44.805 10.955 44.820 ;
        RECT 10.060 44.780 10.955 44.805 ;
        RECT 9.565 44.310 9.895 44.735 ;
        RECT 9.645 44.285 9.895 44.310 ;
        RECT 8.825 43.775 9.085 44.255 ;
        RECT 9.255 43.605 9.505 44.145 ;
        RECT 9.675 43.825 9.895 44.285 ;
        RECT 10.065 44.710 10.955 44.780 ;
        RECT 10.065 43.985 10.235 44.710 ;
        RECT 10.405 44.155 10.955 44.540 ;
        RECT 11.140 44.515 11.435 44.845 ;
        RECT 11.615 44.515 12.030 44.845 ;
        RECT 10.065 43.815 10.955 43.985 ;
        RECT 11.135 43.605 11.435 44.335 ;
        RECT 11.615 43.895 11.845 44.515 ;
        RECT 12.200 44.345 12.375 45.015 ;
        RECT 12.045 44.165 12.375 44.345 ;
        RECT 12.545 44.195 12.785 44.845 ;
        RECT 12.965 44.375 14.175 44.895 ;
        RECT 14.345 44.545 15.555 45.065 ;
        RECT 16.370 45.185 16.760 45.360 ;
        RECT 17.245 45.355 17.575 46.155 ;
        RECT 17.745 45.365 18.280 45.985 ;
        RECT 16.370 45.015 17.795 45.185 ;
        RECT 12.045 43.785 12.270 44.165 ;
        RECT 12.440 43.605 12.770 43.995 ;
        RECT 12.965 43.605 15.555 44.375 ;
        RECT 16.245 44.285 16.600 44.845 ;
        RECT 16.770 44.115 16.940 45.015 ;
        RECT 17.110 44.285 17.375 44.845 ;
        RECT 17.625 44.515 17.795 45.015 ;
        RECT 17.965 44.345 18.280 45.365 ;
        RECT 18.485 44.990 18.775 46.155 ;
        RECT 18.950 45.645 20.605 45.935 ;
        RECT 18.950 45.305 20.540 45.475 ;
        RECT 20.775 45.355 21.055 46.155 ;
        RECT 18.950 45.015 19.270 45.305 ;
        RECT 20.370 45.185 20.540 45.305 ;
        RECT 16.350 43.605 16.590 44.115 ;
        RECT 16.770 43.785 17.050 44.115 ;
        RECT 17.280 43.605 17.495 44.115 ;
        RECT 17.665 43.775 18.280 44.345 ;
        RECT 18.485 43.605 18.775 44.330 ;
        RECT 18.950 44.275 19.300 44.845 ;
        RECT 19.470 44.515 20.180 45.135 ;
        RECT 20.370 45.015 21.095 45.185 ;
        RECT 21.265 45.015 21.535 45.985 ;
        RECT 20.925 44.845 21.095 45.015 ;
        RECT 20.350 44.515 20.755 44.845 ;
        RECT 20.925 44.515 21.195 44.845 ;
        RECT 20.925 44.345 21.095 44.515 ;
        RECT 19.485 44.175 21.095 44.345 ;
        RECT 21.365 44.280 21.535 45.015 ;
        RECT 18.955 43.605 19.285 44.105 ;
        RECT 19.485 43.825 19.655 44.175 ;
        RECT 19.855 43.605 20.185 44.005 ;
        RECT 20.355 43.825 20.525 44.175 ;
        RECT 20.695 43.605 21.075 44.005 ;
        RECT 21.265 43.935 21.535 44.280 ;
        RECT 22.625 43.885 22.905 45.985 ;
        RECT 23.095 45.395 23.880 46.155 ;
        RECT 24.275 45.325 24.660 45.985 ;
        RECT 24.275 45.225 24.685 45.325 ;
        RECT 23.075 45.015 24.685 45.225 ;
        RECT 24.985 45.135 25.185 45.925 ;
        RECT 23.075 44.415 23.350 45.015 ;
        RECT 24.855 44.965 25.185 45.135 ;
        RECT 25.355 44.975 25.675 46.155 ;
        RECT 26.305 45.320 26.650 46.155 ;
        RECT 26.825 45.150 27.080 45.955 ;
        RECT 27.250 45.320 27.510 46.155 ;
        RECT 27.685 45.150 27.940 45.955 ;
        RECT 28.110 45.320 28.370 46.155 ;
        RECT 28.540 45.150 28.800 45.955 ;
        RECT 28.970 45.320 29.355 46.155 ;
        RECT 29.775 45.425 30.070 46.155 ;
        RECT 30.240 45.255 30.500 45.980 ;
        RECT 30.670 45.425 30.930 46.155 ;
        RECT 31.100 45.255 31.360 45.980 ;
        RECT 31.530 45.425 31.790 46.155 ;
        RECT 31.960 45.255 32.220 45.980 ;
        RECT 32.390 45.425 32.650 46.155 ;
        RECT 32.820 45.255 33.080 45.980 ;
        RECT 26.325 44.980 29.355 45.150 ;
        RECT 24.855 44.845 25.035 44.965 ;
        RECT 23.520 44.595 23.875 44.845 ;
        RECT 24.070 44.795 24.535 44.845 ;
        RECT 24.065 44.625 24.535 44.795 ;
        RECT 24.070 44.595 24.535 44.625 ;
        RECT 24.705 44.595 25.035 44.845 ;
        RECT 25.210 44.595 25.675 44.795 ;
        RECT 26.325 44.415 26.495 44.980 ;
        RECT 26.665 44.585 28.880 44.810 ;
        RECT 29.055 44.415 29.355 44.980 ;
        RECT 23.075 44.235 24.325 44.415 ;
        RECT 23.960 44.165 24.325 44.235 ;
        RECT 24.495 44.215 25.675 44.385 ;
        RECT 26.325 44.245 29.355 44.415 ;
        RECT 29.770 45.015 33.080 45.255 ;
        RECT 33.250 45.045 33.510 46.155 ;
        RECT 29.770 44.425 30.740 45.015 ;
        RECT 33.680 44.845 33.930 45.980 ;
        RECT 34.110 45.045 34.405 46.155 ;
        RECT 34.675 45.485 34.845 45.985 ;
        RECT 35.015 45.655 35.345 46.155 ;
        RECT 34.675 45.315 35.340 45.485 ;
        RECT 30.910 44.595 33.930 44.845 ;
        RECT 29.770 44.255 33.080 44.425 ;
        RECT 23.135 43.605 23.305 44.065 ;
        RECT 24.495 43.995 24.825 44.215 ;
        RECT 23.575 43.815 24.825 43.995 ;
        RECT 24.995 43.605 25.165 44.045 ;
        RECT 25.335 43.800 25.675 44.215 ;
        RECT 26.785 43.605 27.080 44.075 ;
        RECT 27.250 43.800 27.510 44.245 ;
        RECT 27.680 43.605 27.940 44.075 ;
        RECT 28.110 43.800 28.365 44.245 ;
        RECT 28.535 43.605 28.835 44.075 ;
        RECT 29.770 43.605 30.070 44.085 ;
        RECT 30.240 43.800 30.500 44.255 ;
        RECT 30.670 43.605 30.930 44.085 ;
        RECT 31.100 43.800 31.360 44.255 ;
        RECT 31.530 43.605 31.790 44.085 ;
        RECT 31.960 43.800 32.220 44.255 ;
        RECT 32.390 43.605 32.650 44.085 ;
        RECT 32.820 43.800 33.080 44.255 ;
        RECT 33.250 43.605 33.510 44.130 ;
        RECT 33.680 43.785 33.930 44.595 ;
        RECT 34.100 44.235 34.415 44.845 ;
        RECT 34.590 44.495 34.940 45.145 ;
        RECT 35.110 44.325 35.340 45.315 ;
        RECT 34.675 44.155 35.340 44.325 ;
        RECT 34.110 43.605 34.355 44.065 ;
        RECT 34.675 43.865 34.845 44.155 ;
        RECT 35.015 43.605 35.345 43.985 ;
        RECT 35.515 43.865 35.700 45.985 ;
        RECT 35.940 45.695 36.205 46.155 ;
        RECT 36.375 45.560 36.625 45.985 ;
        RECT 36.835 45.710 37.940 45.880 ;
        RECT 36.320 45.430 36.625 45.560 ;
        RECT 35.870 44.235 36.150 45.185 ;
        RECT 36.320 44.325 36.490 45.430 ;
        RECT 36.660 44.645 36.900 45.240 ;
        RECT 37.070 45.175 37.600 45.540 ;
        RECT 37.070 44.475 37.240 45.175 ;
        RECT 37.770 45.095 37.940 45.710 ;
        RECT 38.110 45.355 38.280 46.155 ;
        RECT 38.450 45.655 38.700 45.985 ;
        RECT 38.925 45.685 39.810 45.855 ;
        RECT 37.770 45.005 38.280 45.095 ;
        RECT 36.320 44.195 36.545 44.325 ;
        RECT 36.715 44.255 37.240 44.475 ;
        RECT 37.410 44.835 38.280 45.005 ;
        RECT 35.955 43.605 36.205 44.065 ;
        RECT 36.375 44.055 36.545 44.195 ;
        RECT 37.410 44.055 37.580 44.835 ;
        RECT 38.110 44.765 38.280 44.835 ;
        RECT 37.790 44.585 37.990 44.615 ;
        RECT 38.450 44.585 38.620 45.655 ;
        RECT 38.790 44.765 38.980 45.485 ;
        RECT 37.790 44.285 38.620 44.585 ;
        RECT 39.150 44.555 39.470 45.515 ;
        RECT 36.375 43.885 36.710 44.055 ;
        RECT 36.905 43.885 37.580 44.055 ;
        RECT 37.900 43.605 38.270 44.105 ;
        RECT 38.450 44.055 38.620 44.285 ;
        RECT 39.005 44.225 39.470 44.555 ;
        RECT 39.640 44.845 39.810 45.685 ;
        RECT 39.990 45.655 40.305 46.155 ;
        RECT 40.535 45.425 40.875 45.985 ;
        RECT 39.980 45.050 40.875 45.425 ;
        RECT 41.045 45.145 41.215 46.155 ;
        RECT 40.685 44.845 40.875 45.050 ;
        RECT 41.385 45.095 41.715 45.940 ;
        RECT 41.945 45.600 42.550 46.155 ;
        RECT 42.725 45.645 43.205 45.985 ;
        RECT 43.375 45.610 43.630 46.155 ;
        RECT 41.945 45.500 42.560 45.600 ;
        RECT 42.375 45.475 42.560 45.500 ;
        RECT 41.385 45.015 41.775 45.095 ;
        RECT 41.560 44.965 41.775 45.015 ;
        RECT 39.640 44.515 40.515 44.845 ;
        RECT 40.685 44.515 41.435 44.845 ;
        RECT 39.640 44.055 39.810 44.515 ;
        RECT 40.685 44.345 40.885 44.515 ;
        RECT 41.605 44.385 41.775 44.965 ;
        RECT 41.945 44.880 42.205 45.330 ;
        RECT 42.375 45.230 42.705 45.475 ;
        RECT 42.875 45.155 43.630 45.405 ;
        RECT 43.800 45.285 44.075 45.985 ;
        RECT 42.860 45.120 43.630 45.155 ;
        RECT 42.845 45.110 43.630 45.120 ;
        RECT 42.840 45.095 43.735 45.110 ;
        RECT 42.820 45.080 43.735 45.095 ;
        RECT 42.800 45.070 43.735 45.080 ;
        RECT 42.775 45.060 43.735 45.070 ;
        RECT 42.705 45.030 43.735 45.060 ;
        RECT 42.685 45.000 43.735 45.030 ;
        RECT 42.665 44.970 43.735 45.000 ;
        RECT 42.635 44.945 43.735 44.970 ;
        RECT 42.600 44.910 43.735 44.945 ;
        RECT 42.570 44.905 43.735 44.910 ;
        RECT 42.570 44.900 42.960 44.905 ;
        RECT 42.570 44.890 42.935 44.900 ;
        RECT 42.570 44.885 42.920 44.890 ;
        RECT 42.570 44.880 42.905 44.885 ;
        RECT 41.945 44.875 42.905 44.880 ;
        RECT 41.945 44.865 42.895 44.875 ;
        RECT 41.945 44.860 42.885 44.865 ;
        RECT 41.945 44.850 42.875 44.860 ;
        RECT 41.945 44.840 42.870 44.850 ;
        RECT 41.945 44.835 42.865 44.840 ;
        RECT 41.945 44.820 42.855 44.835 ;
        RECT 41.945 44.805 42.850 44.820 ;
        RECT 41.945 44.780 42.840 44.805 ;
        RECT 41.945 44.710 42.835 44.780 ;
        RECT 41.550 44.345 41.775 44.385 ;
        RECT 38.450 43.885 38.855 44.055 ;
        RECT 39.025 43.885 39.810 44.055 ;
        RECT 40.085 43.605 40.295 44.135 ;
        RECT 40.555 43.820 40.885 44.345 ;
        RECT 41.395 44.260 41.775 44.345 ;
        RECT 41.055 43.605 41.225 44.215 ;
        RECT 41.395 43.825 41.725 44.260 ;
        RECT 41.945 44.155 42.495 44.540 ;
        RECT 42.665 43.985 42.835 44.710 ;
        RECT 41.945 43.815 42.835 43.985 ;
        RECT 43.005 44.310 43.335 44.735 ;
        RECT 43.505 44.510 43.735 44.905 ;
        RECT 43.005 43.825 43.225 44.310 ;
        RECT 43.905 44.255 44.075 45.285 ;
        RECT 44.245 44.990 44.535 46.155 ;
        RECT 44.795 45.485 44.965 45.985 ;
        RECT 45.135 45.655 45.465 46.155 ;
        RECT 44.795 45.315 45.460 45.485 ;
        RECT 44.710 44.495 45.060 45.145 ;
        RECT 43.395 43.605 43.645 44.145 ;
        RECT 43.815 43.775 44.075 44.255 ;
        RECT 44.245 43.605 44.535 44.330 ;
        RECT 45.230 44.325 45.460 45.315 ;
        RECT 44.795 44.155 45.460 44.325 ;
        RECT 44.795 43.865 44.965 44.155 ;
        RECT 45.135 43.605 45.465 43.985 ;
        RECT 45.635 43.865 45.820 45.985 ;
        RECT 46.060 45.695 46.325 46.155 ;
        RECT 46.495 45.560 46.745 45.985 ;
        RECT 46.955 45.710 48.060 45.880 ;
        RECT 46.440 45.430 46.745 45.560 ;
        RECT 45.990 44.235 46.270 45.185 ;
        RECT 46.440 44.325 46.610 45.430 ;
        RECT 46.780 44.645 47.020 45.240 ;
        RECT 47.190 45.175 47.720 45.540 ;
        RECT 47.190 44.475 47.360 45.175 ;
        RECT 47.890 45.095 48.060 45.710 ;
        RECT 48.230 45.355 48.400 46.155 ;
        RECT 48.570 45.655 48.820 45.985 ;
        RECT 49.045 45.685 49.930 45.855 ;
        RECT 47.890 45.005 48.400 45.095 ;
        RECT 46.440 44.195 46.665 44.325 ;
        RECT 46.835 44.255 47.360 44.475 ;
        RECT 47.530 44.835 48.400 45.005 ;
        RECT 46.075 43.605 46.325 44.065 ;
        RECT 46.495 44.055 46.665 44.195 ;
        RECT 47.530 44.055 47.700 44.835 ;
        RECT 48.230 44.765 48.400 44.835 ;
        RECT 47.910 44.585 48.110 44.615 ;
        RECT 48.570 44.585 48.740 45.655 ;
        RECT 48.910 44.765 49.100 45.485 ;
        RECT 47.910 44.285 48.740 44.585 ;
        RECT 49.270 44.555 49.590 45.515 ;
        RECT 46.495 43.885 46.830 44.055 ;
        RECT 47.025 43.885 47.700 44.055 ;
        RECT 48.020 43.605 48.390 44.105 ;
        RECT 48.570 44.055 48.740 44.285 ;
        RECT 49.125 44.225 49.590 44.555 ;
        RECT 49.760 44.845 49.930 45.685 ;
        RECT 50.110 45.655 50.425 46.155 ;
        RECT 50.655 45.425 50.995 45.985 ;
        RECT 50.100 45.050 50.995 45.425 ;
        RECT 51.165 45.145 51.335 46.155 ;
        RECT 50.805 44.845 50.995 45.050 ;
        RECT 51.505 45.095 51.835 45.940 ;
        RECT 52.315 45.425 52.610 46.155 ;
        RECT 52.780 45.255 53.040 45.980 ;
        RECT 53.210 45.425 53.470 46.155 ;
        RECT 53.640 45.255 53.900 45.980 ;
        RECT 54.070 45.425 54.330 46.155 ;
        RECT 54.500 45.255 54.760 45.980 ;
        RECT 54.930 45.425 55.190 46.155 ;
        RECT 55.360 45.255 55.620 45.980 ;
        RECT 51.505 45.015 51.895 45.095 ;
        RECT 51.680 44.965 51.895 45.015 ;
        RECT 49.760 44.515 50.635 44.845 ;
        RECT 50.805 44.515 51.555 44.845 ;
        RECT 49.760 44.055 49.930 44.515 ;
        RECT 50.805 44.345 51.005 44.515 ;
        RECT 51.725 44.385 51.895 44.965 ;
        RECT 51.670 44.345 51.895 44.385 ;
        RECT 48.570 43.885 48.975 44.055 ;
        RECT 49.145 43.885 49.930 44.055 ;
        RECT 50.205 43.605 50.415 44.135 ;
        RECT 50.675 43.820 51.005 44.345 ;
        RECT 51.515 44.260 51.895 44.345 ;
        RECT 52.310 45.015 55.620 45.255 ;
        RECT 55.790 45.045 56.050 46.155 ;
        RECT 52.310 44.425 53.280 45.015 ;
        RECT 56.220 44.845 56.470 45.980 ;
        RECT 56.650 45.045 56.945 46.155 ;
        RECT 57.130 45.015 57.465 45.985 ;
        RECT 57.635 45.015 57.805 46.155 ;
        RECT 57.975 45.815 60.005 45.985 ;
        RECT 53.450 44.595 56.470 44.845 ;
        RECT 51.175 43.605 51.345 44.215 ;
        RECT 51.515 43.825 51.845 44.260 ;
        RECT 52.310 44.255 55.620 44.425 ;
        RECT 52.310 43.605 52.610 44.085 ;
        RECT 52.780 43.800 53.040 44.255 ;
        RECT 53.210 43.605 53.470 44.085 ;
        RECT 53.640 43.800 53.900 44.255 ;
        RECT 54.070 43.605 54.330 44.085 ;
        RECT 54.500 43.800 54.760 44.255 ;
        RECT 54.930 43.605 55.190 44.085 ;
        RECT 55.360 43.800 55.620 44.255 ;
        RECT 55.790 43.605 56.050 44.130 ;
        RECT 56.220 43.785 56.470 44.595 ;
        RECT 56.640 44.235 56.955 44.845 ;
        RECT 57.130 44.345 57.300 45.015 ;
        RECT 57.975 44.845 58.145 45.815 ;
        RECT 57.470 44.515 57.725 44.845 ;
        RECT 57.950 44.515 58.145 44.845 ;
        RECT 58.315 45.475 59.440 45.645 ;
        RECT 57.555 44.345 57.725 44.515 ;
        RECT 58.315 44.345 58.485 45.475 ;
        RECT 56.650 43.605 56.895 44.065 ;
        RECT 57.130 43.775 57.385 44.345 ;
        RECT 57.555 44.175 58.485 44.345 ;
        RECT 58.655 45.135 59.665 45.305 ;
        RECT 58.655 44.335 58.825 45.135 ;
        RECT 59.030 44.455 59.305 44.935 ;
        RECT 59.025 44.285 59.305 44.455 ;
        RECT 58.310 44.140 58.485 44.175 ;
        RECT 57.555 43.605 57.885 44.005 ;
        RECT 58.310 43.775 58.840 44.140 ;
        RECT 59.030 43.775 59.305 44.285 ;
        RECT 59.475 43.775 59.665 45.135 ;
        RECT 59.835 45.150 60.005 45.815 ;
        RECT 60.175 45.395 60.345 46.155 ;
        RECT 60.580 45.395 61.095 45.805 ;
        RECT 62.435 45.425 62.730 46.155 ;
        RECT 59.835 44.960 60.585 45.150 ;
        RECT 60.755 44.585 61.095 45.395 ;
        RECT 62.900 45.255 63.160 45.980 ;
        RECT 63.330 45.425 63.590 46.155 ;
        RECT 63.760 45.255 64.020 45.980 ;
        RECT 64.190 45.425 64.450 46.155 ;
        RECT 64.620 45.255 64.880 45.980 ;
        RECT 65.050 45.425 65.310 46.155 ;
        RECT 65.480 45.255 65.740 45.980 ;
        RECT 59.865 44.415 61.095 44.585 ;
        RECT 62.430 45.015 65.740 45.255 ;
        RECT 65.910 45.045 66.170 46.155 ;
        RECT 62.430 44.425 63.400 45.015 ;
        RECT 66.340 44.845 66.590 45.980 ;
        RECT 66.770 45.045 67.065 46.155 ;
        RECT 67.245 45.645 68.435 45.935 ;
        RECT 67.265 45.305 68.435 45.475 ;
        RECT 68.605 45.355 68.885 46.155 ;
        RECT 67.265 45.015 67.590 45.305 ;
        RECT 68.265 45.185 68.435 45.305 ;
        RECT 67.760 44.845 67.955 45.135 ;
        RECT 68.265 45.015 68.925 45.185 ;
        RECT 69.095 45.015 69.370 45.985 ;
        RECT 68.755 44.845 68.925 45.015 ;
        RECT 63.570 44.595 66.590 44.845 ;
        RECT 59.845 43.605 60.355 44.140 ;
        RECT 60.575 43.810 60.820 44.415 ;
        RECT 62.430 44.255 65.740 44.425 ;
        RECT 62.430 43.605 62.730 44.085 ;
        RECT 62.900 43.800 63.160 44.255 ;
        RECT 63.330 43.605 63.590 44.085 ;
        RECT 63.760 43.800 64.020 44.255 ;
        RECT 64.190 43.605 64.450 44.085 ;
        RECT 64.620 43.800 64.880 44.255 ;
        RECT 65.050 43.605 65.310 44.085 ;
        RECT 65.480 43.800 65.740 44.255 ;
        RECT 65.910 43.605 66.170 44.130 ;
        RECT 66.340 43.785 66.590 44.595 ;
        RECT 66.760 44.235 67.075 44.845 ;
        RECT 67.245 44.515 67.590 44.845 ;
        RECT 67.760 44.515 68.585 44.845 ;
        RECT 68.755 44.515 69.030 44.845 ;
        RECT 68.755 44.345 68.925 44.515 ;
        RECT 67.260 44.175 68.925 44.345 ;
        RECT 69.200 44.280 69.370 45.015 ;
        RECT 70.005 44.990 70.295 46.155 ;
        RECT 70.500 45.365 71.035 45.985 ;
        RECT 70.500 44.345 70.815 45.365 ;
        RECT 71.205 45.355 71.535 46.155 ;
        RECT 72.020 45.185 72.410 45.360 ;
        RECT 70.985 45.015 72.410 45.185 ;
        RECT 72.765 45.065 73.975 46.155 ;
        RECT 70.985 44.515 71.155 45.015 ;
        RECT 66.770 43.605 67.015 44.065 ;
        RECT 67.260 43.825 67.515 44.175 ;
        RECT 67.685 43.605 68.015 44.005 ;
        RECT 68.185 43.825 68.355 44.175 ;
        RECT 68.525 43.605 68.905 44.005 ;
        RECT 69.095 43.935 69.370 44.280 ;
        RECT 70.005 43.605 70.295 44.330 ;
        RECT 70.500 43.775 71.115 44.345 ;
        RECT 71.405 44.285 71.670 44.845 ;
        RECT 71.840 44.115 72.010 45.015 ;
        RECT 72.180 44.285 72.535 44.845 ;
        RECT 72.765 44.355 73.285 44.895 ;
        RECT 73.455 44.525 73.975 45.065 ;
        RECT 74.145 45.015 74.485 45.985 ;
        RECT 74.655 45.015 74.825 46.155 ;
        RECT 75.095 45.355 75.345 46.155 ;
        RECT 75.990 45.185 76.320 45.985 ;
        RECT 76.620 45.355 76.950 46.155 ;
        RECT 77.120 45.185 77.450 45.985 ;
        RECT 75.015 45.015 77.450 45.185 ;
        RECT 77.860 45.365 78.395 45.985 ;
        RECT 74.145 44.405 74.320 45.015 ;
        RECT 75.015 44.765 75.185 45.015 ;
        RECT 74.490 44.595 75.185 44.765 ;
        RECT 75.360 44.595 75.780 44.795 ;
        RECT 75.950 44.595 76.280 44.795 ;
        RECT 76.450 44.595 76.780 44.795 ;
        RECT 71.285 43.605 71.500 44.115 ;
        RECT 71.730 43.785 72.010 44.115 ;
        RECT 72.190 43.605 72.430 44.115 ;
        RECT 72.765 43.605 73.975 44.355 ;
        RECT 74.145 43.775 74.485 44.405 ;
        RECT 74.655 43.605 74.905 44.405 ;
        RECT 75.095 44.255 76.320 44.425 ;
        RECT 75.095 43.775 75.425 44.255 ;
        RECT 75.595 43.605 75.820 44.065 ;
        RECT 75.990 43.775 76.320 44.255 ;
        RECT 76.950 44.385 77.120 45.015 ;
        RECT 77.305 44.595 77.655 44.845 ;
        RECT 76.950 43.775 77.450 44.385 ;
        RECT 77.860 44.345 78.175 45.365 ;
        RECT 78.565 45.355 78.895 46.155 ;
        RECT 79.380 45.185 79.770 45.360 ;
        RECT 78.345 45.015 79.770 45.185 ;
        RECT 80.215 45.225 80.385 45.985 ;
        RECT 80.600 45.395 80.930 46.155 ;
        RECT 80.215 45.055 80.930 45.225 ;
        RECT 81.100 45.080 81.355 45.985 ;
        RECT 78.345 44.515 78.515 45.015 ;
        RECT 77.860 43.775 78.475 44.345 ;
        RECT 78.765 44.285 79.030 44.845 ;
        RECT 79.200 44.115 79.370 45.015 ;
        RECT 79.540 44.285 79.895 44.845 ;
        RECT 80.125 44.505 80.480 44.875 ;
        RECT 80.760 44.845 80.930 45.055 ;
        RECT 80.760 44.515 81.015 44.845 ;
        RECT 80.760 44.325 80.930 44.515 ;
        RECT 81.185 44.350 81.355 45.080 ;
        RECT 81.530 45.005 81.790 46.155 ;
        RECT 81.965 45.065 83.175 46.155 ;
        RECT 81.965 44.525 82.485 45.065 ;
        RECT 80.215 44.155 80.930 44.325 ;
        RECT 78.645 43.605 78.860 44.115 ;
        RECT 79.090 43.785 79.370 44.115 ;
        RECT 79.550 43.605 79.790 44.115 ;
        RECT 80.215 43.775 80.385 44.155 ;
        RECT 80.600 43.605 80.930 43.985 ;
        RECT 81.100 43.775 81.355 44.350 ;
        RECT 81.530 43.605 81.790 44.445 ;
        RECT 82.655 44.355 83.175 44.895 ;
        RECT 81.965 43.605 83.175 44.355 ;
        RECT 5.520 43.435 83.260 43.605 ;
        RECT 5.605 42.685 6.815 43.435 ;
        RECT 7.035 42.780 7.365 43.215 ;
        RECT 7.535 42.825 7.705 43.435 ;
        RECT 6.985 42.695 7.365 42.780 ;
        RECT 7.875 42.695 8.205 43.220 ;
        RECT 8.465 42.905 8.675 43.435 ;
        RECT 8.950 42.985 9.735 43.155 ;
        RECT 9.905 42.985 10.310 43.155 ;
        RECT 5.605 42.145 6.125 42.685 ;
        RECT 6.985 42.655 7.210 42.695 ;
        RECT 6.295 41.975 6.815 42.515 ;
        RECT 5.605 40.885 6.815 41.975 ;
        RECT 6.985 42.075 7.155 42.655 ;
        RECT 7.875 42.525 8.075 42.695 ;
        RECT 8.950 42.525 9.120 42.985 ;
        RECT 7.325 42.195 8.075 42.525 ;
        RECT 8.245 42.195 9.120 42.525 ;
        RECT 6.985 42.025 7.200 42.075 ;
        RECT 6.985 41.945 7.375 42.025 ;
        RECT 7.045 41.100 7.375 41.945 ;
        RECT 7.885 41.990 8.075 42.195 ;
        RECT 7.545 40.885 7.715 41.895 ;
        RECT 7.885 41.615 8.780 41.990 ;
        RECT 7.885 41.055 8.225 41.615 ;
        RECT 8.455 40.885 8.770 41.385 ;
        RECT 8.950 41.355 9.120 42.195 ;
        RECT 9.290 42.485 9.755 42.815 ;
        RECT 10.140 42.755 10.310 42.985 ;
        RECT 10.490 42.935 10.860 43.435 ;
        RECT 11.180 42.985 11.855 43.155 ;
        RECT 12.050 42.985 12.385 43.155 ;
        RECT 9.290 41.525 9.610 42.485 ;
        RECT 10.140 42.455 10.970 42.755 ;
        RECT 9.780 41.555 9.970 42.275 ;
        RECT 10.140 41.385 10.310 42.455 ;
        RECT 10.770 42.425 10.970 42.455 ;
        RECT 10.480 42.205 10.650 42.275 ;
        RECT 11.180 42.205 11.350 42.985 ;
        RECT 12.215 42.845 12.385 42.985 ;
        RECT 12.555 42.975 12.805 43.435 ;
        RECT 10.480 42.035 11.350 42.205 ;
        RECT 11.520 42.565 12.045 42.785 ;
        RECT 12.215 42.715 12.440 42.845 ;
        RECT 10.480 41.945 10.990 42.035 ;
        RECT 8.950 41.185 9.835 41.355 ;
        RECT 10.060 41.055 10.310 41.385 ;
        RECT 10.480 40.885 10.650 41.685 ;
        RECT 10.820 41.330 10.990 41.945 ;
        RECT 11.520 41.865 11.690 42.565 ;
        RECT 11.160 41.500 11.690 41.865 ;
        RECT 11.860 41.800 12.100 42.395 ;
        RECT 12.270 41.610 12.440 42.715 ;
        RECT 12.610 41.855 12.890 42.805 ;
        RECT 12.135 41.480 12.440 41.610 ;
        RECT 10.820 41.160 11.925 41.330 ;
        RECT 12.135 41.055 12.385 41.480 ;
        RECT 12.555 40.885 12.820 41.345 ;
        RECT 13.060 41.055 13.245 43.175 ;
        RECT 13.415 43.055 13.745 43.435 ;
        RECT 13.915 42.885 14.085 43.175 ;
        RECT 14.345 43.055 15.235 43.225 ;
        RECT 13.420 42.715 14.085 42.885 ;
        RECT 13.420 41.725 13.650 42.715 ;
        RECT 13.820 41.895 14.170 42.545 ;
        RECT 14.345 42.500 14.895 42.885 ;
        RECT 15.065 42.330 15.235 43.055 ;
        RECT 14.345 42.260 15.235 42.330 ;
        RECT 15.405 42.730 15.625 43.215 ;
        RECT 15.795 42.895 16.045 43.435 ;
        RECT 16.215 42.785 16.475 43.265 ;
        RECT 15.405 42.305 15.735 42.730 ;
        RECT 14.345 42.235 15.240 42.260 ;
        RECT 14.345 42.220 15.250 42.235 ;
        RECT 14.345 42.205 15.255 42.220 ;
        RECT 14.345 42.200 15.265 42.205 ;
        RECT 14.345 42.190 15.270 42.200 ;
        RECT 14.345 42.180 15.275 42.190 ;
        RECT 14.345 42.175 15.285 42.180 ;
        RECT 14.345 42.165 15.295 42.175 ;
        RECT 14.345 42.160 15.305 42.165 ;
        RECT 13.420 41.555 14.085 41.725 ;
        RECT 14.345 41.710 14.605 42.160 ;
        RECT 14.970 42.155 15.305 42.160 ;
        RECT 14.970 42.150 15.320 42.155 ;
        RECT 14.970 42.140 15.335 42.150 ;
        RECT 14.970 42.135 15.360 42.140 ;
        RECT 15.905 42.135 16.135 42.530 ;
        RECT 14.970 42.130 16.135 42.135 ;
        RECT 15.000 42.095 16.135 42.130 ;
        RECT 15.035 42.070 16.135 42.095 ;
        RECT 15.065 42.040 16.135 42.070 ;
        RECT 15.085 42.010 16.135 42.040 ;
        RECT 15.105 41.980 16.135 42.010 ;
        RECT 15.175 41.970 16.135 41.980 ;
        RECT 15.200 41.960 16.135 41.970 ;
        RECT 15.220 41.945 16.135 41.960 ;
        RECT 15.240 41.930 16.135 41.945 ;
        RECT 15.245 41.920 16.030 41.930 ;
        RECT 15.260 41.885 16.030 41.920 ;
        RECT 13.415 40.885 13.745 41.385 ;
        RECT 13.915 41.055 14.085 41.555 ;
        RECT 14.775 41.565 15.105 41.810 ;
        RECT 15.275 41.635 16.030 41.885 ;
        RECT 16.305 41.755 16.475 42.785 ;
        RECT 16.665 42.625 16.905 43.435 ;
        RECT 17.075 42.625 17.405 43.265 ;
        RECT 17.575 42.625 17.845 43.435 ;
        RECT 18.025 42.665 21.535 43.435 ;
        RECT 21.740 42.695 22.355 43.265 ;
        RECT 22.525 42.925 22.740 43.435 ;
        RECT 22.970 42.925 23.250 43.255 ;
        RECT 23.430 42.925 23.670 43.435 ;
        RECT 24.005 43.055 24.895 43.225 ;
        RECT 16.645 42.195 16.995 42.445 ;
        RECT 17.165 42.025 17.335 42.625 ;
        RECT 17.505 42.195 17.855 42.445 ;
        RECT 18.025 42.145 19.675 42.665 ;
        RECT 14.775 41.540 14.960 41.565 ;
        RECT 14.345 41.440 14.960 41.540 ;
        RECT 14.345 40.885 14.950 41.440 ;
        RECT 15.125 41.055 15.605 41.395 ;
        RECT 15.775 40.885 16.030 41.430 ;
        RECT 16.200 41.055 16.475 41.755 ;
        RECT 16.655 41.855 17.335 42.025 ;
        RECT 16.655 41.070 16.985 41.855 ;
        RECT 17.515 40.885 17.845 42.025 ;
        RECT 19.845 41.975 21.535 42.495 ;
        RECT 18.025 40.885 21.535 41.975 ;
        RECT 21.740 41.675 22.055 42.695 ;
        RECT 22.225 42.025 22.395 42.525 ;
        RECT 22.645 42.195 22.910 42.755 ;
        RECT 23.080 42.025 23.250 42.925 ;
        RECT 23.420 42.195 23.775 42.755 ;
        RECT 24.005 42.500 24.555 42.885 ;
        RECT 24.725 42.330 24.895 43.055 ;
        RECT 24.005 42.260 24.895 42.330 ;
        RECT 25.065 42.730 25.285 43.215 ;
        RECT 25.455 42.895 25.705 43.435 ;
        RECT 25.875 42.785 26.135 43.265 ;
        RECT 25.065 42.305 25.395 42.730 ;
        RECT 24.005 42.235 24.900 42.260 ;
        RECT 24.005 42.220 24.910 42.235 ;
        RECT 24.005 42.205 24.915 42.220 ;
        RECT 24.005 42.200 24.925 42.205 ;
        RECT 24.005 42.190 24.930 42.200 ;
        RECT 24.005 42.180 24.935 42.190 ;
        RECT 24.005 42.175 24.945 42.180 ;
        RECT 24.005 42.165 24.955 42.175 ;
        RECT 24.005 42.160 24.965 42.165 ;
        RECT 22.225 41.855 23.650 42.025 ;
        RECT 21.740 41.055 22.275 41.675 ;
        RECT 22.445 40.885 22.775 41.685 ;
        RECT 23.260 41.680 23.650 41.855 ;
        RECT 24.005 41.710 24.265 42.160 ;
        RECT 24.630 42.155 24.965 42.160 ;
        RECT 24.630 42.150 24.980 42.155 ;
        RECT 24.630 42.140 24.995 42.150 ;
        RECT 24.630 42.135 25.020 42.140 ;
        RECT 25.565 42.135 25.795 42.530 ;
        RECT 24.630 42.130 25.795 42.135 ;
        RECT 24.660 42.095 25.795 42.130 ;
        RECT 24.695 42.070 25.795 42.095 ;
        RECT 24.725 42.040 25.795 42.070 ;
        RECT 24.745 42.010 25.795 42.040 ;
        RECT 24.765 41.980 25.795 42.010 ;
        RECT 24.835 41.970 25.795 41.980 ;
        RECT 24.860 41.960 25.795 41.970 ;
        RECT 24.880 41.945 25.795 41.960 ;
        RECT 24.900 41.930 25.795 41.945 ;
        RECT 24.905 41.920 25.690 41.930 ;
        RECT 24.920 41.885 25.690 41.920 ;
        RECT 24.435 41.565 24.765 41.810 ;
        RECT 24.935 41.635 25.690 41.885 ;
        RECT 25.965 41.755 26.135 42.785 ;
        RECT 24.435 41.540 24.620 41.565 ;
        RECT 24.005 41.440 24.620 41.540 ;
        RECT 24.005 40.885 24.610 41.440 ;
        RECT 24.785 41.055 25.265 41.395 ;
        RECT 25.435 40.885 25.690 41.430 ;
        RECT 25.860 41.055 26.135 41.755 ;
        RECT 26.305 42.695 26.745 43.255 ;
        RECT 26.915 42.695 27.365 43.435 ;
        RECT 27.535 42.865 27.705 43.265 ;
        RECT 27.875 43.035 28.295 43.435 ;
        RECT 28.465 42.865 28.695 43.265 ;
        RECT 27.535 42.695 28.695 42.865 ;
        RECT 28.865 42.695 29.355 43.265 ;
        RECT 26.305 41.685 26.615 42.695 ;
        RECT 26.785 42.075 26.955 42.525 ;
        RECT 27.125 42.245 27.515 42.525 ;
        RECT 27.700 42.195 27.945 42.525 ;
        RECT 26.785 41.905 27.575 42.075 ;
        RECT 26.305 41.055 26.745 41.685 ;
        RECT 26.920 40.885 27.235 41.735 ;
        RECT 27.405 41.225 27.575 41.905 ;
        RECT 27.745 41.395 27.945 42.195 ;
        RECT 28.145 41.395 28.395 42.525 ;
        RECT 28.610 42.195 29.015 42.525 ;
        RECT 29.185 42.025 29.355 42.695 ;
        RECT 29.525 42.665 31.195 43.435 ;
        RECT 31.365 42.710 31.655 43.435 ;
        RECT 31.825 42.975 32.385 43.265 ;
        RECT 32.555 42.975 32.805 43.435 ;
        RECT 29.525 42.145 30.275 42.665 ;
        RECT 28.585 41.855 29.355 42.025 ;
        RECT 30.445 41.975 31.195 42.495 ;
        RECT 28.585 41.225 28.835 41.855 ;
        RECT 27.405 41.055 28.835 41.225 ;
        RECT 29.015 40.885 29.345 41.685 ;
        RECT 29.525 40.885 31.195 41.975 ;
        RECT 31.365 40.885 31.655 42.050 ;
        RECT 31.825 41.605 32.075 42.975 ;
        RECT 33.425 42.805 33.755 43.165 ;
        RECT 32.365 42.615 33.755 42.805 ;
        RECT 34.675 42.885 34.845 43.175 ;
        RECT 35.015 43.055 35.345 43.435 ;
        RECT 34.675 42.715 35.340 42.885 ;
        RECT 32.365 42.525 32.535 42.615 ;
        RECT 32.245 42.195 32.535 42.525 ;
        RECT 32.705 42.195 33.045 42.445 ;
        RECT 33.265 42.195 33.940 42.445 ;
        RECT 32.365 41.945 32.535 42.195 ;
        RECT 32.365 41.775 33.305 41.945 ;
        RECT 33.675 41.835 33.940 42.195 ;
        RECT 34.590 41.895 34.940 42.545 ;
        RECT 31.825 41.055 32.285 41.605 ;
        RECT 32.475 40.885 32.805 41.605 ;
        RECT 33.005 41.225 33.305 41.775 ;
        RECT 35.110 41.725 35.340 42.715 ;
        RECT 34.675 41.555 35.340 41.725 ;
        RECT 33.475 40.885 33.755 41.555 ;
        RECT 34.675 41.055 34.845 41.555 ;
        RECT 35.015 40.885 35.345 41.385 ;
        RECT 35.515 41.055 35.700 43.175 ;
        RECT 35.955 42.975 36.205 43.435 ;
        RECT 36.375 42.985 36.710 43.155 ;
        RECT 36.905 42.985 37.580 43.155 ;
        RECT 36.375 42.845 36.545 42.985 ;
        RECT 35.870 41.855 36.150 42.805 ;
        RECT 36.320 42.715 36.545 42.845 ;
        RECT 36.320 41.610 36.490 42.715 ;
        RECT 36.715 42.565 37.240 42.785 ;
        RECT 36.660 41.800 36.900 42.395 ;
        RECT 37.070 41.865 37.240 42.565 ;
        RECT 37.410 42.205 37.580 42.985 ;
        RECT 37.900 42.935 38.270 43.435 ;
        RECT 38.450 42.985 38.855 43.155 ;
        RECT 39.025 42.985 39.810 43.155 ;
        RECT 38.450 42.755 38.620 42.985 ;
        RECT 37.790 42.455 38.620 42.755 ;
        RECT 39.005 42.485 39.470 42.815 ;
        RECT 37.790 42.425 37.990 42.455 ;
        RECT 38.110 42.205 38.280 42.275 ;
        RECT 37.410 42.035 38.280 42.205 ;
        RECT 37.770 41.945 38.280 42.035 ;
        RECT 36.320 41.480 36.625 41.610 ;
        RECT 37.070 41.500 37.600 41.865 ;
        RECT 35.940 40.885 36.205 41.345 ;
        RECT 36.375 41.055 36.625 41.480 ;
        RECT 37.770 41.330 37.940 41.945 ;
        RECT 36.835 41.160 37.940 41.330 ;
        RECT 38.110 40.885 38.280 41.685 ;
        RECT 38.450 41.385 38.620 42.455 ;
        RECT 38.790 41.555 38.980 42.275 ;
        RECT 39.150 41.525 39.470 42.485 ;
        RECT 39.640 42.525 39.810 42.985 ;
        RECT 40.085 42.905 40.295 43.435 ;
        RECT 40.555 42.695 40.885 43.220 ;
        RECT 41.055 42.825 41.225 43.435 ;
        RECT 41.395 42.780 41.725 43.215 ;
        RECT 42.035 42.885 42.205 43.175 ;
        RECT 42.375 43.055 42.705 43.435 ;
        RECT 41.395 42.695 41.775 42.780 ;
        RECT 42.035 42.715 42.700 42.885 ;
        RECT 40.685 42.525 40.885 42.695 ;
        RECT 41.550 42.655 41.775 42.695 ;
        RECT 39.640 42.195 40.515 42.525 ;
        RECT 40.685 42.195 41.435 42.525 ;
        RECT 38.450 41.055 38.700 41.385 ;
        RECT 39.640 41.355 39.810 42.195 ;
        RECT 40.685 41.990 40.875 42.195 ;
        RECT 41.605 42.075 41.775 42.655 ;
        RECT 41.560 42.025 41.775 42.075 ;
        RECT 39.980 41.615 40.875 41.990 ;
        RECT 41.385 41.945 41.775 42.025 ;
        RECT 38.925 41.185 39.810 41.355 ;
        RECT 39.990 40.885 40.305 41.385 ;
        RECT 40.535 41.055 40.875 41.615 ;
        RECT 41.045 40.885 41.215 41.895 ;
        RECT 41.385 41.100 41.715 41.945 ;
        RECT 41.950 41.895 42.300 42.545 ;
        RECT 42.470 41.725 42.700 42.715 ;
        RECT 42.035 41.555 42.700 41.725 ;
        RECT 42.035 41.055 42.205 41.555 ;
        RECT 42.375 40.885 42.705 41.385 ;
        RECT 42.875 41.055 43.060 43.175 ;
        RECT 43.315 42.975 43.565 43.435 ;
        RECT 43.735 42.985 44.070 43.155 ;
        RECT 44.265 42.985 44.940 43.155 ;
        RECT 43.735 42.845 43.905 42.985 ;
        RECT 43.230 41.855 43.510 42.805 ;
        RECT 43.680 42.715 43.905 42.845 ;
        RECT 43.680 41.610 43.850 42.715 ;
        RECT 44.075 42.565 44.600 42.785 ;
        RECT 44.020 41.800 44.260 42.395 ;
        RECT 44.430 41.865 44.600 42.565 ;
        RECT 44.770 42.205 44.940 42.985 ;
        RECT 45.260 42.935 45.630 43.435 ;
        RECT 45.810 42.985 46.215 43.155 ;
        RECT 46.385 42.985 47.170 43.155 ;
        RECT 45.810 42.755 45.980 42.985 ;
        RECT 45.150 42.455 45.980 42.755 ;
        RECT 46.365 42.485 46.830 42.815 ;
        RECT 45.150 42.425 45.350 42.455 ;
        RECT 45.470 42.205 45.640 42.275 ;
        RECT 44.770 42.035 45.640 42.205 ;
        RECT 45.130 41.945 45.640 42.035 ;
        RECT 43.680 41.480 43.985 41.610 ;
        RECT 44.430 41.500 44.960 41.865 ;
        RECT 43.300 40.885 43.565 41.345 ;
        RECT 43.735 41.055 43.985 41.480 ;
        RECT 45.130 41.330 45.300 41.945 ;
        RECT 44.195 41.160 45.300 41.330 ;
        RECT 45.470 40.885 45.640 41.685 ;
        RECT 45.810 41.385 45.980 42.455 ;
        RECT 46.150 41.555 46.340 42.275 ;
        RECT 46.510 41.525 46.830 42.485 ;
        RECT 47.000 42.525 47.170 42.985 ;
        RECT 47.445 42.905 47.655 43.435 ;
        RECT 47.915 42.695 48.245 43.220 ;
        RECT 48.415 42.825 48.585 43.435 ;
        RECT 48.755 42.780 49.085 43.215 ;
        RECT 49.315 42.945 49.645 43.435 ;
        RECT 49.815 42.840 50.435 43.265 ;
        RECT 48.755 42.695 49.135 42.780 ;
        RECT 48.045 42.525 48.245 42.695 ;
        RECT 48.910 42.655 49.135 42.695 ;
        RECT 47.000 42.195 47.875 42.525 ;
        RECT 48.045 42.195 48.795 42.525 ;
        RECT 45.810 41.055 46.060 41.385 ;
        RECT 47.000 41.355 47.170 42.195 ;
        RECT 48.045 41.990 48.235 42.195 ;
        RECT 48.965 42.075 49.135 42.655 ;
        RECT 49.305 42.195 49.645 42.775 ;
        RECT 49.815 42.505 50.175 42.840 ;
        RECT 50.895 42.745 51.225 43.435 ;
        RECT 52.070 42.695 52.325 43.265 ;
        RECT 52.495 43.035 52.825 43.435 ;
        RECT 53.250 42.900 53.780 43.265 ;
        RECT 53.970 43.095 54.245 43.265 ;
        RECT 53.965 42.925 54.245 43.095 ;
        RECT 53.250 42.865 53.425 42.900 ;
        RECT 52.495 42.695 53.425 42.865 ;
        RECT 49.815 42.225 51.235 42.505 ;
        RECT 48.920 42.025 49.135 42.075 ;
        RECT 47.340 41.615 48.235 41.990 ;
        RECT 48.745 41.945 49.135 42.025 ;
        RECT 46.285 41.185 47.170 41.355 ;
        RECT 47.350 40.885 47.665 41.385 ;
        RECT 47.895 41.055 48.235 41.615 ;
        RECT 48.405 40.885 48.575 41.895 ;
        RECT 48.745 41.100 49.075 41.945 ;
        RECT 49.315 40.885 49.645 42.025 ;
        RECT 49.815 41.055 50.175 42.225 ;
        RECT 50.375 40.885 50.705 42.055 ;
        RECT 50.905 41.055 51.235 42.225 ;
        RECT 51.435 40.885 51.765 42.055 ;
        RECT 52.070 42.025 52.240 42.695 ;
        RECT 52.495 42.525 52.665 42.695 ;
        RECT 52.410 42.195 52.665 42.525 ;
        RECT 52.890 42.195 53.085 42.525 ;
        RECT 52.070 41.055 52.405 42.025 ;
        RECT 52.575 40.885 52.745 42.025 ;
        RECT 52.915 41.225 53.085 42.195 ;
        RECT 53.255 41.565 53.425 42.695 ;
        RECT 53.595 41.905 53.765 42.705 ;
        RECT 53.970 42.105 54.245 42.925 ;
        RECT 54.415 41.905 54.605 43.265 ;
        RECT 54.785 42.900 55.295 43.435 ;
        RECT 55.515 42.625 55.760 43.230 ;
        RECT 57.125 42.710 57.415 43.435 ;
        RECT 58.510 42.695 58.765 43.265 ;
        RECT 58.935 43.035 59.265 43.435 ;
        RECT 59.690 42.900 60.220 43.265 ;
        RECT 59.690 42.865 59.865 42.900 ;
        RECT 58.935 42.695 59.865 42.865 ;
        RECT 54.805 42.455 56.035 42.625 ;
        RECT 53.595 41.735 54.605 41.905 ;
        RECT 54.775 41.890 55.525 42.080 ;
        RECT 53.255 41.395 54.380 41.565 ;
        RECT 54.775 41.225 54.945 41.890 ;
        RECT 55.695 41.645 56.035 42.455 ;
        RECT 52.915 41.055 54.945 41.225 ;
        RECT 55.115 40.885 55.285 41.645 ;
        RECT 55.520 41.235 56.035 41.645 ;
        RECT 57.125 40.885 57.415 42.050 ;
        RECT 58.510 42.025 58.680 42.695 ;
        RECT 58.935 42.525 59.105 42.695 ;
        RECT 58.850 42.195 59.105 42.525 ;
        RECT 59.330 42.195 59.525 42.525 ;
        RECT 58.510 41.055 58.845 42.025 ;
        RECT 59.015 40.885 59.185 42.025 ;
        RECT 59.355 41.225 59.525 42.195 ;
        RECT 59.695 41.565 59.865 42.695 ;
        RECT 60.035 41.905 60.205 42.705 ;
        RECT 60.410 42.415 60.685 43.265 ;
        RECT 60.405 42.245 60.685 42.415 ;
        RECT 60.410 42.105 60.685 42.245 ;
        RECT 60.855 41.905 61.045 43.265 ;
        RECT 61.225 42.900 61.735 43.435 ;
        RECT 61.955 42.625 62.200 43.230 ;
        RECT 62.650 42.695 62.905 43.265 ;
        RECT 63.075 43.035 63.405 43.435 ;
        RECT 63.830 42.900 64.360 43.265 ;
        RECT 63.830 42.865 64.005 42.900 ;
        RECT 63.075 42.695 64.005 42.865 ;
        RECT 61.245 42.455 62.475 42.625 ;
        RECT 60.035 41.735 61.045 41.905 ;
        RECT 61.215 41.890 61.965 42.080 ;
        RECT 59.695 41.395 60.820 41.565 ;
        RECT 61.215 41.225 61.385 41.890 ;
        RECT 62.135 41.645 62.475 42.455 ;
        RECT 59.355 41.055 61.385 41.225 ;
        RECT 61.555 40.885 61.725 41.645 ;
        RECT 61.960 41.235 62.475 41.645 ;
        RECT 62.650 42.025 62.820 42.695 ;
        RECT 63.075 42.525 63.245 42.695 ;
        RECT 62.990 42.195 63.245 42.525 ;
        RECT 63.470 42.195 63.665 42.525 ;
        RECT 62.650 41.055 62.985 42.025 ;
        RECT 63.155 40.885 63.325 42.025 ;
        RECT 63.495 41.225 63.665 42.195 ;
        RECT 63.835 41.565 64.005 42.695 ;
        RECT 64.175 41.905 64.345 42.705 ;
        RECT 64.550 42.415 64.825 43.265 ;
        RECT 64.545 42.245 64.825 42.415 ;
        RECT 64.550 42.105 64.825 42.245 ;
        RECT 64.995 41.905 65.185 43.265 ;
        RECT 65.365 42.900 65.875 43.435 ;
        RECT 66.095 42.625 66.340 43.230 ;
        RECT 66.785 42.635 67.125 43.265 ;
        RECT 67.295 42.635 67.545 43.435 ;
        RECT 67.735 42.785 68.065 43.265 ;
        RECT 68.235 42.975 68.460 43.435 ;
        RECT 68.630 42.785 68.960 43.265 ;
        RECT 65.385 42.455 66.615 42.625 ;
        RECT 64.175 41.735 65.185 41.905 ;
        RECT 65.355 41.890 66.105 42.080 ;
        RECT 63.835 41.395 64.960 41.565 ;
        RECT 65.355 41.225 65.525 41.890 ;
        RECT 66.275 41.645 66.615 42.455 ;
        RECT 63.495 41.055 65.525 41.225 ;
        RECT 65.695 40.885 65.865 41.645 ;
        RECT 66.100 41.235 66.615 41.645 ;
        RECT 66.785 42.025 66.960 42.635 ;
        RECT 67.735 42.615 68.960 42.785 ;
        RECT 69.590 42.655 70.090 43.265 ;
        RECT 71.130 42.655 71.630 43.265 ;
        RECT 67.130 42.275 67.825 42.445 ;
        RECT 67.655 42.025 67.825 42.275 ;
        RECT 68.000 42.245 68.420 42.445 ;
        RECT 68.590 42.245 68.920 42.445 ;
        RECT 69.090 42.245 69.420 42.445 ;
        RECT 69.590 42.025 69.760 42.655 ;
        RECT 69.945 42.195 70.295 42.445 ;
        RECT 70.925 42.195 71.275 42.445 ;
        RECT 71.460 42.025 71.630 42.655 ;
        RECT 72.260 42.785 72.590 43.265 ;
        RECT 72.760 42.975 72.985 43.435 ;
        RECT 73.155 42.785 73.485 43.265 ;
        RECT 72.260 42.615 73.485 42.785 ;
        RECT 73.675 42.635 73.925 43.435 ;
        RECT 74.095 42.635 74.435 43.265 ;
        RECT 74.695 42.885 74.865 43.175 ;
        RECT 75.035 43.055 75.365 43.435 ;
        RECT 74.695 42.715 75.360 42.885 ;
        RECT 71.800 42.245 72.130 42.445 ;
        RECT 72.300 42.245 72.630 42.445 ;
        RECT 72.800 42.245 73.220 42.445 ;
        RECT 73.395 42.275 74.090 42.445 ;
        RECT 73.395 42.025 73.565 42.275 ;
        RECT 74.260 42.025 74.435 42.635 ;
        RECT 66.785 41.055 67.125 42.025 ;
        RECT 67.295 40.885 67.465 42.025 ;
        RECT 67.655 41.855 70.090 42.025 ;
        RECT 67.735 40.885 67.985 41.685 ;
        RECT 68.630 41.055 68.960 41.855 ;
        RECT 69.260 40.885 69.590 41.685 ;
        RECT 69.760 41.055 70.090 41.855 ;
        RECT 71.130 41.855 73.565 42.025 ;
        RECT 71.130 41.055 71.460 41.855 ;
        RECT 71.630 40.885 71.960 41.685 ;
        RECT 72.260 41.055 72.590 41.855 ;
        RECT 73.235 40.885 73.485 41.685 ;
        RECT 73.755 40.885 73.925 42.025 ;
        RECT 74.095 41.055 74.435 42.025 ;
        RECT 74.610 41.895 74.960 42.545 ;
        RECT 75.130 41.725 75.360 42.715 ;
        RECT 74.695 41.555 75.360 41.725 ;
        RECT 74.695 41.055 74.865 41.555 ;
        RECT 75.035 40.885 75.365 41.385 ;
        RECT 75.535 41.055 75.720 43.175 ;
        RECT 75.975 42.975 76.225 43.435 ;
        RECT 76.395 42.985 76.730 43.155 ;
        RECT 76.925 42.985 77.600 43.155 ;
        RECT 76.395 42.845 76.565 42.985 ;
        RECT 75.890 41.855 76.170 42.805 ;
        RECT 76.340 42.715 76.565 42.845 ;
        RECT 76.340 41.610 76.510 42.715 ;
        RECT 76.735 42.565 77.260 42.785 ;
        RECT 76.680 41.800 76.920 42.395 ;
        RECT 77.090 41.865 77.260 42.565 ;
        RECT 77.430 42.205 77.600 42.985 ;
        RECT 77.920 42.935 78.290 43.435 ;
        RECT 78.470 42.985 78.875 43.155 ;
        RECT 79.045 42.985 79.830 43.155 ;
        RECT 78.470 42.755 78.640 42.985 ;
        RECT 77.810 42.455 78.640 42.755 ;
        RECT 79.025 42.485 79.490 42.815 ;
        RECT 77.810 42.425 78.010 42.455 ;
        RECT 78.130 42.205 78.300 42.275 ;
        RECT 77.430 42.035 78.300 42.205 ;
        RECT 77.790 41.945 78.300 42.035 ;
        RECT 76.340 41.480 76.645 41.610 ;
        RECT 77.090 41.500 77.620 41.865 ;
        RECT 75.960 40.885 76.225 41.345 ;
        RECT 76.395 41.055 76.645 41.480 ;
        RECT 77.790 41.330 77.960 41.945 ;
        RECT 76.855 41.160 77.960 41.330 ;
        RECT 78.130 40.885 78.300 41.685 ;
        RECT 78.470 41.385 78.640 42.455 ;
        RECT 78.810 41.555 79.000 42.275 ;
        RECT 79.170 41.525 79.490 42.485 ;
        RECT 79.660 42.525 79.830 42.985 ;
        RECT 80.105 42.905 80.315 43.435 ;
        RECT 80.575 42.695 80.905 43.220 ;
        RECT 81.075 42.825 81.245 43.435 ;
        RECT 81.415 42.780 81.745 43.215 ;
        RECT 81.415 42.695 81.795 42.780 ;
        RECT 80.705 42.525 80.905 42.695 ;
        RECT 81.570 42.655 81.795 42.695 ;
        RECT 81.965 42.685 83.175 43.435 ;
        RECT 79.660 42.195 80.535 42.525 ;
        RECT 80.705 42.195 81.455 42.525 ;
        RECT 78.470 41.055 78.720 41.385 ;
        RECT 79.660 41.355 79.830 42.195 ;
        RECT 80.705 41.990 80.895 42.195 ;
        RECT 81.625 42.075 81.795 42.655 ;
        RECT 81.580 42.025 81.795 42.075 ;
        RECT 80.000 41.615 80.895 41.990 ;
        RECT 81.405 41.945 81.795 42.025 ;
        RECT 81.965 41.975 82.485 42.515 ;
        RECT 82.655 42.145 83.175 42.685 ;
        RECT 78.945 41.185 79.830 41.355 ;
        RECT 80.010 40.885 80.325 41.385 ;
        RECT 80.555 41.055 80.895 41.615 ;
        RECT 81.065 40.885 81.235 41.895 ;
        RECT 81.405 41.100 81.735 41.945 ;
        RECT 81.965 40.885 83.175 41.975 ;
        RECT 5.520 40.715 83.260 40.885 ;
        RECT 5.605 39.625 6.815 40.715 ;
        RECT 7.995 40.045 8.165 40.545 ;
        RECT 8.335 40.215 8.665 40.715 ;
        RECT 7.995 39.875 8.660 40.045 ;
        RECT 5.605 38.915 6.125 39.455 ;
        RECT 6.295 39.085 6.815 39.625 ;
        RECT 7.910 39.055 8.260 39.705 ;
        RECT 5.605 38.165 6.815 38.915 ;
        RECT 8.430 38.885 8.660 39.875 ;
        RECT 7.995 38.715 8.660 38.885 ;
        RECT 7.995 38.425 8.165 38.715 ;
        RECT 8.335 38.165 8.665 38.545 ;
        RECT 8.835 38.425 9.020 40.545 ;
        RECT 9.260 40.255 9.525 40.715 ;
        RECT 9.695 40.120 9.945 40.545 ;
        RECT 10.155 40.270 11.260 40.440 ;
        RECT 9.640 39.990 9.945 40.120 ;
        RECT 9.190 38.795 9.470 39.745 ;
        RECT 9.640 38.885 9.810 39.990 ;
        RECT 9.980 39.205 10.220 39.800 ;
        RECT 10.390 39.735 10.920 40.100 ;
        RECT 10.390 39.035 10.560 39.735 ;
        RECT 11.090 39.655 11.260 40.270 ;
        RECT 11.430 39.915 11.600 40.715 ;
        RECT 11.770 40.215 12.020 40.545 ;
        RECT 12.245 40.245 13.130 40.415 ;
        RECT 11.090 39.565 11.600 39.655 ;
        RECT 9.640 38.755 9.865 38.885 ;
        RECT 10.035 38.815 10.560 39.035 ;
        RECT 10.730 39.395 11.600 39.565 ;
        RECT 9.275 38.165 9.525 38.625 ;
        RECT 9.695 38.615 9.865 38.755 ;
        RECT 10.730 38.615 10.900 39.395 ;
        RECT 11.430 39.325 11.600 39.395 ;
        RECT 11.110 39.145 11.310 39.175 ;
        RECT 11.770 39.145 11.940 40.215 ;
        RECT 12.110 39.325 12.300 40.045 ;
        RECT 11.110 38.845 11.940 39.145 ;
        RECT 12.470 39.115 12.790 40.075 ;
        RECT 9.695 38.445 10.030 38.615 ;
        RECT 10.225 38.445 10.900 38.615 ;
        RECT 11.220 38.165 11.590 38.665 ;
        RECT 11.770 38.615 11.940 38.845 ;
        RECT 12.325 38.785 12.790 39.115 ;
        RECT 12.960 39.405 13.130 40.245 ;
        RECT 13.310 40.215 13.625 40.715 ;
        RECT 13.855 39.985 14.195 40.545 ;
        RECT 13.300 39.610 14.195 39.985 ;
        RECT 14.365 39.705 14.535 40.715 ;
        RECT 14.005 39.405 14.195 39.610 ;
        RECT 14.705 39.655 15.035 40.500 ;
        RECT 15.265 40.285 15.605 40.545 ;
        RECT 14.705 39.575 15.095 39.655 ;
        RECT 14.880 39.525 15.095 39.575 ;
        RECT 12.960 39.075 13.835 39.405 ;
        RECT 14.005 39.075 14.755 39.405 ;
        RECT 12.960 38.615 13.130 39.075 ;
        RECT 14.005 38.905 14.205 39.075 ;
        RECT 14.925 38.945 15.095 39.525 ;
        RECT 14.870 38.905 15.095 38.945 ;
        RECT 11.770 38.445 12.175 38.615 ;
        RECT 12.345 38.445 13.130 38.615 ;
        RECT 13.405 38.165 13.615 38.695 ;
        RECT 13.875 38.380 14.205 38.905 ;
        RECT 14.715 38.820 15.095 38.905 ;
        RECT 15.265 38.885 15.525 40.285 ;
        RECT 15.775 39.915 16.105 40.715 ;
        RECT 16.570 39.745 16.820 40.545 ;
        RECT 17.005 39.995 17.335 40.715 ;
        RECT 17.555 39.745 17.805 40.545 ;
        RECT 17.975 40.335 18.310 40.715 ;
        RECT 15.715 39.575 17.905 39.745 ;
        RECT 15.715 39.405 16.030 39.575 ;
        RECT 15.700 39.155 16.030 39.405 ;
        RECT 14.375 38.165 14.545 38.775 ;
        RECT 14.715 38.385 15.045 38.820 ;
        RECT 15.265 38.375 15.605 38.885 ;
        RECT 15.775 38.165 16.045 38.965 ;
        RECT 16.225 38.435 16.505 39.405 ;
        RECT 16.685 38.435 16.985 39.405 ;
        RECT 17.165 38.440 17.515 39.405 ;
        RECT 17.735 38.665 17.905 39.575 ;
        RECT 18.075 38.845 18.315 40.155 ;
        RECT 18.485 39.550 18.775 40.715 ;
        RECT 18.955 40.105 19.285 40.535 ;
        RECT 19.465 40.275 19.660 40.715 ;
        RECT 19.830 40.105 20.160 40.535 ;
        RECT 18.955 39.935 20.160 40.105 ;
        RECT 18.955 39.605 19.850 39.935 ;
        RECT 20.330 39.765 20.605 40.535 ;
        RECT 20.020 39.575 20.605 39.765 ;
        RECT 20.795 39.745 21.125 40.530 ;
        RECT 20.795 39.575 21.475 39.745 ;
        RECT 21.655 39.575 21.985 40.715 ;
        RECT 22.165 39.625 25.675 40.715 ;
        RECT 18.960 39.075 19.255 39.405 ;
        RECT 19.435 39.075 19.850 39.405 ;
        RECT 17.735 38.335 18.230 38.665 ;
        RECT 18.485 38.165 18.775 38.890 ;
        RECT 18.955 38.165 19.255 38.895 ;
        RECT 19.435 38.455 19.665 39.075 ;
        RECT 20.020 38.905 20.195 39.575 ;
        RECT 19.865 38.725 20.195 38.905 ;
        RECT 20.365 38.755 20.605 39.405 ;
        RECT 20.785 39.155 21.135 39.405 ;
        RECT 21.305 38.975 21.475 39.575 ;
        RECT 21.645 39.155 21.995 39.405 ;
        RECT 19.865 38.345 20.090 38.725 ;
        RECT 20.260 38.165 20.590 38.555 ;
        RECT 20.805 38.165 21.045 38.975 ;
        RECT 21.215 38.335 21.545 38.975 ;
        RECT 21.715 38.165 21.985 38.975 ;
        RECT 22.165 38.935 23.815 39.455 ;
        RECT 23.985 39.105 25.675 39.625 ;
        RECT 25.845 39.845 26.120 40.545 ;
        RECT 26.330 40.170 26.545 40.715 ;
        RECT 26.715 40.205 27.190 40.545 ;
        RECT 27.360 40.210 27.975 40.715 ;
        RECT 27.360 40.035 27.555 40.210 ;
        RECT 22.165 38.165 25.675 38.935 ;
        RECT 25.845 38.815 26.015 39.845 ;
        RECT 26.290 39.675 27.005 39.970 ;
        RECT 27.225 39.845 27.555 40.035 ;
        RECT 27.725 39.675 27.975 40.040 ;
        RECT 26.185 39.505 27.975 39.675 ;
        RECT 26.185 39.075 26.415 39.505 ;
        RECT 25.845 38.335 26.105 38.815 ;
        RECT 26.585 38.805 26.995 39.325 ;
        RECT 26.275 38.165 26.605 38.625 ;
        RECT 26.795 38.385 26.995 38.805 ;
        RECT 27.165 38.650 27.420 39.505 ;
        RECT 28.215 39.325 28.385 40.545 ;
        RECT 28.635 40.205 28.895 40.715 ;
        RECT 29.065 40.285 29.405 40.545 ;
        RECT 27.590 39.075 28.385 39.325 ;
        RECT 28.555 39.155 28.895 40.035 ;
        RECT 28.135 38.985 28.385 39.075 ;
        RECT 27.165 38.385 27.955 38.650 ;
        RECT 28.135 38.565 28.465 38.985 ;
        RECT 28.635 38.165 28.895 38.985 ;
        RECT 29.065 38.885 29.325 40.285 ;
        RECT 29.575 39.915 29.905 40.715 ;
        RECT 30.370 39.745 30.620 40.545 ;
        RECT 30.805 39.995 31.135 40.715 ;
        RECT 31.355 39.745 31.605 40.545 ;
        RECT 31.775 40.335 32.110 40.715 ;
        RECT 29.515 39.575 31.705 39.745 ;
        RECT 29.515 39.405 29.830 39.575 ;
        RECT 29.500 39.155 29.830 39.405 ;
        RECT 29.065 38.375 29.405 38.885 ;
        RECT 29.575 38.165 29.845 38.965 ;
        RECT 30.025 38.435 30.305 39.405 ;
        RECT 30.485 38.435 30.785 39.405 ;
        RECT 30.965 38.440 31.315 39.405 ;
        RECT 31.535 38.665 31.705 39.575 ;
        RECT 31.875 38.845 32.115 40.155 ;
        RECT 32.295 39.655 32.625 40.505 ;
        RECT 32.295 38.890 32.485 39.655 ;
        RECT 32.795 39.575 33.045 40.715 ;
        RECT 33.235 40.075 33.485 40.495 ;
        RECT 33.715 40.245 34.045 40.715 ;
        RECT 34.275 40.075 34.525 40.495 ;
        RECT 33.235 39.905 34.525 40.075 ;
        RECT 34.705 40.075 35.035 40.505 ;
        RECT 34.705 39.905 35.160 40.075 ;
        RECT 33.225 39.405 33.440 39.735 ;
        RECT 32.655 39.075 32.965 39.405 ;
        RECT 33.135 39.075 33.440 39.405 ;
        RECT 33.615 39.075 33.900 39.735 ;
        RECT 34.095 39.075 34.360 39.735 ;
        RECT 34.575 39.075 34.820 39.735 ;
        RECT 32.795 38.905 32.965 39.075 ;
        RECT 34.990 38.905 35.160 39.905 ;
        RECT 31.535 38.335 32.030 38.665 ;
        RECT 32.295 38.380 32.625 38.890 ;
        RECT 32.795 38.735 35.160 38.905 ;
        RECT 35.540 39.925 36.075 40.545 ;
        RECT 35.540 38.905 35.855 39.925 ;
        RECT 36.245 39.915 36.575 40.715 ;
        RECT 37.060 39.745 37.450 39.920 ;
        RECT 36.025 39.575 37.450 39.745 ;
        RECT 37.805 39.625 39.015 40.715 ;
        RECT 36.025 39.075 36.195 39.575 ;
        RECT 32.795 38.165 33.125 38.565 ;
        RECT 34.175 38.395 34.505 38.735 ;
        RECT 34.675 38.165 35.005 38.565 ;
        RECT 35.540 38.335 36.155 38.905 ;
        RECT 36.445 38.845 36.710 39.405 ;
        RECT 36.880 38.675 37.050 39.575 ;
        RECT 37.220 38.845 37.575 39.405 ;
        RECT 37.805 38.915 38.325 39.455 ;
        RECT 38.495 39.085 39.015 39.625 ;
        RECT 39.185 39.575 39.465 40.715 ;
        RECT 39.635 39.565 39.965 40.545 ;
        RECT 40.135 39.575 40.395 40.715 ;
        RECT 40.565 39.575 40.950 40.545 ;
        RECT 41.120 40.255 41.445 40.715 ;
        RECT 41.965 40.085 42.245 40.545 ;
        RECT 41.120 39.865 42.245 40.085 ;
        RECT 39.195 39.135 39.530 39.405 ;
        RECT 39.700 38.965 39.870 39.565 ;
        RECT 40.040 39.155 40.375 39.405 ;
        RECT 36.325 38.165 36.540 38.675 ;
        RECT 36.770 38.345 37.050 38.675 ;
        RECT 37.230 38.165 37.470 38.675 ;
        RECT 37.805 38.165 39.015 38.915 ;
        RECT 39.185 38.165 39.495 38.965 ;
        RECT 39.700 38.335 40.395 38.965 ;
        RECT 40.565 38.905 40.845 39.575 ;
        RECT 41.120 39.405 41.570 39.865 ;
        RECT 42.435 39.695 42.835 40.545 ;
        RECT 43.235 40.255 43.505 40.715 ;
        RECT 43.675 40.085 43.960 40.545 ;
        RECT 41.015 39.075 41.570 39.405 ;
        RECT 41.740 39.135 42.835 39.695 ;
        RECT 41.120 38.965 41.570 39.075 ;
        RECT 40.565 38.335 40.950 38.905 ;
        RECT 41.120 38.795 42.245 38.965 ;
        RECT 41.120 38.165 41.445 38.625 ;
        RECT 41.965 38.335 42.245 38.795 ;
        RECT 42.435 38.335 42.835 39.135 ;
        RECT 43.005 39.865 43.960 40.085 ;
        RECT 43.005 38.965 43.215 39.865 ;
        RECT 43.385 39.135 44.075 39.695 ;
        RECT 44.245 39.550 44.535 40.715 ;
        RECT 44.710 39.575 44.985 40.545 ;
        RECT 45.195 39.915 45.475 40.715 ;
        RECT 45.645 40.205 46.835 40.495 ;
        RECT 45.645 39.865 46.815 40.035 ;
        RECT 45.645 39.745 45.815 39.865 ;
        RECT 45.155 39.575 45.815 39.745 ;
        RECT 43.005 38.795 43.960 38.965 ;
        RECT 43.235 38.165 43.505 38.625 ;
        RECT 43.675 38.335 43.960 38.795 ;
        RECT 44.245 38.165 44.535 38.890 ;
        RECT 44.710 38.840 44.880 39.575 ;
        RECT 45.155 39.405 45.325 39.575 ;
        RECT 46.125 39.405 46.320 39.695 ;
        RECT 46.490 39.575 46.815 39.865 ;
        RECT 47.525 39.655 47.855 40.500 ;
        RECT 48.025 39.705 48.195 40.715 ;
        RECT 48.365 39.985 48.705 40.545 ;
        RECT 48.935 40.215 49.250 40.715 ;
        RECT 49.430 40.245 50.315 40.415 ;
        RECT 47.465 39.575 47.855 39.655 ;
        RECT 48.365 39.610 49.260 39.985 ;
        RECT 47.465 39.525 47.680 39.575 ;
        RECT 45.050 39.075 45.325 39.405 ;
        RECT 45.495 39.075 46.320 39.405 ;
        RECT 46.490 39.075 46.835 39.405 ;
        RECT 45.155 38.905 45.325 39.075 ;
        RECT 47.465 38.945 47.635 39.525 ;
        RECT 48.365 39.405 48.555 39.610 ;
        RECT 49.430 39.405 49.600 40.245 ;
        RECT 50.540 40.215 50.790 40.545 ;
        RECT 47.805 39.075 48.555 39.405 ;
        RECT 48.725 39.075 49.600 39.405 ;
        RECT 47.465 38.905 47.690 38.945 ;
        RECT 48.355 38.905 48.555 39.075 ;
        RECT 44.710 38.495 44.985 38.840 ;
        RECT 45.155 38.735 46.820 38.905 ;
        RECT 47.465 38.820 47.845 38.905 ;
        RECT 45.175 38.165 45.555 38.565 ;
        RECT 45.725 38.385 45.895 38.735 ;
        RECT 46.065 38.165 46.395 38.565 ;
        RECT 46.565 38.385 46.820 38.735 ;
        RECT 47.515 38.385 47.845 38.820 ;
        RECT 48.015 38.165 48.185 38.775 ;
        RECT 48.355 38.380 48.685 38.905 ;
        RECT 48.945 38.165 49.155 38.695 ;
        RECT 49.430 38.615 49.600 39.075 ;
        RECT 49.770 39.115 50.090 40.075 ;
        RECT 50.260 39.325 50.450 40.045 ;
        RECT 50.620 39.145 50.790 40.215 ;
        RECT 50.960 39.915 51.130 40.715 ;
        RECT 51.300 40.270 52.405 40.440 ;
        RECT 51.300 39.655 51.470 40.270 ;
        RECT 52.615 40.120 52.865 40.545 ;
        RECT 53.035 40.255 53.300 40.715 ;
        RECT 51.640 39.735 52.170 40.100 ;
        RECT 52.615 39.990 52.920 40.120 ;
        RECT 50.960 39.565 51.470 39.655 ;
        RECT 50.960 39.395 51.830 39.565 ;
        RECT 50.960 39.325 51.130 39.395 ;
        RECT 51.250 39.145 51.450 39.175 ;
        RECT 49.770 38.785 50.235 39.115 ;
        RECT 50.620 38.845 51.450 39.145 ;
        RECT 50.620 38.615 50.790 38.845 ;
        RECT 49.430 38.445 50.215 38.615 ;
        RECT 50.385 38.445 50.790 38.615 ;
        RECT 50.970 38.165 51.340 38.665 ;
        RECT 51.660 38.615 51.830 39.395 ;
        RECT 52.000 39.035 52.170 39.735 ;
        RECT 52.340 39.205 52.580 39.800 ;
        RECT 52.000 38.815 52.525 39.035 ;
        RECT 52.750 38.885 52.920 39.990 ;
        RECT 52.695 38.755 52.920 38.885 ;
        RECT 53.090 38.795 53.370 39.745 ;
        RECT 52.695 38.615 52.865 38.755 ;
        RECT 51.660 38.445 52.335 38.615 ;
        RECT 52.530 38.445 52.865 38.615 ;
        RECT 53.035 38.165 53.285 38.625 ;
        RECT 53.540 38.425 53.725 40.545 ;
        RECT 53.895 40.215 54.225 40.715 ;
        RECT 54.395 40.045 54.565 40.545 ;
        RECT 54.825 40.205 56.020 40.495 ;
        RECT 53.900 39.875 54.565 40.045 ;
        RECT 53.900 38.885 54.130 39.875 ;
        RECT 54.845 39.865 56.010 40.035 ;
        RECT 56.190 39.915 56.470 40.715 ;
        RECT 54.300 39.055 54.650 39.705 ;
        RECT 54.845 39.575 55.175 39.865 ;
        RECT 55.840 39.745 56.010 39.865 ;
        RECT 55.345 39.405 55.570 39.695 ;
        RECT 55.840 39.575 56.510 39.745 ;
        RECT 56.680 39.575 56.955 40.545 ;
        RECT 56.340 39.405 56.510 39.575 ;
        RECT 54.825 39.075 55.175 39.405 ;
        RECT 55.345 39.075 56.170 39.405 ;
        RECT 56.340 39.075 56.615 39.405 ;
        RECT 56.340 38.905 56.510 39.075 ;
        RECT 53.900 38.715 54.565 38.885 ;
        RECT 53.895 38.165 54.225 38.545 ;
        RECT 54.395 38.425 54.565 38.715 ;
        RECT 54.845 38.735 56.510 38.905 ;
        RECT 56.785 38.840 56.955 39.575 ;
        RECT 57.125 39.510 57.415 40.715 ;
        RECT 57.675 40.045 57.845 40.545 ;
        RECT 58.015 40.215 58.345 40.715 ;
        RECT 57.675 39.875 58.340 40.045 ;
        RECT 57.590 39.055 57.940 39.705 ;
        RECT 54.845 38.385 55.100 38.735 ;
        RECT 55.270 38.165 55.600 38.565 ;
        RECT 55.770 38.385 55.940 38.735 ;
        RECT 56.110 38.165 56.490 38.565 ;
        RECT 56.680 38.495 56.955 38.840 ;
        RECT 57.125 38.165 57.415 38.995 ;
        RECT 58.110 38.885 58.340 39.875 ;
        RECT 57.675 38.715 58.340 38.885 ;
        RECT 57.675 38.425 57.845 38.715 ;
        RECT 58.015 38.165 58.345 38.545 ;
        RECT 58.515 38.425 58.700 40.545 ;
        RECT 58.940 40.255 59.205 40.715 ;
        RECT 59.375 40.120 59.625 40.545 ;
        RECT 59.835 40.270 60.940 40.440 ;
        RECT 59.320 39.990 59.625 40.120 ;
        RECT 58.870 38.795 59.150 39.745 ;
        RECT 59.320 38.885 59.490 39.990 ;
        RECT 59.660 39.205 59.900 39.800 ;
        RECT 60.070 39.735 60.600 40.100 ;
        RECT 60.070 39.035 60.240 39.735 ;
        RECT 60.770 39.655 60.940 40.270 ;
        RECT 61.110 39.915 61.280 40.715 ;
        RECT 61.450 40.215 61.700 40.545 ;
        RECT 61.925 40.245 62.810 40.415 ;
        RECT 60.770 39.565 61.280 39.655 ;
        RECT 59.320 38.755 59.545 38.885 ;
        RECT 59.715 38.815 60.240 39.035 ;
        RECT 60.410 39.395 61.280 39.565 ;
        RECT 58.955 38.165 59.205 38.625 ;
        RECT 59.375 38.615 59.545 38.755 ;
        RECT 60.410 38.615 60.580 39.395 ;
        RECT 61.110 39.325 61.280 39.395 ;
        RECT 60.790 39.145 60.990 39.175 ;
        RECT 61.450 39.145 61.620 40.215 ;
        RECT 61.790 39.325 61.980 40.045 ;
        RECT 60.790 38.845 61.620 39.145 ;
        RECT 62.150 39.115 62.470 40.075 ;
        RECT 59.375 38.445 59.710 38.615 ;
        RECT 59.905 38.445 60.580 38.615 ;
        RECT 60.900 38.165 61.270 38.665 ;
        RECT 61.450 38.615 61.620 38.845 ;
        RECT 62.005 38.785 62.470 39.115 ;
        RECT 62.640 39.405 62.810 40.245 ;
        RECT 62.990 40.215 63.305 40.715 ;
        RECT 63.535 39.985 63.875 40.545 ;
        RECT 62.980 39.610 63.875 39.985 ;
        RECT 64.045 39.705 64.215 40.715 ;
        RECT 63.685 39.405 63.875 39.610 ;
        RECT 64.385 39.655 64.715 40.500 ;
        RECT 64.885 39.800 65.055 40.715 ;
        RECT 64.385 39.575 64.775 39.655 ;
        RECT 64.560 39.525 64.775 39.575 ;
        RECT 62.640 39.075 63.515 39.405 ;
        RECT 63.685 39.075 64.435 39.405 ;
        RECT 62.640 38.615 62.810 39.075 ;
        RECT 63.685 38.905 63.885 39.075 ;
        RECT 64.605 38.945 64.775 39.525 ;
        RECT 64.550 38.905 64.775 38.945 ;
        RECT 61.450 38.445 61.855 38.615 ;
        RECT 62.025 38.445 62.810 38.615 ;
        RECT 63.085 38.165 63.295 38.695 ;
        RECT 63.555 38.380 63.885 38.905 ;
        RECT 64.395 38.820 64.775 38.905 ;
        RECT 65.405 39.575 65.680 40.545 ;
        RECT 65.890 39.915 66.170 40.715 ;
        RECT 66.340 40.205 67.955 40.535 ;
        RECT 66.340 39.865 67.515 40.035 ;
        RECT 66.340 39.745 66.510 39.865 ;
        RECT 65.850 39.575 66.510 39.745 ;
        RECT 65.405 38.840 65.575 39.575 ;
        RECT 65.850 39.405 66.020 39.575 ;
        RECT 66.770 39.405 67.015 39.695 ;
        RECT 67.185 39.575 67.515 39.865 ;
        RECT 67.775 39.405 67.945 39.965 ;
        RECT 68.195 39.575 68.455 40.715 ;
        RECT 68.625 39.625 69.835 40.715 ;
        RECT 65.745 39.075 66.020 39.405 ;
        RECT 66.190 39.075 67.015 39.405 ;
        RECT 67.230 39.075 67.945 39.405 ;
        RECT 68.115 39.155 68.450 39.405 ;
        RECT 65.850 38.905 66.020 39.075 ;
        RECT 67.695 38.985 67.945 39.075 ;
        RECT 64.055 38.165 64.225 38.775 ;
        RECT 64.395 38.385 64.725 38.820 ;
        RECT 64.895 38.165 65.065 38.680 ;
        RECT 65.405 38.495 65.680 38.840 ;
        RECT 65.850 38.735 67.515 38.905 ;
        RECT 65.870 38.165 66.245 38.565 ;
        RECT 66.415 38.385 66.585 38.735 ;
        RECT 66.755 38.165 67.085 38.565 ;
        RECT 67.255 38.335 67.515 38.735 ;
        RECT 67.695 38.565 68.025 38.985 ;
        RECT 68.195 38.165 68.455 38.985 ;
        RECT 68.625 38.915 69.145 39.455 ;
        RECT 69.315 39.085 69.835 39.625 ;
        RECT 70.005 39.550 70.295 40.715 ;
        RECT 70.670 39.745 71.000 40.545 ;
        RECT 71.170 39.915 71.500 40.715 ;
        RECT 71.800 39.745 72.130 40.545 ;
        RECT 72.775 39.915 73.025 40.715 ;
        RECT 70.670 39.575 73.105 39.745 ;
        RECT 73.295 39.575 73.465 40.715 ;
        RECT 73.635 39.575 73.975 40.545 ;
        RECT 74.695 40.045 74.865 40.545 ;
        RECT 75.035 40.215 75.365 40.715 ;
        RECT 74.695 39.875 75.360 40.045 ;
        RECT 70.465 39.155 70.815 39.405 ;
        RECT 71.000 38.945 71.170 39.575 ;
        RECT 71.340 39.155 71.670 39.355 ;
        RECT 71.840 39.155 72.170 39.355 ;
        RECT 72.340 39.155 72.760 39.355 ;
        RECT 72.935 39.325 73.105 39.575 ;
        RECT 72.935 39.155 73.630 39.325 ;
        RECT 68.625 38.165 69.835 38.915 ;
        RECT 70.005 38.165 70.295 38.890 ;
        RECT 70.670 38.335 71.170 38.945 ;
        RECT 71.800 38.815 73.025 38.985 ;
        RECT 73.800 38.965 73.975 39.575 ;
        RECT 74.610 39.055 74.960 39.705 ;
        RECT 71.800 38.335 72.130 38.815 ;
        RECT 72.300 38.165 72.525 38.625 ;
        RECT 72.695 38.335 73.025 38.815 ;
        RECT 73.215 38.165 73.465 38.965 ;
        RECT 73.635 38.335 73.975 38.965 ;
        RECT 75.130 38.885 75.360 39.875 ;
        RECT 74.695 38.715 75.360 38.885 ;
        RECT 74.695 38.425 74.865 38.715 ;
        RECT 75.035 38.165 75.365 38.545 ;
        RECT 75.535 38.425 75.720 40.545 ;
        RECT 75.960 40.255 76.225 40.715 ;
        RECT 76.395 40.120 76.645 40.545 ;
        RECT 76.855 40.270 77.960 40.440 ;
        RECT 76.340 39.990 76.645 40.120 ;
        RECT 75.890 38.795 76.170 39.745 ;
        RECT 76.340 38.885 76.510 39.990 ;
        RECT 76.680 39.205 76.920 39.800 ;
        RECT 77.090 39.735 77.620 40.100 ;
        RECT 77.090 39.035 77.260 39.735 ;
        RECT 77.790 39.655 77.960 40.270 ;
        RECT 78.130 39.915 78.300 40.715 ;
        RECT 78.470 40.215 78.720 40.545 ;
        RECT 78.945 40.245 79.830 40.415 ;
        RECT 77.790 39.565 78.300 39.655 ;
        RECT 76.340 38.755 76.565 38.885 ;
        RECT 76.735 38.815 77.260 39.035 ;
        RECT 77.430 39.395 78.300 39.565 ;
        RECT 75.975 38.165 76.225 38.625 ;
        RECT 76.395 38.615 76.565 38.755 ;
        RECT 77.430 38.615 77.600 39.395 ;
        RECT 78.130 39.325 78.300 39.395 ;
        RECT 77.810 39.145 78.010 39.175 ;
        RECT 78.470 39.145 78.640 40.215 ;
        RECT 78.810 39.325 79.000 40.045 ;
        RECT 77.810 38.845 78.640 39.145 ;
        RECT 79.170 39.115 79.490 40.075 ;
        RECT 76.395 38.445 76.730 38.615 ;
        RECT 76.925 38.445 77.600 38.615 ;
        RECT 77.920 38.165 78.290 38.665 ;
        RECT 78.470 38.615 78.640 38.845 ;
        RECT 79.025 38.785 79.490 39.115 ;
        RECT 79.660 39.405 79.830 40.245 ;
        RECT 80.010 40.215 80.325 40.715 ;
        RECT 80.555 39.985 80.895 40.545 ;
        RECT 80.000 39.610 80.895 39.985 ;
        RECT 81.065 39.705 81.235 40.715 ;
        RECT 80.705 39.405 80.895 39.610 ;
        RECT 81.405 39.655 81.735 40.500 ;
        RECT 81.405 39.575 81.795 39.655 ;
        RECT 81.580 39.525 81.795 39.575 ;
        RECT 79.660 39.075 80.535 39.405 ;
        RECT 80.705 39.075 81.455 39.405 ;
        RECT 79.660 38.615 79.830 39.075 ;
        RECT 80.705 38.905 80.905 39.075 ;
        RECT 81.625 38.945 81.795 39.525 ;
        RECT 81.965 39.625 83.175 40.715 ;
        RECT 81.965 39.085 82.485 39.625 ;
        RECT 81.570 38.905 81.795 38.945 ;
        RECT 82.655 38.915 83.175 39.455 ;
        RECT 78.470 38.445 78.875 38.615 ;
        RECT 79.045 38.445 79.830 38.615 ;
        RECT 80.105 38.165 80.315 38.695 ;
        RECT 80.575 38.380 80.905 38.905 ;
        RECT 81.415 38.820 81.795 38.905 ;
        RECT 81.075 38.165 81.245 38.775 ;
        RECT 81.415 38.385 81.745 38.820 ;
        RECT 81.965 38.165 83.175 38.915 ;
        RECT 5.520 37.995 83.260 38.165 ;
        RECT 5.605 37.245 6.815 37.995 ;
        RECT 5.605 36.705 6.125 37.245 ;
        RECT 6.995 37.185 7.265 37.995 ;
        RECT 7.435 37.185 7.765 37.825 ;
        RECT 7.935 37.185 8.175 37.995 ;
        RECT 8.455 37.445 8.625 37.735 ;
        RECT 8.795 37.615 9.125 37.995 ;
        RECT 8.455 37.275 9.120 37.445 ;
        RECT 6.295 36.535 6.815 37.075 ;
        RECT 6.985 36.755 7.335 37.005 ;
        RECT 7.505 36.585 7.675 37.185 ;
        RECT 7.845 36.755 8.195 37.005 ;
        RECT 5.605 35.445 6.815 36.535 ;
        RECT 6.995 35.445 7.325 36.585 ;
        RECT 7.505 36.415 8.185 36.585 ;
        RECT 8.370 36.455 8.720 37.105 ;
        RECT 7.855 35.630 8.185 36.415 ;
        RECT 8.890 36.285 9.120 37.275 ;
        RECT 8.455 36.115 9.120 36.285 ;
        RECT 8.455 35.615 8.625 36.115 ;
        RECT 8.795 35.445 9.125 35.945 ;
        RECT 9.295 35.615 9.480 37.735 ;
        RECT 9.735 37.535 9.985 37.995 ;
        RECT 10.155 37.545 10.490 37.715 ;
        RECT 10.685 37.545 11.360 37.715 ;
        RECT 10.155 37.405 10.325 37.545 ;
        RECT 9.650 36.415 9.930 37.365 ;
        RECT 10.100 37.275 10.325 37.405 ;
        RECT 10.100 36.170 10.270 37.275 ;
        RECT 10.495 37.125 11.020 37.345 ;
        RECT 10.440 36.360 10.680 36.955 ;
        RECT 10.850 36.425 11.020 37.125 ;
        RECT 11.190 36.765 11.360 37.545 ;
        RECT 11.680 37.495 12.050 37.995 ;
        RECT 12.230 37.545 12.635 37.715 ;
        RECT 12.805 37.545 13.590 37.715 ;
        RECT 12.230 37.315 12.400 37.545 ;
        RECT 11.570 37.015 12.400 37.315 ;
        RECT 12.785 37.045 13.250 37.375 ;
        RECT 11.570 36.985 11.770 37.015 ;
        RECT 11.890 36.765 12.060 36.835 ;
        RECT 11.190 36.595 12.060 36.765 ;
        RECT 11.550 36.505 12.060 36.595 ;
        RECT 10.100 36.040 10.405 36.170 ;
        RECT 10.850 36.060 11.380 36.425 ;
        RECT 9.720 35.445 9.985 35.905 ;
        RECT 10.155 35.615 10.405 36.040 ;
        RECT 11.550 35.890 11.720 36.505 ;
        RECT 10.615 35.720 11.720 35.890 ;
        RECT 11.890 35.445 12.060 36.245 ;
        RECT 12.230 35.945 12.400 37.015 ;
        RECT 12.570 36.115 12.760 36.835 ;
        RECT 12.930 36.085 13.250 37.045 ;
        RECT 13.420 37.085 13.590 37.545 ;
        RECT 13.865 37.465 14.075 37.995 ;
        RECT 14.335 37.255 14.665 37.780 ;
        RECT 14.835 37.385 15.005 37.995 ;
        RECT 15.175 37.340 15.505 37.775 ;
        RECT 15.725 37.345 15.985 37.825 ;
        RECT 16.155 37.455 16.405 37.995 ;
        RECT 15.175 37.255 15.555 37.340 ;
        RECT 14.465 37.085 14.665 37.255 ;
        RECT 15.330 37.215 15.555 37.255 ;
        RECT 13.420 36.755 14.295 37.085 ;
        RECT 14.465 36.755 15.215 37.085 ;
        RECT 12.230 35.615 12.480 35.945 ;
        RECT 13.420 35.915 13.590 36.755 ;
        RECT 14.465 36.550 14.655 36.755 ;
        RECT 15.385 36.635 15.555 37.215 ;
        RECT 15.340 36.585 15.555 36.635 ;
        RECT 13.760 36.175 14.655 36.550 ;
        RECT 15.165 36.505 15.555 36.585 ;
        RECT 12.705 35.745 13.590 35.915 ;
        RECT 13.770 35.445 14.085 35.945 ;
        RECT 14.315 35.615 14.655 36.175 ;
        RECT 14.825 35.445 14.995 36.455 ;
        RECT 15.165 35.660 15.495 36.505 ;
        RECT 15.725 36.315 15.895 37.345 ;
        RECT 16.575 37.290 16.795 37.775 ;
        RECT 16.065 36.695 16.295 37.090 ;
        RECT 16.465 36.865 16.795 37.290 ;
        RECT 16.965 37.615 17.855 37.785 ;
        RECT 16.965 36.890 17.135 37.615 ;
        RECT 17.305 37.060 17.855 37.445 ;
        RECT 18.690 37.215 19.190 37.825 ;
        RECT 16.965 36.820 17.855 36.890 ;
        RECT 16.960 36.795 17.855 36.820 ;
        RECT 16.950 36.780 17.855 36.795 ;
        RECT 16.945 36.765 17.855 36.780 ;
        RECT 16.935 36.760 17.855 36.765 ;
        RECT 16.930 36.750 17.855 36.760 ;
        RECT 18.485 36.755 18.835 37.005 ;
        RECT 16.925 36.740 17.855 36.750 ;
        RECT 16.915 36.735 17.855 36.740 ;
        RECT 16.905 36.725 17.855 36.735 ;
        RECT 16.895 36.720 17.855 36.725 ;
        RECT 16.895 36.715 17.230 36.720 ;
        RECT 16.880 36.710 17.230 36.715 ;
        RECT 16.865 36.700 17.230 36.710 ;
        RECT 16.840 36.695 17.230 36.700 ;
        RECT 16.065 36.690 17.230 36.695 ;
        RECT 16.065 36.655 17.200 36.690 ;
        RECT 16.065 36.630 17.165 36.655 ;
        RECT 16.065 36.600 17.135 36.630 ;
        RECT 16.065 36.570 17.115 36.600 ;
        RECT 16.065 36.540 17.095 36.570 ;
        RECT 16.065 36.530 17.025 36.540 ;
        RECT 16.065 36.520 17.000 36.530 ;
        RECT 16.065 36.505 16.980 36.520 ;
        RECT 16.065 36.490 16.960 36.505 ;
        RECT 16.170 36.480 16.955 36.490 ;
        RECT 16.170 36.445 16.940 36.480 ;
        RECT 15.725 35.615 16.000 36.315 ;
        RECT 16.170 36.195 16.925 36.445 ;
        RECT 17.095 36.125 17.425 36.370 ;
        RECT 17.595 36.270 17.855 36.720 ;
        RECT 19.020 36.585 19.190 37.215 ;
        RECT 19.820 37.345 20.150 37.825 ;
        RECT 20.320 37.535 20.545 37.995 ;
        RECT 20.715 37.345 21.045 37.825 ;
        RECT 19.820 37.175 21.045 37.345 ;
        RECT 21.235 37.195 21.485 37.995 ;
        RECT 21.655 37.195 21.995 37.825 ;
        RECT 22.170 37.505 22.425 37.995 ;
        RECT 22.595 37.485 23.825 37.825 ;
        RECT 19.360 36.805 19.690 37.005 ;
        RECT 19.860 36.805 20.190 37.005 ;
        RECT 20.360 36.805 20.780 37.005 ;
        RECT 20.955 36.835 21.650 37.005 ;
        RECT 20.955 36.585 21.125 36.835 ;
        RECT 21.820 36.585 21.995 37.195 ;
        RECT 22.190 36.755 22.410 37.335 ;
        RECT 22.595 36.585 22.775 37.485 ;
        RECT 22.945 36.755 23.320 37.315 ;
        RECT 23.495 37.255 23.825 37.485 ;
        RECT 24.095 37.445 24.265 37.735 ;
        RECT 24.435 37.615 24.765 37.995 ;
        RECT 24.095 37.275 24.760 37.445 ;
        RECT 23.525 36.755 23.835 37.085 ;
        RECT 18.690 36.415 21.125 36.585 ;
        RECT 17.240 36.100 17.425 36.125 ;
        RECT 17.240 36.000 17.855 36.100 ;
        RECT 16.170 35.445 16.425 35.990 ;
        RECT 16.595 35.615 17.075 35.955 ;
        RECT 17.250 35.445 17.855 36.000 ;
        RECT 18.690 35.615 19.020 36.415 ;
        RECT 19.190 35.445 19.520 36.245 ;
        RECT 19.820 35.615 20.150 36.415 ;
        RECT 20.795 35.445 21.045 36.245 ;
        RECT 21.315 35.445 21.485 36.585 ;
        RECT 21.655 35.615 21.995 36.585 ;
        RECT 22.170 35.445 22.425 36.585 ;
        RECT 22.595 36.415 23.825 36.585 ;
        RECT 24.010 36.455 24.360 37.105 ;
        RECT 22.595 35.615 22.925 36.415 ;
        RECT 23.095 35.445 23.325 36.245 ;
        RECT 23.495 35.615 23.825 36.415 ;
        RECT 24.530 36.285 24.760 37.275 ;
        RECT 24.095 36.115 24.760 36.285 ;
        RECT 24.095 35.615 24.265 36.115 ;
        RECT 24.435 35.445 24.765 35.945 ;
        RECT 24.935 35.615 25.120 37.735 ;
        RECT 25.375 37.535 25.625 37.995 ;
        RECT 25.795 37.545 26.130 37.715 ;
        RECT 26.325 37.545 27.000 37.715 ;
        RECT 25.795 37.405 25.965 37.545 ;
        RECT 25.290 36.415 25.570 37.365 ;
        RECT 25.740 37.275 25.965 37.405 ;
        RECT 25.740 36.170 25.910 37.275 ;
        RECT 26.135 37.125 26.660 37.345 ;
        RECT 26.080 36.360 26.320 36.955 ;
        RECT 26.490 36.425 26.660 37.125 ;
        RECT 26.830 36.765 27.000 37.545 ;
        RECT 27.320 37.495 27.690 37.995 ;
        RECT 27.870 37.545 28.275 37.715 ;
        RECT 28.445 37.545 29.230 37.715 ;
        RECT 27.870 37.315 28.040 37.545 ;
        RECT 27.210 37.015 28.040 37.315 ;
        RECT 28.425 37.045 28.890 37.375 ;
        RECT 27.210 36.985 27.410 37.015 ;
        RECT 27.530 36.765 27.700 36.835 ;
        RECT 26.830 36.595 27.700 36.765 ;
        RECT 27.190 36.505 27.700 36.595 ;
        RECT 25.740 36.040 26.045 36.170 ;
        RECT 26.490 36.060 27.020 36.425 ;
        RECT 25.360 35.445 25.625 35.905 ;
        RECT 25.795 35.615 26.045 36.040 ;
        RECT 27.190 35.890 27.360 36.505 ;
        RECT 26.255 35.720 27.360 35.890 ;
        RECT 27.530 35.445 27.700 36.245 ;
        RECT 27.870 35.945 28.040 37.015 ;
        RECT 28.210 36.115 28.400 36.835 ;
        RECT 28.570 36.085 28.890 37.045 ;
        RECT 29.060 37.085 29.230 37.545 ;
        RECT 29.505 37.465 29.715 37.995 ;
        RECT 29.975 37.255 30.305 37.780 ;
        RECT 30.475 37.385 30.645 37.995 ;
        RECT 30.815 37.340 31.145 37.775 ;
        RECT 30.815 37.255 31.195 37.340 ;
        RECT 31.365 37.270 31.655 37.995 ;
        RECT 31.915 37.445 32.085 37.735 ;
        RECT 32.255 37.615 32.585 37.995 ;
        RECT 31.915 37.275 32.580 37.445 ;
        RECT 30.105 37.085 30.305 37.255 ;
        RECT 30.970 37.215 31.195 37.255 ;
        RECT 29.060 36.755 29.935 37.085 ;
        RECT 30.105 36.755 30.855 37.085 ;
        RECT 27.870 35.615 28.120 35.945 ;
        RECT 29.060 35.915 29.230 36.755 ;
        RECT 30.105 36.550 30.295 36.755 ;
        RECT 31.025 36.635 31.195 37.215 ;
        RECT 30.980 36.585 31.195 36.635 ;
        RECT 29.400 36.175 30.295 36.550 ;
        RECT 30.805 36.505 31.195 36.585 ;
        RECT 28.345 35.745 29.230 35.915 ;
        RECT 29.410 35.445 29.725 35.945 ;
        RECT 29.955 35.615 30.295 36.175 ;
        RECT 30.465 35.445 30.635 36.455 ;
        RECT 30.805 35.660 31.135 36.505 ;
        RECT 31.365 35.445 31.655 36.610 ;
        RECT 31.830 36.455 32.180 37.105 ;
        RECT 32.350 36.285 32.580 37.275 ;
        RECT 31.915 36.115 32.580 36.285 ;
        RECT 31.915 35.615 32.085 36.115 ;
        RECT 32.255 35.445 32.585 35.945 ;
        RECT 32.755 35.615 32.940 37.735 ;
        RECT 33.195 37.535 33.445 37.995 ;
        RECT 33.615 37.545 33.950 37.715 ;
        RECT 34.145 37.545 34.820 37.715 ;
        RECT 33.615 37.405 33.785 37.545 ;
        RECT 33.110 36.415 33.390 37.365 ;
        RECT 33.560 37.275 33.785 37.405 ;
        RECT 33.560 36.170 33.730 37.275 ;
        RECT 33.955 37.125 34.480 37.345 ;
        RECT 33.900 36.360 34.140 36.955 ;
        RECT 34.310 36.425 34.480 37.125 ;
        RECT 34.650 36.765 34.820 37.545 ;
        RECT 35.140 37.495 35.510 37.995 ;
        RECT 35.690 37.545 36.095 37.715 ;
        RECT 36.265 37.545 37.050 37.715 ;
        RECT 35.690 37.315 35.860 37.545 ;
        RECT 35.030 37.015 35.860 37.315 ;
        RECT 36.245 37.045 36.710 37.375 ;
        RECT 35.030 36.985 35.230 37.015 ;
        RECT 35.350 36.765 35.520 36.835 ;
        RECT 34.650 36.595 35.520 36.765 ;
        RECT 35.010 36.505 35.520 36.595 ;
        RECT 33.560 36.040 33.865 36.170 ;
        RECT 34.310 36.060 34.840 36.425 ;
        RECT 33.180 35.445 33.445 35.905 ;
        RECT 33.615 35.615 33.865 36.040 ;
        RECT 35.010 35.890 35.180 36.505 ;
        RECT 34.075 35.720 35.180 35.890 ;
        RECT 35.350 35.445 35.520 36.245 ;
        RECT 35.690 35.945 35.860 37.015 ;
        RECT 36.030 36.115 36.220 36.835 ;
        RECT 36.390 36.085 36.710 37.045 ;
        RECT 36.880 37.085 37.050 37.545 ;
        RECT 37.325 37.465 37.535 37.995 ;
        RECT 37.795 37.255 38.125 37.780 ;
        RECT 38.295 37.385 38.465 37.995 ;
        RECT 38.635 37.340 38.965 37.775 ;
        RECT 39.190 37.465 39.480 37.815 ;
        RECT 39.675 37.635 40.005 37.995 ;
        RECT 40.175 37.465 40.405 37.770 ;
        RECT 38.635 37.255 39.015 37.340 ;
        RECT 39.190 37.295 40.405 37.465 ;
        RECT 40.595 37.655 40.765 37.690 ;
        RECT 40.595 37.485 40.795 37.655 ;
        RECT 37.925 37.085 38.125 37.255 ;
        RECT 38.790 37.215 39.015 37.255 ;
        RECT 36.880 36.755 37.755 37.085 ;
        RECT 37.925 36.755 38.675 37.085 ;
        RECT 35.690 35.615 35.940 35.945 ;
        RECT 36.880 35.915 37.050 36.755 ;
        RECT 37.925 36.550 38.115 36.755 ;
        RECT 38.845 36.635 39.015 37.215 ;
        RECT 40.595 37.125 40.765 37.485 ;
        RECT 39.250 36.975 39.510 37.085 ;
        RECT 39.245 36.805 39.510 36.975 ;
        RECT 39.250 36.755 39.510 36.805 ;
        RECT 39.690 36.755 40.075 37.085 ;
        RECT 40.245 36.955 40.765 37.125 ;
        RECT 41.025 37.255 41.490 37.800 ;
        RECT 38.800 36.585 39.015 36.635 ;
        RECT 37.220 36.175 38.115 36.550 ;
        RECT 38.625 36.505 39.015 36.585 ;
        RECT 36.165 35.745 37.050 35.915 ;
        RECT 37.230 35.445 37.545 35.945 ;
        RECT 37.775 35.615 38.115 36.175 ;
        RECT 38.285 35.445 38.455 36.455 ;
        RECT 38.625 35.660 38.955 36.505 ;
        RECT 39.190 35.445 39.510 36.585 ;
        RECT 39.690 35.705 39.885 36.755 ;
        RECT 40.245 36.575 40.415 36.955 ;
        RECT 40.065 36.295 40.415 36.575 ;
        RECT 40.605 36.425 40.850 36.785 ;
        RECT 41.025 36.295 41.195 37.255 ;
        RECT 41.995 37.175 42.165 37.995 ;
        RECT 42.335 37.345 42.665 37.825 ;
        RECT 42.835 37.605 43.185 37.995 ;
        RECT 43.355 37.425 43.585 37.825 ;
        RECT 43.075 37.345 43.585 37.425 ;
        RECT 42.335 37.255 43.585 37.345 ;
        RECT 43.755 37.255 44.075 37.735 ;
        RECT 45.255 37.445 45.425 37.735 ;
        RECT 45.595 37.615 45.925 37.995 ;
        RECT 45.255 37.275 45.920 37.445 ;
        RECT 42.335 37.175 43.245 37.255 ;
        RECT 41.365 36.635 41.610 37.085 ;
        RECT 41.870 36.805 42.565 37.005 ;
        RECT 42.735 36.835 43.335 37.005 ;
        RECT 42.735 36.635 42.905 36.835 ;
        RECT 43.565 36.665 43.735 37.085 ;
        RECT 41.365 36.465 42.905 36.635 ;
        RECT 43.075 36.495 43.735 36.665 ;
        RECT 43.075 36.295 43.245 36.495 ;
        RECT 43.905 36.325 44.075 37.255 ;
        RECT 45.170 36.455 45.520 37.105 ;
        RECT 40.065 35.615 40.395 36.295 ;
        RECT 40.595 35.445 40.850 36.245 ;
        RECT 41.025 36.125 43.245 36.295 ;
        RECT 43.415 36.125 44.075 36.325 ;
        RECT 45.690 36.285 45.920 37.275 ;
        RECT 41.025 35.445 41.325 35.955 ;
        RECT 41.495 35.615 41.825 36.125 ;
        RECT 43.415 35.955 43.585 36.125 ;
        RECT 45.255 36.115 45.920 36.285 ;
        RECT 41.995 35.445 42.625 35.955 ;
        RECT 43.205 35.785 43.585 35.955 ;
        RECT 43.755 35.445 44.055 35.955 ;
        RECT 45.255 35.615 45.425 36.115 ;
        RECT 45.595 35.445 45.925 35.945 ;
        RECT 46.095 35.615 46.280 37.735 ;
        RECT 46.535 37.535 46.785 37.995 ;
        RECT 46.955 37.545 47.290 37.715 ;
        RECT 47.485 37.545 48.160 37.715 ;
        RECT 46.955 37.405 47.125 37.545 ;
        RECT 46.450 36.415 46.730 37.365 ;
        RECT 46.900 37.275 47.125 37.405 ;
        RECT 46.900 36.170 47.070 37.275 ;
        RECT 47.295 37.125 47.820 37.345 ;
        RECT 47.240 36.360 47.480 36.955 ;
        RECT 47.650 36.425 47.820 37.125 ;
        RECT 47.990 36.765 48.160 37.545 ;
        RECT 48.480 37.495 48.850 37.995 ;
        RECT 49.030 37.545 49.435 37.715 ;
        RECT 49.605 37.545 50.390 37.715 ;
        RECT 49.030 37.315 49.200 37.545 ;
        RECT 48.370 37.015 49.200 37.315 ;
        RECT 49.585 37.045 50.050 37.375 ;
        RECT 48.370 36.985 48.570 37.015 ;
        RECT 48.690 36.765 48.860 36.835 ;
        RECT 47.990 36.595 48.860 36.765 ;
        RECT 48.350 36.505 48.860 36.595 ;
        RECT 46.900 36.040 47.205 36.170 ;
        RECT 47.650 36.060 48.180 36.425 ;
        RECT 46.520 35.445 46.785 35.905 ;
        RECT 46.955 35.615 47.205 36.040 ;
        RECT 48.350 35.890 48.520 36.505 ;
        RECT 47.415 35.720 48.520 35.890 ;
        RECT 48.690 35.445 48.860 36.245 ;
        RECT 49.030 35.945 49.200 37.015 ;
        RECT 49.370 36.115 49.560 36.835 ;
        RECT 49.730 36.085 50.050 37.045 ;
        RECT 50.220 37.085 50.390 37.545 ;
        RECT 50.665 37.465 50.875 37.995 ;
        RECT 51.135 37.255 51.465 37.780 ;
        RECT 51.635 37.385 51.805 37.995 ;
        RECT 51.975 37.340 52.305 37.775 ;
        RECT 51.975 37.255 52.355 37.340 ;
        RECT 51.265 37.085 51.465 37.255 ;
        RECT 52.130 37.215 52.355 37.255 ;
        RECT 50.220 36.755 51.095 37.085 ;
        RECT 51.265 36.755 52.015 37.085 ;
        RECT 49.030 35.615 49.280 35.945 ;
        RECT 50.220 35.915 50.390 36.755 ;
        RECT 51.265 36.550 51.455 36.755 ;
        RECT 52.185 36.635 52.355 37.215 ;
        RECT 52.140 36.585 52.355 36.635 ;
        RECT 50.560 36.175 51.455 36.550 ;
        RECT 51.965 36.505 52.355 36.585 ;
        RECT 52.525 37.255 52.910 37.825 ;
        RECT 53.080 37.535 53.405 37.995 ;
        RECT 53.925 37.365 54.205 37.825 ;
        RECT 52.525 36.585 52.805 37.255 ;
        RECT 53.080 37.195 54.205 37.365 ;
        RECT 53.080 37.085 53.530 37.195 ;
        RECT 52.975 36.755 53.530 37.085 ;
        RECT 54.395 37.025 54.795 37.825 ;
        RECT 55.195 37.535 55.465 37.995 ;
        RECT 55.635 37.365 55.920 37.825 ;
        RECT 49.505 35.745 50.390 35.915 ;
        RECT 50.570 35.445 50.885 35.945 ;
        RECT 51.115 35.615 51.455 36.175 ;
        RECT 51.625 35.445 51.795 36.455 ;
        RECT 51.965 35.660 52.295 36.505 ;
        RECT 52.525 35.615 52.910 36.585 ;
        RECT 53.080 36.295 53.530 36.755 ;
        RECT 53.700 36.465 54.795 37.025 ;
        RECT 53.080 36.075 54.205 36.295 ;
        RECT 53.080 35.445 53.405 35.905 ;
        RECT 53.925 35.615 54.205 36.075 ;
        RECT 54.395 35.615 54.795 36.465 ;
        RECT 54.965 37.195 55.920 37.365 ;
        RECT 57.125 37.270 57.415 37.995 ;
        RECT 57.675 37.445 57.845 37.735 ;
        RECT 58.015 37.615 58.345 37.995 ;
        RECT 57.675 37.275 58.340 37.445 ;
        RECT 54.965 36.295 55.175 37.195 ;
        RECT 55.345 36.465 56.035 37.025 ;
        RECT 54.965 36.075 55.920 36.295 ;
        RECT 55.195 35.445 55.465 35.905 ;
        RECT 55.635 35.615 55.920 36.075 ;
        RECT 57.125 35.445 57.415 36.610 ;
        RECT 57.590 36.455 57.940 37.105 ;
        RECT 58.110 36.285 58.340 37.275 ;
        RECT 57.675 36.115 58.340 36.285 ;
        RECT 57.675 35.615 57.845 36.115 ;
        RECT 58.015 35.445 58.345 35.945 ;
        RECT 58.515 35.615 58.700 37.735 ;
        RECT 58.955 37.535 59.205 37.995 ;
        RECT 59.375 37.545 59.710 37.715 ;
        RECT 59.905 37.545 60.580 37.715 ;
        RECT 59.375 37.405 59.545 37.545 ;
        RECT 58.870 36.415 59.150 37.365 ;
        RECT 59.320 37.275 59.545 37.405 ;
        RECT 59.320 36.170 59.490 37.275 ;
        RECT 59.715 37.125 60.240 37.345 ;
        RECT 59.660 36.360 59.900 36.955 ;
        RECT 60.070 36.425 60.240 37.125 ;
        RECT 60.410 36.765 60.580 37.545 ;
        RECT 60.900 37.495 61.270 37.995 ;
        RECT 61.450 37.545 61.855 37.715 ;
        RECT 62.025 37.545 62.810 37.715 ;
        RECT 61.450 37.315 61.620 37.545 ;
        RECT 60.790 37.015 61.620 37.315 ;
        RECT 62.005 37.045 62.470 37.375 ;
        RECT 60.790 36.985 60.990 37.015 ;
        RECT 61.110 36.765 61.280 36.835 ;
        RECT 60.410 36.595 61.280 36.765 ;
        RECT 60.770 36.505 61.280 36.595 ;
        RECT 59.320 36.040 59.625 36.170 ;
        RECT 60.070 36.060 60.600 36.425 ;
        RECT 58.940 35.445 59.205 35.905 ;
        RECT 59.375 35.615 59.625 36.040 ;
        RECT 60.770 35.890 60.940 36.505 ;
        RECT 59.835 35.720 60.940 35.890 ;
        RECT 61.110 35.445 61.280 36.245 ;
        RECT 61.450 35.945 61.620 37.015 ;
        RECT 61.790 36.115 61.980 36.835 ;
        RECT 62.150 36.085 62.470 37.045 ;
        RECT 62.640 37.085 62.810 37.545 ;
        RECT 63.085 37.465 63.295 37.995 ;
        RECT 63.555 37.255 63.885 37.780 ;
        RECT 64.055 37.385 64.225 37.995 ;
        RECT 64.395 37.340 64.725 37.775 ;
        RECT 64.895 37.480 65.065 37.995 ;
        RECT 65.495 37.445 65.665 37.735 ;
        RECT 65.835 37.615 66.165 37.995 ;
        RECT 64.395 37.255 64.775 37.340 ;
        RECT 65.495 37.275 66.160 37.445 ;
        RECT 63.685 37.085 63.885 37.255 ;
        RECT 64.550 37.215 64.775 37.255 ;
        RECT 62.640 36.755 63.515 37.085 ;
        RECT 63.685 36.755 64.435 37.085 ;
        RECT 61.450 35.615 61.700 35.945 ;
        RECT 62.640 35.915 62.810 36.755 ;
        RECT 63.685 36.550 63.875 36.755 ;
        RECT 64.605 36.635 64.775 37.215 ;
        RECT 64.560 36.585 64.775 36.635 ;
        RECT 62.980 36.175 63.875 36.550 ;
        RECT 64.385 36.505 64.775 36.585 ;
        RECT 61.925 35.745 62.810 35.915 ;
        RECT 62.990 35.445 63.305 35.945 ;
        RECT 63.535 35.615 63.875 36.175 ;
        RECT 64.045 35.445 64.215 36.455 ;
        RECT 64.385 35.660 64.715 36.505 ;
        RECT 65.410 36.455 65.760 37.105 ;
        RECT 64.885 35.445 65.055 36.360 ;
        RECT 65.930 36.285 66.160 37.275 ;
        RECT 65.495 36.115 66.160 36.285 ;
        RECT 65.495 35.615 65.665 36.115 ;
        RECT 65.835 35.445 66.165 35.945 ;
        RECT 66.335 35.615 66.520 37.735 ;
        RECT 66.775 37.535 67.025 37.995 ;
        RECT 67.195 37.545 67.530 37.715 ;
        RECT 67.725 37.545 68.400 37.715 ;
        RECT 67.195 37.405 67.365 37.545 ;
        RECT 66.690 36.415 66.970 37.365 ;
        RECT 67.140 37.275 67.365 37.405 ;
        RECT 67.140 36.170 67.310 37.275 ;
        RECT 67.535 37.125 68.060 37.345 ;
        RECT 67.480 36.360 67.720 36.955 ;
        RECT 67.890 36.425 68.060 37.125 ;
        RECT 68.230 36.765 68.400 37.545 ;
        RECT 68.720 37.495 69.090 37.995 ;
        RECT 69.270 37.545 69.675 37.715 ;
        RECT 69.845 37.545 70.630 37.715 ;
        RECT 69.270 37.315 69.440 37.545 ;
        RECT 68.610 37.015 69.440 37.315 ;
        RECT 69.825 37.045 70.290 37.375 ;
        RECT 68.610 36.985 68.810 37.015 ;
        RECT 68.930 36.765 69.100 36.835 ;
        RECT 68.230 36.595 69.100 36.765 ;
        RECT 68.590 36.505 69.100 36.595 ;
        RECT 67.140 36.040 67.445 36.170 ;
        RECT 67.890 36.060 68.420 36.425 ;
        RECT 66.760 35.445 67.025 35.905 ;
        RECT 67.195 35.615 67.445 36.040 ;
        RECT 68.590 35.890 68.760 36.505 ;
        RECT 67.655 35.720 68.760 35.890 ;
        RECT 68.930 35.445 69.100 36.245 ;
        RECT 69.270 35.945 69.440 37.015 ;
        RECT 69.610 36.115 69.800 36.835 ;
        RECT 69.970 36.085 70.290 37.045 ;
        RECT 70.460 37.085 70.630 37.545 ;
        RECT 70.905 37.465 71.115 37.995 ;
        RECT 71.375 37.255 71.705 37.780 ;
        RECT 71.875 37.385 72.045 37.995 ;
        RECT 72.215 37.340 72.545 37.775 ;
        RECT 72.815 37.340 73.145 37.775 ;
        RECT 73.315 37.385 73.485 37.995 ;
        RECT 72.215 37.255 72.595 37.340 ;
        RECT 71.505 37.085 71.705 37.255 ;
        RECT 72.370 37.215 72.595 37.255 ;
        RECT 70.460 36.755 71.335 37.085 ;
        RECT 71.505 36.755 72.255 37.085 ;
        RECT 69.270 35.615 69.520 35.945 ;
        RECT 70.460 35.915 70.630 36.755 ;
        RECT 71.505 36.550 71.695 36.755 ;
        RECT 72.425 36.635 72.595 37.215 ;
        RECT 72.380 36.585 72.595 36.635 ;
        RECT 70.800 36.175 71.695 36.550 ;
        RECT 72.205 36.505 72.595 36.585 ;
        RECT 72.765 37.255 73.145 37.340 ;
        RECT 73.655 37.255 73.985 37.780 ;
        RECT 74.245 37.465 74.455 37.995 ;
        RECT 74.730 37.545 75.515 37.715 ;
        RECT 75.685 37.545 76.090 37.715 ;
        RECT 72.765 37.215 72.990 37.255 ;
        RECT 72.765 36.635 72.935 37.215 ;
        RECT 73.655 37.085 73.855 37.255 ;
        RECT 74.730 37.085 74.900 37.545 ;
        RECT 73.105 36.755 73.855 37.085 ;
        RECT 74.025 36.755 74.900 37.085 ;
        RECT 72.765 36.585 72.980 36.635 ;
        RECT 72.765 36.505 73.155 36.585 ;
        RECT 69.745 35.745 70.630 35.915 ;
        RECT 70.810 35.445 71.125 35.945 ;
        RECT 71.355 35.615 71.695 36.175 ;
        RECT 71.865 35.445 72.035 36.455 ;
        RECT 72.205 35.660 72.535 36.505 ;
        RECT 72.825 35.660 73.155 36.505 ;
        RECT 73.665 36.550 73.855 36.755 ;
        RECT 73.325 35.445 73.495 36.455 ;
        RECT 73.665 36.175 74.560 36.550 ;
        RECT 73.665 35.615 74.005 36.175 ;
        RECT 74.235 35.445 74.550 35.945 ;
        RECT 74.730 35.915 74.900 36.755 ;
        RECT 75.070 37.045 75.535 37.375 ;
        RECT 75.920 37.315 76.090 37.545 ;
        RECT 76.270 37.495 76.640 37.995 ;
        RECT 76.960 37.545 77.635 37.715 ;
        RECT 77.830 37.545 78.165 37.715 ;
        RECT 75.070 36.085 75.390 37.045 ;
        RECT 75.920 37.015 76.750 37.315 ;
        RECT 75.560 36.115 75.750 36.835 ;
        RECT 75.920 35.945 76.090 37.015 ;
        RECT 76.550 36.985 76.750 37.015 ;
        RECT 76.260 36.765 76.430 36.835 ;
        RECT 76.960 36.765 77.130 37.545 ;
        RECT 77.995 37.405 78.165 37.545 ;
        RECT 78.335 37.535 78.585 37.995 ;
        RECT 76.260 36.595 77.130 36.765 ;
        RECT 77.300 37.125 77.825 37.345 ;
        RECT 77.995 37.275 78.220 37.405 ;
        RECT 76.260 36.505 76.770 36.595 ;
        RECT 74.730 35.745 75.615 35.915 ;
        RECT 75.840 35.615 76.090 35.945 ;
        RECT 76.260 35.445 76.430 36.245 ;
        RECT 76.600 35.890 76.770 36.505 ;
        RECT 77.300 36.425 77.470 37.125 ;
        RECT 76.940 36.060 77.470 36.425 ;
        RECT 77.640 36.360 77.880 36.955 ;
        RECT 78.050 36.170 78.220 37.275 ;
        RECT 78.390 36.415 78.670 37.365 ;
        RECT 77.915 36.040 78.220 36.170 ;
        RECT 76.600 35.720 77.705 35.890 ;
        RECT 77.915 35.615 78.165 36.040 ;
        RECT 78.335 35.445 78.600 35.905 ;
        RECT 78.840 35.615 79.025 37.735 ;
        RECT 79.195 37.615 79.525 37.995 ;
        RECT 79.695 37.445 79.865 37.735 ;
        RECT 79.200 37.275 79.865 37.445 ;
        RECT 80.215 37.445 80.385 37.825 ;
        RECT 80.600 37.615 80.930 37.995 ;
        RECT 80.215 37.275 80.930 37.445 ;
        RECT 79.200 36.285 79.430 37.275 ;
        RECT 79.600 36.455 79.950 37.105 ;
        RECT 80.125 36.725 80.480 37.095 ;
        RECT 80.760 37.085 80.930 37.275 ;
        RECT 81.100 37.250 81.355 37.825 ;
        RECT 80.760 36.755 81.015 37.085 ;
        RECT 80.760 36.545 80.930 36.755 ;
        RECT 80.215 36.375 80.930 36.545 ;
        RECT 81.185 36.520 81.355 37.250 ;
        RECT 81.530 37.155 81.790 37.995 ;
        RECT 81.965 37.245 83.175 37.995 ;
        RECT 79.200 36.115 79.865 36.285 ;
        RECT 79.195 35.445 79.525 35.945 ;
        RECT 79.695 35.615 79.865 36.115 ;
        RECT 80.215 35.615 80.385 36.375 ;
        RECT 80.600 35.445 80.930 36.205 ;
        RECT 81.100 35.615 81.355 36.520 ;
        RECT 81.530 35.445 81.790 36.595 ;
        RECT 81.965 36.535 82.485 37.075 ;
        RECT 82.655 36.705 83.175 37.245 ;
        RECT 81.965 35.445 83.175 36.535 ;
        RECT 5.520 35.275 83.260 35.445 ;
        RECT 5.605 34.185 6.815 35.275 ;
        RECT 5.605 33.475 6.125 34.015 ;
        RECT 6.295 33.645 6.815 34.185 ;
        RECT 7.445 34.425 7.825 35.105 ;
        RECT 8.415 34.425 8.585 35.275 ;
        RECT 8.755 34.595 9.085 35.105 ;
        RECT 9.255 34.765 9.425 35.275 ;
        RECT 9.595 34.595 9.995 35.105 ;
        RECT 8.755 34.425 9.995 34.595 ;
        RECT 5.605 32.725 6.815 33.475 ;
        RECT 7.445 33.465 7.615 34.425 ;
        RECT 7.785 34.085 9.090 34.255 ;
        RECT 10.175 34.175 10.495 35.105 ;
        RECT 10.665 34.720 11.270 35.275 ;
        RECT 11.445 34.765 11.925 35.105 ;
        RECT 12.095 34.730 12.350 35.275 ;
        RECT 10.665 34.620 11.280 34.720 ;
        RECT 11.095 34.595 11.280 34.620 ;
        RECT 7.785 33.635 8.030 34.085 ;
        RECT 8.200 33.715 8.750 33.915 ;
        RECT 8.920 33.885 9.090 34.085 ;
        RECT 9.865 34.005 10.495 34.175 ;
        RECT 8.920 33.715 9.295 33.885 ;
        RECT 9.465 33.465 9.695 33.965 ;
        RECT 7.445 33.295 9.695 33.465 ;
        RECT 7.495 32.725 7.825 33.115 ;
        RECT 7.995 32.975 8.165 33.295 ;
        RECT 9.865 33.125 10.035 34.005 ;
        RECT 10.665 34.000 10.925 34.450 ;
        RECT 11.095 34.350 11.425 34.595 ;
        RECT 11.595 34.275 12.350 34.525 ;
        RECT 12.520 34.405 12.795 35.105 ;
        RECT 13.885 34.720 14.490 35.275 ;
        RECT 14.665 34.765 15.145 35.105 ;
        RECT 15.315 34.730 15.570 35.275 ;
        RECT 13.885 34.620 14.500 34.720 ;
        RECT 14.315 34.595 14.500 34.620 ;
        RECT 11.580 34.240 12.350 34.275 ;
        RECT 11.565 34.230 12.350 34.240 ;
        RECT 11.560 34.215 12.455 34.230 ;
        RECT 11.540 34.200 12.455 34.215 ;
        RECT 11.520 34.190 12.455 34.200 ;
        RECT 11.495 34.180 12.455 34.190 ;
        RECT 11.425 34.150 12.455 34.180 ;
        RECT 11.405 34.120 12.455 34.150 ;
        RECT 11.385 34.090 12.455 34.120 ;
        RECT 11.355 34.065 12.455 34.090 ;
        RECT 11.320 34.030 12.455 34.065 ;
        RECT 11.290 34.025 12.455 34.030 ;
        RECT 11.290 34.020 11.680 34.025 ;
        RECT 11.290 34.010 11.655 34.020 ;
        RECT 11.290 34.005 11.640 34.010 ;
        RECT 11.290 34.000 11.625 34.005 ;
        RECT 10.665 33.995 11.625 34.000 ;
        RECT 10.665 33.985 11.615 33.995 ;
        RECT 10.665 33.980 11.605 33.985 ;
        RECT 10.665 33.970 11.595 33.980 ;
        RECT 10.665 33.960 11.590 33.970 ;
        RECT 10.665 33.955 11.585 33.960 ;
        RECT 10.665 33.940 11.575 33.955 ;
        RECT 10.665 33.925 11.570 33.940 ;
        RECT 10.665 33.900 11.560 33.925 ;
        RECT 10.665 33.830 11.555 33.900 ;
        RECT 8.335 32.725 8.665 33.115 ;
        RECT 9.080 32.955 10.035 33.125 ;
        RECT 10.205 32.725 10.495 33.560 ;
        RECT 10.665 33.275 11.215 33.660 ;
        RECT 11.385 33.105 11.555 33.830 ;
        RECT 10.665 32.935 11.555 33.105 ;
        RECT 11.725 33.430 12.055 33.855 ;
        RECT 12.225 33.630 12.455 34.025 ;
        RECT 11.725 32.945 11.945 33.430 ;
        RECT 12.625 33.375 12.795 34.405 ;
        RECT 13.885 34.000 14.145 34.450 ;
        RECT 14.315 34.350 14.645 34.595 ;
        RECT 14.815 34.275 15.570 34.525 ;
        RECT 15.740 34.405 16.015 35.105 ;
        RECT 16.185 34.720 16.790 35.275 ;
        RECT 16.965 34.765 17.445 35.105 ;
        RECT 17.615 34.730 17.870 35.275 ;
        RECT 16.185 34.620 16.800 34.720 ;
        RECT 16.615 34.595 16.800 34.620 ;
        RECT 14.800 34.240 15.570 34.275 ;
        RECT 14.785 34.230 15.570 34.240 ;
        RECT 14.780 34.215 15.675 34.230 ;
        RECT 14.760 34.200 15.675 34.215 ;
        RECT 14.740 34.190 15.675 34.200 ;
        RECT 14.715 34.180 15.675 34.190 ;
        RECT 14.645 34.150 15.675 34.180 ;
        RECT 14.625 34.120 15.675 34.150 ;
        RECT 14.605 34.090 15.675 34.120 ;
        RECT 14.575 34.065 15.675 34.090 ;
        RECT 14.540 34.030 15.675 34.065 ;
        RECT 14.510 34.025 15.675 34.030 ;
        RECT 14.510 34.020 14.900 34.025 ;
        RECT 14.510 34.010 14.875 34.020 ;
        RECT 14.510 34.005 14.860 34.010 ;
        RECT 14.510 34.000 14.845 34.005 ;
        RECT 13.885 33.995 14.845 34.000 ;
        RECT 13.885 33.985 14.835 33.995 ;
        RECT 13.885 33.980 14.825 33.985 ;
        RECT 13.885 33.970 14.815 33.980 ;
        RECT 13.885 33.960 14.810 33.970 ;
        RECT 13.885 33.955 14.805 33.960 ;
        RECT 13.885 33.940 14.795 33.955 ;
        RECT 13.885 33.925 14.790 33.940 ;
        RECT 13.885 33.900 14.780 33.925 ;
        RECT 13.885 33.830 14.775 33.900 ;
        RECT 12.115 32.725 12.365 33.265 ;
        RECT 12.535 32.895 12.795 33.375 ;
        RECT 13.885 33.275 14.435 33.660 ;
        RECT 14.605 33.105 14.775 33.830 ;
        RECT 13.885 32.935 14.775 33.105 ;
        RECT 14.945 33.430 15.275 33.855 ;
        RECT 15.445 33.630 15.675 34.025 ;
        RECT 14.945 32.945 15.165 33.430 ;
        RECT 15.845 33.375 16.015 34.405 ;
        RECT 16.185 34.000 16.445 34.450 ;
        RECT 16.615 34.350 16.945 34.595 ;
        RECT 17.115 34.275 17.870 34.525 ;
        RECT 18.040 34.405 18.315 35.105 ;
        RECT 17.100 34.240 17.870 34.275 ;
        RECT 17.085 34.230 17.870 34.240 ;
        RECT 17.080 34.215 17.975 34.230 ;
        RECT 17.060 34.200 17.975 34.215 ;
        RECT 17.040 34.190 17.975 34.200 ;
        RECT 17.015 34.180 17.975 34.190 ;
        RECT 16.945 34.150 17.975 34.180 ;
        RECT 16.925 34.120 17.975 34.150 ;
        RECT 16.905 34.090 17.975 34.120 ;
        RECT 16.875 34.065 17.975 34.090 ;
        RECT 16.840 34.030 17.975 34.065 ;
        RECT 16.810 34.025 17.975 34.030 ;
        RECT 16.810 34.020 17.200 34.025 ;
        RECT 16.810 34.010 17.175 34.020 ;
        RECT 16.810 34.005 17.160 34.010 ;
        RECT 16.810 34.000 17.145 34.005 ;
        RECT 16.185 33.995 17.145 34.000 ;
        RECT 16.185 33.985 17.135 33.995 ;
        RECT 16.185 33.980 17.125 33.985 ;
        RECT 16.185 33.970 17.115 33.980 ;
        RECT 16.185 33.960 17.110 33.970 ;
        RECT 16.185 33.955 17.105 33.960 ;
        RECT 16.185 33.940 17.095 33.955 ;
        RECT 16.185 33.925 17.090 33.940 ;
        RECT 16.185 33.900 17.080 33.925 ;
        RECT 16.185 33.830 17.075 33.900 ;
        RECT 15.335 32.725 15.585 33.265 ;
        RECT 15.755 32.895 16.015 33.375 ;
        RECT 16.185 33.275 16.735 33.660 ;
        RECT 16.905 33.105 17.075 33.830 ;
        RECT 16.185 32.935 17.075 33.105 ;
        RECT 17.245 33.430 17.575 33.855 ;
        RECT 17.745 33.630 17.975 34.025 ;
        RECT 17.245 32.945 17.465 33.430 ;
        RECT 18.145 33.375 18.315 34.405 ;
        RECT 18.485 34.110 18.775 35.275 ;
        RECT 19.035 34.605 19.205 35.105 ;
        RECT 19.375 34.775 19.705 35.275 ;
        RECT 19.035 34.435 19.700 34.605 ;
        RECT 18.950 33.615 19.300 34.265 ;
        RECT 17.635 32.725 17.885 33.265 ;
        RECT 18.055 32.895 18.315 33.375 ;
        RECT 18.485 32.725 18.775 33.450 ;
        RECT 19.470 33.445 19.700 34.435 ;
        RECT 19.035 33.275 19.700 33.445 ;
        RECT 19.035 32.985 19.205 33.275 ;
        RECT 19.375 32.725 19.705 33.105 ;
        RECT 19.875 32.985 20.060 35.105 ;
        RECT 20.300 34.815 20.565 35.275 ;
        RECT 20.735 34.680 20.985 35.105 ;
        RECT 21.195 34.830 22.300 35.000 ;
        RECT 20.680 34.550 20.985 34.680 ;
        RECT 20.230 33.355 20.510 34.305 ;
        RECT 20.680 33.445 20.850 34.550 ;
        RECT 21.020 33.765 21.260 34.360 ;
        RECT 21.430 34.295 21.960 34.660 ;
        RECT 21.430 33.595 21.600 34.295 ;
        RECT 22.130 34.215 22.300 34.830 ;
        RECT 22.470 34.475 22.640 35.275 ;
        RECT 22.810 34.775 23.060 35.105 ;
        RECT 23.285 34.805 24.170 34.975 ;
        RECT 22.130 34.125 22.640 34.215 ;
        RECT 20.680 33.315 20.905 33.445 ;
        RECT 21.075 33.375 21.600 33.595 ;
        RECT 21.770 33.955 22.640 34.125 ;
        RECT 20.315 32.725 20.565 33.185 ;
        RECT 20.735 33.175 20.905 33.315 ;
        RECT 21.770 33.175 21.940 33.955 ;
        RECT 22.470 33.885 22.640 33.955 ;
        RECT 22.150 33.705 22.350 33.735 ;
        RECT 22.810 33.705 22.980 34.775 ;
        RECT 23.150 33.885 23.340 34.605 ;
        RECT 22.150 33.405 22.980 33.705 ;
        RECT 23.510 33.675 23.830 34.635 ;
        RECT 20.735 33.005 21.070 33.175 ;
        RECT 21.265 33.005 21.940 33.175 ;
        RECT 22.260 32.725 22.630 33.225 ;
        RECT 22.810 33.175 22.980 33.405 ;
        RECT 23.365 33.345 23.830 33.675 ;
        RECT 24.000 33.965 24.170 34.805 ;
        RECT 24.350 34.775 24.665 35.275 ;
        RECT 24.895 34.545 25.235 35.105 ;
        RECT 24.340 34.170 25.235 34.545 ;
        RECT 25.405 34.265 25.575 35.275 ;
        RECT 25.045 33.965 25.235 34.170 ;
        RECT 25.745 34.215 26.075 35.060 ;
        RECT 26.315 34.305 26.645 35.090 ;
        RECT 25.745 34.135 26.135 34.215 ;
        RECT 26.315 34.135 26.995 34.305 ;
        RECT 27.175 34.135 27.505 35.275 ;
        RECT 27.775 34.605 27.945 35.105 ;
        RECT 28.115 34.775 28.445 35.275 ;
        RECT 27.775 34.435 28.440 34.605 ;
        RECT 25.920 34.085 26.135 34.135 ;
        RECT 24.000 33.635 24.875 33.965 ;
        RECT 25.045 33.635 25.795 33.965 ;
        RECT 24.000 33.175 24.170 33.635 ;
        RECT 25.045 33.465 25.245 33.635 ;
        RECT 25.965 33.505 26.135 34.085 ;
        RECT 26.305 33.715 26.655 33.965 ;
        RECT 26.825 33.535 26.995 34.135 ;
        RECT 27.165 33.715 27.515 33.965 ;
        RECT 27.690 33.615 28.040 34.265 ;
        RECT 25.910 33.465 26.135 33.505 ;
        RECT 22.810 33.005 23.215 33.175 ;
        RECT 23.385 33.005 24.170 33.175 ;
        RECT 24.445 32.725 24.655 33.255 ;
        RECT 24.915 32.940 25.245 33.465 ;
        RECT 25.755 33.380 26.135 33.465 ;
        RECT 25.415 32.725 25.585 33.335 ;
        RECT 25.755 32.945 26.085 33.380 ;
        RECT 26.325 32.725 26.565 33.535 ;
        RECT 26.735 32.895 27.065 33.535 ;
        RECT 27.235 32.725 27.505 33.535 ;
        RECT 28.210 33.445 28.440 34.435 ;
        RECT 27.775 33.275 28.440 33.445 ;
        RECT 27.775 32.985 27.945 33.275 ;
        RECT 28.115 32.725 28.445 33.105 ;
        RECT 28.615 32.985 28.800 35.105 ;
        RECT 29.040 34.815 29.305 35.275 ;
        RECT 29.475 34.680 29.725 35.105 ;
        RECT 29.935 34.830 31.040 35.000 ;
        RECT 29.420 34.550 29.725 34.680 ;
        RECT 28.970 33.355 29.250 34.305 ;
        RECT 29.420 33.445 29.590 34.550 ;
        RECT 29.760 33.765 30.000 34.360 ;
        RECT 30.170 34.295 30.700 34.660 ;
        RECT 30.170 33.595 30.340 34.295 ;
        RECT 30.870 34.215 31.040 34.830 ;
        RECT 31.210 34.475 31.380 35.275 ;
        RECT 31.550 34.775 31.800 35.105 ;
        RECT 32.025 34.805 32.910 34.975 ;
        RECT 30.870 34.125 31.380 34.215 ;
        RECT 29.420 33.315 29.645 33.445 ;
        RECT 29.815 33.375 30.340 33.595 ;
        RECT 30.510 33.955 31.380 34.125 ;
        RECT 29.055 32.725 29.305 33.185 ;
        RECT 29.475 33.175 29.645 33.315 ;
        RECT 30.510 33.175 30.680 33.955 ;
        RECT 31.210 33.885 31.380 33.955 ;
        RECT 30.890 33.705 31.090 33.735 ;
        RECT 31.550 33.705 31.720 34.775 ;
        RECT 31.890 33.885 32.080 34.605 ;
        RECT 30.890 33.405 31.720 33.705 ;
        RECT 32.250 33.675 32.570 34.635 ;
        RECT 29.475 33.005 29.810 33.175 ;
        RECT 30.005 33.005 30.680 33.175 ;
        RECT 31.000 32.725 31.370 33.225 ;
        RECT 31.550 33.175 31.720 33.405 ;
        RECT 32.105 33.345 32.570 33.675 ;
        RECT 32.740 33.965 32.910 34.805 ;
        RECT 33.090 34.775 33.405 35.275 ;
        RECT 33.635 34.545 33.975 35.105 ;
        RECT 33.080 34.170 33.975 34.545 ;
        RECT 34.145 34.265 34.315 35.275 ;
        RECT 33.785 33.965 33.975 34.170 ;
        RECT 34.485 34.215 34.815 35.060 ;
        RECT 35.045 34.405 35.320 35.105 ;
        RECT 35.490 34.730 35.745 35.275 ;
        RECT 35.915 34.765 36.395 35.105 ;
        RECT 36.570 34.720 37.175 35.275 ;
        RECT 36.560 34.620 37.175 34.720 ;
        RECT 36.560 34.595 36.745 34.620 ;
        RECT 34.485 34.135 34.875 34.215 ;
        RECT 34.660 34.085 34.875 34.135 ;
        RECT 32.740 33.635 33.615 33.965 ;
        RECT 33.785 33.635 34.535 33.965 ;
        RECT 32.740 33.175 32.910 33.635 ;
        RECT 33.785 33.465 33.985 33.635 ;
        RECT 34.705 33.505 34.875 34.085 ;
        RECT 34.650 33.465 34.875 33.505 ;
        RECT 31.550 33.005 31.955 33.175 ;
        RECT 32.125 33.005 32.910 33.175 ;
        RECT 33.185 32.725 33.395 33.255 ;
        RECT 33.655 32.940 33.985 33.465 ;
        RECT 34.495 33.380 34.875 33.465 ;
        RECT 34.155 32.725 34.325 33.335 ;
        RECT 34.495 32.945 34.825 33.380 ;
        RECT 35.045 33.375 35.215 34.405 ;
        RECT 35.490 34.275 36.245 34.525 ;
        RECT 36.415 34.350 36.745 34.595 ;
        RECT 35.490 34.240 36.260 34.275 ;
        RECT 35.490 34.230 36.275 34.240 ;
        RECT 35.385 34.215 36.280 34.230 ;
        RECT 35.385 34.200 36.300 34.215 ;
        RECT 35.385 34.190 36.320 34.200 ;
        RECT 35.385 34.180 36.345 34.190 ;
        RECT 35.385 34.150 36.415 34.180 ;
        RECT 35.385 34.120 36.435 34.150 ;
        RECT 35.385 34.090 36.455 34.120 ;
        RECT 35.385 34.065 36.485 34.090 ;
        RECT 35.385 34.030 36.520 34.065 ;
        RECT 35.385 34.025 36.550 34.030 ;
        RECT 35.385 33.630 35.615 34.025 ;
        RECT 36.160 34.020 36.550 34.025 ;
        RECT 36.185 34.010 36.550 34.020 ;
        RECT 36.200 34.005 36.550 34.010 ;
        RECT 36.215 34.000 36.550 34.005 ;
        RECT 36.915 34.000 37.175 34.450 ;
        RECT 37.345 34.185 39.015 35.275 ;
        RECT 36.215 33.995 37.175 34.000 ;
        RECT 36.225 33.985 37.175 33.995 ;
        RECT 36.235 33.980 37.175 33.985 ;
        RECT 36.245 33.970 37.175 33.980 ;
        RECT 36.250 33.960 37.175 33.970 ;
        RECT 36.255 33.955 37.175 33.960 ;
        RECT 36.265 33.940 37.175 33.955 ;
        RECT 36.270 33.925 37.175 33.940 ;
        RECT 36.280 33.900 37.175 33.925 ;
        RECT 35.785 33.430 36.115 33.855 ;
        RECT 35.865 33.405 36.115 33.430 ;
        RECT 35.045 32.895 35.305 33.375 ;
        RECT 35.475 32.725 35.725 33.265 ;
        RECT 35.895 32.945 36.115 33.405 ;
        RECT 36.285 33.830 37.175 33.900 ;
        RECT 36.285 33.105 36.455 33.830 ;
        RECT 36.625 33.275 37.175 33.660 ;
        RECT 37.345 33.495 38.095 34.015 ;
        RECT 38.265 33.665 39.015 34.185 ;
        RECT 39.185 34.135 39.445 35.275 ;
        RECT 39.615 34.125 39.945 35.105 ;
        RECT 40.115 34.135 40.395 35.275 ;
        RECT 40.565 34.185 44.075 35.275 ;
        RECT 39.205 33.715 39.540 33.965 ;
        RECT 39.710 33.575 39.880 34.125 ;
        RECT 40.050 33.695 40.385 33.965 ;
        RECT 39.705 33.525 39.880 33.575 ;
        RECT 36.285 32.935 37.175 33.105 ;
        RECT 37.345 32.725 39.015 33.495 ;
        RECT 39.185 32.895 39.880 33.525 ;
        RECT 40.085 32.725 40.395 33.525 ;
        RECT 40.565 33.495 42.215 34.015 ;
        RECT 42.385 33.665 44.075 34.185 ;
        RECT 44.245 34.110 44.535 35.275 ;
        RECT 44.705 34.185 45.915 35.275 ;
        RECT 40.565 32.725 44.075 33.495 ;
        RECT 44.705 33.475 45.225 34.015 ;
        RECT 45.395 33.645 45.915 34.185 ;
        RECT 46.085 34.135 46.470 35.105 ;
        RECT 46.640 34.815 46.965 35.275 ;
        RECT 47.485 34.645 47.765 35.105 ;
        RECT 46.640 34.425 47.765 34.645 ;
        RECT 44.245 32.725 44.535 33.450 ;
        RECT 44.705 32.725 45.915 33.475 ;
        RECT 46.085 33.465 46.365 34.135 ;
        RECT 46.640 33.965 47.090 34.425 ;
        RECT 47.955 34.255 48.355 35.105 ;
        RECT 48.755 34.815 49.025 35.275 ;
        RECT 49.195 34.645 49.480 35.105 ;
        RECT 46.535 33.635 47.090 33.965 ;
        RECT 47.260 33.695 48.355 34.255 ;
        RECT 46.640 33.525 47.090 33.635 ;
        RECT 46.085 32.895 46.470 33.465 ;
        RECT 46.640 33.355 47.765 33.525 ;
        RECT 46.640 32.725 46.965 33.185 ;
        RECT 47.485 32.895 47.765 33.355 ;
        RECT 47.955 32.895 48.355 33.695 ;
        RECT 48.525 34.425 49.480 34.645 ;
        RECT 48.525 33.525 48.735 34.425 ;
        RECT 48.905 33.695 49.595 34.255 ;
        RECT 49.765 34.135 50.150 35.105 ;
        RECT 50.320 34.815 50.645 35.275 ;
        RECT 51.165 34.645 51.445 35.105 ;
        RECT 50.320 34.425 51.445 34.645 ;
        RECT 48.525 33.355 49.480 33.525 ;
        RECT 48.755 32.725 49.025 33.185 ;
        RECT 49.195 32.895 49.480 33.355 ;
        RECT 49.765 33.465 50.045 34.135 ;
        RECT 50.320 33.965 50.770 34.425 ;
        RECT 51.635 34.255 52.035 35.105 ;
        RECT 52.435 34.815 52.705 35.275 ;
        RECT 52.875 34.645 53.160 35.105 ;
        RECT 50.215 33.635 50.770 33.965 ;
        RECT 50.940 33.695 52.035 34.255 ;
        RECT 50.320 33.525 50.770 33.635 ;
        RECT 49.765 32.895 50.150 33.465 ;
        RECT 50.320 33.355 51.445 33.525 ;
        RECT 50.320 32.725 50.645 33.185 ;
        RECT 51.165 32.895 51.445 33.355 ;
        RECT 51.635 32.895 52.035 33.695 ;
        RECT 52.205 34.425 53.160 34.645 ;
        RECT 53.530 34.655 53.705 35.105 ;
        RECT 53.875 34.835 54.205 35.275 ;
        RECT 54.510 34.685 54.680 35.105 ;
        RECT 54.915 34.865 55.585 35.275 ;
        RECT 55.800 34.685 55.970 35.105 ;
        RECT 56.170 34.865 56.500 35.275 ;
        RECT 53.530 34.485 54.160 34.655 ;
        RECT 52.205 33.525 52.415 34.425 ;
        RECT 52.585 33.695 53.275 34.255 ;
        RECT 53.445 33.635 53.810 34.315 ;
        RECT 53.990 33.965 54.160 34.485 ;
        RECT 54.510 34.515 56.525 34.685 ;
        RECT 53.990 33.635 54.340 33.965 ;
        RECT 52.205 33.355 53.160 33.525 ;
        RECT 53.990 33.465 54.160 33.635 ;
        RECT 52.435 32.725 52.705 33.185 ;
        RECT 52.875 32.895 53.160 33.355 ;
        RECT 53.530 33.295 54.160 33.465 ;
        RECT 53.530 32.895 53.705 33.295 ;
        RECT 54.510 33.225 54.680 34.515 ;
        RECT 53.875 32.725 54.205 33.105 ;
        RECT 54.450 32.895 54.680 33.225 ;
        RECT 54.880 33.060 55.160 34.335 ;
        RECT 55.385 33.575 55.655 34.335 ;
        RECT 55.345 33.405 55.655 33.575 ;
        RECT 55.385 33.060 55.655 33.405 ;
        RECT 55.845 33.305 56.185 34.335 ;
        RECT 56.355 33.965 56.525 34.515 ;
        RECT 56.695 34.135 56.955 35.105 ;
        RECT 56.355 33.635 56.615 33.965 ;
        RECT 56.785 33.445 56.955 34.135 ;
        RECT 56.115 32.725 56.445 33.105 ;
        RECT 56.615 32.980 56.955 33.445 ;
        RECT 57.590 34.135 57.925 35.105 ;
        RECT 58.095 34.135 58.265 35.275 ;
        RECT 58.435 34.935 60.465 35.105 ;
        RECT 57.590 33.465 57.760 34.135 ;
        RECT 58.435 33.965 58.605 34.935 ;
        RECT 57.930 33.635 58.185 33.965 ;
        RECT 58.410 33.635 58.605 33.965 ;
        RECT 58.775 34.595 59.900 34.765 ;
        RECT 58.015 33.465 58.185 33.635 ;
        RECT 58.775 33.465 58.945 34.595 ;
        RECT 56.615 32.935 56.950 32.980 ;
        RECT 57.590 32.895 57.845 33.465 ;
        RECT 58.015 33.295 58.945 33.465 ;
        RECT 59.115 34.255 60.125 34.425 ;
        RECT 59.115 33.455 59.285 34.255 ;
        RECT 58.770 33.260 58.945 33.295 ;
        RECT 58.015 32.725 58.345 33.125 ;
        RECT 58.770 32.895 59.300 33.260 ;
        RECT 59.490 33.235 59.765 34.055 ;
        RECT 59.485 33.065 59.765 33.235 ;
        RECT 59.490 32.895 59.765 33.065 ;
        RECT 59.935 32.895 60.125 34.255 ;
        RECT 60.295 34.270 60.465 34.935 ;
        RECT 60.635 34.515 60.805 35.275 ;
        RECT 61.040 34.515 61.555 34.925 ;
        RECT 60.295 34.080 61.045 34.270 ;
        RECT 61.215 33.705 61.555 34.515 ;
        RECT 61.725 34.185 62.935 35.275 ;
        RECT 60.325 33.535 61.555 33.705 ;
        RECT 60.305 32.725 60.815 33.260 ;
        RECT 61.035 32.930 61.280 33.535 ;
        RECT 61.725 33.475 62.245 34.015 ;
        RECT 62.415 33.645 62.935 34.185 ;
        RECT 63.110 34.125 63.370 35.275 ;
        RECT 63.545 34.200 63.800 35.105 ;
        RECT 63.970 34.515 64.300 35.275 ;
        RECT 64.515 34.345 64.685 35.105 ;
        RECT 61.725 32.725 62.935 33.475 ;
        RECT 63.110 32.725 63.370 33.565 ;
        RECT 63.545 33.470 63.715 34.200 ;
        RECT 63.970 34.175 64.685 34.345 ;
        RECT 63.970 33.965 64.140 34.175 ;
        RECT 64.945 34.135 65.285 35.105 ;
        RECT 65.455 34.135 65.625 35.275 ;
        RECT 65.895 34.475 66.145 35.275 ;
        RECT 66.790 34.305 67.120 35.105 ;
        RECT 67.420 34.475 67.750 35.275 ;
        RECT 67.920 34.305 68.250 35.105 ;
        RECT 65.815 34.135 68.250 34.305 ;
        RECT 68.625 34.185 69.835 35.275 ;
        RECT 63.885 33.635 64.140 33.965 ;
        RECT 63.545 32.895 63.800 33.470 ;
        RECT 63.970 33.445 64.140 33.635 ;
        RECT 64.420 33.625 64.775 33.995 ;
        RECT 64.945 33.525 65.120 34.135 ;
        RECT 65.815 33.885 65.985 34.135 ;
        RECT 65.290 33.715 65.985 33.885 ;
        RECT 66.160 33.715 66.580 33.915 ;
        RECT 66.750 33.715 67.080 33.915 ;
        RECT 67.250 33.715 67.580 33.915 ;
        RECT 63.970 33.275 64.685 33.445 ;
        RECT 63.970 32.725 64.300 33.105 ;
        RECT 64.515 32.895 64.685 33.275 ;
        RECT 64.945 32.895 65.285 33.525 ;
        RECT 65.455 32.725 65.705 33.525 ;
        RECT 65.895 33.375 67.120 33.545 ;
        RECT 65.895 32.895 66.225 33.375 ;
        RECT 66.395 32.725 66.620 33.185 ;
        RECT 66.790 32.895 67.120 33.375 ;
        RECT 67.750 33.505 67.920 34.135 ;
        RECT 68.105 33.715 68.455 33.965 ;
        RECT 67.750 32.895 68.250 33.505 ;
        RECT 68.625 33.475 69.145 34.015 ;
        RECT 69.315 33.645 69.835 34.185 ;
        RECT 70.005 34.110 70.295 35.275 ;
        RECT 70.470 34.885 70.805 35.105 ;
        RECT 71.810 34.895 72.165 35.275 ;
        RECT 70.470 34.265 70.725 34.885 ;
        RECT 70.975 34.725 71.205 34.765 ;
        RECT 72.335 34.725 72.585 35.105 ;
        RECT 70.975 34.525 72.585 34.725 ;
        RECT 70.975 34.435 71.160 34.525 ;
        RECT 71.750 34.515 72.585 34.525 ;
        RECT 72.835 34.495 73.085 35.275 ;
        RECT 73.255 34.425 73.515 35.105 ;
        RECT 74.695 34.605 74.865 35.105 ;
        RECT 75.035 34.775 75.365 35.275 ;
        RECT 74.695 34.435 75.360 34.605 ;
        RECT 71.315 34.325 71.645 34.355 ;
        RECT 71.315 34.265 73.115 34.325 ;
        RECT 70.470 34.155 73.175 34.265 ;
        RECT 70.470 34.095 71.645 34.155 ;
        RECT 72.975 34.120 73.175 34.155 ;
        RECT 70.465 33.715 70.955 33.915 ;
        RECT 71.145 33.715 71.620 33.925 ;
        RECT 68.625 32.725 69.835 33.475 ;
        RECT 70.005 32.725 70.295 33.450 ;
        RECT 70.470 32.725 70.925 33.490 ;
        RECT 71.400 33.315 71.620 33.715 ;
        RECT 71.865 33.715 72.195 33.925 ;
        RECT 71.865 33.315 72.075 33.715 ;
        RECT 72.365 33.680 72.775 33.985 ;
        RECT 73.005 33.545 73.175 34.120 ;
        RECT 72.905 33.425 73.175 33.545 ;
        RECT 72.330 33.380 73.175 33.425 ;
        RECT 72.330 33.255 73.085 33.380 ;
        RECT 72.330 33.105 72.500 33.255 ;
        RECT 73.345 33.225 73.515 34.425 ;
        RECT 74.610 33.615 74.960 34.265 ;
        RECT 75.130 33.445 75.360 34.435 ;
        RECT 71.200 32.895 72.500 33.105 ;
        RECT 72.755 32.725 73.085 33.085 ;
        RECT 73.255 32.895 73.515 33.225 ;
        RECT 74.695 33.275 75.360 33.445 ;
        RECT 74.695 32.985 74.865 33.275 ;
        RECT 75.035 32.725 75.365 33.105 ;
        RECT 75.535 32.985 75.720 35.105 ;
        RECT 75.960 34.815 76.225 35.275 ;
        RECT 76.395 34.680 76.645 35.105 ;
        RECT 76.855 34.830 77.960 35.000 ;
        RECT 76.340 34.550 76.645 34.680 ;
        RECT 75.890 33.355 76.170 34.305 ;
        RECT 76.340 33.445 76.510 34.550 ;
        RECT 76.680 33.765 76.920 34.360 ;
        RECT 77.090 34.295 77.620 34.660 ;
        RECT 77.090 33.595 77.260 34.295 ;
        RECT 77.790 34.215 77.960 34.830 ;
        RECT 78.130 34.475 78.300 35.275 ;
        RECT 78.470 34.775 78.720 35.105 ;
        RECT 78.945 34.805 79.830 34.975 ;
        RECT 77.790 34.125 78.300 34.215 ;
        RECT 76.340 33.315 76.565 33.445 ;
        RECT 76.735 33.375 77.260 33.595 ;
        RECT 77.430 33.955 78.300 34.125 ;
        RECT 75.975 32.725 76.225 33.185 ;
        RECT 76.395 33.175 76.565 33.315 ;
        RECT 77.430 33.175 77.600 33.955 ;
        RECT 78.130 33.885 78.300 33.955 ;
        RECT 77.810 33.705 78.010 33.735 ;
        RECT 78.470 33.705 78.640 34.775 ;
        RECT 78.810 33.885 79.000 34.605 ;
        RECT 77.810 33.405 78.640 33.705 ;
        RECT 79.170 33.675 79.490 34.635 ;
        RECT 76.395 33.005 76.730 33.175 ;
        RECT 76.925 33.005 77.600 33.175 ;
        RECT 77.920 32.725 78.290 33.225 ;
        RECT 78.470 33.175 78.640 33.405 ;
        RECT 79.025 33.345 79.490 33.675 ;
        RECT 79.660 33.965 79.830 34.805 ;
        RECT 80.010 34.775 80.325 35.275 ;
        RECT 80.555 34.545 80.895 35.105 ;
        RECT 80.000 34.170 80.895 34.545 ;
        RECT 81.065 34.265 81.235 35.275 ;
        RECT 80.705 33.965 80.895 34.170 ;
        RECT 81.405 34.215 81.735 35.060 ;
        RECT 81.405 34.135 81.795 34.215 ;
        RECT 81.580 34.085 81.795 34.135 ;
        RECT 79.660 33.635 80.535 33.965 ;
        RECT 80.705 33.635 81.455 33.965 ;
        RECT 79.660 33.175 79.830 33.635 ;
        RECT 80.705 33.465 80.905 33.635 ;
        RECT 81.625 33.505 81.795 34.085 ;
        RECT 81.965 34.185 83.175 35.275 ;
        RECT 81.965 33.645 82.485 34.185 ;
        RECT 81.570 33.465 81.795 33.505 ;
        RECT 82.655 33.475 83.175 34.015 ;
        RECT 78.470 33.005 78.875 33.175 ;
        RECT 79.045 33.005 79.830 33.175 ;
        RECT 80.105 32.725 80.315 33.255 ;
        RECT 80.575 32.940 80.905 33.465 ;
        RECT 81.415 33.380 81.795 33.465 ;
        RECT 81.075 32.725 81.245 33.335 ;
        RECT 81.415 32.945 81.745 33.380 ;
        RECT 81.965 32.725 83.175 33.475 ;
        RECT 5.520 32.555 83.260 32.725 ;
        RECT 5.605 31.805 6.815 32.555 ;
        RECT 6.985 32.010 12.330 32.555 ;
        RECT 13.015 32.165 13.345 32.555 ;
        RECT 5.605 31.265 6.125 31.805 ;
        RECT 6.295 31.095 6.815 31.635 ;
        RECT 8.570 31.180 8.910 32.010 ;
        RECT 13.515 31.985 13.685 32.305 ;
        RECT 13.855 32.165 14.185 32.555 ;
        RECT 14.600 32.155 15.555 32.325 ;
        RECT 12.965 31.815 15.215 31.985 ;
        RECT 5.605 30.005 6.815 31.095 ;
        RECT 10.390 30.440 10.740 31.690 ;
        RECT 12.965 30.855 13.135 31.815 ;
        RECT 13.305 31.195 13.550 31.645 ;
        RECT 13.720 31.365 14.270 31.565 ;
        RECT 14.440 31.395 14.815 31.565 ;
        RECT 14.440 31.195 14.610 31.395 ;
        RECT 14.985 31.315 15.215 31.815 ;
        RECT 13.305 31.025 14.610 31.195 ;
        RECT 15.385 31.275 15.555 32.155 ;
        RECT 15.725 31.720 16.015 32.555 ;
        RECT 16.275 32.005 16.445 32.295 ;
        RECT 16.615 32.175 16.945 32.555 ;
        RECT 16.275 31.835 16.940 32.005 ;
        RECT 15.385 31.105 16.015 31.275 ;
        RECT 6.985 30.005 12.330 30.440 ;
        RECT 12.965 30.175 13.345 30.855 ;
        RECT 13.935 30.005 14.105 30.855 ;
        RECT 14.275 30.685 15.515 30.855 ;
        RECT 14.275 30.175 14.605 30.685 ;
        RECT 14.775 30.005 14.945 30.515 ;
        RECT 15.115 30.175 15.515 30.685 ;
        RECT 15.695 30.175 16.015 31.105 ;
        RECT 16.190 31.015 16.540 31.665 ;
        RECT 16.710 30.845 16.940 31.835 ;
        RECT 16.275 30.675 16.940 30.845 ;
        RECT 16.275 30.175 16.445 30.675 ;
        RECT 16.615 30.005 16.945 30.505 ;
        RECT 17.115 30.175 17.300 32.295 ;
        RECT 17.555 32.095 17.805 32.555 ;
        RECT 17.975 32.105 18.310 32.275 ;
        RECT 18.505 32.105 19.180 32.275 ;
        RECT 17.975 31.965 18.145 32.105 ;
        RECT 17.470 30.975 17.750 31.925 ;
        RECT 17.920 31.835 18.145 31.965 ;
        RECT 17.920 30.730 18.090 31.835 ;
        RECT 18.315 31.685 18.840 31.905 ;
        RECT 18.260 30.920 18.500 31.515 ;
        RECT 18.670 30.985 18.840 31.685 ;
        RECT 19.010 31.325 19.180 32.105 ;
        RECT 19.500 32.055 19.870 32.555 ;
        RECT 20.050 32.105 20.455 32.275 ;
        RECT 20.625 32.105 21.410 32.275 ;
        RECT 20.050 31.875 20.220 32.105 ;
        RECT 19.390 31.575 20.220 31.875 ;
        RECT 20.605 31.605 21.070 31.935 ;
        RECT 19.390 31.545 19.590 31.575 ;
        RECT 19.710 31.325 19.880 31.395 ;
        RECT 19.010 31.155 19.880 31.325 ;
        RECT 19.370 31.065 19.880 31.155 ;
        RECT 17.920 30.600 18.225 30.730 ;
        RECT 18.670 30.620 19.200 30.985 ;
        RECT 17.540 30.005 17.805 30.465 ;
        RECT 17.975 30.175 18.225 30.600 ;
        RECT 19.370 30.450 19.540 31.065 ;
        RECT 18.435 30.280 19.540 30.450 ;
        RECT 19.710 30.005 19.880 30.805 ;
        RECT 20.050 30.505 20.220 31.575 ;
        RECT 20.390 30.675 20.580 31.395 ;
        RECT 20.750 30.645 21.070 31.605 ;
        RECT 21.240 31.645 21.410 32.105 ;
        RECT 21.685 32.025 21.895 32.555 ;
        RECT 22.155 31.815 22.485 32.340 ;
        RECT 22.655 31.945 22.825 32.555 ;
        RECT 22.995 31.900 23.325 32.335 ;
        RECT 23.545 31.905 23.805 32.385 ;
        RECT 23.975 32.015 24.225 32.555 ;
        RECT 22.995 31.815 23.375 31.900 ;
        RECT 22.285 31.645 22.485 31.815 ;
        RECT 23.150 31.775 23.375 31.815 ;
        RECT 21.240 31.315 22.115 31.645 ;
        RECT 22.285 31.315 23.035 31.645 ;
        RECT 20.050 30.175 20.300 30.505 ;
        RECT 21.240 30.475 21.410 31.315 ;
        RECT 22.285 31.110 22.475 31.315 ;
        RECT 23.205 31.195 23.375 31.775 ;
        RECT 23.160 31.145 23.375 31.195 ;
        RECT 21.580 30.735 22.475 31.110 ;
        RECT 22.985 31.065 23.375 31.145 ;
        RECT 20.525 30.305 21.410 30.475 ;
        RECT 21.590 30.005 21.905 30.505 ;
        RECT 22.135 30.175 22.475 30.735 ;
        RECT 22.645 30.005 22.815 31.015 ;
        RECT 22.985 30.220 23.315 31.065 ;
        RECT 23.545 30.875 23.715 31.905 ;
        RECT 24.395 31.875 24.615 32.335 ;
        RECT 24.365 31.850 24.615 31.875 ;
        RECT 23.885 31.255 24.115 31.650 ;
        RECT 24.285 31.425 24.615 31.850 ;
        RECT 24.785 32.175 25.675 32.345 ;
        RECT 24.785 31.450 24.955 32.175 ;
        RECT 25.125 31.620 25.675 32.005 ;
        RECT 25.845 31.805 27.055 32.555 ;
        RECT 27.245 31.865 27.485 32.385 ;
        RECT 27.655 32.060 28.050 32.555 ;
        RECT 28.615 32.225 28.785 32.370 ;
        RECT 28.410 32.030 28.785 32.225 ;
        RECT 24.785 31.380 25.675 31.450 ;
        RECT 24.780 31.355 25.675 31.380 ;
        RECT 24.770 31.340 25.675 31.355 ;
        RECT 24.765 31.325 25.675 31.340 ;
        RECT 24.755 31.320 25.675 31.325 ;
        RECT 24.750 31.310 25.675 31.320 ;
        RECT 24.745 31.300 25.675 31.310 ;
        RECT 24.735 31.295 25.675 31.300 ;
        RECT 24.725 31.285 25.675 31.295 ;
        RECT 24.715 31.280 25.675 31.285 ;
        RECT 24.715 31.275 25.050 31.280 ;
        RECT 24.700 31.270 25.050 31.275 ;
        RECT 24.685 31.260 25.050 31.270 ;
        RECT 24.660 31.255 25.050 31.260 ;
        RECT 23.885 31.250 25.050 31.255 ;
        RECT 23.885 31.215 25.020 31.250 ;
        RECT 23.885 31.190 24.985 31.215 ;
        RECT 23.885 31.160 24.955 31.190 ;
        RECT 23.885 31.130 24.935 31.160 ;
        RECT 23.885 31.100 24.915 31.130 ;
        RECT 23.885 31.090 24.845 31.100 ;
        RECT 23.885 31.080 24.820 31.090 ;
        RECT 23.885 31.065 24.800 31.080 ;
        RECT 23.885 31.050 24.780 31.065 ;
        RECT 23.990 31.040 24.775 31.050 ;
        RECT 23.990 31.005 24.760 31.040 ;
        RECT 23.545 30.175 23.820 30.875 ;
        RECT 23.990 30.755 24.745 31.005 ;
        RECT 24.915 30.685 25.245 30.930 ;
        RECT 25.415 30.830 25.675 31.280 ;
        RECT 25.845 31.265 26.365 31.805 ;
        RECT 26.535 31.095 27.055 31.635 ;
        RECT 25.060 30.660 25.245 30.685 ;
        RECT 25.060 30.560 25.675 30.660 ;
        RECT 23.990 30.005 24.245 30.550 ;
        RECT 24.415 30.175 24.895 30.515 ;
        RECT 25.070 30.005 25.675 30.560 ;
        RECT 25.845 30.005 27.055 31.095 ;
        RECT 27.245 31.060 27.420 31.865 ;
        RECT 28.410 31.695 28.580 32.030 ;
        RECT 29.065 31.985 29.305 32.360 ;
        RECT 29.475 32.050 29.810 32.555 ;
        RECT 29.065 31.835 29.285 31.985 ;
        RECT 27.595 31.335 28.580 31.695 ;
        RECT 28.750 31.505 29.285 31.835 ;
        RECT 27.595 31.315 28.880 31.335 ;
        RECT 28.020 31.165 28.880 31.315 ;
        RECT 27.245 30.275 27.550 31.060 ;
        RECT 27.725 30.685 28.420 30.995 ;
        RECT 27.730 30.005 28.415 30.475 ;
        RECT 28.595 30.220 28.880 31.165 ;
        RECT 29.050 30.855 29.285 31.505 ;
        RECT 29.455 31.025 29.755 31.875 ;
        RECT 29.985 31.805 31.195 32.555 ;
        RECT 31.365 31.830 31.655 32.555 ;
        RECT 29.985 31.265 30.505 31.805 ;
        RECT 30.675 31.095 31.195 31.635 ;
        RECT 29.050 30.625 29.725 30.855 ;
        RECT 29.055 30.005 29.385 30.455 ;
        RECT 29.555 30.195 29.725 30.625 ;
        RECT 29.985 30.005 31.195 31.095 ;
        RECT 31.365 30.005 31.655 31.170 ;
        RECT 31.835 30.185 32.095 32.375 ;
        RECT 32.355 32.185 33.025 32.555 ;
        RECT 33.205 32.005 33.515 32.375 ;
        RECT 32.285 31.805 33.515 32.005 ;
        RECT 32.285 31.135 32.575 31.805 ;
        RECT 33.695 31.625 33.925 32.265 ;
        RECT 34.105 31.825 34.395 32.555 ;
        RECT 34.585 32.010 39.930 32.555 ;
        RECT 40.105 32.010 45.450 32.555 ;
        RECT 32.755 31.315 33.220 31.625 ;
        RECT 33.400 31.315 33.925 31.625 ;
        RECT 34.105 31.315 34.405 31.645 ;
        RECT 36.170 31.180 36.510 32.010 ;
        RECT 32.285 30.915 33.055 31.135 ;
        RECT 32.265 30.005 32.605 30.735 ;
        RECT 32.785 30.185 33.055 30.915 ;
        RECT 33.235 30.895 34.395 31.135 ;
        RECT 33.235 30.185 33.465 30.895 ;
        RECT 33.635 30.005 33.965 30.715 ;
        RECT 34.135 30.185 34.395 30.895 ;
        RECT 37.990 30.440 38.340 31.690 ;
        RECT 41.690 31.180 42.030 32.010 ;
        RECT 45.625 31.785 47.295 32.555 ;
        RECT 43.510 30.440 43.860 31.690 ;
        RECT 45.625 31.265 46.375 31.785 ;
        RECT 47.465 31.755 48.160 32.385 ;
        RECT 48.365 31.755 48.675 32.555 ;
        RECT 48.850 32.025 49.140 32.375 ;
        RECT 49.335 32.195 49.665 32.555 ;
        RECT 49.835 32.025 50.065 32.330 ;
        RECT 48.850 31.855 50.065 32.025 ;
        RECT 46.545 31.095 47.295 31.615 ;
        RECT 47.485 31.315 47.820 31.565 ;
        RECT 47.990 31.155 48.160 31.755 ;
        RECT 50.255 31.685 50.425 32.250 ;
        RECT 48.330 31.315 48.665 31.585 ;
        RECT 48.910 31.535 49.170 31.645 ;
        RECT 48.905 31.365 49.170 31.535 ;
        RECT 48.910 31.315 49.170 31.365 ;
        RECT 49.350 31.315 49.735 31.645 ;
        RECT 49.905 31.515 50.425 31.685 ;
        RECT 51.605 31.905 51.865 32.385 ;
        RECT 52.035 32.015 52.285 32.555 ;
        RECT 34.585 30.005 39.930 30.440 ;
        RECT 40.105 30.005 45.450 30.440 ;
        RECT 45.625 30.005 47.295 31.095 ;
        RECT 47.465 30.005 47.725 31.145 ;
        RECT 47.895 30.175 48.225 31.155 ;
        RECT 48.395 30.005 48.675 31.145 ;
        RECT 48.850 30.005 49.170 31.145 ;
        RECT 49.350 30.265 49.545 31.315 ;
        RECT 49.905 31.135 50.075 31.515 ;
        RECT 49.725 30.855 50.075 31.135 ;
        RECT 50.265 30.985 50.510 31.345 ;
        RECT 51.605 30.875 51.775 31.905 ;
        RECT 52.455 31.850 52.675 32.335 ;
        RECT 51.945 31.255 52.175 31.650 ;
        RECT 52.345 31.425 52.675 31.850 ;
        RECT 52.845 32.175 53.735 32.345 ;
        RECT 52.845 31.450 53.015 32.175 ;
        RECT 53.185 31.620 53.735 32.005 ;
        RECT 53.905 31.735 54.165 32.555 ;
        RECT 54.335 31.735 54.665 32.155 ;
        RECT 54.845 32.070 55.635 32.335 ;
        RECT 54.415 31.645 54.665 31.735 ;
        RECT 52.845 31.380 53.735 31.450 ;
        RECT 52.840 31.355 53.735 31.380 ;
        RECT 52.830 31.340 53.735 31.355 ;
        RECT 52.825 31.325 53.735 31.340 ;
        RECT 52.815 31.320 53.735 31.325 ;
        RECT 52.810 31.310 53.735 31.320 ;
        RECT 52.805 31.300 53.735 31.310 ;
        RECT 52.795 31.295 53.735 31.300 ;
        RECT 52.785 31.285 53.735 31.295 ;
        RECT 52.775 31.280 53.735 31.285 ;
        RECT 52.775 31.275 53.110 31.280 ;
        RECT 52.760 31.270 53.110 31.275 ;
        RECT 52.745 31.260 53.110 31.270 ;
        RECT 52.720 31.255 53.110 31.260 ;
        RECT 51.945 31.250 53.110 31.255 ;
        RECT 51.945 31.215 53.080 31.250 ;
        RECT 51.945 31.190 53.045 31.215 ;
        RECT 51.945 31.160 53.015 31.190 ;
        RECT 51.945 31.130 52.995 31.160 ;
        RECT 51.945 31.100 52.975 31.130 ;
        RECT 51.945 31.090 52.905 31.100 ;
        RECT 51.945 31.080 52.880 31.090 ;
        RECT 51.945 31.065 52.860 31.080 ;
        RECT 51.945 31.050 52.840 31.065 ;
        RECT 52.050 31.040 52.835 31.050 ;
        RECT 52.050 31.005 52.820 31.040 ;
        RECT 49.725 30.175 50.055 30.855 ;
        RECT 50.255 30.005 50.510 30.805 ;
        RECT 51.605 30.175 51.880 30.875 ;
        RECT 52.050 30.755 52.805 31.005 ;
        RECT 52.975 30.685 53.305 30.930 ;
        RECT 53.475 30.830 53.735 31.280 ;
        RECT 53.905 30.685 54.245 31.565 ;
        RECT 54.415 31.395 55.210 31.645 ;
        RECT 53.120 30.660 53.305 30.685 ;
        RECT 53.120 30.560 53.735 30.660 ;
        RECT 52.050 30.005 52.305 30.550 ;
        RECT 52.475 30.175 52.955 30.515 ;
        RECT 53.130 30.005 53.735 30.560 ;
        RECT 53.905 30.005 54.165 30.515 ;
        RECT 54.415 30.175 54.585 31.395 ;
        RECT 55.380 31.215 55.635 32.070 ;
        RECT 55.805 31.915 56.005 32.335 ;
        RECT 56.195 32.095 56.525 32.555 ;
        RECT 55.805 31.395 56.215 31.915 ;
        RECT 56.695 31.905 56.955 32.385 ;
        RECT 56.385 31.215 56.615 31.645 ;
        RECT 54.825 31.045 56.615 31.215 ;
        RECT 54.825 30.680 55.075 31.045 ;
        RECT 55.245 30.685 55.575 30.875 ;
        RECT 55.795 30.750 56.510 31.045 ;
        RECT 56.785 30.875 56.955 31.905 ;
        RECT 57.125 31.830 57.415 32.555 ;
        RECT 57.585 31.735 57.845 32.555 ;
        RECT 58.015 31.735 58.345 32.155 ;
        RECT 58.525 31.985 58.785 32.385 ;
        RECT 58.955 32.155 59.285 32.555 ;
        RECT 59.455 31.985 59.625 32.335 ;
        RECT 59.795 32.155 60.170 32.555 ;
        RECT 58.525 31.815 60.190 31.985 ;
        RECT 60.360 31.880 60.635 32.225 ;
        RECT 58.095 31.645 58.345 31.735 ;
        RECT 60.020 31.645 60.190 31.815 ;
        RECT 57.590 31.315 57.925 31.565 ;
        RECT 58.095 31.315 58.810 31.645 ;
        RECT 59.025 31.315 59.850 31.645 ;
        RECT 60.020 31.315 60.295 31.645 ;
        RECT 55.245 30.510 55.440 30.685 ;
        RECT 54.825 30.005 55.440 30.510 ;
        RECT 55.610 30.175 56.085 30.515 ;
        RECT 56.255 30.005 56.470 30.550 ;
        RECT 56.680 30.175 56.955 30.875 ;
        RECT 57.125 30.005 57.415 31.170 ;
        RECT 57.585 30.005 57.845 31.145 ;
        RECT 58.095 30.755 58.265 31.315 ;
        RECT 58.525 30.855 58.855 31.145 ;
        RECT 59.025 31.025 59.270 31.315 ;
        RECT 60.020 31.145 60.190 31.315 ;
        RECT 60.465 31.145 60.635 31.880 ;
        RECT 61.730 31.715 61.990 32.555 ;
        RECT 62.165 31.810 62.420 32.385 ;
        RECT 62.590 32.175 62.920 32.555 ;
        RECT 63.135 32.005 63.305 32.385 ;
        RECT 62.590 31.835 63.305 32.005 ;
        RECT 59.530 30.975 60.190 31.145 ;
        RECT 59.530 30.855 59.700 30.975 ;
        RECT 58.525 30.685 59.700 30.855 ;
        RECT 58.085 30.185 59.700 30.515 ;
        RECT 59.870 30.005 60.150 30.805 ;
        RECT 60.360 30.175 60.635 31.145 ;
        RECT 61.730 30.005 61.990 31.155 ;
        RECT 62.165 31.080 62.335 31.810 ;
        RECT 62.590 31.645 62.760 31.835 ;
        RECT 63.570 31.715 63.830 32.555 ;
        RECT 64.005 31.810 64.260 32.385 ;
        RECT 64.430 32.175 64.760 32.555 ;
        RECT 64.975 32.005 65.145 32.385 ;
        RECT 64.430 31.835 65.145 32.005 ;
        RECT 62.505 31.315 62.760 31.645 ;
        RECT 62.590 31.105 62.760 31.315 ;
        RECT 63.040 31.285 63.395 31.655 ;
        RECT 62.165 30.175 62.420 31.080 ;
        RECT 62.590 30.935 63.305 31.105 ;
        RECT 62.590 30.005 62.920 30.765 ;
        RECT 63.135 30.175 63.305 30.935 ;
        RECT 63.570 30.005 63.830 31.155 ;
        RECT 64.005 31.080 64.175 31.810 ;
        RECT 64.430 31.645 64.600 31.835 ;
        RECT 65.440 31.815 66.055 32.385 ;
        RECT 66.225 32.045 66.440 32.555 ;
        RECT 66.670 32.045 66.950 32.375 ;
        RECT 67.130 32.045 67.370 32.555 ;
        RECT 64.345 31.315 64.600 31.645 ;
        RECT 64.430 31.105 64.600 31.315 ;
        RECT 64.880 31.285 65.235 31.655 ;
        RECT 64.005 30.175 64.260 31.080 ;
        RECT 64.430 30.935 65.145 31.105 ;
        RECT 64.430 30.005 64.760 30.765 ;
        RECT 64.975 30.175 65.145 30.935 ;
        RECT 65.440 30.795 65.755 31.815 ;
        RECT 65.925 31.145 66.095 31.645 ;
        RECT 66.345 31.315 66.610 31.875 ;
        RECT 66.780 31.145 66.950 32.045 ;
        RECT 67.120 31.315 67.475 31.875 ;
        RECT 67.740 31.815 68.355 32.385 ;
        RECT 68.525 32.045 68.740 32.555 ;
        RECT 68.970 32.045 69.250 32.375 ;
        RECT 69.430 32.045 69.670 32.555 ;
        RECT 65.925 30.975 67.350 31.145 ;
        RECT 65.440 30.175 65.975 30.795 ;
        RECT 66.145 30.005 66.475 30.805 ;
        RECT 66.960 30.800 67.350 30.975 ;
        RECT 67.740 30.795 68.055 31.815 ;
        RECT 68.225 31.145 68.395 31.645 ;
        RECT 68.645 31.315 68.910 31.875 ;
        RECT 69.080 31.145 69.250 32.045 ;
        RECT 69.420 31.315 69.775 31.875 ;
        RECT 70.500 31.815 71.115 32.385 ;
        RECT 71.285 32.045 71.500 32.555 ;
        RECT 71.730 32.045 72.010 32.375 ;
        RECT 72.190 32.045 72.430 32.555 ;
        RECT 68.225 30.975 69.650 31.145 ;
        RECT 67.740 30.175 68.275 30.795 ;
        RECT 68.445 30.005 68.775 30.805 ;
        RECT 69.260 30.800 69.650 30.975 ;
        RECT 70.500 30.795 70.815 31.815 ;
        RECT 70.985 31.145 71.155 31.645 ;
        RECT 71.405 31.315 71.670 31.875 ;
        RECT 71.840 31.145 72.010 32.045 ;
        RECT 72.855 32.005 73.025 32.385 ;
        RECT 73.240 32.175 73.570 32.555 ;
        RECT 72.180 31.315 72.535 31.875 ;
        RECT 72.855 31.835 73.570 32.005 ;
        RECT 72.765 31.285 73.120 31.655 ;
        RECT 73.400 31.645 73.570 31.835 ;
        RECT 73.740 31.810 73.995 32.385 ;
        RECT 73.400 31.315 73.655 31.645 ;
        RECT 70.985 30.975 72.410 31.145 ;
        RECT 73.400 31.105 73.570 31.315 ;
        RECT 70.500 30.175 71.035 30.795 ;
        RECT 71.205 30.005 71.535 30.805 ;
        RECT 72.020 30.800 72.410 30.975 ;
        RECT 72.855 30.935 73.570 31.105 ;
        RECT 73.825 31.080 73.995 31.810 ;
        RECT 74.170 31.715 74.430 32.555 ;
        RECT 74.810 31.775 75.310 32.385 ;
        RECT 74.605 31.315 74.955 31.565 ;
        RECT 72.855 30.175 73.025 30.935 ;
        RECT 73.240 30.005 73.570 30.765 ;
        RECT 73.740 30.175 73.995 31.080 ;
        RECT 74.170 30.005 74.430 31.155 ;
        RECT 75.140 31.145 75.310 31.775 ;
        RECT 75.940 31.905 76.270 32.385 ;
        RECT 76.440 32.095 76.665 32.555 ;
        RECT 76.835 31.905 77.165 32.385 ;
        RECT 75.940 31.735 77.165 31.905 ;
        RECT 77.355 31.755 77.605 32.555 ;
        RECT 77.775 31.755 78.115 32.385 ;
        RECT 75.480 31.365 75.810 31.565 ;
        RECT 75.980 31.365 76.310 31.565 ;
        RECT 76.480 31.535 76.900 31.565 ;
        RECT 76.480 31.365 76.905 31.535 ;
        RECT 77.075 31.395 77.770 31.565 ;
        RECT 77.075 31.145 77.245 31.395 ;
        RECT 77.940 31.145 78.115 31.755 ;
        RECT 74.810 30.975 77.245 31.145 ;
        RECT 74.810 30.175 75.140 30.975 ;
        RECT 75.310 30.005 75.640 30.805 ;
        RECT 75.940 30.175 76.270 30.975 ;
        RECT 76.915 30.005 77.165 30.805 ;
        RECT 77.435 30.005 77.605 31.145 ;
        RECT 77.775 30.175 78.115 31.145 ;
        RECT 78.285 32.055 78.545 32.385 ;
        RECT 78.715 32.195 79.045 32.555 ;
        RECT 79.300 32.175 80.600 32.385 ;
        RECT 78.285 32.045 78.515 32.055 ;
        RECT 78.285 30.855 78.455 32.045 ;
        RECT 79.300 32.025 79.470 32.175 ;
        RECT 78.715 31.900 79.470 32.025 ;
        RECT 78.625 31.855 79.470 31.900 ;
        RECT 78.625 31.735 78.895 31.855 ;
        RECT 78.625 31.160 78.795 31.735 ;
        RECT 79.025 31.295 79.435 31.600 ;
        RECT 79.725 31.565 79.935 31.965 ;
        RECT 79.605 31.355 79.935 31.565 ;
        RECT 80.180 31.565 80.400 31.965 ;
        RECT 80.875 31.790 81.330 32.555 ;
        RECT 81.965 31.805 83.175 32.555 ;
        RECT 80.180 31.355 80.655 31.565 ;
        RECT 80.845 31.365 81.335 31.565 ;
        RECT 78.625 31.125 78.825 31.160 ;
        RECT 80.155 31.125 81.330 31.185 ;
        RECT 78.625 31.015 81.330 31.125 ;
        RECT 78.685 30.955 80.485 31.015 ;
        RECT 80.155 30.925 80.485 30.955 ;
        RECT 78.285 30.175 78.545 30.855 ;
        RECT 78.715 30.005 78.965 30.785 ;
        RECT 79.215 30.755 80.050 30.765 ;
        RECT 80.640 30.755 80.825 30.845 ;
        RECT 79.215 30.555 80.825 30.755 ;
        RECT 79.215 30.175 79.465 30.555 ;
        RECT 80.595 30.515 80.825 30.555 ;
        RECT 81.075 30.395 81.330 31.015 ;
        RECT 79.635 30.005 79.990 30.385 ;
        RECT 80.995 30.175 81.330 30.395 ;
        RECT 81.965 31.095 82.485 31.635 ;
        RECT 82.655 31.265 83.175 31.805 ;
        RECT 81.965 30.005 83.175 31.095 ;
        RECT 5.520 29.835 83.260 30.005 ;
        RECT 5.605 28.745 6.815 29.835 ;
        RECT 6.985 29.400 12.330 29.835 ;
        RECT 12.505 29.400 17.850 29.835 ;
        RECT 5.605 28.035 6.125 28.575 ;
        RECT 6.295 28.205 6.815 28.745 ;
        RECT 5.605 27.285 6.815 28.035 ;
        RECT 8.570 27.830 8.910 28.660 ;
        RECT 10.390 28.150 10.740 29.400 ;
        RECT 14.090 27.830 14.430 28.660 ;
        RECT 15.910 28.150 16.260 29.400 ;
        RECT 18.485 28.670 18.775 29.835 ;
        RECT 19.005 28.775 19.335 29.620 ;
        RECT 19.505 28.825 19.675 29.835 ;
        RECT 19.845 29.105 20.185 29.665 ;
        RECT 20.415 29.335 20.730 29.835 ;
        RECT 20.910 29.365 21.795 29.535 ;
        RECT 18.945 28.695 19.335 28.775 ;
        RECT 19.845 28.730 20.740 29.105 ;
        RECT 18.945 28.645 19.160 28.695 ;
        RECT 18.945 28.065 19.115 28.645 ;
        RECT 19.845 28.525 20.035 28.730 ;
        RECT 20.910 28.525 21.080 29.365 ;
        RECT 22.020 29.335 22.270 29.665 ;
        RECT 19.285 28.195 20.035 28.525 ;
        RECT 20.205 28.195 21.080 28.525 ;
        RECT 18.945 28.025 19.170 28.065 ;
        RECT 19.835 28.025 20.035 28.195 ;
        RECT 6.985 27.285 12.330 27.830 ;
        RECT 12.505 27.285 17.850 27.830 ;
        RECT 18.485 27.285 18.775 28.010 ;
        RECT 18.945 27.940 19.325 28.025 ;
        RECT 18.995 27.505 19.325 27.940 ;
        RECT 19.495 27.285 19.665 27.895 ;
        RECT 19.835 27.500 20.165 28.025 ;
        RECT 20.425 27.285 20.635 27.815 ;
        RECT 20.910 27.735 21.080 28.195 ;
        RECT 21.250 28.235 21.570 29.195 ;
        RECT 21.740 28.445 21.930 29.165 ;
        RECT 22.100 28.265 22.270 29.335 ;
        RECT 22.440 29.035 22.610 29.835 ;
        RECT 22.780 29.390 23.885 29.560 ;
        RECT 22.780 28.775 22.950 29.390 ;
        RECT 24.095 29.240 24.345 29.665 ;
        RECT 24.515 29.375 24.780 29.835 ;
        RECT 23.120 28.855 23.650 29.220 ;
        RECT 24.095 29.110 24.400 29.240 ;
        RECT 22.440 28.685 22.950 28.775 ;
        RECT 22.440 28.515 23.310 28.685 ;
        RECT 22.440 28.445 22.610 28.515 ;
        RECT 22.730 28.265 22.930 28.295 ;
        RECT 21.250 27.905 21.715 28.235 ;
        RECT 22.100 27.965 22.930 28.265 ;
        RECT 22.100 27.735 22.270 27.965 ;
        RECT 20.910 27.565 21.695 27.735 ;
        RECT 21.865 27.565 22.270 27.735 ;
        RECT 22.450 27.285 22.820 27.785 ;
        RECT 23.140 27.735 23.310 28.515 ;
        RECT 23.480 28.155 23.650 28.855 ;
        RECT 23.820 28.325 24.060 28.920 ;
        RECT 23.480 27.935 24.005 28.155 ;
        RECT 24.230 28.005 24.400 29.110 ;
        RECT 24.175 27.875 24.400 28.005 ;
        RECT 24.570 27.915 24.850 28.865 ;
        RECT 24.175 27.735 24.345 27.875 ;
        RECT 23.140 27.565 23.815 27.735 ;
        RECT 24.010 27.565 24.345 27.735 ;
        RECT 24.515 27.285 24.765 27.745 ;
        RECT 25.020 27.545 25.205 29.665 ;
        RECT 25.375 29.335 25.705 29.835 ;
        RECT 25.875 29.165 26.045 29.665 ;
        RECT 25.380 28.995 26.045 29.165 ;
        RECT 26.395 29.165 26.565 29.665 ;
        RECT 26.735 29.335 27.065 29.835 ;
        RECT 26.395 28.995 27.060 29.165 ;
        RECT 25.380 28.005 25.610 28.995 ;
        RECT 25.780 28.175 26.130 28.825 ;
        RECT 26.310 28.175 26.660 28.825 ;
        RECT 26.830 28.005 27.060 28.995 ;
        RECT 25.380 27.835 26.045 28.005 ;
        RECT 25.375 27.285 25.705 27.665 ;
        RECT 25.875 27.545 26.045 27.835 ;
        RECT 26.395 27.835 27.060 28.005 ;
        RECT 26.395 27.545 26.565 27.835 ;
        RECT 26.735 27.285 27.065 27.665 ;
        RECT 27.235 27.545 27.420 29.665 ;
        RECT 27.660 29.375 27.925 29.835 ;
        RECT 28.095 29.240 28.345 29.665 ;
        RECT 28.555 29.390 29.660 29.560 ;
        RECT 28.040 29.110 28.345 29.240 ;
        RECT 27.590 27.915 27.870 28.865 ;
        RECT 28.040 28.005 28.210 29.110 ;
        RECT 28.380 28.325 28.620 28.920 ;
        RECT 28.790 28.855 29.320 29.220 ;
        RECT 28.790 28.155 28.960 28.855 ;
        RECT 29.490 28.775 29.660 29.390 ;
        RECT 29.830 29.035 30.000 29.835 ;
        RECT 30.170 29.335 30.420 29.665 ;
        RECT 30.645 29.365 31.530 29.535 ;
        RECT 29.490 28.685 30.000 28.775 ;
        RECT 28.040 27.875 28.265 28.005 ;
        RECT 28.435 27.935 28.960 28.155 ;
        RECT 29.130 28.515 30.000 28.685 ;
        RECT 27.675 27.285 27.925 27.745 ;
        RECT 28.095 27.735 28.265 27.875 ;
        RECT 29.130 27.735 29.300 28.515 ;
        RECT 29.830 28.445 30.000 28.515 ;
        RECT 29.510 28.265 29.710 28.295 ;
        RECT 30.170 28.265 30.340 29.335 ;
        RECT 30.510 28.445 30.700 29.165 ;
        RECT 29.510 27.965 30.340 28.265 ;
        RECT 30.870 28.235 31.190 29.195 ;
        RECT 28.095 27.565 28.430 27.735 ;
        RECT 28.625 27.565 29.300 27.735 ;
        RECT 29.620 27.285 29.990 27.785 ;
        RECT 30.170 27.735 30.340 27.965 ;
        RECT 30.725 27.905 31.190 28.235 ;
        RECT 31.360 28.525 31.530 29.365 ;
        RECT 31.710 29.335 32.025 29.835 ;
        RECT 32.255 29.105 32.595 29.665 ;
        RECT 31.700 28.730 32.595 29.105 ;
        RECT 32.765 28.825 32.935 29.835 ;
        RECT 32.405 28.525 32.595 28.730 ;
        RECT 33.105 28.775 33.435 29.620 ;
        RECT 33.665 29.400 39.010 29.835 ;
        RECT 33.105 28.695 33.495 28.775 ;
        RECT 33.280 28.645 33.495 28.695 ;
        RECT 31.360 28.195 32.235 28.525 ;
        RECT 32.405 28.195 33.155 28.525 ;
        RECT 31.360 27.735 31.530 28.195 ;
        RECT 32.405 28.025 32.605 28.195 ;
        RECT 33.325 28.065 33.495 28.645 ;
        RECT 33.270 28.025 33.495 28.065 ;
        RECT 30.170 27.565 30.575 27.735 ;
        RECT 30.745 27.565 31.530 27.735 ;
        RECT 31.805 27.285 32.015 27.815 ;
        RECT 32.275 27.500 32.605 28.025 ;
        RECT 33.115 27.940 33.495 28.025 ;
        RECT 32.775 27.285 32.945 27.895 ;
        RECT 33.115 27.505 33.445 27.940 ;
        RECT 35.250 27.830 35.590 28.660 ;
        RECT 37.070 28.150 37.420 29.400 ;
        RECT 39.185 28.745 42.695 29.835 ;
        RECT 42.865 28.745 44.075 29.835 ;
        RECT 39.185 28.055 40.835 28.575 ;
        RECT 41.005 28.225 42.695 28.745 ;
        RECT 33.665 27.285 39.010 27.830 ;
        RECT 39.185 27.285 42.695 28.055 ;
        RECT 42.865 28.035 43.385 28.575 ;
        RECT 43.555 28.205 44.075 28.745 ;
        RECT 44.245 28.670 44.535 29.835 ;
        RECT 44.705 29.400 50.050 29.835 ;
        RECT 42.865 27.285 44.075 28.035 ;
        RECT 44.245 27.285 44.535 28.010 ;
        RECT 46.290 27.830 46.630 28.660 ;
        RECT 48.110 28.150 48.460 29.400 ;
        RECT 50.225 28.745 51.895 29.835 ;
        RECT 50.225 28.055 50.975 28.575 ;
        RECT 51.145 28.225 51.895 28.745 ;
        RECT 52.525 28.695 52.805 29.835 ;
        RECT 52.975 28.685 53.305 29.665 ;
        RECT 53.475 28.695 53.735 29.835 ;
        RECT 53.915 28.865 54.245 29.650 ;
        RECT 53.915 28.695 54.595 28.865 ;
        RECT 54.775 28.695 55.105 29.835 ;
        RECT 55.285 28.745 56.495 29.835 ;
        RECT 52.535 28.255 52.870 28.525 ;
        RECT 53.040 28.085 53.210 28.685 ;
        RECT 53.380 28.275 53.715 28.525 ;
        RECT 53.905 28.275 54.255 28.525 ;
        RECT 54.425 28.095 54.595 28.695 ;
        RECT 54.765 28.275 55.115 28.525 ;
        RECT 44.705 27.285 50.050 27.830 ;
        RECT 50.225 27.285 51.895 28.055 ;
        RECT 52.525 27.285 52.835 28.085 ;
        RECT 53.040 27.455 53.735 28.085 ;
        RECT 53.925 27.285 54.165 28.095 ;
        RECT 54.335 27.455 54.665 28.095 ;
        RECT 54.835 27.285 55.105 28.095 ;
        RECT 55.285 28.035 55.805 28.575 ;
        RECT 55.975 28.205 56.495 28.745 ;
        RECT 56.705 28.695 56.935 29.835 ;
        RECT 57.105 28.685 57.435 29.665 ;
        RECT 57.605 28.695 57.815 29.835 ;
        RECT 58.045 28.745 59.255 29.835 ;
        RECT 56.685 28.275 57.015 28.525 ;
        RECT 55.285 27.285 56.495 28.035 ;
        RECT 56.705 27.285 56.935 28.105 ;
        RECT 57.185 28.085 57.435 28.685 ;
        RECT 57.105 27.455 57.435 28.085 ;
        RECT 57.605 27.285 57.815 28.105 ;
        RECT 58.045 28.035 58.565 28.575 ;
        RECT 58.735 28.205 59.255 28.745 ;
        RECT 59.430 28.685 59.690 29.835 ;
        RECT 59.865 28.760 60.120 29.665 ;
        RECT 60.290 29.075 60.620 29.835 ;
        RECT 60.835 28.905 61.005 29.665 ;
        RECT 58.045 27.285 59.255 28.035 ;
        RECT 59.430 27.285 59.690 28.125 ;
        RECT 59.865 28.030 60.035 28.760 ;
        RECT 60.290 28.735 61.005 28.905 ;
        RECT 60.290 28.525 60.460 28.735 ;
        RECT 61.270 28.685 61.530 29.835 ;
        RECT 61.705 28.760 61.960 29.665 ;
        RECT 62.130 29.075 62.460 29.835 ;
        RECT 62.675 28.905 62.845 29.665 ;
        RECT 60.205 28.195 60.460 28.525 ;
        RECT 59.865 27.455 60.120 28.030 ;
        RECT 60.290 28.005 60.460 28.195 ;
        RECT 60.740 28.185 61.095 28.555 ;
        RECT 60.290 27.835 61.005 28.005 ;
        RECT 60.290 27.285 60.620 27.665 ;
        RECT 60.835 27.455 61.005 27.835 ;
        RECT 61.270 27.285 61.530 28.125 ;
        RECT 61.705 28.030 61.875 28.760 ;
        RECT 62.130 28.735 62.845 28.905 ;
        RECT 63.140 29.045 63.675 29.665 ;
        RECT 62.130 28.525 62.300 28.735 ;
        RECT 62.045 28.195 62.300 28.525 ;
        RECT 61.705 27.455 61.960 28.030 ;
        RECT 62.130 28.005 62.300 28.195 ;
        RECT 62.580 28.185 62.935 28.555 ;
        RECT 63.140 28.025 63.455 29.045 ;
        RECT 63.845 29.035 64.175 29.835 ;
        RECT 64.660 28.865 65.050 29.040 ;
        RECT 63.625 28.695 65.050 28.865 ;
        RECT 65.590 28.865 65.980 29.040 ;
        RECT 66.465 29.035 66.795 29.835 ;
        RECT 66.965 29.045 67.500 29.665 ;
        RECT 65.590 28.695 67.015 28.865 ;
        RECT 63.625 28.195 63.795 28.695 ;
        RECT 62.130 27.835 62.845 28.005 ;
        RECT 62.130 27.285 62.460 27.665 ;
        RECT 62.675 27.455 62.845 27.835 ;
        RECT 63.140 27.455 63.755 28.025 ;
        RECT 64.045 27.965 64.310 28.525 ;
        RECT 64.480 27.795 64.650 28.695 ;
        RECT 64.820 27.965 65.175 28.525 ;
        RECT 65.465 27.965 65.820 28.525 ;
        RECT 65.990 27.795 66.160 28.695 ;
        RECT 66.330 27.965 66.595 28.525 ;
        RECT 66.845 28.195 67.015 28.695 ;
        RECT 67.185 28.025 67.500 29.045 ;
        RECT 67.890 28.865 68.280 29.040 ;
        RECT 68.765 29.035 69.095 29.835 ;
        RECT 69.265 29.045 69.800 29.665 ;
        RECT 67.890 28.695 69.315 28.865 ;
        RECT 63.925 27.285 64.140 27.795 ;
        RECT 64.370 27.465 64.650 27.795 ;
        RECT 64.830 27.285 65.070 27.795 ;
        RECT 65.570 27.285 65.810 27.795 ;
        RECT 65.990 27.465 66.270 27.795 ;
        RECT 66.500 27.285 66.715 27.795 ;
        RECT 66.885 27.455 67.500 28.025 ;
        RECT 67.765 27.965 68.120 28.525 ;
        RECT 68.290 27.795 68.460 28.695 ;
        RECT 68.630 27.965 68.895 28.525 ;
        RECT 69.145 28.195 69.315 28.695 ;
        RECT 69.485 28.025 69.800 29.045 ;
        RECT 70.005 28.670 70.295 29.835 ;
        RECT 70.470 29.445 70.805 29.665 ;
        RECT 71.810 29.455 72.165 29.835 ;
        RECT 70.470 28.825 70.725 29.445 ;
        RECT 70.975 29.285 71.205 29.325 ;
        RECT 72.335 29.285 72.585 29.665 ;
        RECT 70.975 29.085 72.585 29.285 ;
        RECT 70.975 28.995 71.160 29.085 ;
        RECT 71.750 29.075 72.585 29.085 ;
        RECT 72.835 29.055 73.085 29.835 ;
        RECT 73.255 28.985 73.515 29.665 ;
        RECT 71.315 28.885 71.645 28.915 ;
        RECT 71.315 28.825 73.115 28.885 ;
        RECT 70.470 28.715 73.175 28.825 ;
        RECT 70.470 28.655 71.645 28.715 ;
        RECT 72.975 28.680 73.175 28.715 ;
        RECT 70.465 28.275 70.955 28.475 ;
        RECT 71.145 28.275 71.620 28.485 ;
        RECT 67.870 27.285 68.110 27.795 ;
        RECT 68.290 27.465 68.570 27.795 ;
        RECT 68.800 27.285 69.015 27.795 ;
        RECT 69.185 27.455 69.800 28.025 ;
        RECT 70.005 27.285 70.295 28.010 ;
        RECT 70.470 27.285 70.925 28.050 ;
        RECT 71.400 27.875 71.620 28.275 ;
        RECT 71.865 28.275 72.195 28.485 ;
        RECT 71.865 27.875 72.075 28.275 ;
        RECT 72.365 28.240 72.775 28.545 ;
        RECT 73.005 28.105 73.175 28.680 ;
        RECT 72.905 27.985 73.175 28.105 ;
        RECT 72.330 27.940 73.175 27.985 ;
        RECT 72.330 27.815 73.085 27.940 ;
        RECT 72.330 27.665 72.500 27.815 ;
        RECT 73.345 27.795 73.515 28.985 ;
        RECT 73.285 27.785 73.515 27.795 ;
        RECT 71.200 27.455 72.500 27.665 ;
        RECT 72.755 27.285 73.085 27.645 ;
        RECT 73.255 27.455 73.515 27.785 ;
        RECT 73.685 28.985 73.945 29.665 ;
        RECT 74.115 29.055 74.365 29.835 ;
        RECT 74.615 29.285 74.865 29.665 ;
        RECT 75.035 29.455 75.390 29.835 ;
        RECT 76.395 29.445 76.730 29.665 ;
        RECT 75.995 29.285 76.225 29.325 ;
        RECT 74.615 29.085 76.225 29.285 ;
        RECT 74.615 29.075 75.450 29.085 ;
        RECT 76.040 28.995 76.225 29.085 ;
        RECT 73.685 27.785 73.855 28.985 ;
        RECT 75.555 28.885 75.885 28.915 ;
        RECT 74.085 28.825 75.885 28.885 ;
        RECT 76.475 28.825 76.730 29.445 ;
        RECT 74.025 28.715 76.730 28.825 ;
        RECT 74.025 28.680 74.225 28.715 ;
        RECT 74.025 28.105 74.195 28.680 ;
        RECT 75.555 28.655 76.730 28.715 ;
        RECT 77.365 28.695 77.705 29.665 ;
        RECT 77.875 28.695 78.045 29.835 ;
        RECT 78.315 29.035 78.565 29.835 ;
        RECT 79.210 28.865 79.540 29.665 ;
        RECT 79.840 29.035 80.170 29.835 ;
        RECT 80.340 28.865 80.670 29.665 ;
        RECT 78.235 28.695 80.670 28.865 ;
        RECT 81.965 28.745 83.175 29.835 ;
        RECT 74.425 28.240 74.835 28.545 ;
        RECT 75.005 28.275 75.335 28.485 ;
        RECT 74.025 27.985 74.295 28.105 ;
        RECT 74.025 27.940 74.870 27.985 ;
        RECT 74.115 27.815 74.870 27.940 ;
        RECT 75.125 27.875 75.335 28.275 ;
        RECT 75.580 28.275 76.055 28.485 ;
        RECT 76.245 28.275 76.735 28.475 ;
        RECT 75.580 27.875 75.800 28.275 ;
        RECT 77.365 28.085 77.540 28.695 ;
        RECT 78.235 28.445 78.405 28.695 ;
        RECT 77.710 28.275 78.405 28.445 ;
        RECT 78.580 28.275 79.000 28.475 ;
        RECT 79.170 28.275 79.500 28.475 ;
        RECT 79.670 28.275 80.000 28.475 ;
        RECT 73.685 27.455 73.945 27.785 ;
        RECT 74.700 27.665 74.870 27.815 ;
        RECT 74.115 27.285 74.445 27.645 ;
        RECT 74.700 27.455 76.000 27.665 ;
        RECT 76.275 27.285 76.730 28.050 ;
        RECT 77.365 27.455 77.705 28.085 ;
        RECT 77.875 27.285 78.125 28.085 ;
        RECT 78.315 27.935 79.540 28.105 ;
        RECT 78.315 27.455 78.645 27.935 ;
        RECT 78.815 27.285 79.040 27.745 ;
        RECT 79.210 27.455 79.540 27.935 ;
        RECT 80.170 28.065 80.340 28.695 ;
        RECT 80.525 28.275 80.875 28.525 ;
        RECT 81.965 28.205 82.485 28.745 ;
        RECT 80.170 27.455 80.670 28.065 ;
        RECT 82.655 28.035 83.175 28.575 ;
        RECT 81.965 27.285 83.175 28.035 ;
        RECT 5.520 27.115 83.260 27.285 ;
        RECT 5.605 26.365 6.815 27.115 ;
        RECT 6.985 26.570 12.330 27.115 ;
        RECT 12.505 26.570 17.850 27.115 ;
        RECT 18.025 26.570 23.370 27.115 ;
        RECT 23.545 26.570 28.890 27.115 ;
        RECT 5.605 25.825 6.125 26.365 ;
        RECT 6.295 25.655 6.815 26.195 ;
        RECT 8.570 25.740 8.910 26.570 ;
        RECT 5.605 24.565 6.815 25.655 ;
        RECT 10.390 25.000 10.740 26.250 ;
        RECT 14.090 25.740 14.430 26.570 ;
        RECT 15.910 25.000 16.260 26.250 ;
        RECT 19.610 25.740 19.950 26.570 ;
        RECT 21.430 25.000 21.780 26.250 ;
        RECT 25.130 25.740 25.470 26.570 ;
        RECT 29.065 26.345 30.735 27.115 ;
        RECT 31.365 26.390 31.655 27.115 ;
        RECT 31.825 26.570 37.170 27.115 ;
        RECT 37.345 26.570 42.690 27.115 ;
        RECT 42.865 26.570 48.210 27.115 ;
        RECT 26.950 25.000 27.300 26.250 ;
        RECT 29.065 25.825 29.815 26.345 ;
        RECT 29.985 25.655 30.735 26.175 ;
        RECT 33.410 25.740 33.750 26.570 ;
        RECT 6.985 24.565 12.330 25.000 ;
        RECT 12.505 24.565 17.850 25.000 ;
        RECT 18.025 24.565 23.370 25.000 ;
        RECT 23.545 24.565 28.890 25.000 ;
        RECT 29.065 24.565 30.735 25.655 ;
        RECT 31.365 24.565 31.655 25.730 ;
        RECT 35.230 25.000 35.580 26.250 ;
        RECT 38.930 25.740 39.270 26.570 ;
        RECT 40.750 25.000 41.100 26.250 ;
        RECT 44.450 25.740 44.790 26.570 ;
        RECT 48.385 26.365 49.595 27.115 ;
        RECT 46.270 25.000 46.620 26.250 ;
        RECT 48.385 25.825 48.905 26.365 ;
        RECT 49.765 26.315 50.460 26.945 ;
        RECT 50.665 26.315 50.975 27.115 ;
        RECT 51.180 26.375 51.795 26.945 ;
        RECT 51.965 26.605 52.180 27.115 ;
        RECT 52.410 26.605 52.690 26.935 ;
        RECT 52.870 26.605 53.110 27.115 ;
        RECT 49.075 25.655 49.595 26.195 ;
        RECT 49.785 25.875 50.120 26.125 ;
        RECT 50.290 25.715 50.460 26.315 ;
        RECT 50.630 25.875 50.965 26.145 ;
        RECT 31.825 24.565 37.170 25.000 ;
        RECT 37.345 24.565 42.690 25.000 ;
        RECT 42.865 24.565 48.210 25.000 ;
        RECT 48.385 24.565 49.595 25.655 ;
        RECT 49.765 24.565 50.025 25.705 ;
        RECT 50.195 24.735 50.525 25.715 ;
        RECT 50.695 24.565 50.975 25.705 ;
        RECT 51.180 25.355 51.495 26.375 ;
        RECT 51.665 25.705 51.835 26.205 ;
        RECT 52.085 25.875 52.350 26.435 ;
        RECT 52.520 25.705 52.690 26.605 ;
        RECT 52.860 25.875 53.215 26.435 ;
        RECT 53.905 26.295 54.165 27.115 ;
        RECT 54.335 26.295 54.665 26.715 ;
        RECT 54.845 26.545 55.105 26.945 ;
        RECT 55.275 26.715 55.605 27.115 ;
        RECT 55.775 26.545 55.945 26.895 ;
        RECT 56.115 26.715 56.490 27.115 ;
        RECT 54.845 26.375 56.510 26.545 ;
        RECT 56.680 26.440 56.955 26.785 ;
        RECT 54.415 26.205 54.665 26.295 ;
        RECT 56.340 26.205 56.510 26.375 ;
        RECT 53.910 25.875 54.245 26.125 ;
        RECT 54.415 25.875 55.130 26.205 ;
        RECT 55.345 25.875 56.170 26.205 ;
        RECT 56.340 25.875 56.615 26.205 ;
        RECT 51.665 25.535 53.090 25.705 ;
        RECT 51.180 24.735 51.715 25.355 ;
        RECT 51.885 24.565 52.215 25.365 ;
        RECT 52.700 25.360 53.090 25.535 ;
        RECT 53.905 24.565 54.165 25.705 ;
        RECT 54.415 25.315 54.585 25.875 ;
        RECT 54.845 25.415 55.175 25.705 ;
        RECT 55.345 25.585 55.590 25.875 ;
        RECT 56.340 25.705 56.510 25.875 ;
        RECT 56.785 25.705 56.955 26.440 ;
        RECT 57.125 26.390 57.415 27.115 ;
        RECT 58.050 26.375 58.305 26.945 ;
        RECT 58.475 26.715 58.805 27.115 ;
        RECT 59.230 26.580 59.760 26.945 ;
        RECT 59.950 26.775 60.225 26.945 ;
        RECT 59.945 26.605 60.225 26.775 ;
        RECT 59.230 26.545 59.405 26.580 ;
        RECT 58.475 26.375 59.405 26.545 ;
        RECT 55.850 25.535 56.510 25.705 ;
        RECT 55.850 25.415 56.020 25.535 ;
        RECT 54.845 25.245 56.020 25.415 ;
        RECT 54.405 24.745 56.020 25.075 ;
        RECT 56.190 24.565 56.470 25.365 ;
        RECT 56.680 24.735 56.955 25.705 ;
        RECT 57.125 24.565 57.415 25.730 ;
        RECT 58.050 25.705 58.220 26.375 ;
        RECT 58.475 26.205 58.645 26.375 ;
        RECT 58.390 25.875 58.645 26.205 ;
        RECT 58.870 25.875 59.065 26.205 ;
        RECT 58.050 24.735 58.385 25.705 ;
        RECT 58.555 24.565 58.725 25.705 ;
        RECT 58.895 24.905 59.065 25.875 ;
        RECT 59.235 25.245 59.405 26.375 ;
        RECT 59.575 25.585 59.745 26.385 ;
        RECT 59.950 25.785 60.225 26.605 ;
        RECT 60.395 25.585 60.585 26.945 ;
        RECT 60.765 26.580 61.275 27.115 ;
        RECT 61.495 26.305 61.740 26.910 ;
        RECT 62.190 26.375 62.445 26.945 ;
        RECT 62.615 26.715 62.945 27.115 ;
        RECT 63.370 26.580 63.900 26.945 ;
        RECT 64.090 26.775 64.365 26.945 ;
        RECT 64.085 26.605 64.365 26.775 ;
        RECT 63.370 26.545 63.545 26.580 ;
        RECT 62.615 26.375 63.545 26.545 ;
        RECT 60.785 26.135 62.015 26.305 ;
        RECT 59.575 25.415 60.585 25.585 ;
        RECT 60.755 25.570 61.505 25.760 ;
        RECT 59.235 25.075 60.360 25.245 ;
        RECT 60.755 24.905 60.925 25.570 ;
        RECT 61.675 25.325 62.015 26.135 ;
        RECT 58.895 24.735 60.925 24.905 ;
        RECT 61.095 24.565 61.265 25.325 ;
        RECT 61.500 24.915 62.015 25.325 ;
        RECT 62.190 25.705 62.360 26.375 ;
        RECT 62.615 26.205 62.785 26.375 ;
        RECT 62.530 25.875 62.785 26.205 ;
        RECT 63.010 25.875 63.205 26.205 ;
        RECT 62.190 24.735 62.525 25.705 ;
        RECT 62.695 24.565 62.865 25.705 ;
        RECT 63.035 24.905 63.205 25.875 ;
        RECT 63.375 25.245 63.545 26.375 ;
        RECT 63.715 25.585 63.885 26.385 ;
        RECT 64.090 25.785 64.365 26.605 ;
        RECT 64.535 25.585 64.725 26.945 ;
        RECT 64.905 26.580 65.415 27.115 ;
        RECT 65.635 26.305 65.880 26.910 ;
        RECT 66.325 26.315 66.665 26.945 ;
        RECT 66.835 26.315 67.085 27.115 ;
        RECT 67.275 26.465 67.605 26.945 ;
        RECT 67.775 26.655 68.000 27.115 ;
        RECT 68.170 26.465 68.500 26.945 ;
        RECT 64.925 26.135 66.155 26.305 ;
        RECT 63.715 25.415 64.725 25.585 ;
        RECT 64.895 25.570 65.645 25.760 ;
        RECT 63.375 25.075 64.500 25.245 ;
        RECT 64.895 24.905 65.065 25.570 ;
        RECT 65.815 25.325 66.155 26.135 ;
        RECT 63.035 24.735 65.065 24.905 ;
        RECT 65.235 24.565 65.405 25.325 ;
        RECT 65.640 24.915 66.155 25.325 ;
        RECT 66.325 25.705 66.500 26.315 ;
        RECT 67.275 26.295 68.500 26.465 ;
        RECT 69.130 26.335 69.630 26.945 ;
        RECT 70.005 26.375 70.390 26.945 ;
        RECT 70.560 26.655 70.885 27.115 ;
        RECT 71.405 26.485 71.685 26.945 ;
        RECT 66.670 25.955 67.365 26.125 ;
        RECT 67.195 25.705 67.365 25.955 ;
        RECT 67.540 25.925 67.960 26.125 ;
        RECT 68.130 25.925 68.460 26.125 ;
        RECT 68.630 25.925 68.960 26.125 ;
        RECT 69.130 25.705 69.300 26.335 ;
        RECT 69.485 25.875 69.835 26.125 ;
        RECT 70.005 25.705 70.285 26.375 ;
        RECT 70.560 26.315 71.685 26.485 ;
        RECT 70.560 26.205 71.010 26.315 ;
        RECT 70.455 25.875 71.010 26.205 ;
        RECT 71.875 26.145 72.275 26.945 ;
        RECT 72.675 26.655 72.945 27.115 ;
        RECT 73.115 26.485 73.400 26.945 ;
        RECT 66.325 24.735 66.665 25.705 ;
        RECT 66.835 24.565 67.005 25.705 ;
        RECT 67.195 25.535 69.630 25.705 ;
        RECT 67.275 24.565 67.525 25.365 ;
        RECT 68.170 24.735 68.500 25.535 ;
        RECT 68.800 24.565 69.130 25.365 ;
        RECT 69.300 24.735 69.630 25.535 ;
        RECT 70.005 24.735 70.390 25.705 ;
        RECT 70.560 25.415 71.010 25.875 ;
        RECT 71.180 25.585 72.275 26.145 ;
        RECT 70.560 25.195 71.685 25.415 ;
        RECT 70.560 24.565 70.885 25.025 ;
        RECT 71.405 24.735 71.685 25.195 ;
        RECT 71.875 24.735 72.275 25.585 ;
        RECT 72.445 26.315 73.400 26.485 ;
        RECT 73.685 26.315 74.025 26.945 ;
        RECT 74.195 26.315 74.445 27.115 ;
        RECT 74.635 26.465 74.965 26.945 ;
        RECT 75.135 26.655 75.360 27.115 ;
        RECT 75.530 26.465 75.860 26.945 ;
        RECT 72.445 25.415 72.655 26.315 ;
        RECT 72.825 25.585 73.515 26.145 ;
        RECT 73.685 25.705 73.860 26.315 ;
        RECT 74.635 26.295 75.860 26.465 ;
        RECT 76.490 26.335 76.990 26.945 ;
        RECT 74.030 25.955 74.725 26.125 ;
        RECT 74.555 25.705 74.725 25.955 ;
        RECT 74.900 25.925 75.320 26.125 ;
        RECT 75.490 25.925 75.820 26.125 ;
        RECT 75.990 25.925 76.320 26.125 ;
        RECT 76.490 25.705 76.660 26.335 ;
        RECT 77.365 26.315 77.705 26.945 ;
        RECT 77.875 26.315 78.125 27.115 ;
        RECT 78.315 26.465 78.645 26.945 ;
        RECT 78.815 26.655 79.040 27.115 ;
        RECT 79.210 26.465 79.540 26.945 ;
        RECT 76.845 25.875 77.195 26.125 ;
        RECT 77.365 25.705 77.540 26.315 ;
        RECT 78.315 26.295 79.540 26.465 ;
        RECT 80.170 26.335 80.670 26.945 ;
        RECT 81.965 26.365 83.175 27.115 ;
        RECT 77.710 25.955 78.405 26.125 ;
        RECT 78.235 25.705 78.405 25.955 ;
        RECT 78.580 25.925 79.000 26.125 ;
        RECT 79.170 25.925 79.500 26.125 ;
        RECT 79.670 25.925 80.000 26.125 ;
        RECT 80.170 25.705 80.340 26.335 ;
        RECT 80.525 25.875 80.875 26.125 ;
        RECT 72.445 25.195 73.400 25.415 ;
        RECT 72.675 24.565 72.945 25.025 ;
        RECT 73.115 24.735 73.400 25.195 ;
        RECT 73.685 24.735 74.025 25.705 ;
        RECT 74.195 24.565 74.365 25.705 ;
        RECT 74.555 25.535 76.990 25.705 ;
        RECT 74.635 24.565 74.885 25.365 ;
        RECT 75.530 24.735 75.860 25.535 ;
        RECT 76.160 24.565 76.490 25.365 ;
        RECT 76.660 24.735 76.990 25.535 ;
        RECT 77.365 24.735 77.705 25.705 ;
        RECT 77.875 24.565 78.045 25.705 ;
        RECT 78.235 25.535 80.670 25.705 ;
        RECT 78.315 24.565 78.565 25.365 ;
        RECT 79.210 24.735 79.540 25.535 ;
        RECT 79.840 24.565 80.170 25.365 ;
        RECT 80.340 24.735 80.670 25.535 ;
        RECT 81.965 25.655 82.485 26.195 ;
        RECT 82.655 25.825 83.175 26.365 ;
        RECT 81.965 24.565 83.175 25.655 ;
        RECT 5.520 24.395 83.260 24.565 ;
        RECT 5.605 23.305 6.815 24.395 ;
        RECT 6.985 23.960 12.330 24.395 ;
        RECT 12.505 23.960 17.850 24.395 ;
        RECT 5.605 22.595 6.125 23.135 ;
        RECT 6.295 22.765 6.815 23.305 ;
        RECT 5.605 21.845 6.815 22.595 ;
        RECT 8.570 22.390 8.910 23.220 ;
        RECT 10.390 22.710 10.740 23.960 ;
        RECT 14.090 22.390 14.430 23.220 ;
        RECT 15.910 22.710 16.260 23.960 ;
        RECT 18.485 23.230 18.775 24.395 ;
        RECT 18.945 23.960 24.290 24.395 ;
        RECT 24.465 23.960 29.810 24.395 ;
        RECT 29.985 23.960 35.330 24.395 ;
        RECT 35.505 23.960 40.850 24.395 ;
        RECT 6.985 21.845 12.330 22.390 ;
        RECT 12.505 21.845 17.850 22.390 ;
        RECT 18.485 21.845 18.775 22.570 ;
        RECT 20.530 22.390 20.870 23.220 ;
        RECT 22.350 22.710 22.700 23.960 ;
        RECT 26.050 22.390 26.390 23.220 ;
        RECT 27.870 22.710 28.220 23.960 ;
        RECT 31.570 22.390 31.910 23.220 ;
        RECT 33.390 22.710 33.740 23.960 ;
        RECT 37.090 22.390 37.430 23.220 ;
        RECT 38.910 22.710 39.260 23.960 ;
        RECT 41.025 23.305 43.615 24.395 ;
        RECT 41.025 22.615 42.235 23.135 ;
        RECT 42.405 22.785 43.615 23.305 ;
        RECT 44.245 23.230 44.535 24.395 ;
        RECT 44.710 23.255 45.030 24.395 ;
        RECT 45.210 23.085 45.405 24.135 ;
        RECT 45.585 23.545 45.915 24.225 ;
        RECT 46.115 23.595 46.370 24.395 ;
        RECT 46.745 23.725 47.025 24.395 ;
        RECT 45.585 23.265 45.935 23.545 ;
        RECT 47.195 23.505 47.495 24.055 ;
        RECT 47.695 23.675 48.025 24.395 ;
        RECT 48.215 23.675 48.675 24.225 ;
        RECT 44.770 23.035 45.030 23.085 ;
        RECT 44.765 22.865 45.030 23.035 ;
        RECT 44.770 22.755 45.030 22.865 ;
        RECT 45.210 22.755 45.595 23.085 ;
        RECT 45.765 22.885 45.935 23.265 ;
        RECT 46.125 23.055 46.370 23.415 ;
        RECT 46.560 23.085 46.825 23.445 ;
        RECT 47.195 23.335 48.135 23.505 ;
        RECT 47.965 23.085 48.135 23.335 ;
        RECT 45.765 22.715 46.285 22.885 ;
        RECT 46.560 22.835 47.235 23.085 ;
        RECT 47.455 22.835 47.795 23.085 ;
        RECT 18.945 21.845 24.290 22.390 ;
        RECT 24.465 21.845 29.810 22.390 ;
        RECT 29.985 21.845 35.330 22.390 ;
        RECT 35.505 21.845 40.850 22.390 ;
        RECT 41.025 21.845 43.615 22.615 ;
        RECT 44.245 21.845 44.535 22.570 ;
        RECT 44.710 22.375 45.925 22.545 ;
        RECT 44.710 22.025 45.000 22.375 ;
        RECT 45.195 21.845 45.525 22.205 ;
        RECT 45.695 22.070 45.925 22.375 ;
        RECT 46.115 22.355 46.285 22.715 ;
        RECT 47.965 22.755 48.255 23.085 ;
        RECT 47.965 22.665 48.135 22.755 ;
        RECT 46.745 22.475 48.135 22.665 ;
        RECT 46.115 22.185 46.315 22.355 ;
        RECT 46.115 22.150 46.285 22.185 ;
        RECT 46.745 22.115 47.075 22.475 ;
        RECT 48.425 22.305 48.675 23.675 ;
        RECT 48.935 23.725 49.105 24.225 ;
        RECT 49.275 23.895 49.605 24.395 ;
        RECT 48.935 23.555 49.600 23.725 ;
        RECT 48.850 22.735 49.200 23.385 ;
        RECT 49.370 22.565 49.600 23.555 ;
        RECT 47.695 21.845 47.945 22.305 ;
        RECT 48.115 22.015 48.675 22.305 ;
        RECT 48.935 22.395 49.600 22.565 ;
        RECT 48.935 22.105 49.105 22.395 ;
        RECT 49.275 21.845 49.605 22.225 ;
        RECT 49.775 22.105 49.960 24.225 ;
        RECT 50.200 23.935 50.465 24.395 ;
        RECT 50.635 23.800 50.885 24.225 ;
        RECT 51.095 23.950 52.200 24.120 ;
        RECT 50.580 23.670 50.885 23.800 ;
        RECT 50.130 22.475 50.410 23.425 ;
        RECT 50.580 22.565 50.750 23.670 ;
        RECT 50.920 22.885 51.160 23.480 ;
        RECT 51.330 23.415 51.860 23.780 ;
        RECT 51.330 22.715 51.500 23.415 ;
        RECT 52.030 23.335 52.200 23.950 ;
        RECT 52.370 23.595 52.540 24.395 ;
        RECT 52.710 23.895 52.960 24.225 ;
        RECT 53.185 23.925 54.070 24.095 ;
        RECT 52.030 23.245 52.540 23.335 ;
        RECT 50.580 22.435 50.805 22.565 ;
        RECT 50.975 22.495 51.500 22.715 ;
        RECT 51.670 23.075 52.540 23.245 ;
        RECT 50.215 21.845 50.465 22.305 ;
        RECT 50.635 22.295 50.805 22.435 ;
        RECT 51.670 22.295 51.840 23.075 ;
        RECT 52.370 23.005 52.540 23.075 ;
        RECT 52.050 22.825 52.250 22.855 ;
        RECT 52.710 22.825 52.880 23.895 ;
        RECT 53.050 23.005 53.240 23.725 ;
        RECT 52.050 22.525 52.880 22.825 ;
        RECT 53.410 22.795 53.730 23.755 ;
        RECT 50.635 22.125 50.970 22.295 ;
        RECT 51.165 22.125 51.840 22.295 ;
        RECT 52.160 21.845 52.530 22.345 ;
        RECT 52.710 22.295 52.880 22.525 ;
        RECT 53.265 22.465 53.730 22.795 ;
        RECT 53.900 23.085 54.070 23.925 ;
        RECT 54.250 23.895 54.565 24.395 ;
        RECT 54.795 23.665 55.135 24.225 ;
        RECT 54.240 23.290 55.135 23.665 ;
        RECT 55.305 23.385 55.475 24.395 ;
        RECT 54.945 23.085 55.135 23.290 ;
        RECT 55.645 23.335 55.975 24.180 ;
        RECT 57.215 23.725 57.385 24.225 ;
        RECT 57.555 23.895 57.885 24.395 ;
        RECT 57.215 23.555 57.880 23.725 ;
        RECT 55.645 23.255 56.035 23.335 ;
        RECT 55.820 23.205 56.035 23.255 ;
        RECT 53.900 22.755 54.775 23.085 ;
        RECT 54.945 22.755 55.695 23.085 ;
        RECT 53.900 22.295 54.070 22.755 ;
        RECT 54.945 22.585 55.145 22.755 ;
        RECT 55.865 22.625 56.035 23.205 ;
        RECT 57.130 22.735 57.480 23.385 ;
        RECT 55.810 22.585 56.035 22.625 ;
        RECT 52.710 22.125 53.115 22.295 ;
        RECT 53.285 22.125 54.070 22.295 ;
        RECT 54.345 21.845 54.555 22.375 ;
        RECT 54.815 22.060 55.145 22.585 ;
        RECT 55.655 22.500 56.035 22.585 ;
        RECT 57.650 22.565 57.880 23.555 ;
        RECT 55.315 21.845 55.485 22.455 ;
        RECT 55.655 22.065 55.985 22.500 ;
        RECT 57.215 22.395 57.880 22.565 ;
        RECT 57.215 22.105 57.385 22.395 ;
        RECT 57.555 21.845 57.885 22.225 ;
        RECT 58.055 22.105 58.240 24.225 ;
        RECT 58.480 23.935 58.745 24.395 ;
        RECT 58.915 23.800 59.165 24.225 ;
        RECT 59.375 23.950 60.480 24.120 ;
        RECT 58.860 23.670 59.165 23.800 ;
        RECT 58.410 22.475 58.690 23.425 ;
        RECT 58.860 22.565 59.030 23.670 ;
        RECT 59.200 22.885 59.440 23.480 ;
        RECT 59.610 23.415 60.140 23.780 ;
        RECT 59.610 22.715 59.780 23.415 ;
        RECT 60.310 23.335 60.480 23.950 ;
        RECT 60.650 23.595 60.820 24.395 ;
        RECT 60.990 23.895 61.240 24.225 ;
        RECT 61.465 23.925 62.350 24.095 ;
        RECT 60.310 23.245 60.820 23.335 ;
        RECT 58.860 22.435 59.085 22.565 ;
        RECT 59.255 22.495 59.780 22.715 ;
        RECT 59.950 23.075 60.820 23.245 ;
        RECT 58.495 21.845 58.745 22.305 ;
        RECT 58.915 22.295 59.085 22.435 ;
        RECT 59.950 22.295 60.120 23.075 ;
        RECT 60.650 23.005 60.820 23.075 ;
        RECT 60.330 22.825 60.530 22.855 ;
        RECT 60.990 22.825 61.160 23.895 ;
        RECT 61.330 23.005 61.520 23.725 ;
        RECT 60.330 22.525 61.160 22.825 ;
        RECT 61.690 22.795 62.010 23.755 ;
        RECT 58.915 22.125 59.250 22.295 ;
        RECT 59.445 22.125 60.120 22.295 ;
        RECT 60.440 21.845 60.810 22.345 ;
        RECT 60.990 22.295 61.160 22.525 ;
        RECT 61.545 22.465 62.010 22.795 ;
        RECT 62.180 23.085 62.350 23.925 ;
        RECT 62.530 23.895 62.845 24.395 ;
        RECT 63.075 23.665 63.415 24.225 ;
        RECT 62.520 23.290 63.415 23.665 ;
        RECT 63.585 23.385 63.755 24.395 ;
        RECT 63.225 23.085 63.415 23.290 ;
        RECT 63.925 23.335 64.255 24.180 ;
        RECT 64.425 23.480 64.595 24.395 ;
        RECT 63.925 23.255 64.315 23.335 ;
        RECT 64.100 23.205 64.315 23.255 ;
        RECT 62.180 22.755 63.055 23.085 ;
        RECT 63.225 22.755 63.975 23.085 ;
        RECT 62.180 22.295 62.350 22.755 ;
        RECT 63.225 22.585 63.425 22.755 ;
        RECT 64.145 22.625 64.315 23.205 ;
        RECT 64.090 22.585 64.315 22.625 ;
        RECT 60.990 22.125 61.395 22.295 ;
        RECT 61.565 22.125 62.350 22.295 ;
        RECT 62.625 21.845 62.835 22.375 ;
        RECT 63.095 22.060 63.425 22.585 ;
        RECT 63.935 22.500 64.315 22.585 ;
        RECT 64.950 23.255 65.285 24.225 ;
        RECT 65.455 23.255 65.625 24.395 ;
        RECT 65.795 24.055 67.825 24.225 ;
        RECT 64.950 22.585 65.120 23.255 ;
        RECT 65.795 23.085 65.965 24.055 ;
        RECT 65.290 22.755 65.545 23.085 ;
        RECT 65.770 22.755 65.965 23.085 ;
        RECT 66.135 23.715 67.260 23.885 ;
        RECT 65.375 22.585 65.545 22.755 ;
        RECT 66.135 22.585 66.305 23.715 ;
        RECT 63.595 21.845 63.765 22.455 ;
        RECT 63.935 22.065 64.265 22.500 ;
        RECT 64.435 21.845 64.605 22.360 ;
        RECT 64.950 22.015 65.205 22.585 ;
        RECT 65.375 22.415 66.305 22.585 ;
        RECT 66.475 23.375 67.485 23.545 ;
        RECT 66.475 22.575 66.645 23.375 ;
        RECT 66.850 22.695 67.125 23.175 ;
        RECT 66.845 22.525 67.125 22.695 ;
        RECT 66.130 22.380 66.305 22.415 ;
        RECT 65.375 21.845 65.705 22.245 ;
        RECT 66.130 22.015 66.660 22.380 ;
        RECT 66.850 22.015 67.125 22.525 ;
        RECT 67.295 22.015 67.485 23.375 ;
        RECT 67.655 23.390 67.825 24.055 ;
        RECT 67.995 23.635 68.165 24.395 ;
        RECT 68.400 23.635 68.915 24.045 ;
        RECT 67.655 23.200 68.405 23.390 ;
        RECT 68.575 22.825 68.915 23.635 ;
        RECT 70.005 23.230 70.295 24.395 ;
        RECT 70.525 23.335 70.855 24.180 ;
        RECT 71.025 23.385 71.195 24.395 ;
        RECT 71.365 23.665 71.705 24.225 ;
        RECT 71.935 23.895 72.250 24.395 ;
        RECT 72.430 23.925 73.315 24.095 ;
        RECT 70.465 23.255 70.855 23.335 ;
        RECT 71.365 23.290 72.260 23.665 ;
        RECT 67.685 22.655 68.915 22.825 ;
        RECT 70.465 23.205 70.680 23.255 ;
        RECT 67.665 21.845 68.175 22.380 ;
        RECT 68.395 22.050 68.640 22.655 ;
        RECT 70.465 22.625 70.635 23.205 ;
        RECT 71.365 23.085 71.555 23.290 ;
        RECT 72.430 23.085 72.600 23.925 ;
        RECT 73.540 23.895 73.790 24.225 ;
        RECT 70.805 22.755 71.555 23.085 ;
        RECT 71.725 22.755 72.600 23.085 ;
        RECT 70.465 22.585 70.690 22.625 ;
        RECT 71.355 22.585 71.555 22.755 ;
        RECT 70.005 21.845 70.295 22.570 ;
        RECT 70.465 22.500 70.845 22.585 ;
        RECT 70.515 22.065 70.845 22.500 ;
        RECT 71.015 21.845 71.185 22.455 ;
        RECT 71.355 22.060 71.685 22.585 ;
        RECT 71.945 21.845 72.155 22.375 ;
        RECT 72.430 22.295 72.600 22.755 ;
        RECT 72.770 22.795 73.090 23.755 ;
        RECT 73.260 23.005 73.450 23.725 ;
        RECT 73.620 22.825 73.790 23.895 ;
        RECT 73.960 23.595 74.130 24.395 ;
        RECT 74.300 23.950 75.405 24.120 ;
        RECT 74.300 23.335 74.470 23.950 ;
        RECT 75.615 23.800 75.865 24.225 ;
        RECT 76.035 23.935 76.300 24.395 ;
        RECT 74.640 23.415 75.170 23.780 ;
        RECT 75.615 23.670 75.920 23.800 ;
        RECT 73.960 23.245 74.470 23.335 ;
        RECT 73.960 23.075 74.830 23.245 ;
        RECT 73.960 23.005 74.130 23.075 ;
        RECT 74.250 22.825 74.450 22.855 ;
        RECT 72.770 22.465 73.235 22.795 ;
        RECT 73.620 22.525 74.450 22.825 ;
        RECT 73.620 22.295 73.790 22.525 ;
        RECT 72.430 22.125 73.215 22.295 ;
        RECT 73.385 22.125 73.790 22.295 ;
        RECT 73.970 21.845 74.340 22.345 ;
        RECT 74.660 22.295 74.830 23.075 ;
        RECT 75.000 22.715 75.170 23.415 ;
        RECT 75.340 22.885 75.580 23.480 ;
        RECT 75.000 22.495 75.525 22.715 ;
        RECT 75.750 22.565 75.920 23.670 ;
        RECT 75.695 22.435 75.920 22.565 ;
        RECT 76.090 22.475 76.370 23.425 ;
        RECT 75.695 22.295 75.865 22.435 ;
        RECT 74.660 22.125 75.335 22.295 ;
        RECT 75.530 22.125 75.865 22.295 ;
        RECT 76.035 21.845 76.285 22.305 ;
        RECT 76.540 22.105 76.725 24.225 ;
        RECT 76.895 23.895 77.225 24.395 ;
        RECT 77.395 23.725 77.565 24.225 ;
        RECT 76.900 23.555 77.565 23.725 ;
        RECT 76.900 22.565 77.130 23.555 ;
        RECT 77.300 22.735 77.650 23.385 ;
        RECT 77.825 23.255 78.165 24.225 ;
        RECT 78.335 23.255 78.505 24.395 ;
        RECT 78.775 23.595 79.025 24.395 ;
        RECT 79.670 23.425 80.000 24.225 ;
        RECT 80.300 23.595 80.630 24.395 ;
        RECT 80.800 23.425 81.130 24.225 ;
        RECT 78.695 23.255 81.130 23.425 ;
        RECT 81.965 23.305 83.175 24.395 ;
        RECT 77.825 22.645 78.000 23.255 ;
        RECT 78.695 23.005 78.865 23.255 ;
        RECT 78.170 22.835 78.865 23.005 ;
        RECT 79.040 22.835 79.460 23.035 ;
        RECT 79.630 22.835 79.960 23.035 ;
        RECT 80.130 22.835 80.460 23.035 ;
        RECT 76.900 22.395 77.565 22.565 ;
        RECT 76.895 21.845 77.225 22.225 ;
        RECT 77.395 22.105 77.565 22.395 ;
        RECT 77.825 22.015 78.165 22.645 ;
        RECT 78.335 21.845 78.585 22.645 ;
        RECT 78.775 22.495 80.000 22.665 ;
        RECT 78.775 22.015 79.105 22.495 ;
        RECT 79.275 21.845 79.500 22.305 ;
        RECT 79.670 22.015 80.000 22.495 ;
        RECT 80.630 22.625 80.800 23.255 ;
        RECT 80.985 22.835 81.335 23.085 ;
        RECT 81.965 22.765 82.485 23.305 ;
        RECT 80.630 22.015 81.130 22.625 ;
        RECT 82.655 22.595 83.175 23.135 ;
        RECT 81.965 21.845 83.175 22.595 ;
        RECT 5.520 21.675 83.260 21.845 ;
        RECT 5.605 20.925 6.815 21.675 ;
        RECT 6.985 21.130 12.330 21.675 ;
        RECT 12.505 21.130 17.850 21.675 ;
        RECT 18.025 21.130 23.370 21.675 ;
        RECT 23.545 21.130 28.890 21.675 ;
        RECT 5.605 20.385 6.125 20.925 ;
        RECT 6.295 20.215 6.815 20.755 ;
        RECT 8.570 20.300 8.910 21.130 ;
        RECT 5.605 19.125 6.815 20.215 ;
        RECT 10.390 19.560 10.740 20.810 ;
        RECT 14.090 20.300 14.430 21.130 ;
        RECT 15.910 19.560 16.260 20.810 ;
        RECT 19.610 20.300 19.950 21.130 ;
        RECT 21.430 19.560 21.780 20.810 ;
        RECT 25.130 20.300 25.470 21.130 ;
        RECT 29.065 20.905 30.735 21.675 ;
        RECT 31.365 20.950 31.655 21.675 ;
        RECT 31.825 21.130 37.170 21.675 ;
        RECT 26.950 19.560 27.300 20.810 ;
        RECT 29.065 20.385 29.815 20.905 ;
        RECT 29.985 20.215 30.735 20.735 ;
        RECT 33.410 20.300 33.750 21.130 ;
        RECT 37.345 20.905 39.935 21.675 ;
        RECT 40.140 20.935 40.755 21.505 ;
        RECT 40.925 21.165 41.140 21.675 ;
        RECT 41.370 21.165 41.650 21.495 ;
        RECT 41.830 21.165 42.070 21.675 ;
        RECT 42.405 21.215 42.965 21.505 ;
        RECT 43.135 21.215 43.385 21.675 ;
        RECT 6.985 19.125 12.330 19.560 ;
        RECT 12.505 19.125 17.850 19.560 ;
        RECT 18.025 19.125 23.370 19.560 ;
        RECT 23.545 19.125 28.890 19.560 ;
        RECT 29.065 19.125 30.735 20.215 ;
        RECT 31.365 19.125 31.655 20.290 ;
        RECT 35.230 19.560 35.580 20.810 ;
        RECT 37.345 20.385 38.555 20.905 ;
        RECT 38.725 20.215 39.935 20.735 ;
        RECT 31.825 19.125 37.170 19.560 ;
        RECT 37.345 19.125 39.935 20.215 ;
        RECT 40.140 19.915 40.455 20.935 ;
        RECT 40.625 20.265 40.795 20.765 ;
        RECT 41.045 20.435 41.310 20.995 ;
        RECT 41.480 20.265 41.650 21.165 ;
        RECT 41.820 20.435 42.175 20.995 ;
        RECT 40.625 20.095 42.050 20.265 ;
        RECT 40.140 19.295 40.675 19.915 ;
        RECT 40.845 19.125 41.175 19.925 ;
        RECT 41.660 19.920 42.050 20.095 ;
        RECT 42.405 19.845 42.655 21.215 ;
        RECT 44.005 21.045 44.335 21.405 ;
        RECT 42.945 20.855 44.335 21.045 ;
        RECT 44.710 21.200 45.045 21.460 ;
        RECT 45.215 21.275 45.545 21.675 ;
        RECT 45.715 21.275 47.330 21.445 ;
        RECT 42.945 20.765 43.115 20.855 ;
        RECT 42.825 20.435 43.115 20.765 ;
        RECT 43.285 20.435 43.625 20.685 ;
        RECT 43.845 20.435 44.520 20.685 ;
        RECT 42.945 20.185 43.115 20.435 ;
        RECT 42.945 20.015 43.885 20.185 ;
        RECT 44.255 20.075 44.520 20.435 ;
        RECT 42.405 19.295 42.865 19.845 ;
        RECT 43.055 19.125 43.385 19.845 ;
        RECT 43.585 19.465 43.885 20.015 ;
        RECT 44.710 19.845 44.965 21.200 ;
        RECT 45.715 21.105 45.885 21.275 ;
        RECT 45.325 20.935 45.885 21.105 ;
        RECT 46.150 20.995 46.420 21.095 ;
        RECT 46.610 20.995 46.900 21.095 ;
        RECT 45.325 20.765 45.495 20.935 ;
        RECT 46.145 20.825 46.420 20.995 ;
        RECT 46.605 20.825 46.900 20.995 ;
        RECT 45.190 20.435 45.495 20.765 ;
        RECT 45.690 20.655 45.940 20.765 ;
        RECT 45.685 20.485 45.940 20.655 ;
        RECT 45.690 20.435 45.940 20.485 ;
        RECT 46.150 20.435 46.420 20.825 ;
        RECT 46.610 20.435 46.900 20.825 ;
        RECT 47.070 20.435 47.490 21.100 ;
        RECT 47.875 20.955 48.205 21.675 ;
        RECT 49.395 21.125 49.565 21.415 ;
        RECT 49.735 21.295 50.065 21.675 ;
        RECT 49.395 20.955 50.060 21.125 ;
        RECT 47.800 20.655 48.150 20.765 ;
        RECT 47.800 20.485 48.155 20.655 ;
        RECT 47.800 20.435 48.150 20.485 ;
        RECT 45.325 20.265 45.495 20.435 ;
        RECT 45.325 20.095 47.695 20.265 ;
        RECT 47.945 20.145 48.150 20.435 ;
        RECT 49.310 20.135 49.660 20.785 ;
        RECT 44.055 19.125 44.335 19.795 ;
        RECT 44.710 19.335 45.045 19.845 ;
        RECT 45.295 19.125 45.625 19.925 ;
        RECT 45.870 19.715 47.295 19.885 ;
        RECT 45.870 19.295 46.155 19.715 ;
        RECT 46.410 19.125 46.740 19.545 ;
        RECT 46.965 19.465 47.295 19.715 ;
        RECT 47.525 19.635 47.695 20.095 ;
        RECT 49.830 19.965 50.060 20.955 ;
        RECT 47.955 19.465 48.125 19.965 ;
        RECT 46.965 19.295 48.125 19.465 ;
        RECT 49.395 19.795 50.060 19.965 ;
        RECT 49.395 19.295 49.565 19.795 ;
        RECT 49.735 19.125 50.065 19.625 ;
        RECT 50.235 19.295 50.420 21.415 ;
        RECT 50.675 21.215 50.925 21.675 ;
        RECT 51.095 21.225 51.430 21.395 ;
        RECT 51.625 21.225 52.300 21.395 ;
        RECT 51.095 21.085 51.265 21.225 ;
        RECT 50.590 20.095 50.870 21.045 ;
        RECT 51.040 20.955 51.265 21.085 ;
        RECT 51.040 19.850 51.210 20.955 ;
        RECT 51.435 20.805 51.960 21.025 ;
        RECT 51.380 20.040 51.620 20.635 ;
        RECT 51.790 20.105 51.960 20.805 ;
        RECT 52.130 20.445 52.300 21.225 ;
        RECT 52.620 21.175 52.990 21.675 ;
        RECT 53.170 21.225 53.575 21.395 ;
        RECT 53.745 21.225 54.530 21.395 ;
        RECT 53.170 20.995 53.340 21.225 ;
        RECT 52.510 20.695 53.340 20.995 ;
        RECT 53.725 20.725 54.190 21.055 ;
        RECT 52.510 20.665 52.710 20.695 ;
        RECT 52.830 20.445 53.000 20.515 ;
        RECT 52.130 20.275 53.000 20.445 ;
        RECT 52.490 20.185 53.000 20.275 ;
        RECT 51.040 19.720 51.345 19.850 ;
        RECT 51.790 19.740 52.320 20.105 ;
        RECT 50.660 19.125 50.925 19.585 ;
        RECT 51.095 19.295 51.345 19.720 ;
        RECT 52.490 19.570 52.660 20.185 ;
        RECT 51.555 19.400 52.660 19.570 ;
        RECT 52.830 19.125 53.000 19.925 ;
        RECT 53.170 19.625 53.340 20.695 ;
        RECT 53.510 19.795 53.700 20.515 ;
        RECT 53.870 19.765 54.190 20.725 ;
        RECT 54.360 20.765 54.530 21.225 ;
        RECT 54.805 21.145 55.015 21.675 ;
        RECT 55.275 20.935 55.605 21.460 ;
        RECT 55.775 21.065 55.945 21.675 ;
        RECT 56.115 21.020 56.445 21.455 ;
        RECT 56.615 21.160 56.785 21.675 ;
        RECT 56.115 20.935 56.495 21.020 ;
        RECT 57.125 20.950 57.415 21.675 ;
        RECT 57.755 21.160 57.925 21.675 ;
        RECT 58.095 21.020 58.425 21.455 ;
        RECT 58.595 21.065 58.765 21.675 ;
        RECT 55.405 20.765 55.605 20.935 ;
        RECT 56.270 20.895 56.495 20.935 ;
        RECT 54.360 20.435 55.235 20.765 ;
        RECT 55.405 20.435 56.155 20.765 ;
        RECT 53.170 19.295 53.420 19.625 ;
        RECT 54.360 19.595 54.530 20.435 ;
        RECT 55.405 20.230 55.595 20.435 ;
        RECT 56.325 20.315 56.495 20.895 ;
        RECT 56.280 20.265 56.495 20.315 ;
        RECT 58.045 20.935 58.425 21.020 ;
        RECT 58.935 20.935 59.265 21.460 ;
        RECT 59.525 21.145 59.735 21.675 ;
        RECT 60.010 21.225 60.795 21.395 ;
        RECT 60.965 21.225 61.370 21.395 ;
        RECT 58.045 20.895 58.270 20.935 ;
        RECT 58.045 20.315 58.215 20.895 ;
        RECT 58.935 20.765 59.135 20.935 ;
        RECT 60.010 20.765 60.180 21.225 ;
        RECT 58.385 20.435 59.135 20.765 ;
        RECT 59.305 20.435 60.180 20.765 ;
        RECT 54.700 19.855 55.595 20.230 ;
        RECT 56.105 20.185 56.495 20.265 ;
        RECT 53.645 19.425 54.530 19.595 ;
        RECT 54.710 19.125 55.025 19.625 ;
        RECT 55.255 19.295 55.595 19.855 ;
        RECT 55.765 19.125 55.935 20.135 ;
        RECT 56.105 19.340 56.435 20.185 ;
        RECT 56.605 19.125 56.775 20.040 ;
        RECT 57.125 19.125 57.415 20.290 ;
        RECT 58.045 20.265 58.260 20.315 ;
        RECT 58.045 20.185 58.435 20.265 ;
        RECT 57.765 19.125 57.935 20.040 ;
        RECT 58.105 19.340 58.435 20.185 ;
        RECT 58.945 20.230 59.135 20.435 ;
        RECT 58.605 19.125 58.775 20.135 ;
        RECT 58.945 19.855 59.840 20.230 ;
        RECT 58.945 19.295 59.285 19.855 ;
        RECT 59.515 19.125 59.830 19.625 ;
        RECT 60.010 19.595 60.180 20.435 ;
        RECT 60.350 20.725 60.815 21.055 ;
        RECT 61.200 20.995 61.370 21.225 ;
        RECT 61.550 21.175 61.920 21.675 ;
        RECT 62.240 21.225 62.915 21.395 ;
        RECT 63.110 21.225 63.445 21.395 ;
        RECT 60.350 19.765 60.670 20.725 ;
        RECT 61.200 20.695 62.030 20.995 ;
        RECT 60.840 19.795 61.030 20.515 ;
        RECT 61.200 19.625 61.370 20.695 ;
        RECT 61.830 20.665 62.030 20.695 ;
        RECT 61.540 20.445 61.710 20.515 ;
        RECT 62.240 20.445 62.410 21.225 ;
        RECT 63.275 21.085 63.445 21.225 ;
        RECT 63.615 21.215 63.865 21.675 ;
        RECT 61.540 20.275 62.410 20.445 ;
        RECT 62.580 20.805 63.105 21.025 ;
        RECT 63.275 20.955 63.500 21.085 ;
        RECT 61.540 20.185 62.050 20.275 ;
        RECT 60.010 19.425 60.895 19.595 ;
        RECT 61.120 19.295 61.370 19.625 ;
        RECT 61.540 19.125 61.710 19.925 ;
        RECT 61.880 19.570 62.050 20.185 ;
        RECT 62.580 20.105 62.750 20.805 ;
        RECT 62.220 19.740 62.750 20.105 ;
        RECT 62.920 20.040 63.160 20.635 ;
        RECT 63.330 19.850 63.500 20.955 ;
        RECT 63.670 20.095 63.950 21.045 ;
        RECT 63.195 19.720 63.500 19.850 ;
        RECT 61.880 19.400 62.985 19.570 ;
        RECT 63.195 19.295 63.445 19.720 ;
        RECT 63.615 19.125 63.880 19.585 ;
        RECT 64.120 19.295 64.305 21.415 ;
        RECT 64.475 21.295 64.805 21.675 ;
        RECT 64.975 21.125 65.145 21.415 ;
        RECT 64.480 20.955 65.145 21.125 ;
        RECT 65.495 21.125 65.665 21.415 ;
        RECT 65.835 21.295 66.165 21.675 ;
        RECT 65.495 20.955 66.160 21.125 ;
        RECT 64.480 19.965 64.710 20.955 ;
        RECT 64.880 20.135 65.230 20.785 ;
        RECT 65.410 20.135 65.760 20.785 ;
        RECT 65.930 19.965 66.160 20.955 ;
        RECT 64.480 19.795 65.145 19.965 ;
        RECT 64.475 19.125 64.805 19.625 ;
        RECT 64.975 19.295 65.145 19.795 ;
        RECT 65.495 19.795 66.160 19.965 ;
        RECT 65.495 19.295 65.665 19.795 ;
        RECT 65.835 19.125 66.165 19.625 ;
        RECT 66.335 19.295 66.520 21.415 ;
        RECT 66.775 21.215 67.025 21.675 ;
        RECT 67.195 21.225 67.530 21.395 ;
        RECT 67.725 21.225 68.400 21.395 ;
        RECT 67.195 21.085 67.365 21.225 ;
        RECT 66.690 20.095 66.970 21.045 ;
        RECT 67.140 20.955 67.365 21.085 ;
        RECT 67.140 19.850 67.310 20.955 ;
        RECT 67.535 20.805 68.060 21.025 ;
        RECT 67.480 20.040 67.720 20.635 ;
        RECT 67.890 20.105 68.060 20.805 ;
        RECT 68.230 20.445 68.400 21.225 ;
        RECT 68.720 21.175 69.090 21.675 ;
        RECT 69.270 21.225 69.675 21.395 ;
        RECT 69.845 21.225 70.630 21.395 ;
        RECT 69.270 20.995 69.440 21.225 ;
        RECT 68.610 20.695 69.440 20.995 ;
        RECT 69.825 20.725 70.290 21.055 ;
        RECT 68.610 20.665 68.810 20.695 ;
        RECT 68.930 20.445 69.100 20.515 ;
        RECT 68.230 20.275 69.100 20.445 ;
        RECT 68.590 20.185 69.100 20.275 ;
        RECT 67.140 19.720 67.445 19.850 ;
        RECT 67.890 19.740 68.420 20.105 ;
        RECT 66.760 19.125 67.025 19.585 ;
        RECT 67.195 19.295 67.445 19.720 ;
        RECT 68.590 19.570 68.760 20.185 ;
        RECT 67.655 19.400 68.760 19.570 ;
        RECT 68.930 19.125 69.100 19.925 ;
        RECT 69.270 19.625 69.440 20.695 ;
        RECT 69.610 19.795 69.800 20.515 ;
        RECT 69.970 19.765 70.290 20.725 ;
        RECT 70.460 20.765 70.630 21.225 ;
        RECT 70.905 21.145 71.115 21.675 ;
        RECT 71.375 20.935 71.705 21.460 ;
        RECT 71.875 21.065 72.045 21.675 ;
        RECT 72.215 21.020 72.545 21.455 ;
        RECT 73.275 21.020 73.605 21.455 ;
        RECT 73.775 21.065 73.945 21.675 ;
        RECT 72.215 20.935 72.595 21.020 ;
        RECT 71.505 20.765 71.705 20.935 ;
        RECT 72.370 20.895 72.595 20.935 ;
        RECT 70.460 20.435 71.335 20.765 ;
        RECT 71.505 20.435 72.255 20.765 ;
        RECT 69.270 19.295 69.520 19.625 ;
        RECT 70.460 19.595 70.630 20.435 ;
        RECT 71.505 20.230 71.695 20.435 ;
        RECT 72.425 20.315 72.595 20.895 ;
        RECT 72.380 20.265 72.595 20.315 ;
        RECT 70.800 19.855 71.695 20.230 ;
        RECT 72.205 20.185 72.595 20.265 ;
        RECT 73.225 20.935 73.605 21.020 ;
        RECT 74.115 20.935 74.445 21.460 ;
        RECT 74.705 21.145 74.915 21.675 ;
        RECT 75.190 21.225 75.975 21.395 ;
        RECT 76.145 21.225 76.550 21.395 ;
        RECT 73.225 20.895 73.450 20.935 ;
        RECT 73.225 20.315 73.395 20.895 ;
        RECT 74.115 20.765 74.315 20.935 ;
        RECT 75.190 20.765 75.360 21.225 ;
        RECT 73.565 20.435 74.315 20.765 ;
        RECT 74.485 20.435 75.360 20.765 ;
        RECT 73.225 20.265 73.440 20.315 ;
        RECT 73.225 20.185 73.615 20.265 ;
        RECT 69.745 19.425 70.630 19.595 ;
        RECT 70.810 19.125 71.125 19.625 ;
        RECT 71.355 19.295 71.695 19.855 ;
        RECT 71.865 19.125 72.035 20.135 ;
        RECT 72.205 19.340 72.535 20.185 ;
        RECT 73.285 19.340 73.615 20.185 ;
        RECT 74.125 20.230 74.315 20.435 ;
        RECT 73.785 19.125 73.955 20.135 ;
        RECT 74.125 19.855 75.020 20.230 ;
        RECT 74.125 19.295 74.465 19.855 ;
        RECT 74.695 19.125 75.010 19.625 ;
        RECT 75.190 19.595 75.360 20.435 ;
        RECT 75.530 20.725 75.995 21.055 ;
        RECT 76.380 20.995 76.550 21.225 ;
        RECT 76.730 21.175 77.100 21.675 ;
        RECT 77.420 21.225 78.095 21.395 ;
        RECT 78.290 21.225 78.625 21.395 ;
        RECT 75.530 19.765 75.850 20.725 ;
        RECT 76.380 20.695 77.210 20.995 ;
        RECT 76.020 19.795 76.210 20.515 ;
        RECT 76.380 19.625 76.550 20.695 ;
        RECT 77.010 20.665 77.210 20.695 ;
        RECT 76.720 20.445 76.890 20.515 ;
        RECT 77.420 20.445 77.590 21.225 ;
        RECT 78.455 21.085 78.625 21.225 ;
        RECT 78.795 21.215 79.045 21.675 ;
        RECT 76.720 20.275 77.590 20.445 ;
        RECT 77.760 20.805 78.285 21.025 ;
        RECT 78.455 20.955 78.680 21.085 ;
        RECT 76.720 20.185 77.230 20.275 ;
        RECT 75.190 19.425 76.075 19.595 ;
        RECT 76.300 19.295 76.550 19.625 ;
        RECT 76.720 19.125 76.890 19.925 ;
        RECT 77.060 19.570 77.230 20.185 ;
        RECT 77.760 20.105 77.930 20.805 ;
        RECT 77.400 19.740 77.930 20.105 ;
        RECT 78.100 20.040 78.340 20.635 ;
        RECT 78.510 19.850 78.680 20.955 ;
        RECT 78.850 20.095 79.130 21.045 ;
        RECT 78.375 19.720 78.680 19.850 ;
        RECT 77.060 19.400 78.165 19.570 ;
        RECT 78.375 19.295 78.625 19.720 ;
        RECT 78.795 19.125 79.060 19.585 ;
        RECT 79.300 19.295 79.485 21.415 ;
        RECT 79.655 21.295 79.985 21.675 ;
        RECT 80.155 21.125 80.325 21.415 ;
        RECT 79.660 20.955 80.325 21.125 ;
        RECT 79.660 19.965 79.890 20.955 ;
        RECT 80.585 20.925 81.795 21.675 ;
        RECT 81.965 20.925 83.175 21.675 ;
        RECT 80.060 20.135 80.410 20.785 ;
        RECT 80.585 20.385 81.105 20.925 ;
        RECT 81.275 20.215 81.795 20.755 ;
        RECT 79.660 19.795 80.325 19.965 ;
        RECT 79.655 19.125 79.985 19.625 ;
        RECT 80.155 19.295 80.325 19.795 ;
        RECT 80.585 19.125 81.795 20.215 ;
        RECT 81.965 20.215 82.485 20.755 ;
        RECT 82.655 20.385 83.175 20.925 ;
        RECT 81.965 19.125 83.175 20.215 ;
        RECT 5.520 18.955 83.260 19.125 ;
        RECT 5.605 17.865 6.815 18.955 ;
        RECT 6.985 18.520 12.330 18.955 ;
        RECT 12.505 18.520 17.850 18.955 ;
        RECT 5.605 17.155 6.125 17.695 ;
        RECT 6.295 17.325 6.815 17.865 ;
        RECT 5.605 16.405 6.815 17.155 ;
        RECT 8.570 16.950 8.910 17.780 ;
        RECT 10.390 17.270 10.740 18.520 ;
        RECT 14.090 16.950 14.430 17.780 ;
        RECT 15.910 17.270 16.260 18.520 ;
        RECT 18.485 17.790 18.775 18.955 ;
        RECT 18.945 18.520 24.290 18.955 ;
        RECT 24.465 18.520 29.810 18.955 ;
        RECT 29.985 18.520 35.330 18.955 ;
        RECT 35.505 18.520 40.850 18.955 ;
        RECT 6.985 16.405 12.330 16.950 ;
        RECT 12.505 16.405 17.850 16.950 ;
        RECT 18.485 16.405 18.775 17.130 ;
        RECT 20.530 16.950 20.870 17.780 ;
        RECT 22.350 17.270 22.700 18.520 ;
        RECT 26.050 16.950 26.390 17.780 ;
        RECT 27.870 17.270 28.220 18.520 ;
        RECT 31.570 16.950 31.910 17.780 ;
        RECT 33.390 17.270 33.740 18.520 ;
        RECT 37.090 16.950 37.430 17.780 ;
        RECT 38.910 17.270 39.260 18.520 ;
        RECT 41.025 17.865 42.695 18.955 ;
        RECT 41.025 17.175 41.775 17.695 ;
        RECT 41.945 17.345 42.695 17.865 ;
        RECT 42.865 17.880 43.135 18.785 ;
        RECT 43.305 18.195 43.635 18.955 ;
        RECT 43.815 18.025 43.985 18.785 ;
        RECT 18.945 16.405 24.290 16.950 ;
        RECT 24.465 16.405 29.810 16.950 ;
        RECT 29.985 16.405 35.330 16.950 ;
        RECT 35.505 16.405 40.850 16.950 ;
        RECT 41.025 16.405 42.695 17.175 ;
        RECT 42.865 17.080 43.035 17.880 ;
        RECT 43.320 17.855 43.985 18.025 ;
        RECT 43.320 17.710 43.490 17.855 ;
        RECT 44.245 17.790 44.535 18.955 ;
        RECT 45.740 18.325 46.025 18.785 ;
        RECT 46.195 18.495 46.465 18.955 ;
        RECT 45.740 18.105 46.695 18.325 ;
        RECT 43.205 17.380 43.490 17.710 ;
        RECT 43.320 17.125 43.490 17.380 ;
        RECT 43.725 17.305 44.055 17.675 ;
        RECT 45.625 17.375 46.315 17.935 ;
        RECT 46.485 17.205 46.695 18.105 ;
        RECT 42.865 16.575 43.125 17.080 ;
        RECT 43.320 16.955 43.985 17.125 ;
        RECT 43.305 16.405 43.635 16.785 ;
        RECT 43.815 16.575 43.985 16.955 ;
        RECT 44.245 16.405 44.535 17.130 ;
        RECT 45.740 17.035 46.695 17.205 ;
        RECT 46.865 17.935 47.265 18.785 ;
        RECT 47.455 18.325 47.735 18.785 ;
        RECT 48.255 18.495 48.580 18.955 ;
        RECT 47.455 18.105 48.580 18.325 ;
        RECT 46.865 17.375 47.960 17.935 ;
        RECT 48.130 17.645 48.580 18.105 ;
        RECT 48.750 17.815 49.135 18.785 ;
        RECT 49.395 18.285 49.565 18.785 ;
        RECT 49.735 18.455 50.065 18.955 ;
        RECT 49.395 18.115 50.060 18.285 ;
        RECT 45.740 16.575 46.025 17.035 ;
        RECT 46.195 16.405 46.465 16.865 ;
        RECT 46.865 16.575 47.265 17.375 ;
        RECT 48.130 17.315 48.685 17.645 ;
        RECT 48.130 17.205 48.580 17.315 ;
        RECT 47.455 17.035 48.580 17.205 ;
        RECT 48.855 17.145 49.135 17.815 ;
        RECT 49.310 17.295 49.660 17.945 ;
        RECT 47.455 16.575 47.735 17.035 ;
        RECT 48.255 16.405 48.580 16.865 ;
        RECT 48.750 16.575 49.135 17.145 ;
        RECT 49.830 17.125 50.060 18.115 ;
        RECT 49.395 16.955 50.060 17.125 ;
        RECT 49.395 16.665 49.565 16.955 ;
        RECT 49.735 16.405 50.065 16.785 ;
        RECT 50.235 16.665 50.420 18.785 ;
        RECT 50.660 18.495 50.925 18.955 ;
        RECT 51.095 18.360 51.345 18.785 ;
        RECT 51.555 18.510 52.660 18.680 ;
        RECT 51.040 18.230 51.345 18.360 ;
        RECT 50.590 17.035 50.870 17.985 ;
        RECT 51.040 17.125 51.210 18.230 ;
        RECT 51.380 17.445 51.620 18.040 ;
        RECT 51.790 17.975 52.320 18.340 ;
        RECT 51.790 17.275 51.960 17.975 ;
        RECT 52.490 17.895 52.660 18.510 ;
        RECT 52.830 18.155 53.000 18.955 ;
        RECT 53.170 18.455 53.420 18.785 ;
        RECT 53.645 18.485 54.530 18.655 ;
        RECT 52.490 17.805 53.000 17.895 ;
        RECT 51.040 16.995 51.265 17.125 ;
        RECT 51.435 17.055 51.960 17.275 ;
        RECT 52.130 17.635 53.000 17.805 ;
        RECT 50.675 16.405 50.925 16.865 ;
        RECT 51.095 16.855 51.265 16.995 ;
        RECT 52.130 16.855 52.300 17.635 ;
        RECT 52.830 17.565 53.000 17.635 ;
        RECT 52.510 17.385 52.710 17.415 ;
        RECT 53.170 17.385 53.340 18.455 ;
        RECT 53.510 17.565 53.700 18.285 ;
        RECT 52.510 17.085 53.340 17.385 ;
        RECT 53.870 17.355 54.190 18.315 ;
        RECT 51.095 16.685 51.430 16.855 ;
        RECT 51.625 16.685 52.300 16.855 ;
        RECT 52.620 16.405 52.990 16.905 ;
        RECT 53.170 16.855 53.340 17.085 ;
        RECT 53.725 17.025 54.190 17.355 ;
        RECT 54.360 17.645 54.530 18.485 ;
        RECT 54.710 18.455 55.025 18.955 ;
        RECT 55.255 18.225 55.595 18.785 ;
        RECT 54.700 17.850 55.595 18.225 ;
        RECT 55.765 17.945 55.935 18.955 ;
        RECT 55.405 17.645 55.595 17.850 ;
        RECT 56.105 17.895 56.435 18.740 ;
        RECT 56.665 18.400 57.270 18.955 ;
        RECT 57.445 18.445 57.925 18.785 ;
        RECT 58.095 18.410 58.350 18.955 ;
        RECT 56.665 18.300 57.280 18.400 ;
        RECT 57.095 18.275 57.280 18.300 ;
        RECT 56.105 17.815 56.495 17.895 ;
        RECT 56.280 17.765 56.495 17.815 ;
        RECT 54.360 17.315 55.235 17.645 ;
        RECT 55.405 17.315 56.155 17.645 ;
        RECT 54.360 16.855 54.530 17.315 ;
        RECT 55.405 17.145 55.605 17.315 ;
        RECT 56.325 17.185 56.495 17.765 ;
        RECT 56.665 17.680 56.925 18.130 ;
        RECT 57.095 18.030 57.425 18.275 ;
        RECT 57.595 17.955 58.350 18.205 ;
        RECT 58.520 18.085 58.795 18.785 ;
        RECT 59.975 18.285 60.145 18.785 ;
        RECT 60.315 18.455 60.645 18.955 ;
        RECT 59.975 18.115 60.640 18.285 ;
        RECT 57.580 17.920 58.350 17.955 ;
        RECT 57.565 17.910 58.350 17.920 ;
        RECT 57.560 17.895 58.455 17.910 ;
        RECT 57.540 17.880 58.455 17.895 ;
        RECT 57.520 17.870 58.455 17.880 ;
        RECT 57.495 17.860 58.455 17.870 ;
        RECT 57.425 17.830 58.455 17.860 ;
        RECT 57.405 17.800 58.455 17.830 ;
        RECT 57.385 17.770 58.455 17.800 ;
        RECT 57.355 17.745 58.455 17.770 ;
        RECT 57.320 17.710 58.455 17.745 ;
        RECT 57.290 17.705 58.455 17.710 ;
        RECT 57.290 17.700 57.680 17.705 ;
        RECT 57.290 17.690 57.655 17.700 ;
        RECT 57.290 17.685 57.640 17.690 ;
        RECT 57.290 17.680 57.625 17.685 ;
        RECT 56.665 17.675 57.625 17.680 ;
        RECT 56.665 17.665 57.615 17.675 ;
        RECT 56.665 17.660 57.605 17.665 ;
        RECT 56.665 17.650 57.595 17.660 ;
        RECT 56.665 17.640 57.590 17.650 ;
        RECT 56.665 17.635 57.585 17.640 ;
        RECT 56.665 17.620 57.575 17.635 ;
        RECT 56.665 17.605 57.570 17.620 ;
        RECT 56.665 17.580 57.560 17.605 ;
        RECT 56.665 17.510 57.555 17.580 ;
        RECT 56.270 17.145 56.495 17.185 ;
        RECT 53.170 16.685 53.575 16.855 ;
        RECT 53.745 16.685 54.530 16.855 ;
        RECT 54.805 16.405 55.015 16.935 ;
        RECT 55.275 16.620 55.605 17.145 ;
        RECT 56.115 17.060 56.495 17.145 ;
        RECT 55.775 16.405 55.945 17.015 ;
        RECT 56.115 16.625 56.445 17.060 ;
        RECT 56.665 16.955 57.215 17.340 ;
        RECT 57.385 16.785 57.555 17.510 ;
        RECT 56.665 16.615 57.555 16.785 ;
        RECT 57.725 17.110 58.055 17.535 ;
        RECT 58.225 17.310 58.455 17.705 ;
        RECT 57.725 16.625 57.945 17.110 ;
        RECT 58.625 17.055 58.795 18.085 ;
        RECT 59.890 17.295 60.240 17.945 ;
        RECT 60.410 17.125 60.640 18.115 ;
        RECT 58.115 16.405 58.365 16.945 ;
        RECT 58.535 16.575 58.795 17.055 ;
        RECT 59.975 16.955 60.640 17.125 ;
        RECT 59.975 16.665 60.145 16.955 ;
        RECT 60.315 16.405 60.645 16.785 ;
        RECT 60.815 16.665 61.000 18.785 ;
        RECT 61.240 18.495 61.505 18.955 ;
        RECT 61.675 18.360 61.925 18.785 ;
        RECT 62.135 18.510 63.240 18.680 ;
        RECT 61.620 18.230 61.925 18.360 ;
        RECT 61.170 17.035 61.450 17.985 ;
        RECT 61.620 17.125 61.790 18.230 ;
        RECT 61.960 17.445 62.200 18.040 ;
        RECT 62.370 17.975 62.900 18.340 ;
        RECT 62.370 17.275 62.540 17.975 ;
        RECT 63.070 17.895 63.240 18.510 ;
        RECT 63.410 18.155 63.580 18.955 ;
        RECT 63.750 18.455 64.000 18.785 ;
        RECT 64.225 18.485 65.110 18.655 ;
        RECT 63.070 17.805 63.580 17.895 ;
        RECT 61.620 16.995 61.845 17.125 ;
        RECT 62.015 17.055 62.540 17.275 ;
        RECT 62.710 17.635 63.580 17.805 ;
        RECT 61.255 16.405 61.505 16.865 ;
        RECT 61.675 16.855 61.845 16.995 ;
        RECT 62.710 16.855 62.880 17.635 ;
        RECT 63.410 17.565 63.580 17.635 ;
        RECT 63.090 17.385 63.290 17.415 ;
        RECT 63.750 17.385 63.920 18.455 ;
        RECT 64.090 17.565 64.280 18.285 ;
        RECT 63.090 17.085 63.920 17.385 ;
        RECT 64.450 17.355 64.770 18.315 ;
        RECT 61.675 16.685 62.010 16.855 ;
        RECT 62.205 16.685 62.880 16.855 ;
        RECT 63.200 16.405 63.570 16.905 ;
        RECT 63.750 16.855 63.920 17.085 ;
        RECT 64.305 17.025 64.770 17.355 ;
        RECT 64.940 17.645 65.110 18.485 ;
        RECT 65.290 18.455 65.605 18.955 ;
        RECT 65.835 18.225 66.175 18.785 ;
        RECT 65.280 17.850 66.175 18.225 ;
        RECT 66.345 17.945 66.515 18.955 ;
        RECT 65.985 17.645 66.175 17.850 ;
        RECT 66.685 17.895 67.015 18.740 ;
        RECT 67.430 17.985 67.820 18.160 ;
        RECT 68.305 18.155 68.635 18.955 ;
        RECT 68.805 18.165 69.340 18.785 ;
        RECT 66.685 17.815 67.075 17.895 ;
        RECT 67.430 17.815 68.855 17.985 ;
        RECT 66.860 17.765 67.075 17.815 ;
        RECT 64.940 17.315 65.815 17.645 ;
        RECT 65.985 17.315 66.735 17.645 ;
        RECT 64.940 16.855 65.110 17.315 ;
        RECT 65.985 17.145 66.185 17.315 ;
        RECT 66.905 17.185 67.075 17.765 ;
        RECT 66.850 17.145 67.075 17.185 ;
        RECT 63.750 16.685 64.155 16.855 ;
        RECT 64.325 16.685 65.110 16.855 ;
        RECT 65.385 16.405 65.595 16.935 ;
        RECT 65.855 16.620 66.185 17.145 ;
        RECT 66.695 17.060 67.075 17.145 ;
        RECT 67.305 17.085 67.660 17.645 ;
        RECT 66.355 16.405 66.525 17.015 ;
        RECT 66.695 16.625 67.025 17.060 ;
        RECT 67.830 16.915 68.000 17.815 ;
        RECT 68.170 17.085 68.435 17.645 ;
        RECT 68.685 17.315 68.855 17.815 ;
        RECT 69.025 17.145 69.340 18.165 ;
        RECT 70.005 17.790 70.295 18.955 ;
        RECT 70.465 17.815 70.805 18.785 ;
        RECT 70.975 17.815 71.145 18.955 ;
        RECT 71.415 18.155 71.665 18.955 ;
        RECT 72.310 17.985 72.640 18.785 ;
        RECT 72.940 18.155 73.270 18.955 ;
        RECT 73.440 17.985 73.770 18.785 ;
        RECT 74.695 18.285 74.865 18.785 ;
        RECT 75.035 18.455 75.365 18.955 ;
        RECT 74.695 18.115 75.360 18.285 ;
        RECT 71.335 17.815 73.770 17.985 ;
        RECT 67.410 16.405 67.650 16.915 ;
        RECT 67.830 16.585 68.110 16.915 ;
        RECT 68.340 16.405 68.555 16.915 ;
        RECT 68.725 16.575 69.340 17.145 ;
        RECT 70.465 17.205 70.640 17.815 ;
        RECT 71.335 17.565 71.505 17.815 ;
        RECT 70.810 17.395 71.505 17.565 ;
        RECT 71.680 17.395 72.100 17.595 ;
        RECT 72.270 17.395 72.600 17.595 ;
        RECT 72.770 17.395 73.100 17.595 ;
        RECT 70.005 16.405 70.295 17.130 ;
        RECT 70.465 16.575 70.805 17.205 ;
        RECT 70.975 16.405 71.225 17.205 ;
        RECT 71.415 17.055 72.640 17.225 ;
        RECT 71.415 16.575 71.745 17.055 ;
        RECT 71.915 16.405 72.140 16.865 ;
        RECT 72.310 16.575 72.640 17.055 ;
        RECT 73.270 17.185 73.440 17.815 ;
        RECT 73.625 17.395 73.975 17.645 ;
        RECT 74.610 17.295 74.960 17.945 ;
        RECT 73.270 16.575 73.770 17.185 ;
        RECT 75.130 17.125 75.360 18.115 ;
        RECT 74.695 16.955 75.360 17.125 ;
        RECT 74.695 16.665 74.865 16.955 ;
        RECT 75.035 16.405 75.365 16.785 ;
        RECT 75.535 16.665 75.720 18.785 ;
        RECT 75.960 18.495 76.225 18.955 ;
        RECT 76.395 18.360 76.645 18.785 ;
        RECT 76.855 18.510 77.960 18.680 ;
        RECT 76.340 18.230 76.645 18.360 ;
        RECT 75.890 17.035 76.170 17.985 ;
        RECT 76.340 17.125 76.510 18.230 ;
        RECT 76.680 17.445 76.920 18.040 ;
        RECT 77.090 17.975 77.620 18.340 ;
        RECT 77.090 17.275 77.260 17.975 ;
        RECT 77.790 17.895 77.960 18.510 ;
        RECT 78.130 18.155 78.300 18.955 ;
        RECT 78.470 18.455 78.720 18.785 ;
        RECT 78.945 18.485 79.830 18.655 ;
        RECT 77.790 17.805 78.300 17.895 ;
        RECT 76.340 16.995 76.565 17.125 ;
        RECT 76.735 17.055 77.260 17.275 ;
        RECT 77.430 17.635 78.300 17.805 ;
        RECT 75.975 16.405 76.225 16.865 ;
        RECT 76.395 16.855 76.565 16.995 ;
        RECT 77.430 16.855 77.600 17.635 ;
        RECT 78.130 17.565 78.300 17.635 ;
        RECT 77.810 17.385 78.010 17.415 ;
        RECT 78.470 17.385 78.640 18.455 ;
        RECT 78.810 17.565 79.000 18.285 ;
        RECT 77.810 17.085 78.640 17.385 ;
        RECT 79.170 17.355 79.490 18.315 ;
        RECT 76.395 16.685 76.730 16.855 ;
        RECT 76.925 16.685 77.600 16.855 ;
        RECT 77.920 16.405 78.290 16.905 ;
        RECT 78.470 16.855 78.640 17.085 ;
        RECT 79.025 17.025 79.490 17.355 ;
        RECT 79.660 17.645 79.830 18.485 ;
        RECT 80.010 18.455 80.325 18.955 ;
        RECT 80.555 18.225 80.895 18.785 ;
        RECT 80.000 17.850 80.895 18.225 ;
        RECT 81.065 17.945 81.235 18.955 ;
        RECT 80.705 17.645 80.895 17.850 ;
        RECT 81.405 17.895 81.735 18.740 ;
        RECT 81.405 17.815 81.795 17.895 ;
        RECT 81.580 17.765 81.795 17.815 ;
        RECT 79.660 17.315 80.535 17.645 ;
        RECT 80.705 17.315 81.455 17.645 ;
        RECT 79.660 16.855 79.830 17.315 ;
        RECT 80.705 17.145 80.905 17.315 ;
        RECT 81.625 17.185 81.795 17.765 ;
        RECT 81.965 17.865 83.175 18.955 ;
        RECT 81.965 17.325 82.485 17.865 ;
        RECT 81.570 17.145 81.795 17.185 ;
        RECT 82.655 17.155 83.175 17.695 ;
        RECT 78.470 16.685 78.875 16.855 ;
        RECT 79.045 16.685 79.830 16.855 ;
        RECT 80.105 16.405 80.315 16.935 ;
        RECT 80.575 16.620 80.905 17.145 ;
        RECT 81.415 17.060 81.795 17.145 ;
        RECT 81.075 16.405 81.245 17.015 ;
        RECT 81.415 16.625 81.745 17.060 ;
        RECT 81.965 16.405 83.175 17.155 ;
        RECT 5.520 16.235 83.260 16.405 ;
        RECT 5.605 15.485 6.815 16.235 ;
        RECT 6.985 15.690 12.330 16.235 ;
        RECT 12.505 15.690 17.850 16.235 ;
        RECT 18.025 15.690 23.370 16.235 ;
        RECT 23.545 15.690 28.890 16.235 ;
        RECT 5.605 14.945 6.125 15.485 ;
        RECT 6.295 14.775 6.815 15.315 ;
        RECT 8.570 14.860 8.910 15.690 ;
        RECT 5.605 13.685 6.815 14.775 ;
        RECT 10.390 14.120 10.740 15.370 ;
        RECT 14.090 14.860 14.430 15.690 ;
        RECT 15.910 14.120 16.260 15.370 ;
        RECT 19.610 14.860 19.950 15.690 ;
        RECT 21.430 14.120 21.780 15.370 ;
        RECT 25.130 14.860 25.470 15.690 ;
        RECT 29.065 15.465 30.735 16.235 ;
        RECT 31.365 15.510 31.655 16.235 ;
        RECT 31.825 15.690 37.170 16.235 ;
        RECT 26.950 14.120 27.300 15.370 ;
        RECT 29.065 14.945 29.815 15.465 ;
        RECT 29.985 14.775 30.735 15.295 ;
        RECT 33.410 14.860 33.750 15.690 ;
        RECT 37.345 15.465 39.935 16.235 ;
        RECT 40.195 15.685 40.365 15.975 ;
        RECT 40.535 15.855 40.865 16.235 ;
        RECT 40.195 15.515 40.860 15.685 ;
        RECT 6.985 13.685 12.330 14.120 ;
        RECT 12.505 13.685 17.850 14.120 ;
        RECT 18.025 13.685 23.370 14.120 ;
        RECT 23.545 13.685 28.890 14.120 ;
        RECT 29.065 13.685 30.735 14.775 ;
        RECT 31.365 13.685 31.655 14.850 ;
        RECT 35.230 14.120 35.580 15.370 ;
        RECT 37.345 14.945 38.555 15.465 ;
        RECT 38.725 14.775 39.935 15.295 ;
        RECT 31.825 13.685 37.170 14.120 ;
        RECT 37.345 13.685 39.935 14.775 ;
        RECT 40.110 14.695 40.460 15.345 ;
        RECT 40.630 14.525 40.860 15.515 ;
        RECT 40.195 14.355 40.860 14.525 ;
        RECT 40.195 13.855 40.365 14.355 ;
        RECT 40.535 13.685 40.865 14.185 ;
        RECT 41.035 13.855 41.220 15.975 ;
        RECT 41.475 15.775 41.725 16.235 ;
        RECT 41.895 15.785 42.230 15.955 ;
        RECT 42.425 15.785 43.100 15.955 ;
        RECT 41.895 15.645 42.065 15.785 ;
        RECT 41.390 14.655 41.670 15.605 ;
        RECT 41.840 15.515 42.065 15.645 ;
        RECT 41.840 14.410 42.010 15.515 ;
        RECT 42.235 15.365 42.760 15.585 ;
        RECT 42.180 14.600 42.420 15.195 ;
        RECT 42.590 14.665 42.760 15.365 ;
        RECT 42.930 15.005 43.100 15.785 ;
        RECT 43.420 15.735 43.790 16.235 ;
        RECT 43.970 15.785 44.375 15.955 ;
        RECT 44.545 15.785 45.330 15.955 ;
        RECT 43.970 15.555 44.140 15.785 ;
        RECT 43.310 15.255 44.140 15.555 ;
        RECT 44.525 15.285 44.990 15.615 ;
        RECT 43.310 15.225 43.510 15.255 ;
        RECT 43.630 15.005 43.800 15.075 ;
        RECT 42.930 14.835 43.800 15.005 ;
        RECT 43.290 14.745 43.800 14.835 ;
        RECT 41.840 14.280 42.145 14.410 ;
        RECT 42.590 14.300 43.120 14.665 ;
        RECT 41.460 13.685 41.725 14.145 ;
        RECT 41.895 13.855 42.145 14.280 ;
        RECT 43.290 14.130 43.460 14.745 ;
        RECT 42.355 13.960 43.460 14.130 ;
        RECT 43.630 13.685 43.800 14.485 ;
        RECT 43.970 14.185 44.140 15.255 ;
        RECT 44.310 14.355 44.500 15.075 ;
        RECT 44.670 14.325 44.990 15.285 ;
        RECT 45.160 15.325 45.330 15.785 ;
        RECT 45.605 15.705 45.815 16.235 ;
        RECT 46.075 15.495 46.405 16.020 ;
        RECT 46.575 15.625 46.745 16.235 ;
        RECT 46.915 15.580 47.245 16.015 ;
        RECT 46.915 15.495 47.295 15.580 ;
        RECT 46.205 15.325 46.405 15.495 ;
        RECT 47.070 15.455 47.295 15.495 ;
        RECT 45.160 14.995 46.035 15.325 ;
        RECT 46.205 14.995 46.955 15.325 ;
        RECT 43.970 13.855 44.220 14.185 ;
        RECT 45.160 14.155 45.330 14.995 ;
        RECT 46.205 14.790 46.395 14.995 ;
        RECT 47.125 14.875 47.295 15.455 ;
        RECT 47.465 15.465 50.975 16.235 ;
        RECT 52.070 15.495 52.325 16.065 ;
        RECT 52.495 15.835 52.825 16.235 ;
        RECT 53.250 15.700 53.780 16.065 ;
        RECT 53.970 15.895 54.245 16.065 ;
        RECT 53.965 15.725 54.245 15.895 ;
        RECT 53.250 15.665 53.425 15.700 ;
        RECT 52.495 15.495 53.425 15.665 ;
        RECT 47.465 14.945 49.115 15.465 ;
        RECT 47.080 14.825 47.295 14.875 ;
        RECT 45.500 14.415 46.395 14.790 ;
        RECT 46.905 14.745 47.295 14.825 ;
        RECT 49.285 14.775 50.975 15.295 ;
        RECT 44.445 13.985 45.330 14.155 ;
        RECT 45.510 13.685 45.825 14.185 ;
        RECT 46.055 13.855 46.395 14.415 ;
        RECT 46.565 13.685 46.735 14.695 ;
        RECT 46.905 13.900 47.235 14.745 ;
        RECT 47.465 13.685 50.975 14.775 ;
        RECT 52.070 14.825 52.240 15.495 ;
        RECT 52.495 15.325 52.665 15.495 ;
        RECT 52.410 14.995 52.665 15.325 ;
        RECT 52.890 14.995 53.085 15.325 ;
        RECT 52.070 13.855 52.405 14.825 ;
        RECT 52.575 13.685 52.745 14.825 ;
        RECT 52.915 14.025 53.085 14.995 ;
        RECT 53.255 14.365 53.425 15.495 ;
        RECT 53.595 14.705 53.765 15.505 ;
        RECT 53.970 14.905 54.245 15.725 ;
        RECT 54.415 14.705 54.605 16.065 ;
        RECT 54.785 15.700 55.295 16.235 ;
        RECT 55.515 15.425 55.760 16.030 ;
        RECT 57.125 15.510 57.415 16.235 ;
        RECT 57.585 15.690 62.930 16.235 ;
        RECT 54.805 15.255 56.035 15.425 ;
        RECT 53.595 14.535 54.605 14.705 ;
        RECT 54.775 14.690 55.525 14.880 ;
        RECT 53.255 14.195 54.380 14.365 ;
        RECT 54.775 14.025 54.945 14.690 ;
        RECT 55.695 14.445 56.035 15.255 ;
        RECT 59.170 14.860 59.510 15.690 ;
        RECT 63.655 15.685 63.825 15.975 ;
        RECT 63.995 15.855 64.325 16.235 ;
        RECT 63.655 15.515 64.320 15.685 ;
        RECT 52.915 13.855 54.945 14.025 ;
        RECT 55.115 13.685 55.285 14.445 ;
        RECT 55.520 14.035 56.035 14.445 ;
        RECT 57.125 13.685 57.415 14.850 ;
        RECT 60.990 14.120 61.340 15.370 ;
        RECT 63.570 14.695 63.920 15.345 ;
        RECT 64.090 14.525 64.320 15.515 ;
        RECT 63.655 14.355 64.320 14.525 ;
        RECT 57.585 13.685 62.930 14.120 ;
        RECT 63.655 13.855 63.825 14.355 ;
        RECT 63.995 13.685 64.325 14.185 ;
        RECT 64.495 13.855 64.680 15.975 ;
        RECT 64.935 15.775 65.185 16.235 ;
        RECT 65.355 15.785 65.690 15.955 ;
        RECT 65.885 15.785 66.560 15.955 ;
        RECT 65.355 15.645 65.525 15.785 ;
        RECT 64.850 14.655 65.130 15.605 ;
        RECT 65.300 15.515 65.525 15.645 ;
        RECT 65.300 14.410 65.470 15.515 ;
        RECT 65.695 15.365 66.220 15.585 ;
        RECT 65.640 14.600 65.880 15.195 ;
        RECT 66.050 14.665 66.220 15.365 ;
        RECT 66.390 15.005 66.560 15.785 ;
        RECT 66.880 15.735 67.250 16.235 ;
        RECT 67.430 15.785 67.835 15.955 ;
        RECT 68.005 15.785 68.790 15.955 ;
        RECT 67.430 15.555 67.600 15.785 ;
        RECT 66.770 15.255 67.600 15.555 ;
        RECT 67.985 15.285 68.450 15.615 ;
        RECT 66.770 15.225 66.970 15.255 ;
        RECT 67.090 15.005 67.260 15.075 ;
        RECT 66.390 14.835 67.260 15.005 ;
        RECT 66.750 14.745 67.260 14.835 ;
        RECT 65.300 14.280 65.605 14.410 ;
        RECT 66.050 14.300 66.580 14.665 ;
        RECT 64.920 13.685 65.185 14.145 ;
        RECT 65.355 13.855 65.605 14.280 ;
        RECT 66.750 14.130 66.920 14.745 ;
        RECT 65.815 13.960 66.920 14.130 ;
        RECT 67.090 13.685 67.260 14.485 ;
        RECT 67.430 14.185 67.600 15.255 ;
        RECT 67.770 14.355 67.960 15.075 ;
        RECT 68.130 14.325 68.450 15.285 ;
        RECT 68.620 15.325 68.790 15.785 ;
        RECT 69.065 15.705 69.275 16.235 ;
        RECT 69.535 15.495 69.865 16.020 ;
        RECT 70.035 15.625 70.205 16.235 ;
        RECT 70.375 15.580 70.705 16.015 ;
        RECT 71.015 15.685 71.185 16.065 ;
        RECT 71.365 15.855 71.695 16.235 ;
        RECT 70.375 15.495 70.755 15.580 ;
        RECT 71.015 15.515 71.680 15.685 ;
        RECT 71.875 15.560 72.135 16.065 ;
        RECT 72.470 15.725 72.710 16.235 ;
        RECT 72.890 15.725 73.170 16.055 ;
        RECT 73.400 15.725 73.615 16.235 ;
        RECT 69.665 15.325 69.865 15.495 ;
        RECT 70.530 15.455 70.755 15.495 ;
        RECT 68.620 14.995 69.495 15.325 ;
        RECT 69.665 14.995 70.415 15.325 ;
        RECT 67.430 13.855 67.680 14.185 ;
        RECT 68.620 14.155 68.790 14.995 ;
        RECT 69.665 14.790 69.855 14.995 ;
        RECT 70.585 14.875 70.755 15.455 ;
        RECT 70.945 14.965 71.275 15.335 ;
        RECT 71.510 15.260 71.680 15.515 ;
        RECT 70.540 14.825 70.755 14.875 ;
        RECT 68.960 14.415 69.855 14.790 ;
        RECT 70.365 14.745 70.755 14.825 ;
        RECT 71.510 14.930 71.795 15.260 ;
        RECT 71.510 14.785 71.680 14.930 ;
        RECT 67.905 13.985 68.790 14.155 ;
        RECT 68.970 13.685 69.285 14.185 ;
        RECT 69.515 13.855 69.855 14.415 ;
        RECT 70.025 13.685 70.195 14.695 ;
        RECT 70.365 13.900 70.695 14.745 ;
        RECT 71.015 14.615 71.680 14.785 ;
        RECT 71.965 14.760 72.135 15.560 ;
        RECT 72.365 14.995 72.720 15.555 ;
        RECT 72.890 14.825 73.060 15.725 ;
        RECT 73.230 14.995 73.495 15.555 ;
        RECT 73.785 15.495 74.400 16.065 ;
        RECT 74.695 15.685 74.865 15.975 ;
        RECT 75.035 15.855 75.365 16.235 ;
        RECT 74.695 15.515 75.360 15.685 ;
        RECT 73.745 14.825 73.915 15.325 ;
        RECT 71.015 13.855 71.185 14.615 ;
        RECT 71.365 13.685 71.695 14.445 ;
        RECT 71.865 13.855 72.135 14.760 ;
        RECT 72.490 14.655 73.915 14.825 ;
        RECT 72.490 14.480 72.880 14.655 ;
        RECT 73.365 13.685 73.695 14.485 ;
        RECT 74.085 14.475 74.400 15.495 ;
        RECT 74.610 14.695 74.960 15.345 ;
        RECT 75.130 14.525 75.360 15.515 ;
        RECT 73.865 13.855 74.400 14.475 ;
        RECT 74.695 14.355 75.360 14.525 ;
        RECT 74.695 13.855 74.865 14.355 ;
        RECT 75.035 13.685 75.365 14.185 ;
        RECT 75.535 13.855 75.720 15.975 ;
        RECT 75.975 15.775 76.225 16.235 ;
        RECT 76.395 15.785 76.730 15.955 ;
        RECT 76.925 15.785 77.600 15.955 ;
        RECT 76.395 15.645 76.565 15.785 ;
        RECT 75.890 14.655 76.170 15.605 ;
        RECT 76.340 15.515 76.565 15.645 ;
        RECT 76.340 14.410 76.510 15.515 ;
        RECT 76.735 15.365 77.260 15.585 ;
        RECT 76.680 14.600 76.920 15.195 ;
        RECT 77.090 14.665 77.260 15.365 ;
        RECT 77.430 15.005 77.600 15.785 ;
        RECT 77.920 15.735 78.290 16.235 ;
        RECT 78.470 15.785 78.875 15.955 ;
        RECT 79.045 15.785 79.830 15.955 ;
        RECT 78.470 15.555 78.640 15.785 ;
        RECT 77.810 15.255 78.640 15.555 ;
        RECT 79.025 15.285 79.490 15.615 ;
        RECT 77.810 15.225 78.010 15.255 ;
        RECT 78.130 15.005 78.300 15.075 ;
        RECT 77.430 14.835 78.300 15.005 ;
        RECT 77.790 14.745 78.300 14.835 ;
        RECT 76.340 14.280 76.645 14.410 ;
        RECT 77.090 14.300 77.620 14.665 ;
        RECT 75.960 13.685 76.225 14.145 ;
        RECT 76.395 13.855 76.645 14.280 ;
        RECT 77.790 14.130 77.960 14.745 ;
        RECT 76.855 13.960 77.960 14.130 ;
        RECT 78.130 13.685 78.300 14.485 ;
        RECT 78.470 14.185 78.640 15.255 ;
        RECT 78.810 14.355 79.000 15.075 ;
        RECT 79.170 14.325 79.490 15.285 ;
        RECT 79.660 15.325 79.830 15.785 ;
        RECT 80.105 15.705 80.315 16.235 ;
        RECT 80.575 15.495 80.905 16.020 ;
        RECT 81.075 15.625 81.245 16.235 ;
        RECT 81.415 15.580 81.745 16.015 ;
        RECT 81.415 15.495 81.795 15.580 ;
        RECT 80.705 15.325 80.905 15.495 ;
        RECT 81.570 15.455 81.795 15.495 ;
        RECT 81.965 15.485 83.175 16.235 ;
        RECT 79.660 14.995 80.535 15.325 ;
        RECT 80.705 14.995 81.455 15.325 ;
        RECT 78.470 13.855 78.720 14.185 ;
        RECT 79.660 14.155 79.830 14.995 ;
        RECT 80.705 14.790 80.895 14.995 ;
        RECT 81.625 14.875 81.795 15.455 ;
        RECT 81.580 14.825 81.795 14.875 ;
        RECT 80.000 14.415 80.895 14.790 ;
        RECT 81.405 14.745 81.795 14.825 ;
        RECT 81.965 14.775 82.485 15.315 ;
        RECT 82.655 14.945 83.175 15.485 ;
        RECT 78.945 13.985 79.830 14.155 ;
        RECT 80.010 13.685 80.325 14.185 ;
        RECT 80.555 13.855 80.895 14.415 ;
        RECT 81.065 13.685 81.235 14.695 ;
        RECT 81.405 13.900 81.735 14.745 ;
        RECT 81.965 13.685 83.175 14.775 ;
        RECT 5.520 13.515 83.260 13.685 ;
        RECT 5.605 12.425 6.815 13.515 ;
        RECT 6.985 13.080 12.330 13.515 ;
        RECT 12.505 13.080 17.850 13.515 ;
        RECT 5.605 11.715 6.125 12.255 ;
        RECT 6.295 11.885 6.815 12.425 ;
        RECT 5.605 10.965 6.815 11.715 ;
        RECT 8.570 11.510 8.910 12.340 ;
        RECT 10.390 11.830 10.740 13.080 ;
        RECT 14.090 11.510 14.430 12.340 ;
        RECT 15.910 11.830 16.260 13.080 ;
        RECT 18.485 12.350 18.775 13.515 ;
        RECT 18.945 13.080 24.290 13.515 ;
        RECT 24.465 13.080 29.810 13.515 ;
        RECT 6.985 10.965 12.330 11.510 ;
        RECT 12.505 10.965 17.850 11.510 ;
        RECT 18.485 10.965 18.775 11.690 ;
        RECT 20.530 11.510 20.870 12.340 ;
        RECT 22.350 11.830 22.700 13.080 ;
        RECT 26.050 11.510 26.390 12.340 ;
        RECT 27.870 11.830 28.220 13.080 ;
        RECT 29.985 12.425 31.195 13.515 ;
        RECT 29.985 11.715 30.505 12.255 ;
        RECT 30.675 11.885 31.195 12.425 ;
        RECT 31.365 12.350 31.655 13.515 ;
        RECT 31.825 12.425 35.335 13.515 ;
        RECT 35.965 12.920 36.400 13.345 ;
        RECT 36.570 13.090 36.955 13.515 ;
        RECT 35.965 12.750 36.955 12.920 ;
        RECT 31.825 11.735 33.475 12.255 ;
        RECT 33.645 11.905 35.335 12.425 ;
        RECT 35.965 11.875 36.450 12.580 ;
        RECT 36.620 12.205 36.955 12.750 ;
        RECT 37.125 12.555 37.550 13.345 ;
        RECT 37.720 12.920 37.995 13.345 ;
        RECT 38.165 13.090 38.550 13.515 ;
        RECT 37.720 12.725 38.550 12.920 ;
        RECT 37.125 12.375 38.030 12.555 ;
        RECT 36.620 11.875 37.030 12.205 ;
        RECT 37.200 11.875 38.030 12.375 ;
        RECT 38.200 12.205 38.550 12.725 ;
        RECT 38.720 12.555 38.965 13.345 ;
        RECT 39.155 12.920 39.410 13.345 ;
        RECT 39.580 13.090 39.965 13.515 ;
        RECT 39.155 12.725 39.965 12.920 ;
        RECT 38.720 12.375 39.445 12.555 ;
        RECT 38.200 11.875 38.625 12.205 ;
        RECT 38.795 11.875 39.445 12.375 ;
        RECT 39.615 12.205 39.965 12.725 ;
        RECT 40.135 12.375 40.395 13.345 ;
        RECT 39.615 11.875 40.040 12.205 ;
        RECT 18.945 10.965 24.290 11.510 ;
        RECT 24.465 10.965 29.810 11.510 ;
        RECT 29.985 10.965 31.195 11.715 ;
        RECT 31.365 10.965 31.655 11.690 ;
        RECT 31.825 10.965 35.335 11.735 ;
        RECT 36.620 11.705 36.955 11.875 ;
        RECT 37.200 11.705 37.550 11.875 ;
        RECT 38.200 11.705 38.550 11.875 ;
        RECT 38.795 11.705 38.965 11.875 ;
        RECT 39.615 11.705 39.965 11.875 ;
        RECT 40.210 11.705 40.395 12.375 ;
        RECT 35.965 11.535 36.955 11.705 ;
        RECT 35.965 11.135 36.400 11.535 ;
        RECT 36.570 10.965 36.955 11.365 ;
        RECT 37.125 11.135 37.550 11.705 ;
        RECT 37.740 11.535 38.550 11.705 ;
        RECT 37.740 11.135 37.995 11.535 ;
        RECT 38.165 10.965 38.550 11.365 ;
        RECT 38.720 11.135 38.965 11.705 ;
        RECT 39.155 11.535 39.965 11.705 ;
        RECT 39.155 11.135 39.410 11.535 ;
        RECT 39.580 10.965 39.965 11.365 ;
        RECT 40.135 11.135 40.395 11.705 ;
        RECT 40.565 12.545 40.835 13.315 ;
        RECT 41.005 12.735 41.335 13.515 ;
        RECT 41.540 12.910 41.725 13.315 ;
        RECT 41.895 13.090 42.230 13.515 ;
        RECT 41.540 12.735 42.205 12.910 ;
        RECT 40.565 12.375 41.695 12.545 ;
        RECT 40.565 11.465 40.735 12.375 ;
        RECT 40.905 11.625 41.265 12.205 ;
        RECT 41.445 11.875 41.695 12.375 ;
        RECT 41.865 11.705 42.205 12.735 ;
        RECT 42.410 12.365 42.670 13.515 ;
        RECT 42.845 12.440 43.100 13.345 ;
        RECT 43.270 12.755 43.600 13.515 ;
        RECT 43.815 12.585 43.985 13.345 ;
        RECT 41.520 11.535 42.205 11.705 ;
        RECT 40.565 11.135 40.825 11.465 ;
        RECT 41.035 10.965 41.310 11.445 ;
        RECT 41.520 11.135 41.725 11.535 ;
        RECT 41.895 10.965 42.230 11.365 ;
        RECT 42.410 10.965 42.670 11.805 ;
        RECT 42.845 11.710 43.015 12.440 ;
        RECT 43.270 12.415 43.985 12.585 ;
        RECT 43.270 12.205 43.440 12.415 ;
        RECT 44.245 12.350 44.535 13.515 ;
        RECT 45.630 12.365 45.890 13.515 ;
        RECT 46.065 12.440 46.320 13.345 ;
        RECT 46.490 12.755 46.820 13.515 ;
        RECT 47.035 12.585 47.205 13.345 ;
        RECT 43.185 11.875 43.440 12.205 ;
        RECT 42.845 11.135 43.100 11.710 ;
        RECT 43.270 11.685 43.440 11.875 ;
        RECT 43.720 11.865 44.075 12.235 ;
        RECT 43.270 11.515 43.985 11.685 ;
        RECT 43.270 10.965 43.600 11.345 ;
        RECT 43.815 11.135 43.985 11.515 ;
        RECT 44.245 10.965 44.535 11.690 ;
        RECT 45.630 10.965 45.890 11.805 ;
        RECT 46.065 11.710 46.235 12.440 ;
        RECT 46.490 12.415 47.205 12.585 ;
        RECT 47.465 12.425 48.675 13.515 ;
        RECT 46.490 12.205 46.660 12.415 ;
        RECT 46.405 11.875 46.660 12.205 ;
        RECT 46.065 11.135 46.320 11.710 ;
        RECT 46.490 11.685 46.660 11.875 ;
        RECT 46.940 11.865 47.295 12.235 ;
        RECT 47.465 11.715 47.985 12.255 ;
        RECT 48.155 11.885 48.675 12.425 ;
        RECT 48.845 12.545 49.115 13.315 ;
        RECT 49.285 12.735 49.615 13.515 ;
        RECT 49.820 12.910 50.005 13.315 ;
        RECT 50.175 13.090 50.510 13.515 ;
        RECT 50.685 13.080 56.030 13.515 ;
        RECT 49.820 12.735 50.485 12.910 ;
        RECT 48.845 12.375 49.975 12.545 ;
        RECT 46.490 11.515 47.205 11.685 ;
        RECT 46.490 10.965 46.820 11.345 ;
        RECT 47.035 11.135 47.205 11.515 ;
        RECT 47.465 10.965 48.675 11.715 ;
        RECT 48.845 11.465 49.015 12.375 ;
        RECT 49.185 11.625 49.545 12.205 ;
        RECT 49.725 11.875 49.975 12.375 ;
        RECT 50.145 11.705 50.485 12.735 ;
        RECT 49.800 11.535 50.485 11.705 ;
        RECT 48.845 11.135 49.105 11.465 ;
        RECT 49.315 10.965 49.590 11.445 ;
        RECT 49.800 11.135 50.005 11.535 ;
        RECT 52.270 11.510 52.610 12.340 ;
        RECT 54.090 11.830 54.440 13.080 ;
        RECT 57.125 12.350 57.415 13.515 ;
        RECT 57.585 13.080 62.930 13.515 ;
        RECT 50.175 10.965 50.510 11.365 ;
        RECT 50.685 10.965 56.030 11.510 ;
        RECT 57.125 10.965 57.415 11.690 ;
        RECT 59.170 11.510 59.510 12.340 ;
        RECT 60.990 11.830 61.340 13.080 ;
        RECT 63.105 12.425 64.775 13.515 ;
        RECT 63.105 11.735 63.855 12.255 ;
        RECT 64.025 11.905 64.775 12.425 ;
        RECT 64.950 12.365 65.210 13.515 ;
        RECT 65.385 12.440 65.640 13.345 ;
        RECT 65.810 12.755 66.140 13.515 ;
        RECT 66.355 12.585 66.525 13.345 ;
        RECT 57.585 10.965 62.930 11.510 ;
        RECT 63.105 10.965 64.775 11.735 ;
        RECT 64.950 10.965 65.210 11.805 ;
        RECT 65.385 11.710 65.555 12.440 ;
        RECT 65.810 12.415 66.525 12.585 ;
        RECT 66.785 12.425 67.995 13.515 ;
        RECT 65.810 12.205 65.980 12.415 ;
        RECT 65.725 11.875 65.980 12.205 ;
        RECT 65.385 11.135 65.640 11.710 ;
        RECT 65.810 11.685 65.980 11.875 ;
        RECT 66.260 11.865 66.615 12.235 ;
        RECT 66.785 11.715 67.305 12.255 ;
        RECT 67.475 11.885 67.995 12.425 ;
        RECT 68.170 12.365 68.430 13.515 ;
        RECT 68.605 12.440 68.860 13.345 ;
        RECT 69.030 12.755 69.360 13.515 ;
        RECT 69.575 12.585 69.745 13.345 ;
        RECT 65.810 11.515 66.525 11.685 ;
        RECT 65.810 10.965 66.140 11.345 ;
        RECT 66.355 11.135 66.525 11.515 ;
        RECT 66.785 10.965 67.995 11.715 ;
        RECT 68.170 10.965 68.430 11.805 ;
        RECT 68.605 11.710 68.775 12.440 ;
        RECT 69.030 12.415 69.745 12.585 ;
        RECT 69.030 12.205 69.200 12.415 ;
        RECT 70.005 12.350 70.295 13.515 ;
        RECT 71.390 12.365 71.650 13.515 ;
        RECT 71.825 12.440 72.080 13.345 ;
        RECT 72.250 12.755 72.580 13.515 ;
        RECT 72.795 12.585 72.965 13.345 ;
        RECT 68.945 11.875 69.200 12.205 ;
        RECT 68.605 11.135 68.860 11.710 ;
        RECT 69.030 11.685 69.200 11.875 ;
        RECT 69.480 11.865 69.835 12.235 ;
        RECT 69.030 11.515 69.745 11.685 ;
        RECT 69.030 10.965 69.360 11.345 ;
        RECT 69.575 11.135 69.745 11.515 ;
        RECT 70.005 10.965 70.295 11.690 ;
        RECT 71.390 10.965 71.650 11.805 ;
        RECT 71.825 11.710 71.995 12.440 ;
        RECT 72.250 12.415 72.965 12.585 ;
        RECT 73.315 12.585 73.485 13.345 ;
        RECT 73.700 12.755 74.030 13.515 ;
        RECT 73.315 12.415 74.030 12.585 ;
        RECT 74.200 12.440 74.455 13.345 ;
        RECT 72.250 12.205 72.420 12.415 ;
        RECT 72.165 11.875 72.420 12.205 ;
        RECT 71.825 11.135 72.080 11.710 ;
        RECT 72.250 11.685 72.420 11.875 ;
        RECT 72.700 11.865 73.055 12.235 ;
        RECT 73.225 11.865 73.580 12.235 ;
        RECT 73.860 12.205 74.030 12.415 ;
        RECT 73.860 11.875 74.115 12.205 ;
        RECT 73.860 11.685 74.030 11.875 ;
        RECT 74.285 11.710 74.455 12.440 ;
        RECT 74.630 12.365 74.890 13.515 ;
        RECT 75.155 12.585 75.325 13.345 ;
        RECT 75.540 12.755 75.870 13.515 ;
        RECT 75.155 12.415 75.870 12.585 ;
        RECT 76.040 12.440 76.295 13.345 ;
        RECT 75.065 11.865 75.420 12.235 ;
        RECT 75.700 12.205 75.870 12.415 ;
        RECT 75.700 11.875 75.955 12.205 ;
        RECT 72.250 11.515 72.965 11.685 ;
        RECT 72.250 10.965 72.580 11.345 ;
        RECT 72.795 11.135 72.965 11.515 ;
        RECT 73.315 11.515 74.030 11.685 ;
        RECT 73.315 11.135 73.485 11.515 ;
        RECT 73.700 10.965 74.030 11.345 ;
        RECT 74.200 11.135 74.455 11.710 ;
        RECT 74.630 10.965 74.890 11.805 ;
        RECT 75.700 11.685 75.870 11.875 ;
        RECT 76.125 11.710 76.295 12.440 ;
        RECT 76.470 12.365 76.730 13.515 ;
        RECT 77.090 12.545 77.480 12.720 ;
        RECT 77.965 12.715 78.295 13.515 ;
        RECT 78.465 12.725 79.000 13.345 ;
        RECT 77.090 12.375 78.515 12.545 ;
        RECT 75.155 11.515 75.870 11.685 ;
        RECT 75.155 11.135 75.325 11.515 ;
        RECT 75.540 10.965 75.870 11.345 ;
        RECT 76.040 11.135 76.295 11.710 ;
        RECT 76.470 10.965 76.730 11.805 ;
        RECT 76.965 11.645 77.320 12.205 ;
        RECT 77.490 11.475 77.660 12.375 ;
        RECT 77.830 11.645 78.095 12.205 ;
        RECT 78.345 11.875 78.515 12.375 ;
        RECT 78.685 11.705 79.000 12.725 ;
        RECT 80.215 12.585 80.385 13.345 ;
        RECT 80.600 12.755 80.930 13.515 ;
        RECT 80.215 12.415 80.930 12.585 ;
        RECT 81.100 12.440 81.355 13.345 ;
        RECT 80.125 11.865 80.480 12.235 ;
        RECT 80.760 12.205 80.930 12.415 ;
        RECT 80.760 11.875 81.015 12.205 ;
        RECT 77.070 10.965 77.310 11.475 ;
        RECT 77.490 11.145 77.770 11.475 ;
        RECT 78.000 10.965 78.215 11.475 ;
        RECT 78.385 11.135 79.000 11.705 ;
        RECT 80.760 11.685 80.930 11.875 ;
        RECT 81.185 11.710 81.355 12.440 ;
        RECT 81.530 12.365 81.790 13.515 ;
        RECT 81.965 12.425 83.175 13.515 ;
        RECT 81.965 11.885 82.485 12.425 ;
        RECT 80.215 11.515 80.930 11.685 ;
        RECT 80.215 11.135 80.385 11.515 ;
        RECT 80.600 10.965 80.930 11.345 ;
        RECT 81.100 11.135 81.355 11.710 ;
        RECT 81.530 10.965 81.790 11.805 ;
        RECT 82.655 11.715 83.175 12.255 ;
        RECT 81.965 10.965 83.175 11.715 ;
        RECT 5.520 10.795 83.260 10.965 ;
      LAYER met1 ;
        RECT 5.520 165.680 83.260 166.160 ;
        RECT 38.710 165.480 39.030 165.540 ;
        RECT 39.645 165.480 39.935 165.525 ;
        RECT 38.710 165.340 39.935 165.480 ;
        RECT 38.710 165.280 39.030 165.340 ;
        RECT 39.645 165.295 39.935 165.340 ;
        RECT 58.505 165.480 58.795 165.525 ;
        RECT 64.470 165.480 64.790 165.540 ;
        RECT 58.505 165.340 64.790 165.480 ;
        RECT 58.505 165.295 58.795 165.340 ;
        RECT 64.470 165.280 64.790 165.340 ;
        RECT 64.930 165.480 65.250 165.540 ;
        RECT 68.625 165.480 68.915 165.525 ;
        RECT 74.130 165.480 74.450 165.540 ;
        RECT 64.930 165.340 68.380 165.480 ;
        RECT 64.930 165.280 65.250 165.340 ;
        RECT 55.745 165.140 56.035 165.185 ;
        RECT 67.690 165.140 68.010 165.200 ;
        RECT 55.745 165.000 68.010 165.140 ;
        RECT 68.240 165.140 68.380 165.340 ;
        RECT 68.625 165.340 74.450 165.480 ;
        RECT 68.625 165.295 68.915 165.340 ;
        RECT 74.130 165.280 74.450 165.340 ;
        RECT 76.430 165.480 76.750 165.540 ;
        RECT 82.410 165.480 82.730 165.540 ;
        RECT 76.430 165.340 82.730 165.480 ;
        RECT 76.430 165.280 76.750 165.340 ;
        RECT 82.410 165.280 82.730 165.340 ;
        RECT 68.240 165.000 78.040 165.140 ;
        RECT 55.745 164.955 56.035 165.000 ;
        RECT 67.690 164.940 68.010 165.000 ;
        RECT 77.350 164.800 77.670 164.860 ;
        RECT 60.420 164.660 77.670 164.800 ;
        RECT 40.550 164.260 40.870 164.520 ;
        RECT 52.970 164.260 53.290 164.520 ;
        RECT 54.350 164.460 54.670 164.520 ;
        RECT 54.825 164.460 55.115 164.505 ;
        RECT 54.350 164.320 55.115 164.460 ;
        RECT 54.350 164.260 54.670 164.320 ;
        RECT 54.825 164.275 55.115 164.320 ;
        RECT 56.650 164.260 56.970 164.520 ;
        RECT 57.570 164.260 57.890 164.520 ;
        RECT 52.050 163.580 52.370 163.840 ;
        RECT 53.890 163.580 54.210 163.840 ;
        RECT 59.885 163.780 60.175 163.825 ;
        RECT 60.420 163.780 60.560 164.660 ;
        RECT 77.350 164.600 77.670 164.660 ;
        RECT 60.805 164.275 61.095 164.505 ;
        RECT 63.565 164.460 63.855 164.505 ;
        RECT 63.565 164.320 69.300 164.460 ;
        RECT 63.565 164.275 63.855 164.320 ;
        RECT 60.880 164.120 61.020 164.275 ;
        RECT 62.185 164.120 62.475 164.165 ;
        RECT 62.630 164.120 62.950 164.180 ;
        RECT 60.880 163.980 61.940 164.120 ;
        RECT 59.885 163.640 60.560 163.780 ;
        RECT 59.885 163.595 60.175 163.640 ;
        RECT 61.250 163.580 61.570 163.840 ;
        RECT 61.800 163.780 61.940 163.980 ;
        RECT 62.185 163.980 62.950 164.120 ;
        RECT 62.185 163.935 62.475 163.980 ;
        RECT 62.630 163.920 62.950 163.980 ;
        RECT 63.105 164.120 63.395 164.165 ;
        RECT 64.010 164.120 64.330 164.180 ;
        RECT 63.105 163.980 64.330 164.120 ;
        RECT 63.105 163.935 63.395 163.980 ;
        RECT 64.010 163.920 64.330 163.980 ;
        RECT 64.485 164.120 64.775 164.165 ;
        RECT 64.930 164.120 65.250 164.180 ;
        RECT 64.485 163.980 65.250 164.120 ;
        RECT 64.485 163.935 64.775 163.980 ;
        RECT 64.560 163.780 64.700 163.935 ;
        RECT 64.930 163.920 65.250 163.980 ;
        RECT 65.405 164.120 65.695 164.165 ;
        RECT 65.405 163.980 66.540 164.120 ;
        RECT 65.405 163.935 65.695 163.980 ;
        RECT 61.800 163.640 64.700 163.780 ;
        RECT 65.850 163.580 66.170 163.840 ;
        RECT 66.400 163.780 66.540 163.980 ;
        RECT 66.770 163.920 67.090 164.180 ;
        RECT 67.230 164.120 67.550 164.180 ;
        RECT 67.705 164.120 67.995 164.165 ;
        RECT 67.230 163.980 67.995 164.120 ;
        RECT 69.160 164.120 69.300 164.320 ;
        RECT 69.530 164.260 69.850 164.520 ;
        RECT 74.590 164.460 74.910 164.520 ;
        RECT 70.080 164.320 74.910 164.460 ;
        RECT 70.080 164.120 70.220 164.320 ;
        RECT 74.590 164.260 74.910 164.320 ;
        RECT 75.065 164.460 75.355 164.505 ;
        RECT 76.430 164.460 76.750 164.520 ;
        RECT 75.065 164.320 76.750 164.460 ;
        RECT 75.065 164.275 75.355 164.320 ;
        RECT 76.430 164.260 76.750 164.320 ;
        RECT 76.890 164.460 77.210 164.520 ;
        RECT 77.900 164.505 78.040 165.000 ;
        RECT 77.825 164.460 78.115 164.505 ;
        RECT 76.890 164.320 78.115 164.460 ;
        RECT 76.890 164.260 77.210 164.320 ;
        RECT 77.825 164.275 78.115 164.320 ;
        RECT 79.665 164.460 79.955 164.505 ;
        RECT 80.570 164.460 80.890 164.520 ;
        RECT 79.665 164.320 80.890 164.460 ;
        RECT 79.665 164.275 79.955 164.320 ;
        RECT 80.570 164.260 80.890 164.320 ;
        RECT 69.160 163.980 70.220 164.120 ;
        RECT 70.465 164.120 70.755 164.165 ;
        RECT 70.910 164.120 71.230 164.180 ;
        RECT 70.465 163.980 71.230 164.120 ;
        RECT 67.230 163.920 67.550 163.980 ;
        RECT 67.705 163.935 67.995 163.980 ;
        RECT 70.465 163.935 70.755 163.980 ;
        RECT 70.540 163.780 70.680 163.935 ;
        RECT 70.910 163.920 71.230 163.980 ;
        RECT 71.370 163.920 71.690 164.180 ;
        RECT 71.830 164.120 72.150 164.180 ;
        RECT 72.765 164.120 73.055 164.165 ;
        RECT 71.830 163.980 73.055 164.120 ;
        RECT 71.830 163.920 72.150 163.980 ;
        RECT 72.765 163.935 73.055 163.980 ;
        RECT 73.210 164.120 73.530 164.180 ;
        RECT 73.685 164.120 73.975 164.165 ;
        RECT 73.210 163.980 73.975 164.120 ;
        RECT 73.210 163.920 73.530 163.980 ;
        RECT 73.685 163.935 73.975 163.980 ;
        RECT 75.985 164.120 76.275 164.165 ;
        RECT 78.270 164.120 78.590 164.180 ;
        RECT 75.985 163.980 78.590 164.120 ;
        RECT 75.985 163.935 76.275 163.980 ;
        RECT 78.270 163.920 78.590 163.980 ;
        RECT 78.730 163.920 79.050 164.180 ;
        RECT 79.190 164.120 79.510 164.180 ;
        RECT 81.030 164.120 81.350 164.180 ;
        RECT 79.190 163.980 81.350 164.120 ;
        RECT 79.190 163.920 79.510 163.980 ;
        RECT 81.030 163.920 81.350 163.980 ;
        RECT 66.400 163.640 70.680 163.780 ;
        RECT 72.290 163.580 72.610 163.840 ;
        RECT 74.130 163.780 74.450 163.840 ;
        RECT 74.605 163.780 74.895 163.825 ;
        RECT 74.130 163.640 74.895 163.780 ;
        RECT 74.130 163.580 74.450 163.640 ;
        RECT 74.605 163.595 74.895 163.640 ;
        RECT 76.430 163.780 76.750 163.840 ;
        RECT 76.905 163.780 77.195 163.825 ;
        RECT 76.430 163.640 77.195 163.780 ;
        RECT 76.430 163.580 76.750 163.640 ;
        RECT 76.905 163.595 77.195 163.640 ;
        RECT 77.350 163.780 77.670 163.840 ;
        RECT 80.585 163.780 80.875 163.825 ;
        RECT 77.350 163.640 80.875 163.780 ;
        RECT 77.350 163.580 77.670 163.640 ;
        RECT 80.585 163.595 80.875 163.640 ;
        RECT 5.520 162.960 83.260 163.440 ;
        RECT 56.650 162.760 56.970 162.820 ;
        RECT 62.185 162.760 62.475 162.805 ;
        RECT 66.770 162.760 67.090 162.820 ;
        RECT 56.650 162.620 67.090 162.760 ;
        RECT 56.650 162.560 56.970 162.620 ;
        RECT 62.185 162.575 62.475 162.620 ;
        RECT 66.770 162.560 67.090 162.620 ;
        RECT 67.230 162.760 67.550 162.820 ;
        RECT 71.830 162.760 72.150 162.820 ;
        RECT 67.230 162.620 72.150 162.760 ;
        RECT 67.230 162.560 67.550 162.620 ;
        RECT 71.830 162.560 72.150 162.620 ;
        RECT 72.290 162.560 72.610 162.820 ;
        RECT 73.760 162.620 77.580 162.760 ;
        RECT 53.890 162.220 54.210 162.480 ;
        RECT 69.990 162.420 70.310 162.480 ;
        RECT 72.380 162.420 72.520 162.560 ;
        RECT 69.990 162.280 72.060 162.420 ;
        RECT 72.380 162.280 72.980 162.420 ;
        RECT 69.990 162.220 70.310 162.280 ;
        RECT 34.585 161.895 34.875 162.125 ;
        RECT 34.660 161.740 34.800 161.895 ;
        RECT 35.950 161.880 36.270 162.140 ;
        RECT 36.870 161.880 37.190 162.140 ;
        RECT 37.330 162.080 37.650 162.140 ;
        RECT 44.705 162.080 44.995 162.125 ;
        RECT 37.330 161.940 44.995 162.080 ;
        RECT 37.330 161.880 37.650 161.940 ;
        RECT 44.705 161.895 44.995 161.940 ;
        RECT 45.610 161.880 45.930 162.140 ;
        RECT 52.985 162.080 53.275 162.125 ;
        RECT 53.980 162.080 54.120 162.220 ;
        RECT 67.690 162.125 68.010 162.140 ;
        RECT 52.985 161.940 64.240 162.080 ;
        RECT 52.985 161.895 53.275 161.940 ;
        RECT 38.250 161.740 38.570 161.800 ;
        RECT 34.660 161.600 38.570 161.740 ;
        RECT 38.250 161.540 38.570 161.600 ;
        RECT 53.890 161.540 54.210 161.800 ;
        RECT 54.900 161.600 60.100 161.740 ;
        RECT 35.030 161.200 35.350 161.460 ;
        RECT 35.490 161.200 35.810 161.460 ;
        RECT 52.065 161.400 52.355 161.445 ;
        RECT 54.900 161.400 55.040 161.600 ;
        RECT 52.065 161.260 55.040 161.400 ;
        RECT 55.270 161.400 55.590 161.460 ;
        RECT 57.585 161.400 57.875 161.445 ;
        RECT 55.270 161.260 57.875 161.400 ;
        RECT 59.960 161.400 60.100 161.600 ;
        RECT 60.330 161.540 60.650 161.800 ;
        RECT 63.090 161.400 63.410 161.460 ;
        RECT 59.960 161.260 63.410 161.400 ;
        RECT 52.065 161.215 52.355 161.260 ;
        RECT 55.270 161.200 55.590 161.260 ;
        RECT 57.585 161.215 57.875 161.260 ;
        RECT 63.090 161.200 63.410 161.260 ;
        RECT 33.650 160.860 33.970 161.120 ;
        RECT 41.930 161.060 42.250 161.120 ;
        RECT 45.165 161.060 45.455 161.105 ;
        RECT 41.930 160.920 45.455 161.060 ;
        RECT 41.930 160.860 42.250 160.920 ;
        RECT 45.165 160.875 45.455 160.920 ;
        RECT 56.650 160.860 56.970 161.120 ;
        RECT 64.100 161.060 64.240 161.940 ;
        RECT 67.690 161.895 68.040 162.125 ;
        RECT 68.610 162.080 68.930 162.140 ;
        RECT 71.920 162.125 72.060 162.280 ;
        RECT 68.610 161.940 70.220 162.080 ;
        RECT 67.690 161.880 68.010 161.895 ;
        RECT 68.610 161.880 68.930 161.940 ;
        RECT 64.495 161.740 64.785 161.785 ;
        RECT 67.015 161.740 67.305 161.785 ;
        RECT 68.205 161.740 68.495 161.785 ;
        RECT 64.495 161.600 68.495 161.740 ;
        RECT 64.495 161.555 64.785 161.600 ;
        RECT 67.015 161.555 67.305 161.600 ;
        RECT 68.205 161.555 68.495 161.600 ;
        RECT 69.085 161.740 69.375 161.785 ;
        RECT 69.530 161.740 69.850 161.800 ;
        RECT 69.085 161.600 69.850 161.740 ;
        RECT 70.080 161.740 70.220 161.940 ;
        RECT 71.845 161.895 72.135 162.125 ;
        RECT 72.290 161.880 72.610 162.140 ;
        RECT 72.840 162.125 72.980 162.280 ;
        RECT 73.760 162.125 73.900 162.620 ;
        RECT 74.590 162.420 74.910 162.480 ;
        RECT 74.590 162.280 76.660 162.420 ;
        RECT 74.590 162.220 74.910 162.280 ;
        RECT 72.765 161.895 73.055 162.125 ;
        RECT 73.685 161.895 73.975 162.125 ;
        RECT 75.050 162.080 75.370 162.140 ;
        RECT 76.520 162.125 76.660 162.280 ;
        RECT 77.440 162.125 77.580 162.620 ;
        RECT 78.270 162.420 78.590 162.480 ;
        RECT 79.205 162.420 79.495 162.465 ;
        RECT 78.270 162.280 79.495 162.420 ;
        RECT 78.270 162.220 78.590 162.280 ;
        RECT 79.205 162.235 79.495 162.280 ;
        RECT 75.525 162.080 75.815 162.125 ;
        RECT 75.050 161.940 75.815 162.080 ;
        RECT 73.210 161.740 73.530 161.800 ;
        RECT 70.080 161.600 73.530 161.740 ;
        RECT 69.085 161.555 69.375 161.600 ;
        RECT 69.530 161.540 69.850 161.600 ;
        RECT 73.210 161.540 73.530 161.600 ;
        RECT 73.760 161.740 73.900 161.895 ;
        RECT 75.050 161.880 75.370 161.940 ;
        RECT 75.525 161.895 75.815 161.940 ;
        RECT 75.985 161.895 76.275 162.125 ;
        RECT 76.445 161.895 76.735 162.125 ;
        RECT 77.365 161.895 77.655 162.125 ;
        RECT 78.745 162.080 79.035 162.125 ;
        RECT 78.360 161.940 79.035 162.080 ;
        RECT 74.130 161.740 74.450 161.800 ;
        RECT 73.760 161.600 74.450 161.740 ;
        RECT 64.930 161.400 65.220 161.445 ;
        RECT 66.500 161.400 66.790 161.445 ;
        RECT 68.600 161.400 68.890 161.445 ;
        RECT 73.760 161.400 73.900 161.600 ;
        RECT 74.130 161.540 74.450 161.600 ;
        RECT 64.930 161.260 68.890 161.400 ;
        RECT 64.930 161.215 65.220 161.260 ;
        RECT 66.500 161.215 66.790 161.260 ;
        RECT 68.600 161.215 68.890 161.260 ;
        RECT 70.080 161.260 73.900 161.400 ;
        RECT 75.510 161.400 75.830 161.460 ;
        RECT 76.060 161.400 76.200 161.895 ;
        RECT 78.360 161.800 78.500 161.940 ;
        RECT 78.745 161.895 79.035 161.940 ;
        RECT 79.280 161.800 79.420 162.235 ;
        RECT 79.650 161.880 79.970 162.140 ;
        RECT 80.585 161.895 80.875 162.125 ;
        RECT 78.270 161.540 78.590 161.800 ;
        RECT 79.190 161.540 79.510 161.800 ;
        RECT 80.660 161.400 80.800 161.895 ;
        RECT 75.510 161.260 76.200 161.400 ;
        RECT 76.520 161.260 80.800 161.400 ;
        RECT 70.080 161.060 70.220 161.260 ;
        RECT 75.510 161.200 75.830 161.260 ;
        RECT 64.100 160.920 70.220 161.060 ;
        RECT 70.450 160.860 70.770 161.120 ;
        RECT 71.830 161.060 72.150 161.120 ;
        RECT 74.145 161.060 74.435 161.105 ;
        RECT 71.830 160.920 74.435 161.060 ;
        RECT 71.830 160.860 72.150 160.920 ;
        RECT 74.145 160.875 74.435 160.920 ;
        RECT 74.590 161.060 74.910 161.120 ;
        RECT 76.520 161.060 76.660 161.260 ;
        RECT 74.590 160.920 76.660 161.060 ;
        RECT 74.590 160.860 74.910 160.920 ;
        RECT 77.810 160.860 78.130 161.120 ;
        RECT 5.520 160.240 83.260 160.720 ;
        RECT 39.185 160.040 39.475 160.085 ;
        RECT 40.550 160.040 40.870 160.100 ;
        RECT 39.185 159.900 40.870 160.040 ;
        RECT 39.185 159.855 39.475 159.900 ;
        RECT 40.550 159.840 40.870 159.900 ;
        RECT 44.705 160.040 44.995 160.085 ;
        RECT 45.610 160.040 45.930 160.100 ;
        RECT 44.705 159.900 45.930 160.040 ;
        RECT 44.705 159.855 44.995 159.900 ;
        RECT 32.770 159.700 33.060 159.745 ;
        RECT 34.870 159.700 35.160 159.745 ;
        RECT 36.440 159.700 36.730 159.745 ;
        RECT 32.770 159.560 36.730 159.700 ;
        RECT 32.770 159.515 33.060 159.560 ;
        RECT 34.870 159.515 35.160 159.560 ;
        RECT 36.440 159.515 36.730 159.560 ;
        RECT 33.165 159.360 33.455 159.405 ;
        RECT 34.355 159.360 34.645 159.405 ;
        RECT 36.875 159.360 37.165 159.405 ;
        RECT 33.165 159.220 37.165 159.360 ;
        RECT 33.165 159.175 33.455 159.220 ;
        RECT 34.355 159.175 34.645 159.220 ;
        RECT 36.875 159.175 37.165 159.220 ;
        RECT 41.930 159.160 42.250 159.420 ;
        RECT 32.285 159.020 32.575 159.065 ;
        RECT 32.285 158.880 34.570 159.020 ;
        RECT 32.285 158.835 32.575 158.880 ;
        RECT 34.430 158.740 34.570 158.880 ;
        RECT 40.550 158.820 40.870 159.080 ;
        RECT 42.390 159.020 42.710 159.080 ;
        RECT 42.865 159.020 43.155 159.065 ;
        RECT 42.390 158.880 43.155 159.020 ;
        RECT 42.390 158.820 42.710 158.880 ;
        RECT 42.865 158.835 43.155 158.880 ;
        RECT 43.325 159.020 43.615 159.065 ;
        RECT 44.780 159.020 44.920 159.855 ;
        RECT 45.610 159.840 45.930 159.900 ;
        RECT 57.570 160.040 57.890 160.100 ;
        RECT 60.805 160.040 61.095 160.085 ;
        RECT 68.610 160.040 68.930 160.100 ;
        RECT 57.570 159.900 68.930 160.040 ;
        RECT 57.570 159.840 57.890 159.900 ;
        RECT 60.805 159.855 61.095 159.900 ;
        RECT 68.610 159.840 68.930 159.900 ;
        RECT 69.070 159.840 69.390 160.100 ;
        RECT 76.890 160.040 77.210 160.100 ;
        RECT 77.365 160.040 77.655 160.085 ;
        RECT 76.890 159.900 77.655 160.040 ;
        RECT 76.890 159.840 77.210 159.900 ;
        RECT 77.365 159.855 77.655 159.900 ;
        RECT 48.870 159.700 49.160 159.745 ;
        RECT 50.970 159.700 51.260 159.745 ;
        RECT 52.540 159.700 52.830 159.745 ;
        RECT 48.870 159.560 52.830 159.700 ;
        RECT 48.870 159.515 49.160 159.560 ;
        RECT 50.970 159.515 51.260 159.560 ;
        RECT 52.540 159.515 52.830 159.560 ;
        RECT 53.890 159.700 54.210 159.760 ;
        RECT 54.810 159.700 55.130 159.760 ;
        RECT 55.285 159.700 55.575 159.745 ;
        RECT 53.890 159.560 55.575 159.700 ;
        RECT 53.890 159.500 54.210 159.560 ;
        RECT 54.810 159.500 55.130 159.560 ;
        RECT 55.285 159.515 55.575 159.560 ;
        RECT 55.745 159.515 56.035 159.745 ;
        RECT 63.550 159.700 63.840 159.745 ;
        RECT 65.120 159.700 65.410 159.745 ;
        RECT 67.220 159.700 67.510 159.745 ;
        RECT 63.550 159.560 67.510 159.700 ;
        RECT 63.550 159.515 63.840 159.560 ;
        RECT 65.120 159.515 65.410 159.560 ;
        RECT 67.220 159.515 67.510 159.560 ;
        RECT 70.950 159.700 71.240 159.745 ;
        RECT 73.050 159.700 73.340 159.745 ;
        RECT 74.620 159.700 74.910 159.745 ;
        RECT 70.950 159.560 74.910 159.700 ;
        RECT 70.950 159.515 71.240 159.560 ;
        RECT 73.050 159.515 73.340 159.560 ;
        RECT 74.620 159.515 74.910 159.560 ;
        RECT 80.110 159.700 80.430 159.760 ;
        RECT 81.045 159.700 81.335 159.745 ;
        RECT 80.110 159.560 81.335 159.700 ;
        RECT 49.265 159.360 49.555 159.405 ;
        RECT 50.455 159.360 50.745 159.405 ;
        RECT 52.975 159.360 53.265 159.405 ;
        RECT 49.265 159.220 53.265 159.360 ;
        RECT 49.265 159.175 49.555 159.220 ;
        RECT 50.455 159.175 50.745 159.220 ;
        RECT 52.975 159.175 53.265 159.220 ;
        RECT 43.325 158.880 44.920 159.020 ;
        RECT 46.990 159.020 47.310 159.080 ;
        RECT 47.465 159.020 47.755 159.065 ;
        RECT 46.990 158.880 47.755 159.020 ;
        RECT 43.325 158.835 43.615 158.880 ;
        RECT 46.990 158.820 47.310 158.880 ;
        RECT 47.465 158.835 47.755 158.880 ;
        RECT 48.370 158.820 48.690 159.080 ;
        RECT 49.720 159.020 50.010 159.065 ;
        RECT 55.820 159.020 55.960 159.515 ;
        RECT 80.110 159.500 80.430 159.560 ;
        RECT 81.045 159.515 81.335 159.560 ;
        RECT 56.650 159.360 56.970 159.420 ;
        RECT 58.045 159.360 58.335 159.405 ;
        RECT 56.650 159.220 58.335 159.360 ;
        RECT 56.650 159.160 56.970 159.220 ;
        RECT 58.045 159.175 58.335 159.220 ;
        RECT 58.505 159.175 58.795 159.405 ;
        RECT 63.115 159.360 63.405 159.405 ;
        RECT 65.635 159.360 65.925 159.405 ;
        RECT 66.825 159.360 67.115 159.405 ;
        RECT 71.345 159.360 71.635 159.405 ;
        RECT 72.535 159.360 72.825 159.405 ;
        RECT 75.055 159.360 75.345 159.405 ;
        RECT 79.650 159.360 79.970 159.420 ;
        RECT 81.950 159.360 82.270 159.420 ;
        RECT 63.115 159.220 67.115 159.360 ;
        RECT 63.115 159.175 63.405 159.220 ;
        RECT 65.635 159.175 65.925 159.220 ;
        RECT 66.825 159.175 67.115 159.220 ;
        RECT 67.825 159.220 68.840 159.360 ;
        RECT 58.580 159.020 58.720 159.175 ;
        RECT 67.825 159.065 67.965 159.220 ;
        RECT 68.700 159.080 68.840 159.220 ;
        RECT 71.345 159.220 75.345 159.360 ;
        RECT 71.345 159.175 71.635 159.220 ;
        RECT 72.535 159.175 72.825 159.220 ;
        RECT 75.055 159.175 75.345 159.220 ;
        RECT 79.280 159.220 82.270 159.360 ;
        RECT 49.720 158.880 55.960 159.020 ;
        RECT 56.280 158.880 58.720 159.020 ;
        RECT 49.720 158.835 50.010 158.880 ;
        RECT 33.650 158.725 33.970 158.740 ;
        RECT 33.620 158.495 33.970 158.725 ;
        RECT 34.430 158.540 34.890 158.740 ;
        RECT 33.650 158.480 33.970 158.495 ;
        RECT 34.570 158.480 34.890 158.540 ;
        RECT 41.485 158.680 41.775 158.725 ;
        RECT 44.230 158.680 44.550 158.740 ;
        RECT 41.485 158.540 44.550 158.680 ;
        RECT 41.485 158.495 41.775 158.540 ;
        RECT 44.230 158.480 44.550 158.540 ;
        RECT 53.430 158.680 53.750 158.740 ;
        RECT 56.280 158.680 56.420 158.880 ;
        RECT 67.705 158.835 67.995 159.065 ;
        RECT 68.165 158.835 68.455 159.065 ;
        RECT 68.610 159.020 68.930 159.080 ;
        RECT 69.530 159.020 69.850 159.080 ;
        RECT 70.465 159.020 70.755 159.065 ;
        RECT 74.590 159.020 74.910 159.080 ;
        RECT 75.510 159.020 75.830 159.080 ;
        RECT 68.610 158.880 74.910 159.020 ;
        RECT 53.430 158.540 56.420 158.680 ;
        RECT 65.390 158.680 65.710 158.740 ;
        RECT 66.370 158.680 66.660 158.725 ;
        RECT 65.390 158.540 66.660 158.680 ;
        RECT 53.430 158.480 53.750 158.540 ;
        RECT 65.390 158.480 65.710 158.540 ;
        RECT 66.370 158.495 66.660 158.540 ;
        RECT 68.240 158.400 68.380 158.835 ;
        RECT 68.610 158.820 68.930 158.880 ;
        RECT 69.530 158.820 69.850 158.880 ;
        RECT 70.465 158.835 70.755 158.880 ;
        RECT 74.590 158.820 74.910 158.880 ;
        RECT 75.140 158.880 75.830 159.020 ;
        RECT 71.830 158.725 72.150 158.740 ;
        RECT 71.800 158.495 72.150 158.725 ;
        RECT 71.830 158.480 72.150 158.495 ;
        RECT 72.290 158.680 72.610 158.740 ;
        RECT 75.140 158.680 75.280 158.880 ;
        RECT 75.510 158.820 75.830 158.880 ;
        RECT 75.970 159.020 76.290 159.080 ;
        RECT 79.280 159.065 79.420 159.220 ;
        RECT 79.650 159.160 79.970 159.220 ;
        RECT 81.950 159.160 82.270 159.220 ;
        RECT 78.285 159.020 78.575 159.065 ;
        RECT 75.970 158.880 78.575 159.020 ;
        RECT 75.970 158.820 76.290 158.880 ;
        RECT 78.285 158.835 78.575 158.880 ;
        RECT 79.205 158.835 79.495 159.065 ;
        RECT 80.125 159.020 80.415 159.065 ;
        RECT 80.570 159.020 80.890 159.080 ;
        RECT 80.125 158.880 80.890 159.020 ;
        RECT 80.125 158.835 80.415 158.880 ;
        RECT 80.570 158.820 80.890 158.880 ;
        RECT 72.290 158.540 75.280 158.680 ;
        RECT 72.290 158.480 72.610 158.540 ;
        RECT 79.665 158.495 79.955 158.725 ;
        RECT 39.630 158.140 39.950 158.400 ;
        RECT 41.945 158.340 42.235 158.385 ;
        RECT 42.390 158.340 42.710 158.400 ;
        RECT 41.945 158.200 42.710 158.340 ;
        RECT 41.945 158.155 42.235 158.200 ;
        RECT 42.390 158.140 42.710 158.200 ;
        RECT 57.570 158.140 57.890 158.400 ;
        RECT 68.150 158.140 68.470 158.400 ;
        RECT 79.740 158.340 79.880 158.495 ;
        RECT 80.570 158.340 80.890 158.400 ;
        RECT 79.740 158.200 80.890 158.340 ;
        RECT 80.570 158.140 80.890 158.200 ;
        RECT 5.520 157.520 83.260 158.000 ;
        RECT 36.870 157.320 37.190 157.380 ;
        RECT 37.345 157.320 37.635 157.365 ;
        RECT 36.870 157.180 37.635 157.320 ;
        RECT 36.870 157.120 37.190 157.180 ;
        RECT 37.345 157.135 37.635 157.180 ;
        RECT 55.285 157.320 55.575 157.365 ;
        RECT 56.190 157.320 56.510 157.380 ;
        RECT 60.330 157.320 60.650 157.380 ;
        RECT 55.285 157.180 60.650 157.320 ;
        RECT 55.285 157.135 55.575 157.180 ;
        RECT 56.190 157.120 56.510 157.180 ;
        RECT 60.330 157.120 60.650 157.180 ;
        RECT 71.370 157.320 71.690 157.380 ;
        RECT 74.605 157.320 74.895 157.365 ;
        RECT 71.370 157.180 74.895 157.320 ;
        RECT 71.370 157.120 71.690 157.180 ;
        RECT 74.605 157.135 74.895 157.180 ;
        RECT 39.630 156.980 39.950 157.040 ;
        RECT 40.565 156.980 40.855 157.025 ;
        RECT 68.610 156.980 68.930 157.040 ;
        RECT 39.630 156.840 40.855 156.980 ;
        RECT 39.630 156.780 39.950 156.840 ;
        RECT 40.565 156.795 40.855 156.840 ;
        RECT 64.560 156.840 68.930 156.980 ;
        RECT 35.490 156.640 35.810 156.700 ;
        RECT 37.790 156.640 38.110 156.700 ;
        RECT 42.390 156.685 42.710 156.700 ;
        RECT 38.725 156.640 39.015 156.685 ;
        RECT 42.360 156.640 42.710 156.685 ;
        RECT 35.490 156.500 39.015 156.640 ;
        RECT 42.195 156.500 42.710 156.640 ;
        RECT 35.490 156.440 35.810 156.500 ;
        RECT 37.790 156.440 38.110 156.500 ;
        RECT 38.725 156.455 39.015 156.500 ;
        RECT 42.360 156.455 42.710 156.500 ;
        RECT 42.390 156.440 42.710 156.455 ;
        RECT 48.370 156.440 48.690 156.700 ;
        RECT 49.750 156.685 50.070 156.700 ;
        RECT 49.720 156.455 50.070 156.685 ;
        RECT 49.750 156.440 50.070 156.455 ;
        RECT 61.710 156.640 62.030 156.700 ;
        RECT 64.560 156.685 64.700 156.840 ;
        RECT 63.150 156.640 63.440 156.685 ;
        RECT 61.710 156.500 63.440 156.640 ;
        RECT 61.710 156.440 62.030 156.500 ;
        RECT 63.150 156.455 63.440 156.500 ;
        RECT 64.485 156.455 64.775 156.685 ;
        RECT 64.930 156.440 65.250 156.700 ;
        RECT 67.780 156.685 67.920 156.840 ;
        RECT 68.610 156.780 68.930 156.840 ;
        RECT 70.910 156.980 71.230 157.040 ;
        RECT 75.065 156.980 75.355 157.025 ;
        RECT 70.910 156.840 75.355 156.980 ;
        RECT 70.910 156.780 71.230 156.840 ;
        RECT 75.065 156.795 75.355 156.840 ;
        RECT 66.785 156.455 67.075 156.685 ;
        RECT 67.705 156.455 67.995 156.685 ;
        RECT 30.430 156.300 30.750 156.360 ;
        RECT 36.425 156.300 36.715 156.345 ;
        RECT 30.430 156.160 36.715 156.300 ;
        RECT 30.430 156.100 30.750 156.160 ;
        RECT 36.425 156.115 36.715 156.160 ;
        RECT 38.250 156.100 38.570 156.360 ;
        RECT 40.090 156.100 40.410 156.360 ;
        RECT 41.025 156.115 41.315 156.345 ;
        RECT 41.905 156.300 42.195 156.345 ;
        RECT 43.095 156.300 43.385 156.345 ;
        RECT 45.615 156.300 45.905 156.345 ;
        RECT 41.905 156.160 45.905 156.300 ;
        RECT 41.905 156.115 42.195 156.160 ;
        RECT 43.095 156.115 43.385 156.160 ;
        RECT 45.615 156.115 45.905 156.160 ;
        RECT 49.265 156.300 49.555 156.345 ;
        RECT 50.455 156.300 50.745 156.345 ;
        RECT 52.975 156.300 53.265 156.345 ;
        RECT 49.265 156.160 53.265 156.300 ;
        RECT 49.265 156.115 49.555 156.160 ;
        RECT 50.455 156.115 50.745 156.160 ;
        RECT 52.975 156.115 53.265 156.160 ;
        RECT 59.895 156.300 60.185 156.345 ;
        RECT 62.415 156.300 62.705 156.345 ;
        RECT 63.605 156.300 63.895 156.345 ;
        RECT 59.895 156.160 63.895 156.300 ;
        RECT 66.860 156.300 67.000 156.455 ;
        RECT 68.150 156.440 68.470 156.700 ;
        RECT 69.040 156.640 69.330 156.685 ;
        RECT 70.450 156.640 70.770 156.700 ;
        RECT 69.040 156.500 70.770 156.640 ;
        RECT 69.040 156.455 69.330 156.500 ;
        RECT 70.450 156.440 70.770 156.500 ;
        RECT 75.970 156.440 76.290 156.700 ;
        RECT 81.490 156.440 81.810 156.700 ;
        RECT 68.240 156.300 68.380 156.440 ;
        RECT 66.860 156.160 68.380 156.300 ;
        RECT 68.585 156.300 68.875 156.345 ;
        RECT 69.775 156.300 70.065 156.345 ;
        RECT 72.295 156.300 72.585 156.345 ;
        RECT 68.585 156.160 72.585 156.300 ;
        RECT 59.895 156.115 60.185 156.160 ;
        RECT 62.415 156.115 62.705 156.160 ;
        RECT 63.605 156.115 63.895 156.160 ;
        RECT 68.585 156.115 68.875 156.160 ;
        RECT 69.775 156.115 70.065 156.160 ;
        RECT 72.295 156.115 72.585 156.160 ;
        RECT 76.890 156.300 77.210 156.360 ;
        RECT 80.125 156.300 80.415 156.345 ;
        RECT 76.890 156.160 80.415 156.300 ;
        RECT 34.570 155.960 34.890 156.020 ;
        RECT 41.100 155.960 41.240 156.115 ;
        RECT 76.890 156.100 77.210 156.160 ;
        RECT 80.125 156.115 80.415 156.160 ;
        RECT 34.570 155.820 41.240 155.960 ;
        RECT 41.510 155.960 41.800 156.005 ;
        RECT 43.610 155.960 43.900 156.005 ;
        RECT 45.180 155.960 45.470 156.005 ;
        RECT 41.510 155.820 45.470 155.960 ;
        RECT 34.570 155.760 34.890 155.820 ;
        RECT 41.510 155.775 41.800 155.820 ;
        RECT 43.610 155.775 43.900 155.820 ;
        RECT 45.180 155.775 45.470 155.820 ;
        RECT 48.870 155.960 49.160 156.005 ;
        RECT 50.970 155.960 51.260 156.005 ;
        RECT 52.540 155.960 52.830 156.005 ;
        RECT 48.870 155.820 52.830 155.960 ;
        RECT 48.870 155.775 49.160 155.820 ;
        RECT 50.970 155.775 51.260 155.820 ;
        RECT 52.540 155.775 52.830 155.820 ;
        RECT 60.330 155.960 60.620 156.005 ;
        RECT 61.900 155.960 62.190 156.005 ;
        RECT 64.000 155.960 64.290 156.005 ;
        RECT 68.190 155.960 68.480 156.005 ;
        RECT 70.290 155.960 70.580 156.005 ;
        RECT 71.860 155.960 72.150 156.005 ;
        RECT 79.190 155.960 79.510 156.020 ;
        RECT 81.490 155.960 81.810 156.020 ;
        RECT 60.330 155.820 64.290 155.960 ;
        RECT 60.330 155.775 60.620 155.820 ;
        RECT 61.900 155.775 62.190 155.820 ;
        RECT 64.000 155.775 64.290 155.820 ;
        RECT 65.020 155.820 67.920 155.960 ;
        RECT 33.650 155.420 33.970 155.680 ;
        RECT 46.990 155.620 47.310 155.680 ;
        RECT 47.925 155.620 48.215 155.665 ;
        RECT 46.990 155.480 48.215 155.620 ;
        RECT 46.990 155.420 47.310 155.480 ;
        RECT 47.925 155.435 48.215 155.480 ;
        RECT 57.585 155.620 57.875 155.665 ;
        RECT 59.410 155.620 59.730 155.680 ;
        RECT 57.585 155.480 59.730 155.620 ;
        RECT 57.585 155.435 57.875 155.480 ;
        RECT 59.410 155.420 59.730 155.480 ;
        RECT 59.870 155.620 60.190 155.680 ;
        RECT 65.020 155.620 65.160 155.820 ;
        RECT 59.870 155.480 65.160 155.620 ;
        RECT 67.780 155.620 67.920 155.820 ;
        RECT 68.190 155.820 72.150 155.960 ;
        RECT 68.190 155.775 68.480 155.820 ;
        RECT 70.290 155.775 70.580 155.820 ;
        RECT 71.860 155.775 72.150 155.820 ;
        RECT 76.520 155.820 81.810 155.960 ;
        RECT 76.520 155.620 76.660 155.820 ;
        RECT 79.190 155.760 79.510 155.820 ;
        RECT 81.490 155.760 81.810 155.820 ;
        RECT 67.780 155.480 76.660 155.620 ;
        RECT 76.905 155.620 77.195 155.665 ;
        RECT 78.730 155.620 79.050 155.680 ;
        RECT 76.905 155.480 79.050 155.620 ;
        RECT 59.870 155.420 60.190 155.480 ;
        RECT 76.905 155.435 77.195 155.480 ;
        RECT 78.730 155.420 79.050 155.480 ;
        RECT 5.520 154.800 83.260 155.280 ;
        RECT 30.430 154.400 30.750 154.660 ;
        RECT 40.090 154.600 40.410 154.660 ;
        RECT 44.705 154.600 44.995 154.645 ;
        RECT 40.090 154.460 44.995 154.600 ;
        RECT 40.090 154.400 40.410 154.460 ;
        RECT 44.705 154.415 44.995 154.460 ;
        RECT 49.290 154.400 49.610 154.660 ;
        RECT 49.750 154.600 50.070 154.660 ;
        RECT 50.685 154.600 50.975 154.645 ;
        RECT 49.750 154.460 50.975 154.600 ;
        RECT 49.750 154.400 50.070 154.460 ;
        RECT 50.685 154.415 50.975 154.460 ;
        RECT 59.410 154.600 59.730 154.660 ;
        RECT 59.410 154.460 69.300 154.600 ;
        RECT 59.410 154.400 59.730 154.460 ;
        RECT 33.190 154.260 33.480 154.305 ;
        RECT 34.760 154.260 35.050 154.305 ;
        RECT 36.860 154.260 37.150 154.305 ;
        RECT 42.390 154.260 42.710 154.320 ;
        RECT 33.190 154.120 37.150 154.260 ;
        RECT 33.190 154.075 33.480 154.120 ;
        RECT 34.760 154.075 35.050 154.120 ;
        RECT 36.860 154.075 37.150 154.120 ;
        RECT 38.800 154.120 42.710 154.260 ;
        RECT 32.755 153.920 33.045 153.965 ;
        RECT 35.275 153.920 35.565 153.965 ;
        RECT 36.465 153.920 36.755 153.965 ;
        RECT 32.755 153.780 36.755 153.920 ;
        RECT 32.755 153.735 33.045 153.780 ;
        RECT 35.275 153.735 35.565 153.780 ;
        RECT 36.465 153.735 36.755 153.780 ;
        RECT 32.270 153.580 32.590 153.640 ;
        RECT 34.570 153.580 34.890 153.640 ;
        RECT 37.330 153.580 37.650 153.640 ;
        RECT 38.800 153.625 38.940 154.120 ;
        RECT 42.390 154.060 42.710 154.120 ;
        RECT 48.370 154.260 48.690 154.320 ;
        RECT 55.310 154.260 55.600 154.305 ;
        RECT 57.410 154.260 57.700 154.305 ;
        RECT 58.980 154.260 59.270 154.305 ;
        RECT 48.370 154.120 55.040 154.260 ;
        RECT 48.370 154.060 48.690 154.120 ;
        RECT 41.485 153.920 41.775 153.965 ;
        RECT 41.485 153.780 46.300 153.920 ;
        RECT 41.485 153.735 41.775 153.780 ;
        RECT 46.160 153.640 46.300 153.780 ;
        RECT 49.750 153.720 50.070 153.980 ;
        RECT 51.130 153.920 51.450 153.980 ;
        RECT 53.430 153.920 53.750 153.980 ;
        RECT 54.900 153.965 55.040 154.120 ;
        RECT 55.310 154.120 59.270 154.260 ;
        RECT 55.310 154.075 55.600 154.120 ;
        RECT 57.410 154.075 57.700 154.120 ;
        RECT 58.980 154.075 59.270 154.120 ;
        RECT 62.185 154.075 62.475 154.305 ;
        RECT 51.130 153.780 53.750 153.920 ;
        RECT 51.130 153.720 51.450 153.780 ;
        RECT 53.430 153.720 53.750 153.780 ;
        RECT 54.825 153.735 55.115 153.965 ;
        RECT 55.705 153.920 55.995 153.965 ;
        RECT 56.895 153.920 57.185 153.965 ;
        RECT 59.415 153.920 59.705 153.965 ;
        RECT 55.705 153.780 59.705 153.920 ;
        RECT 55.705 153.735 55.995 153.780 ;
        RECT 56.895 153.735 57.185 153.780 ;
        RECT 59.415 153.735 59.705 153.780 ;
        RECT 32.270 153.440 37.650 153.580 ;
        RECT 32.270 153.380 32.590 153.440 ;
        RECT 34.570 153.380 34.890 153.440 ;
        RECT 37.330 153.380 37.650 153.440 ;
        RECT 38.265 153.395 38.555 153.625 ;
        RECT 38.725 153.395 39.015 153.625 ;
        RECT 39.645 153.580 39.935 153.625 ;
        RECT 41.025 153.580 41.315 153.625 ;
        RECT 39.645 153.440 41.315 153.580 ;
        RECT 39.645 153.395 39.935 153.440 ;
        RECT 41.025 153.395 41.315 153.440 ;
        RECT 35.030 153.240 35.350 153.300 ;
        RECT 36.010 153.240 36.300 153.285 ;
        RECT 35.030 153.100 36.300 153.240 ;
        RECT 38.340 153.240 38.480 153.395 ;
        RECT 41.930 153.380 42.250 153.640 ;
        RECT 42.390 153.380 42.710 153.640 ;
        RECT 43.325 153.580 43.615 153.625 ;
        RECT 44.230 153.580 44.550 153.640 ;
        RECT 43.325 153.440 44.550 153.580 ;
        RECT 43.325 153.395 43.615 153.440 ;
        RECT 44.230 153.380 44.550 153.440 ;
        RECT 45.610 153.380 45.930 153.640 ;
        RECT 46.070 153.380 46.390 153.640 ;
        RECT 47.005 153.395 47.295 153.625 ;
        RECT 42.020 153.240 42.160 153.380 ;
        RECT 47.080 153.240 47.220 153.395 ;
        RECT 47.450 153.380 47.770 153.640 ;
        RECT 48.845 153.580 49.135 153.625 ;
        RECT 50.670 153.580 50.990 153.640 ;
        RECT 48.845 153.440 50.990 153.580 ;
        RECT 48.845 153.395 49.135 153.440 ;
        RECT 50.670 153.380 50.990 153.440 ;
        RECT 52.525 153.580 52.815 153.625 ;
        RECT 62.260 153.580 62.400 154.075 ;
        RECT 63.550 153.920 63.870 153.980 ;
        RECT 69.160 153.965 69.300 154.460 ;
        RECT 81.490 154.400 81.810 154.660 ;
        RECT 72.750 154.060 73.070 154.320 ;
        RECT 75.090 154.260 75.380 154.305 ;
        RECT 77.190 154.260 77.480 154.305 ;
        RECT 78.760 154.260 79.050 154.305 ;
        RECT 75.090 154.120 79.050 154.260 ;
        RECT 75.090 154.075 75.380 154.120 ;
        RECT 77.190 154.075 77.480 154.120 ;
        RECT 78.760 154.075 79.050 154.120 ;
        RECT 64.945 153.920 65.235 153.965 ;
        RECT 63.550 153.780 65.235 153.920 ;
        RECT 63.550 153.720 63.870 153.780 ;
        RECT 64.945 153.735 65.235 153.780 ;
        RECT 69.085 153.735 69.375 153.965 ;
        RECT 72.840 153.920 72.980 154.060 ;
        RECT 75.485 153.920 75.775 153.965 ;
        RECT 76.675 153.920 76.965 153.965 ;
        RECT 79.195 153.920 79.485 153.965 ;
        RECT 69.620 153.780 73.900 153.920 ;
        RECT 52.525 153.440 62.400 153.580 ;
        RECT 63.090 153.580 63.410 153.640 ;
        RECT 69.620 153.580 69.760 153.780 ;
        RECT 63.090 153.440 69.760 153.580 ;
        RECT 69.990 153.580 70.310 153.640 ;
        RECT 71.830 153.580 72.150 153.640 ;
        RECT 69.990 153.440 72.150 153.580 ;
        RECT 52.525 153.395 52.815 153.440 ;
        RECT 63.090 153.380 63.410 153.440 ;
        RECT 69.990 153.380 70.310 153.440 ;
        RECT 71.830 153.380 72.150 153.440 ;
        RECT 72.305 153.395 72.595 153.625 ;
        RECT 72.765 153.580 73.055 153.625 ;
        RECT 73.210 153.580 73.530 153.640 ;
        RECT 73.760 153.625 73.900 153.780 ;
        RECT 75.485 153.780 79.485 153.920 ;
        RECT 75.485 153.735 75.775 153.780 ;
        RECT 76.675 153.735 76.965 153.780 ;
        RECT 79.195 153.735 79.485 153.780 ;
        RECT 72.765 153.440 73.530 153.580 ;
        RECT 72.765 153.395 73.055 153.440 ;
        RECT 38.340 153.100 41.700 153.240 ;
        RECT 42.020 153.100 47.220 153.240 ;
        RECT 50.225 153.240 50.515 153.285 ;
        RECT 52.050 153.240 52.370 153.300 ;
        RECT 50.225 153.100 52.370 153.240 ;
        RECT 35.030 153.040 35.350 153.100 ;
        RECT 36.010 153.055 36.300 153.100 ;
        RECT 40.090 152.700 40.410 152.960 ;
        RECT 41.560 152.900 41.700 153.100 ;
        RECT 50.225 153.055 50.515 153.100 ;
        RECT 52.050 153.040 52.370 153.100 ;
        RECT 52.985 153.240 53.275 153.285 ;
        RECT 55.270 153.240 55.590 153.300 ;
        RECT 52.985 153.100 55.590 153.240 ;
        RECT 52.985 153.055 53.275 153.100 ;
        RECT 55.270 153.040 55.590 153.100 ;
        RECT 56.160 153.240 56.450 153.285 ;
        RECT 58.950 153.240 59.270 153.300 ;
        RECT 64.010 153.240 64.330 153.300 ;
        RECT 56.160 153.100 59.270 153.240 ;
        RECT 56.160 153.055 56.450 153.100 ;
        RECT 58.950 153.040 59.270 153.100 ;
        RECT 61.800 153.100 64.330 153.240 ;
        RECT 46.990 152.900 47.310 152.960 ;
        RECT 41.560 152.760 47.310 152.900 ;
        RECT 46.990 152.700 47.310 152.760 ;
        RECT 47.925 152.900 48.215 152.945 ;
        RECT 48.830 152.900 49.150 152.960 ;
        RECT 61.800 152.945 61.940 153.100 ;
        RECT 64.010 153.040 64.330 153.100 ;
        RECT 65.390 153.240 65.710 153.300 ;
        RECT 70.465 153.240 70.755 153.285 ;
        RECT 65.390 153.100 70.755 153.240 ;
        RECT 65.390 153.040 65.710 153.100 ;
        RECT 70.465 153.055 70.755 153.100 ;
        RECT 71.370 153.240 71.690 153.300 ;
        RECT 72.380 153.240 72.520 153.395 ;
        RECT 73.210 153.380 73.530 153.440 ;
        RECT 73.685 153.395 73.975 153.625 ;
        RECT 74.590 153.380 74.910 153.640 ;
        RECT 71.370 153.100 72.520 153.240 ;
        RECT 74.130 153.240 74.450 153.300 ;
        RECT 75.830 153.240 76.120 153.285 ;
        RECT 74.130 153.100 76.120 153.240 ;
        RECT 71.370 153.040 71.690 153.100 ;
        RECT 74.130 153.040 74.450 153.100 ;
        RECT 75.830 153.055 76.120 153.100 ;
        RECT 47.925 152.760 49.150 152.900 ;
        RECT 47.925 152.715 48.215 152.760 ;
        RECT 48.830 152.700 49.150 152.760 ;
        RECT 61.725 152.715 62.015 152.945 ;
        RECT 62.170 152.900 62.490 152.960 ;
        RECT 64.485 152.900 64.775 152.945 ;
        RECT 62.170 152.760 64.775 152.900 ;
        RECT 62.170 152.700 62.490 152.760 ;
        RECT 64.485 152.715 64.775 152.760 ;
        RECT 66.310 152.700 66.630 152.960 ;
        RECT 5.520 152.080 83.260 152.560 ;
        RECT 30.445 151.880 30.735 151.925 ;
        RECT 33.650 151.880 33.970 151.940 ;
        RECT 30.445 151.740 33.970 151.880 ;
        RECT 30.445 151.695 30.735 151.740 ;
        RECT 33.650 151.680 33.970 151.740 ;
        RECT 34.110 151.680 34.430 151.940 ;
        RECT 42.390 151.880 42.710 151.940 ;
        RECT 46.545 151.880 46.835 151.925 ;
        RECT 47.910 151.880 48.230 151.940 ;
        RECT 42.390 151.740 48.230 151.880 ;
        RECT 42.390 151.680 42.710 151.740 ;
        RECT 46.545 151.695 46.835 151.740 ;
        RECT 47.910 151.680 48.230 151.740 ;
        RECT 49.290 151.880 49.610 151.940 ;
        RECT 54.350 151.880 54.670 151.940 ;
        RECT 49.290 151.740 54.670 151.880 ;
        RECT 49.290 151.680 49.610 151.740 ;
        RECT 54.350 151.680 54.670 151.740 ;
        RECT 57.570 151.680 57.890 151.940 ;
        RECT 59.410 151.680 59.730 151.940 ;
        RECT 61.710 151.680 62.030 151.940 ;
        RECT 63.565 151.880 63.855 151.925 ;
        RECT 66.310 151.880 66.630 151.940 ;
        RECT 63.565 151.740 66.630 151.880 ;
        RECT 63.565 151.695 63.855 151.740 ;
        RECT 66.310 151.680 66.630 151.740 ;
        RECT 81.030 151.880 81.350 151.940 ;
        RECT 81.505 151.880 81.795 151.925 ;
        RECT 81.030 151.740 81.795 151.880 ;
        RECT 81.030 151.680 81.350 151.740 ;
        RECT 81.505 151.695 81.795 151.740 ;
        RECT 32.270 151.540 32.590 151.600 ;
        RECT 27.300 151.400 31.580 151.540 ;
        RECT 27.300 151.245 27.440 151.400 ;
        RECT 27.225 151.015 27.515 151.245 ;
        RECT 28.145 151.015 28.435 151.245 ;
        RECT 28.220 150.860 28.360 151.015 ;
        RECT 29.510 151.000 29.830 151.260 ;
        RECT 30.890 151.000 31.210 151.260 ;
        RECT 30.430 150.860 30.750 150.920 ;
        RECT 28.220 150.720 30.750 150.860 ;
        RECT 31.440 150.860 31.580 151.400 ;
        RECT 31.900 151.400 32.590 151.540 ;
        RECT 31.900 151.245 32.040 151.400 ;
        RECT 32.270 151.340 32.590 151.400 ;
        RECT 33.160 151.540 33.450 151.585 ;
        RECT 34.200 151.540 34.340 151.680 ;
        RECT 33.160 151.400 34.340 151.540 ;
        RECT 40.090 151.540 40.410 151.600 ;
        RECT 40.870 151.540 41.160 151.585 ;
        RECT 40.090 151.400 41.160 151.540 ;
        RECT 33.160 151.355 33.450 151.400 ;
        RECT 40.090 151.340 40.410 151.400 ;
        RECT 40.870 151.355 41.160 151.400 ;
        RECT 47.005 151.540 47.295 151.585 ;
        RECT 50.670 151.540 50.990 151.600 ;
        RECT 47.005 151.400 50.990 151.540 ;
        RECT 47.005 151.355 47.295 151.400 ;
        RECT 50.670 151.340 50.990 151.400 ;
        RECT 51.605 151.540 51.895 151.585 ;
        RECT 53.890 151.540 54.210 151.600 ;
        RECT 51.605 151.400 54.210 151.540 ;
        RECT 51.605 151.355 51.895 151.400 ;
        RECT 53.890 151.340 54.210 151.400 ;
        RECT 64.010 151.540 64.330 151.600 ;
        RECT 67.690 151.540 68.010 151.600 ;
        RECT 69.545 151.540 69.835 151.585 ;
        RECT 64.010 151.400 65.160 151.540 ;
        RECT 64.010 151.340 64.330 151.400 ;
        RECT 31.825 151.015 32.115 151.245 ;
        RECT 37.330 151.200 37.650 151.260 ;
        RECT 39.630 151.200 39.950 151.260 ;
        RECT 32.360 151.060 37.100 151.200 ;
        RECT 32.360 150.860 32.500 151.060 ;
        RECT 31.440 150.720 32.500 150.860 ;
        RECT 32.705 150.860 32.995 150.905 ;
        RECT 33.895 150.860 34.185 150.905 ;
        RECT 36.415 150.860 36.705 150.905 ;
        RECT 32.705 150.720 36.705 150.860 ;
        RECT 36.960 150.860 37.100 151.060 ;
        RECT 37.330 151.060 39.950 151.200 ;
        RECT 37.330 151.000 37.650 151.060 ;
        RECT 39.630 151.000 39.950 151.060 ;
        RECT 49.305 151.200 49.595 151.245 ;
        RECT 50.210 151.200 50.530 151.260 ;
        RECT 49.305 151.060 50.530 151.200 ;
        RECT 49.305 151.015 49.595 151.060 ;
        RECT 50.210 151.000 50.530 151.060 ;
        RECT 52.970 151.200 53.290 151.260 ;
        RECT 65.020 151.200 65.160 151.400 ;
        RECT 67.690 151.400 69.835 151.540 ;
        RECT 67.690 151.340 68.010 151.400 ;
        RECT 69.545 151.355 69.835 151.400 ;
        RECT 68.625 151.200 68.915 151.245 ;
        RECT 52.970 151.060 64.700 151.200 ;
        RECT 65.020 151.060 68.915 151.200 ;
        RECT 52.970 151.000 53.290 151.060 ;
        RECT 40.525 150.860 40.815 150.905 ;
        RECT 41.715 150.860 42.005 150.905 ;
        RECT 44.235 150.860 44.525 150.905 ;
        RECT 36.960 150.720 39.400 150.860 ;
        RECT 30.430 150.660 30.750 150.720 ;
        RECT 32.705 150.675 32.995 150.720 ;
        RECT 33.895 150.675 34.185 150.720 ;
        RECT 36.415 150.675 36.705 150.720 ;
        RECT 32.310 150.520 32.600 150.565 ;
        RECT 34.410 150.520 34.700 150.565 ;
        RECT 35.980 150.520 36.270 150.565 ;
        RECT 32.310 150.380 36.270 150.520 ;
        RECT 32.310 150.335 32.600 150.380 ;
        RECT 34.410 150.335 34.700 150.380 ;
        RECT 35.980 150.335 36.270 150.380 ;
        RECT 27.670 149.980 27.990 150.240 ;
        RECT 28.605 150.180 28.895 150.225 ;
        RECT 35.030 150.180 35.350 150.240 ;
        RECT 28.605 150.040 35.350 150.180 ;
        RECT 28.605 149.995 28.895 150.040 ;
        RECT 35.030 149.980 35.350 150.040 ;
        RECT 38.710 149.980 39.030 150.240 ;
        RECT 39.260 150.180 39.400 150.720 ;
        RECT 40.525 150.720 44.525 150.860 ;
        RECT 40.525 150.675 40.815 150.720 ;
        RECT 41.715 150.675 42.005 150.720 ;
        RECT 44.235 150.675 44.525 150.720 ;
        RECT 48.845 150.860 49.135 150.905 ;
        RECT 53.905 150.860 54.195 150.905 ;
        RECT 56.205 150.860 56.495 150.905 ;
        RECT 48.845 150.720 54.195 150.860 ;
        RECT 48.845 150.675 49.135 150.720 ;
        RECT 53.905 150.675 54.195 150.720 ;
        RECT 54.440 150.720 56.495 150.860 ;
        RECT 40.130 150.520 40.420 150.565 ;
        RECT 42.230 150.520 42.520 150.565 ;
        RECT 43.800 150.520 44.090 150.565 ;
        RECT 50.685 150.520 50.975 150.565 ;
        RECT 40.130 150.380 44.090 150.520 ;
        RECT 40.130 150.335 40.420 150.380 ;
        RECT 42.230 150.335 42.520 150.380 ;
        RECT 43.800 150.335 44.090 150.380 ;
        RECT 48.920 150.380 50.975 150.520 ;
        RECT 44.230 150.180 44.550 150.240 ;
        RECT 48.920 150.225 49.060 150.380 ;
        RECT 50.685 150.335 50.975 150.380 ;
        RECT 53.430 150.320 53.750 150.580 ;
        RECT 39.260 150.040 44.550 150.180 ;
        RECT 44.230 149.980 44.550 150.040 ;
        RECT 48.845 149.995 49.135 150.225 ;
        RECT 49.290 150.180 49.610 150.240 ;
        RECT 50.225 150.180 50.515 150.225 ;
        RECT 49.290 150.040 50.515 150.180 ;
        RECT 49.290 149.980 49.610 150.040 ;
        RECT 50.225 149.995 50.515 150.040 ;
        RECT 51.590 150.180 51.910 150.240 ;
        RECT 54.440 150.180 54.580 150.720 ;
        RECT 56.205 150.675 56.495 150.720 ;
        RECT 56.650 150.860 56.970 150.920 ;
        RECT 59.885 150.860 60.175 150.905 ;
        RECT 56.650 150.720 60.175 150.860 ;
        RECT 56.650 150.660 56.970 150.720 ;
        RECT 59.885 150.675 60.175 150.720 ;
        RECT 60.345 150.860 60.635 150.905 ;
        RECT 63.550 150.860 63.870 150.920 ;
        RECT 60.345 150.720 63.870 150.860 ;
        RECT 60.345 150.675 60.635 150.720 ;
        RECT 54.810 150.320 55.130 150.580 ;
        RECT 55.270 150.520 55.590 150.580 ;
        RECT 60.420 150.520 60.560 150.675 ;
        RECT 63.550 150.660 63.870 150.720 ;
        RECT 64.025 150.675 64.315 150.905 ;
        RECT 55.270 150.380 60.560 150.520 ;
        RECT 61.710 150.520 62.030 150.580 ;
        RECT 64.100 150.520 64.240 150.675 ;
        RECT 61.710 150.380 64.240 150.520 ;
        RECT 64.560 150.520 64.700 151.060 ;
        RECT 68.625 151.015 68.915 151.060 ;
        RECT 70.450 151.200 70.770 151.260 ;
        RECT 70.925 151.200 71.215 151.245 ;
        RECT 70.450 151.060 71.215 151.200 ;
        RECT 70.450 151.000 70.770 151.060 ;
        RECT 70.925 151.015 71.215 151.060 ;
        RECT 71.370 151.000 71.690 151.260 ;
        RECT 71.845 151.015 72.135 151.245 ;
        RECT 64.945 150.860 65.235 150.905 ;
        RECT 65.390 150.860 65.710 150.920 ;
        RECT 64.945 150.720 65.710 150.860 ;
        RECT 64.945 150.675 65.235 150.720 ;
        RECT 65.390 150.660 65.710 150.720 ;
        RECT 65.850 150.860 66.170 150.920 ;
        RECT 71.920 150.860 72.060 151.015 ;
        RECT 72.750 151.000 73.070 151.260 ;
        RECT 74.145 151.015 74.435 151.245 ;
        RECT 65.850 150.720 72.060 150.860 ;
        RECT 72.290 150.860 72.610 150.920 ;
        RECT 74.220 150.860 74.360 151.015 ;
        RECT 74.590 151.000 74.910 151.260 ;
        RECT 75.050 151.000 75.370 151.260 ;
        RECT 75.940 151.200 76.230 151.245 ;
        RECT 77.810 151.200 78.130 151.260 ;
        RECT 75.940 151.060 78.130 151.200 ;
        RECT 75.940 151.015 76.230 151.060 ;
        RECT 77.810 151.000 78.130 151.060 ;
        RECT 75.140 150.860 75.280 151.000 ;
        RECT 72.290 150.720 74.360 150.860 ;
        RECT 74.680 150.720 75.280 150.860 ;
        RECT 75.485 150.860 75.775 150.905 ;
        RECT 76.675 150.860 76.965 150.905 ;
        RECT 79.195 150.860 79.485 150.905 ;
        RECT 75.485 150.720 79.485 150.860 ;
        RECT 65.850 150.660 66.170 150.720 ;
        RECT 72.290 150.660 72.610 150.720 ;
        RECT 73.225 150.520 73.515 150.565 ;
        RECT 64.560 150.380 73.515 150.520 ;
        RECT 55.270 150.320 55.590 150.380 ;
        RECT 61.710 150.320 62.030 150.380 ;
        RECT 73.225 150.335 73.515 150.380 ;
        RECT 51.590 150.040 54.580 150.180 ;
        RECT 60.790 150.180 61.110 150.240 ;
        RECT 65.865 150.180 66.155 150.225 ;
        RECT 60.790 150.040 66.155 150.180 ;
        RECT 51.590 149.980 51.910 150.040 ;
        RECT 60.790 149.980 61.110 150.040 ;
        RECT 65.865 149.995 66.155 150.040 ;
        RECT 70.450 150.180 70.770 150.240 ;
        RECT 74.680 150.180 74.820 150.720 ;
        RECT 75.485 150.675 75.775 150.720 ;
        RECT 76.675 150.675 76.965 150.720 ;
        RECT 79.195 150.675 79.485 150.720 ;
        RECT 75.090 150.520 75.380 150.565 ;
        RECT 77.190 150.520 77.480 150.565 ;
        RECT 78.760 150.520 79.050 150.565 ;
        RECT 75.090 150.380 79.050 150.520 ;
        RECT 75.090 150.335 75.380 150.380 ;
        RECT 77.190 150.335 77.480 150.380 ;
        RECT 78.760 150.335 79.050 150.380 ;
        RECT 79.190 150.180 79.510 150.240 ;
        RECT 70.450 150.040 79.510 150.180 ;
        RECT 70.450 149.980 70.770 150.040 ;
        RECT 79.190 149.980 79.510 150.040 ;
        RECT 5.520 149.360 83.260 149.840 ;
        RECT 30.430 148.960 30.750 149.220 ;
        RECT 35.490 149.160 35.810 149.220 ;
        RECT 36.870 149.160 37.190 149.220 ;
        RECT 39.170 149.160 39.490 149.220 ;
        RECT 35.490 149.020 39.490 149.160 ;
        RECT 35.490 148.960 35.810 149.020 ;
        RECT 36.870 148.960 37.190 149.020 ;
        RECT 39.170 148.960 39.490 149.020 ;
        RECT 46.085 149.160 46.375 149.205 ;
        RECT 47.450 149.160 47.770 149.220 ;
        RECT 46.085 149.020 47.770 149.160 ;
        RECT 46.085 148.975 46.375 149.020 ;
        RECT 47.450 148.960 47.770 149.020 ;
        RECT 49.750 148.960 50.070 149.220 ;
        RECT 50.685 149.160 50.975 149.205 ;
        RECT 51.590 149.160 51.910 149.220 ;
        RECT 50.685 149.020 51.910 149.160 ;
        RECT 50.685 148.975 50.975 149.020 ;
        RECT 33.205 148.820 33.495 148.865 ;
        RECT 35.950 148.820 36.270 148.880 ;
        RECT 29.600 148.680 36.270 148.820 ;
        RECT 29.600 148.140 29.740 148.680 ;
        RECT 33.205 148.635 33.495 148.680 ;
        RECT 35.950 148.620 36.270 148.680 ;
        RECT 47.910 148.820 48.230 148.880 ;
        RECT 50.760 148.820 50.900 148.975 ;
        RECT 51.590 148.960 51.910 149.020 ;
        RECT 52.050 149.160 52.370 149.220 ;
        RECT 52.985 149.160 53.275 149.205 ;
        RECT 64.930 149.160 65.250 149.220 ;
        RECT 70.450 149.160 70.770 149.220 ;
        RECT 52.050 149.020 53.275 149.160 ;
        RECT 52.050 148.960 52.370 149.020 ;
        RECT 52.985 148.975 53.275 149.020 ;
        RECT 56.740 149.020 70.770 149.160 ;
        RECT 53.905 148.820 54.195 148.865 ;
        RECT 56.190 148.820 56.510 148.880 ;
        RECT 47.910 148.680 51.360 148.820 ;
        RECT 47.910 148.620 48.230 148.680 ;
        RECT 29.985 148.480 30.275 148.525 ;
        RECT 38.710 148.480 39.030 148.540 ;
        RECT 39.185 148.480 39.475 148.525 ;
        RECT 29.985 148.340 39.475 148.480 ;
        RECT 29.985 148.295 30.275 148.340 ;
        RECT 38.710 148.280 39.030 148.340 ;
        RECT 39.185 148.295 39.475 148.340 ;
        RECT 40.550 148.480 40.870 148.540 ;
        RECT 49.750 148.480 50.070 148.540 ;
        RECT 50.670 148.480 50.990 148.540 ;
        RECT 40.550 148.340 50.990 148.480 ;
        RECT 51.220 148.480 51.360 148.680 ;
        RECT 53.905 148.680 56.510 148.820 ;
        RECT 53.905 148.635 54.195 148.680 ;
        RECT 56.190 148.620 56.510 148.680 ;
        RECT 55.285 148.480 55.575 148.525 ;
        RECT 55.730 148.480 56.050 148.540 ;
        RECT 51.220 148.340 56.050 148.480 ;
        RECT 40.550 148.280 40.870 148.340 ;
        RECT 49.750 148.280 50.070 148.340 ;
        RECT 50.670 148.280 50.990 148.340 ;
        RECT 55.285 148.295 55.575 148.340 ;
        RECT 55.730 148.280 56.050 148.340 ;
        RECT 30.445 148.140 30.735 148.185 ;
        RECT 29.600 148.000 30.735 148.140 ;
        RECT 30.445 147.955 30.735 148.000 ;
        RECT 30.890 148.140 31.210 148.200 ;
        RECT 30.890 148.000 32.500 148.140 ;
        RECT 30.890 147.940 31.210 148.000 ;
        RECT 31.825 147.615 32.115 147.845 ;
        RECT 32.360 147.800 32.500 148.000 ;
        RECT 34.570 147.940 34.890 148.200 ;
        RECT 35.965 148.190 36.255 148.195 ;
        RECT 35.965 148.050 37.100 148.190 ;
        RECT 35.965 147.965 36.255 148.050 ;
        RECT 35.490 147.800 35.810 147.860 ;
        RECT 32.360 147.660 35.810 147.800 ;
        RECT 36.960 147.800 37.100 148.050 ;
        RECT 44.230 148.140 44.550 148.200 ;
        RECT 44.705 148.140 44.995 148.185 ;
        RECT 44.230 148.000 44.995 148.140 ;
        RECT 44.230 147.940 44.550 148.000 ;
        RECT 44.705 147.955 44.995 148.000 ;
        RECT 45.625 148.140 45.915 148.185 ;
        RECT 46.070 148.140 46.390 148.200 ;
        RECT 45.625 148.000 46.390 148.140 ;
        RECT 45.625 147.955 45.915 148.000 ;
        RECT 45.700 147.800 45.840 147.955 ;
        RECT 46.070 147.940 46.390 148.000 ;
        RECT 46.990 148.140 47.310 148.200 ;
        RECT 47.465 148.140 47.755 148.185 ;
        RECT 46.990 148.000 47.755 148.140 ;
        RECT 46.990 147.940 47.310 148.000 ;
        RECT 47.465 147.955 47.755 148.000 ;
        RECT 36.960 147.660 45.840 147.800 ;
        RECT 47.540 147.800 47.680 147.955 ;
        RECT 47.910 147.940 48.230 148.200 ;
        RECT 48.385 148.140 48.675 148.185 ;
        RECT 48.830 148.140 49.150 148.200 ;
        RECT 48.385 148.000 49.150 148.140 ;
        RECT 48.385 147.955 48.675 148.000 ;
        RECT 48.830 147.940 49.150 148.000 ;
        RECT 49.290 147.940 49.610 148.200 ;
        RECT 52.525 148.140 52.815 148.185 ;
        RECT 53.430 148.140 53.750 148.200 ;
        RECT 56.740 148.185 56.880 149.020 ;
        RECT 64.930 148.960 65.250 149.020 ;
        RECT 70.450 148.960 70.770 149.020 ;
        RECT 74.130 148.960 74.450 149.220 ;
        RECT 77.810 148.960 78.130 149.220 ;
        RECT 58.950 148.620 59.270 148.880 ;
        RECT 61.250 148.820 61.570 148.880 ;
        RECT 61.250 148.680 80.340 148.820 ;
        RECT 61.250 148.620 61.570 148.680 ;
        RECT 61.710 148.480 62.030 148.540 ;
        RECT 59.040 148.340 62.030 148.480 ;
        RECT 52.525 148.000 53.750 148.140 ;
        RECT 52.525 147.955 52.815 148.000 ;
        RECT 52.600 147.800 52.740 147.955 ;
        RECT 53.430 147.940 53.750 148.000 ;
        RECT 56.665 147.955 56.955 148.185 ;
        RECT 57.110 147.940 57.430 148.200 ;
        RECT 58.030 147.940 58.350 148.200 ;
        RECT 58.490 147.940 58.810 148.200 ;
        RECT 47.540 147.660 52.740 147.800 ;
        RECT 55.745 147.800 56.035 147.845 ;
        RECT 59.040 147.800 59.180 148.340 ;
        RECT 61.710 148.280 62.030 148.340 ;
        RECT 62.185 148.480 62.475 148.525 ;
        RECT 63.550 148.480 63.870 148.540 ;
        RECT 65.390 148.480 65.710 148.540 ;
        RECT 65.865 148.480 66.155 148.525 ;
        RECT 62.185 148.340 66.155 148.480 ;
        RECT 62.185 148.295 62.475 148.340 ;
        RECT 63.550 148.280 63.870 148.340 ;
        RECT 65.390 148.280 65.710 148.340 ;
        RECT 65.865 148.295 66.155 148.340 ;
        RECT 66.310 148.480 66.630 148.540 ;
        RECT 71.830 148.480 72.150 148.540 ;
        RECT 78.270 148.480 78.590 148.540 ;
        RECT 66.310 148.340 75.740 148.480 ;
        RECT 66.310 148.280 66.630 148.340 ;
        RECT 71.830 148.280 72.150 148.340 ;
        RECT 60.790 147.940 61.110 148.200 ;
        RECT 64.945 148.140 65.235 148.185 ;
        RECT 70.465 148.140 70.755 148.185 ;
        RECT 64.945 148.000 70.755 148.140 ;
        RECT 64.945 147.955 65.235 148.000 ;
        RECT 70.465 147.955 70.755 148.000 ;
        RECT 73.685 148.140 73.975 148.185 ;
        RECT 74.130 148.140 74.450 148.200 ;
        RECT 75.600 148.185 75.740 148.340 ;
        RECT 76.060 148.340 79.880 148.480 ;
        RECT 76.060 148.185 76.200 148.340 ;
        RECT 78.270 148.280 78.590 148.340 ;
        RECT 73.685 148.000 74.450 148.140 ;
        RECT 73.685 147.955 73.975 148.000 ;
        RECT 55.745 147.660 59.180 147.800 ;
        RECT 61.265 147.800 61.555 147.845 ;
        RECT 67.230 147.800 67.550 147.860 ;
        RECT 61.265 147.660 67.550 147.800 ;
        RECT 28.590 147.260 28.910 147.520 ;
        RECT 30.430 147.460 30.750 147.520 ;
        RECT 31.900 147.460 32.040 147.615 ;
        RECT 35.490 147.600 35.810 147.660 ;
        RECT 55.745 147.615 56.035 147.660 ;
        RECT 61.265 147.615 61.555 147.660 ;
        RECT 67.230 147.600 67.550 147.660 ;
        RECT 67.690 147.600 68.010 147.860 ;
        RECT 68.610 147.600 68.930 147.860 ;
        RECT 73.760 147.800 73.900 147.955 ;
        RECT 74.130 147.940 74.450 148.000 ;
        RECT 75.525 147.955 75.815 148.185 ;
        RECT 75.985 147.955 76.275 148.185 ;
        RECT 76.430 147.940 76.750 148.200 ;
        RECT 77.365 148.140 77.655 148.185 ;
        RECT 76.980 148.000 77.655 148.140 ;
        RECT 69.160 147.660 73.900 147.800 ;
        RECT 76.980 147.800 77.120 148.000 ;
        RECT 77.365 147.955 77.655 148.000 ;
        RECT 79.190 147.940 79.510 148.200 ;
        RECT 79.740 148.185 79.880 148.340 ;
        RECT 80.200 148.185 80.340 148.680 ;
        RECT 79.665 147.955 79.955 148.185 ;
        RECT 80.125 147.955 80.415 148.185 ;
        RECT 81.045 147.955 81.335 148.185 ;
        RECT 81.120 147.800 81.260 147.955 ;
        RECT 76.980 147.660 81.260 147.800 ;
        RECT 30.430 147.320 32.040 147.460 ;
        RECT 32.745 147.460 33.035 147.505 ;
        RECT 33.650 147.460 33.970 147.520 ;
        RECT 32.745 147.320 33.970 147.460 ;
        RECT 30.430 147.260 30.750 147.320 ;
        RECT 32.745 147.275 33.035 147.320 ;
        RECT 33.650 147.260 33.970 147.320 ;
        RECT 34.570 147.460 34.890 147.520 ;
        RECT 36.425 147.460 36.715 147.505 ;
        RECT 34.570 147.320 36.715 147.460 ;
        RECT 34.570 147.260 34.890 147.320 ;
        RECT 36.425 147.275 36.715 147.320 ;
        RECT 43.310 147.260 43.630 147.520 ;
        RECT 45.150 147.260 45.470 147.520 ;
        RECT 50.685 147.460 50.975 147.505 ;
        RECT 51.590 147.460 51.910 147.520 ;
        RECT 50.685 147.320 51.910 147.460 ;
        RECT 50.685 147.275 50.975 147.320 ;
        RECT 51.590 147.260 51.910 147.320 ;
        RECT 52.510 147.460 52.830 147.520 ;
        RECT 62.630 147.460 62.950 147.520 ;
        RECT 52.510 147.320 62.950 147.460 ;
        RECT 52.510 147.260 52.830 147.320 ;
        RECT 62.630 147.260 62.950 147.320 ;
        RECT 63.090 147.260 63.410 147.520 ;
        RECT 64.470 147.460 64.790 147.520 ;
        RECT 65.405 147.460 65.695 147.505 ;
        RECT 66.310 147.460 66.630 147.520 ;
        RECT 64.470 147.320 66.630 147.460 ;
        RECT 64.470 147.260 64.790 147.320 ;
        RECT 65.405 147.275 65.695 147.320 ;
        RECT 66.310 147.260 66.630 147.320 ;
        RECT 68.150 147.460 68.470 147.520 ;
        RECT 69.160 147.460 69.300 147.660 ;
        RECT 68.150 147.320 69.300 147.460 ;
        RECT 69.545 147.460 69.835 147.505 ;
        RECT 71.370 147.460 71.690 147.520 ;
        RECT 69.545 147.320 71.690 147.460 ;
        RECT 68.150 147.260 68.470 147.320 ;
        RECT 69.545 147.275 69.835 147.320 ;
        RECT 71.370 147.260 71.690 147.320 ;
        RECT 72.750 147.460 73.070 147.520 ;
        RECT 76.980 147.460 77.120 147.660 ;
        RECT 72.750 147.320 77.120 147.460 ;
        RECT 72.750 147.260 73.070 147.320 ;
        RECT 5.520 146.640 83.260 147.120 ;
        RECT 32.745 146.440 33.035 146.485 ;
        RECT 33.190 146.440 33.510 146.500 ;
        RECT 32.745 146.300 33.510 146.440 ;
        RECT 32.745 146.255 33.035 146.300 ;
        RECT 33.190 146.240 33.510 146.300 ;
        RECT 33.650 146.440 33.970 146.500 ;
        RECT 41.930 146.440 42.250 146.500 ;
        RECT 33.650 146.300 42.250 146.440 ;
        RECT 33.650 146.240 33.970 146.300 ;
        RECT 41.930 146.240 42.250 146.300 ;
        RECT 43.310 146.440 43.630 146.500 ;
        RECT 45.625 146.440 45.915 146.485 ;
        RECT 43.310 146.300 45.915 146.440 ;
        RECT 43.310 146.240 43.630 146.300 ;
        RECT 45.625 146.255 45.915 146.300 ;
        RECT 54.350 146.440 54.670 146.500 ;
        RECT 54.825 146.440 55.115 146.485 ;
        RECT 54.350 146.300 55.115 146.440 ;
        RECT 54.350 146.240 54.670 146.300 ;
        RECT 54.825 146.255 55.115 146.300 ;
        RECT 55.665 146.440 55.955 146.485 ;
        RECT 58.030 146.440 58.350 146.500 ;
        RECT 55.665 146.300 58.350 146.440 ;
        RECT 55.665 146.255 55.955 146.300 ;
        RECT 58.030 146.240 58.350 146.300 ;
        RECT 68.150 146.240 68.470 146.500 ;
        RECT 70.450 146.440 70.770 146.500 ;
        RECT 73.210 146.440 73.530 146.500 ;
        RECT 79.650 146.440 79.970 146.500 ;
        RECT 80.585 146.440 80.875 146.485 ;
        RECT 70.450 146.300 78.500 146.440 ;
        RECT 70.450 146.240 70.770 146.300 ;
        RECT 73.210 146.240 73.530 146.300 ;
        RECT 29.510 146.100 29.830 146.160 ;
        RECT 34.110 146.100 34.430 146.160 ;
        RECT 39.630 146.100 39.950 146.160 ;
        RECT 45.150 146.100 45.470 146.160 ;
        RECT 53.430 146.100 53.750 146.160 ;
        RECT 56.665 146.100 56.955 146.145 ;
        RECT 29.510 145.960 35.260 146.100 ;
        RECT 29.510 145.900 29.830 145.960 ;
        RECT 34.110 145.900 34.430 145.960 ;
        RECT 27.670 145.760 27.990 145.820 ;
        RECT 33.190 145.760 33.510 145.820 ;
        RECT 27.670 145.620 34.340 145.760 ;
        RECT 27.670 145.560 27.990 145.620 ;
        RECT 33.190 145.560 33.510 145.620 ;
        RECT 34.200 145.465 34.340 145.620 ;
        RECT 34.570 145.560 34.890 145.820 ;
        RECT 35.120 145.805 35.260 145.960 ;
        RECT 39.630 145.960 43.540 146.100 ;
        RECT 39.630 145.900 39.950 145.960 ;
        RECT 43.400 145.805 43.540 145.960 ;
        RECT 45.150 145.960 46.300 146.100 ;
        RECT 45.150 145.900 45.470 145.960 ;
        RECT 35.045 145.575 35.335 145.805 ;
        RECT 42.045 145.760 42.335 145.805 ;
        RECT 42.045 145.620 43.080 145.760 ;
        RECT 42.045 145.575 42.335 145.620 ;
        RECT 33.665 145.235 33.955 145.465 ;
        RECT 34.125 145.235 34.415 145.465 ;
        RECT 38.735 145.420 39.025 145.465 ;
        RECT 41.255 145.420 41.545 145.465 ;
        RECT 42.445 145.420 42.735 145.465 ;
        RECT 38.735 145.280 42.735 145.420 ;
        RECT 42.940 145.420 43.080 145.620 ;
        RECT 43.325 145.575 43.615 145.805 ;
        RECT 44.690 145.560 45.010 145.820 ;
        RECT 46.160 145.805 46.300 145.960 ;
        RECT 53.430 145.960 56.955 146.100 ;
        RECT 53.430 145.900 53.750 145.960 ;
        RECT 56.665 145.915 56.955 145.960 ;
        RECT 62.600 146.100 62.890 146.145 ;
        RECT 63.090 146.100 63.410 146.160 ;
        RECT 62.600 145.960 63.410 146.100 ;
        RECT 62.600 145.915 62.890 145.960 ;
        RECT 63.090 145.900 63.410 145.960 ;
        RECT 66.770 146.100 67.090 146.160 ;
        RECT 77.350 146.100 77.670 146.160 ;
        RECT 66.770 145.960 73.900 146.100 ;
        RECT 66.770 145.900 67.090 145.960 ;
        RECT 46.085 145.575 46.375 145.805 ;
        RECT 47.465 145.760 47.755 145.805 ;
        RECT 47.910 145.760 48.230 145.820 ;
        RECT 47.465 145.620 48.230 145.760 ;
        RECT 47.465 145.575 47.755 145.620 ;
        RECT 47.910 145.560 48.230 145.620 ;
        RECT 48.800 145.760 49.090 145.805 ;
        RECT 50.670 145.760 50.990 145.820 ;
        RECT 48.800 145.620 50.990 145.760 ;
        RECT 48.800 145.575 49.090 145.620 ;
        RECT 50.670 145.560 50.990 145.620 ;
        RECT 71.845 145.760 72.135 145.805 ;
        RECT 72.290 145.760 72.610 145.820 ;
        RECT 71.845 145.620 72.610 145.760 ;
        RECT 71.845 145.575 72.135 145.620 ;
        RECT 72.290 145.560 72.610 145.620 ;
        RECT 73.210 145.560 73.530 145.820 ;
        RECT 73.760 145.805 73.900 145.960 ;
        RECT 74.680 145.960 77.670 146.100 ;
        RECT 74.680 145.805 74.820 145.960 ;
        RECT 77.350 145.900 77.670 145.960 ;
        RECT 73.685 145.575 73.975 145.805 ;
        RECT 74.605 145.575 74.895 145.805 ;
        RECT 75.050 145.560 75.370 145.820 ;
        RECT 75.525 145.780 75.815 145.805 ;
        RECT 76.430 145.780 76.750 145.820 ;
        RECT 78.360 145.805 78.500 146.300 ;
        RECT 79.650 146.300 80.875 146.440 ;
        RECT 79.650 146.240 79.970 146.300 ;
        RECT 80.585 146.255 80.875 146.300 ;
        RECT 75.525 145.640 76.750 145.780 ;
        RECT 75.525 145.575 75.815 145.640 ;
        RECT 76.430 145.560 76.750 145.640 ;
        RECT 78.285 145.575 78.575 145.805 ;
        RECT 78.745 145.575 79.035 145.805 ;
        RECT 43.785 145.420 44.075 145.465 ;
        RECT 42.940 145.280 44.075 145.420 ;
        RECT 38.735 145.235 39.025 145.280 ;
        RECT 41.255 145.235 41.545 145.280 ;
        RECT 42.445 145.235 42.735 145.280 ;
        RECT 43.785 145.235 44.075 145.280 ;
        RECT 48.345 145.420 48.635 145.465 ;
        RECT 49.535 145.420 49.825 145.465 ;
        RECT 52.055 145.420 52.345 145.465 ;
        RECT 48.345 145.280 52.345 145.420 ;
        RECT 48.345 145.235 48.635 145.280 ;
        RECT 49.535 145.235 49.825 145.280 ;
        RECT 52.055 145.235 52.345 145.280 ;
        RECT 60.345 145.235 60.635 145.465 ;
        RECT 33.740 145.080 33.880 145.235 ;
        RECT 35.950 145.080 36.270 145.140 ;
        RECT 33.740 144.940 36.270 145.080 ;
        RECT 35.950 144.880 36.270 144.940 ;
        RECT 36.410 144.880 36.730 145.140 ;
        RECT 39.170 145.080 39.460 145.125 ;
        RECT 40.740 145.080 41.030 145.125 ;
        RECT 42.840 145.080 43.130 145.125 ;
        RECT 39.170 144.940 43.130 145.080 ;
        RECT 39.170 144.895 39.460 144.940 ;
        RECT 40.740 144.895 41.030 144.940 ;
        RECT 42.840 144.895 43.130 144.940 ;
        RECT 47.950 145.080 48.240 145.125 ;
        RECT 50.050 145.080 50.340 145.125 ;
        RECT 51.620 145.080 51.910 145.125 ;
        RECT 47.950 144.940 51.910 145.080 ;
        RECT 47.950 144.895 48.240 144.940 ;
        RECT 50.050 144.895 50.340 144.940 ;
        RECT 51.620 144.895 51.910 144.940 ;
        RECT 53.890 145.080 54.210 145.140 ;
        RECT 54.365 145.080 54.655 145.125 ;
        RECT 60.420 145.080 60.560 145.235 ;
        RECT 61.250 145.220 61.570 145.480 ;
        RECT 62.145 145.420 62.435 145.465 ;
        RECT 63.335 145.420 63.625 145.465 ;
        RECT 65.855 145.420 66.145 145.465 ;
        RECT 62.145 145.280 66.145 145.420 ;
        RECT 62.145 145.235 62.435 145.280 ;
        RECT 63.335 145.235 63.625 145.280 ;
        RECT 65.855 145.235 66.145 145.280 ;
        RECT 68.610 145.420 68.930 145.480 ;
        RECT 77.350 145.420 77.670 145.480 ;
        RECT 78.820 145.420 78.960 145.575 ;
        RECT 79.650 145.560 79.970 145.820 ;
        RECT 80.110 145.560 80.430 145.820 ;
        RECT 81.490 145.560 81.810 145.820 ;
        RECT 68.610 145.280 78.960 145.420 ;
        RECT 68.610 145.220 68.930 145.280 ;
        RECT 77.350 145.220 77.670 145.280 ;
        RECT 53.890 144.940 60.560 145.080 ;
        RECT 61.750 145.080 62.040 145.125 ;
        RECT 63.850 145.080 64.140 145.125 ;
        RECT 65.420 145.080 65.710 145.125 ;
        RECT 61.750 144.940 65.710 145.080 ;
        RECT 53.890 144.880 54.210 144.940 ;
        RECT 54.365 144.895 54.655 144.940 ;
        RECT 61.750 144.895 62.040 144.940 ;
        RECT 63.850 144.895 64.140 144.940 ;
        RECT 65.420 144.895 65.710 144.940 ;
        RECT 67.230 145.080 67.550 145.140 ;
        RECT 74.130 145.080 74.450 145.140 ;
        RECT 75.970 145.080 76.290 145.140 ;
        RECT 67.230 144.940 69.300 145.080 ;
        RECT 67.230 144.880 67.550 144.940 ;
        RECT 45.150 144.740 45.470 144.800 ;
        RECT 47.450 144.740 47.770 144.800 ;
        RECT 45.150 144.600 47.770 144.740 ;
        RECT 45.150 144.540 45.470 144.600 ;
        RECT 47.450 144.540 47.770 144.600 ;
        RECT 55.730 144.540 56.050 144.800 ;
        RECT 57.570 144.540 57.890 144.800 ;
        RECT 68.610 144.540 68.930 144.800 ;
        RECT 69.160 144.740 69.300 144.940 ;
        RECT 74.130 144.940 76.290 145.080 ;
        RECT 74.130 144.880 74.450 144.940 ;
        RECT 75.970 144.880 76.290 144.940 ;
        RECT 76.445 145.080 76.735 145.125 ;
        RECT 76.890 145.080 77.210 145.140 ;
        RECT 76.445 144.940 77.210 145.080 ;
        RECT 76.445 144.895 76.735 144.940 ;
        RECT 76.890 144.880 77.210 144.940 ;
        RECT 72.305 144.740 72.595 144.785 ;
        RECT 69.160 144.600 72.595 144.740 ;
        RECT 72.305 144.555 72.595 144.600 ;
        RECT 72.750 144.740 73.070 144.800 ;
        RECT 77.365 144.740 77.655 144.785 ;
        RECT 72.750 144.600 77.655 144.740 ;
        RECT 72.750 144.540 73.070 144.600 ;
        RECT 77.365 144.555 77.655 144.600 ;
        RECT 5.520 143.920 83.260 144.400 ;
        RECT 34.110 143.520 34.430 143.780 ;
        RECT 35.505 143.720 35.795 143.765 ;
        RECT 44.690 143.720 45.010 143.780 ;
        RECT 35.505 143.580 45.010 143.720 ;
        RECT 35.505 143.535 35.795 143.580 ;
        RECT 44.690 143.520 45.010 143.580 ;
        RECT 45.150 143.720 45.470 143.780 ;
        RECT 45.625 143.720 45.915 143.765 ;
        RECT 45.150 143.580 45.915 143.720 ;
        RECT 45.150 143.520 45.470 143.580 ;
        RECT 45.625 143.535 45.915 143.580 ;
        RECT 46.545 143.720 46.835 143.765 ;
        RECT 50.210 143.720 50.530 143.780 ;
        RECT 46.545 143.580 50.530 143.720 ;
        RECT 46.545 143.535 46.835 143.580 ;
        RECT 50.210 143.520 50.530 143.580 ;
        RECT 50.670 143.520 50.990 143.780 ;
        RECT 68.625 143.720 68.915 143.765 ;
        RECT 72.290 143.720 72.610 143.780 ;
        RECT 68.625 143.580 72.610 143.720 ;
        RECT 68.625 143.535 68.915 143.580 ;
        RECT 72.290 143.520 72.610 143.580 ;
        RECT 76.430 143.720 76.750 143.780 ;
        RECT 81.505 143.720 81.795 143.765 ;
        RECT 76.430 143.580 81.795 143.720 ;
        RECT 76.430 143.520 76.750 143.580 ;
        RECT 81.505 143.535 81.795 143.580 ;
        RECT 43.785 143.380 44.075 143.425 ;
        RECT 46.070 143.380 46.390 143.440 ;
        RECT 43.785 143.240 46.390 143.380 ;
        RECT 43.785 143.195 44.075 143.240 ;
        RECT 46.070 143.180 46.390 143.240 ;
        RECT 49.305 143.380 49.595 143.425 ;
        RECT 62.210 143.380 62.500 143.425 ;
        RECT 64.310 143.380 64.600 143.425 ;
        RECT 65.880 143.380 66.170 143.425 ;
        RECT 49.305 143.240 55.960 143.380 ;
        RECT 49.305 143.195 49.595 143.240 ;
        RECT 38.250 143.040 38.570 143.100 ;
        RECT 40.565 143.040 40.855 143.085 ;
        RECT 38.250 142.900 40.855 143.040 ;
        RECT 38.250 142.840 38.570 142.900 ;
        RECT 40.565 142.855 40.855 142.900 ;
        RECT 51.130 143.040 51.450 143.100 ;
        RECT 53.445 143.040 53.735 143.085 ;
        RECT 51.130 142.900 53.735 143.040 ;
        RECT 55.820 143.040 55.960 143.240 ;
        RECT 62.210 143.240 66.170 143.380 ;
        RECT 62.210 143.195 62.500 143.240 ;
        RECT 64.310 143.195 64.600 143.240 ;
        RECT 65.880 143.195 66.170 143.240 ;
        RECT 66.770 143.380 67.090 143.440 ;
        RECT 72.750 143.380 73.070 143.440 ;
        RECT 66.770 143.240 73.070 143.380 ;
        RECT 66.770 143.180 67.090 143.240 ;
        RECT 72.750 143.180 73.070 143.240 ;
        RECT 75.090 143.380 75.380 143.425 ;
        RECT 77.190 143.380 77.480 143.425 ;
        RECT 78.760 143.380 79.050 143.425 ;
        RECT 75.090 143.240 79.050 143.380 ;
        RECT 75.090 143.195 75.380 143.240 ;
        RECT 77.190 143.195 77.480 143.240 ;
        RECT 78.760 143.195 79.050 143.240 ;
        RECT 62.605 143.040 62.895 143.085 ;
        RECT 63.795 143.040 64.085 143.085 ;
        RECT 66.315 143.040 66.605 143.085 ;
        RECT 73.210 143.040 73.530 143.100 ;
        RECT 74.130 143.040 74.450 143.100 ;
        RECT 55.820 142.900 62.400 143.040 ;
        RECT 51.130 142.840 51.450 142.900 ;
        RECT 53.445 142.855 53.735 142.900 ;
        RECT 28.590 142.700 28.910 142.760 ;
        RECT 33.665 142.700 33.955 142.745 ;
        RECT 28.590 142.560 33.955 142.700 ;
        RECT 28.590 142.500 28.910 142.560 ;
        RECT 33.665 142.515 33.955 142.560 ;
        RECT 34.110 142.700 34.430 142.760 ;
        RECT 35.045 142.700 35.335 142.745 ;
        RECT 34.110 142.560 35.335 142.700 ;
        RECT 34.110 142.500 34.430 142.560 ;
        RECT 35.045 142.515 35.335 142.560 ;
        RECT 35.950 142.500 36.270 142.760 ;
        RECT 42.865 142.515 43.155 142.745 ;
        RECT 43.785 142.700 44.075 142.745 ;
        RECT 45.150 142.700 45.470 142.760 ;
        RECT 43.785 142.560 45.470 142.700 ;
        RECT 43.785 142.515 44.075 142.560 ;
        RECT 14.790 142.360 15.110 142.420 ;
        RECT 16.645 142.360 16.935 142.405 ;
        RECT 14.790 142.220 16.935 142.360 ;
        RECT 14.790 142.160 15.110 142.220 ;
        RECT 16.645 142.175 16.935 142.220 ;
        RECT 17.565 142.360 17.855 142.405 ;
        RECT 41.010 142.360 41.330 142.420 ;
        RECT 17.565 142.220 41.330 142.360 ;
        RECT 42.940 142.360 43.080 142.515 ;
        RECT 45.150 142.500 45.470 142.560 ;
        RECT 50.225 142.700 50.515 142.745 ;
        RECT 52.510 142.700 52.830 142.760 ;
        RECT 50.225 142.560 52.830 142.700 ;
        RECT 50.225 142.515 50.515 142.560 ;
        RECT 52.510 142.500 52.830 142.560 ;
        RECT 52.985 142.700 53.275 142.745 ;
        RECT 57.570 142.700 57.890 142.760 ;
        RECT 52.985 142.560 57.890 142.700 ;
        RECT 52.985 142.515 53.275 142.560 ;
        RECT 57.570 142.500 57.890 142.560 ;
        RECT 58.030 142.500 58.350 142.760 ;
        RECT 61.250 142.700 61.570 142.760 ;
        RECT 61.725 142.700 62.015 142.745 ;
        RECT 61.250 142.560 62.015 142.700 ;
        RECT 62.260 142.700 62.400 142.900 ;
        RECT 62.605 142.900 66.605 143.040 ;
        RECT 62.605 142.855 62.895 142.900 ;
        RECT 63.795 142.855 64.085 142.900 ;
        RECT 66.315 142.855 66.605 142.900 ;
        RECT 70.540 142.900 74.450 143.040 ;
        RECT 70.540 142.745 70.680 142.900 ;
        RECT 73.210 142.840 73.530 142.900 ;
        RECT 74.130 142.840 74.450 142.900 ;
        RECT 74.590 142.840 74.910 143.100 ;
        RECT 75.485 143.040 75.775 143.085 ;
        RECT 76.675 143.040 76.965 143.085 ;
        RECT 79.195 143.040 79.485 143.085 ;
        RECT 75.485 142.900 79.485 143.040 ;
        RECT 75.485 142.855 75.775 142.900 ;
        RECT 76.675 142.855 76.965 142.900 ;
        RECT 79.195 142.855 79.485 142.900 ;
        RECT 62.260 142.560 65.620 142.700 ;
        RECT 61.250 142.500 61.570 142.560 ;
        RECT 61.725 142.515 62.015 142.560 ;
        RECT 44.705 142.360 44.995 142.405 ;
        RECT 46.990 142.360 47.310 142.420 ;
        RECT 42.940 142.220 47.310 142.360 ;
        RECT 17.565 142.175 17.855 142.220 ;
        RECT 41.010 142.160 41.330 142.220 ;
        RECT 44.705 142.175 44.995 142.220 ;
        RECT 46.990 142.160 47.310 142.220 ;
        RECT 48.370 142.360 48.690 142.420 ;
        RECT 54.825 142.360 55.115 142.405 ;
        RECT 61.800 142.360 61.940 142.515 ;
        RECT 48.370 142.220 61.940 142.360 ;
        RECT 63.060 142.360 63.350 142.405 ;
        RECT 64.930 142.360 65.250 142.420 ;
        RECT 63.060 142.220 65.250 142.360 ;
        RECT 65.480 142.360 65.620 142.560 ;
        RECT 70.465 142.515 70.755 142.745 ;
        RECT 71.370 142.500 71.690 142.760 ;
        RECT 71.830 142.500 72.150 142.760 ;
        RECT 72.305 142.700 72.595 142.745 ;
        RECT 77.810 142.700 78.130 142.760 ;
        RECT 72.305 142.560 78.130 142.700 ;
        RECT 72.305 142.515 72.595 142.560 ;
        RECT 77.810 142.500 78.130 142.560 ;
        RECT 75.940 142.360 76.230 142.405 ;
        RECT 76.430 142.360 76.750 142.420 ;
        RECT 65.480 142.220 74.360 142.360 ;
        RECT 48.370 142.160 48.690 142.220 ;
        RECT 54.825 142.175 55.115 142.220 ;
        RECT 63.060 142.175 63.350 142.220 ;
        RECT 64.930 142.160 65.250 142.220 ;
        RECT 37.790 141.820 38.110 142.080 ;
        RECT 44.230 142.020 44.550 142.080 ;
        RECT 45.705 142.020 45.995 142.065 ;
        RECT 44.230 141.880 45.995 142.020 ;
        RECT 44.230 141.820 44.550 141.880 ;
        RECT 45.705 141.835 45.995 141.880 ;
        RECT 52.510 141.820 52.830 142.080 ;
        RECT 61.265 142.020 61.555 142.065 ;
        RECT 64.010 142.020 64.330 142.080 ;
        RECT 61.265 141.880 64.330 142.020 ;
        RECT 61.265 141.835 61.555 141.880 ;
        RECT 64.010 141.820 64.330 141.880 ;
        RECT 73.670 141.820 73.990 142.080 ;
        RECT 74.220 142.020 74.360 142.220 ;
        RECT 75.940 142.220 76.750 142.360 ;
        RECT 75.940 142.175 76.230 142.220 ;
        RECT 76.430 142.160 76.750 142.220 ;
        RECT 76.890 142.020 77.210 142.080 ;
        RECT 74.220 141.880 77.210 142.020 ;
        RECT 76.890 141.820 77.210 141.880 ;
        RECT 5.520 141.200 83.260 141.680 ;
        RECT 38.725 141.000 39.015 141.045 ;
        RECT 39.170 141.000 39.490 141.060 ;
        RECT 38.725 140.860 39.490 141.000 ;
        RECT 38.725 140.815 39.015 140.860 ;
        RECT 39.170 140.800 39.490 140.860 ;
        RECT 43.785 141.000 44.075 141.045 ;
        RECT 45.610 141.000 45.930 141.060 ;
        RECT 43.785 140.860 45.930 141.000 ;
        RECT 43.785 140.815 44.075 140.860 ;
        RECT 45.610 140.800 45.930 140.860 ;
        RECT 52.510 141.000 52.830 141.060 ;
        RECT 52.985 141.000 53.275 141.045 ;
        RECT 52.510 140.860 53.275 141.000 ;
        RECT 52.510 140.800 52.830 140.860 ;
        RECT 52.985 140.815 53.275 140.860 ;
        RECT 54.825 141.000 55.115 141.045 ;
        RECT 57.585 141.000 57.875 141.045 ;
        RECT 54.825 140.860 57.875 141.000 ;
        RECT 54.825 140.815 55.115 140.860 ;
        RECT 57.585 140.815 57.875 140.860 ;
        RECT 59.870 141.000 60.190 141.060 ;
        RECT 59.870 140.860 64.700 141.000 ;
        RECT 34.125 140.660 34.415 140.705 ;
        RECT 35.030 140.660 35.350 140.720 ;
        RECT 40.565 140.660 40.855 140.705 ;
        RECT 34.125 140.520 35.350 140.660 ;
        RECT 34.125 140.475 34.415 140.520 ;
        RECT 35.030 140.460 35.350 140.520 ;
        RECT 36.500 140.520 40.855 140.660 ;
        RECT 36.500 140.380 36.640 140.520 ;
        RECT 40.565 140.475 40.855 140.520 ;
        RECT 12.950 140.320 13.270 140.380 ;
        RECT 15.165 140.320 15.455 140.365 ;
        RECT 12.950 140.180 15.455 140.320 ;
        RECT 12.950 140.120 13.270 140.180 ;
        RECT 15.165 140.135 15.455 140.180 ;
        RECT 17.090 140.320 17.410 140.380 ;
        RECT 21.245 140.320 21.535 140.365 ;
        RECT 17.090 140.180 21.535 140.320 ;
        RECT 17.090 140.120 17.410 140.180 ;
        RECT 21.245 140.135 21.535 140.180 ;
        RECT 22.165 140.320 22.455 140.365 ;
        RECT 23.530 140.320 23.850 140.380 ;
        RECT 22.165 140.180 23.850 140.320 ;
        RECT 22.165 140.135 22.455 140.180 ;
        RECT 23.530 140.120 23.850 140.180 ;
        RECT 33.650 140.120 33.970 140.380 ;
        RECT 34.585 140.320 34.875 140.365 ;
        RECT 35.490 140.320 35.810 140.380 ;
        RECT 34.585 140.180 35.810 140.320 ;
        RECT 34.585 140.135 34.875 140.180 ;
        RECT 35.490 140.120 35.810 140.180 ;
        RECT 36.410 140.120 36.730 140.380 ;
        RECT 37.805 140.320 38.095 140.365 ;
        RECT 39.170 140.320 39.490 140.380 ;
        RECT 39.645 140.320 39.935 140.365 ;
        RECT 37.805 140.180 38.940 140.320 ;
        RECT 37.805 140.135 38.095 140.180 ;
        RECT 13.870 139.780 14.190 140.040 ;
        RECT 14.765 139.980 15.055 140.025 ;
        RECT 15.955 139.980 16.245 140.025 ;
        RECT 18.475 139.980 18.765 140.025 ;
        RECT 14.765 139.840 18.765 139.980 ;
        RECT 14.765 139.795 15.055 139.840 ;
        RECT 15.955 139.795 16.245 139.840 ;
        RECT 18.475 139.795 18.765 139.840 ;
        RECT 35.950 139.780 36.270 140.040 ;
        RECT 14.370 139.640 14.660 139.685 ;
        RECT 16.470 139.640 16.760 139.685 ;
        RECT 18.040 139.640 18.330 139.685 ;
        RECT 14.370 139.500 18.330 139.640 ;
        RECT 14.370 139.455 14.660 139.500 ;
        RECT 16.470 139.455 16.760 139.500 ;
        RECT 18.040 139.455 18.330 139.500 ;
        RECT 18.930 139.640 19.250 139.700 ;
        RECT 21.245 139.640 21.535 139.685 ;
        RECT 18.930 139.500 21.535 139.640 ;
        RECT 18.930 139.440 19.250 139.500 ;
        RECT 21.245 139.455 21.535 139.500 ;
        RECT 29.050 139.640 29.370 139.700 ;
        RECT 37.880 139.640 38.020 140.135 ;
        RECT 38.265 139.795 38.555 140.025 ;
        RECT 38.800 139.980 38.940 140.180 ;
        RECT 39.170 140.180 39.935 140.320 ;
        RECT 39.170 140.120 39.490 140.180 ;
        RECT 39.645 140.135 39.935 140.180 ;
        RECT 41.010 140.320 41.330 140.380 ;
        RECT 41.945 140.320 42.235 140.365 ;
        RECT 41.010 140.180 42.235 140.320 ;
        RECT 41.010 140.120 41.330 140.180 ;
        RECT 41.945 140.135 42.235 140.180 ;
        RECT 43.770 140.320 44.090 140.380 ;
        RECT 45.625 140.320 45.915 140.365 ;
        RECT 43.770 140.180 45.915 140.320 ;
        RECT 43.770 140.120 44.090 140.180 ;
        RECT 45.625 140.135 45.915 140.180 ;
        RECT 38.800 139.840 41.240 139.980 ;
        RECT 29.050 139.500 38.020 139.640 ;
        RECT 29.050 139.440 29.370 139.500 ;
        RECT 19.850 139.300 20.170 139.360 ;
        RECT 20.785 139.300 21.075 139.345 ;
        RECT 19.850 139.160 21.075 139.300 ;
        RECT 19.850 139.100 20.170 139.160 ;
        RECT 20.785 139.115 21.075 139.160 ;
        RECT 34.570 139.300 34.890 139.360 ;
        RECT 35.045 139.300 35.335 139.345 ;
        RECT 34.570 139.160 35.335 139.300 ;
        RECT 38.340 139.300 38.480 139.795 ;
        RECT 41.100 139.685 41.240 139.840 ;
        RECT 46.070 139.780 46.390 140.040 ;
        RECT 47.005 139.980 47.295 140.025 ;
        RECT 49.750 139.980 50.070 140.040 ;
        RECT 47.005 139.840 50.070 139.980 ;
        RECT 47.005 139.795 47.295 139.840 ;
        RECT 49.750 139.780 50.070 139.840 ;
        RECT 54.350 139.980 54.670 140.040 ;
        RECT 55.285 139.980 55.575 140.025 ;
        RECT 54.350 139.840 55.575 139.980 ;
        RECT 54.350 139.780 54.670 139.840 ;
        RECT 55.285 139.795 55.575 139.840 ;
        RECT 55.730 139.780 56.050 140.040 ;
        RECT 41.025 139.455 41.315 139.685 ;
        RECT 51.130 139.300 51.450 139.360 ;
        RECT 38.340 139.160 51.450 139.300 ;
        RECT 57.660 139.300 57.800 140.815 ;
        RECT 59.870 140.800 60.190 140.860 ;
        RECT 61.250 140.660 61.570 140.720 ;
        RECT 64.560 140.660 64.700 140.860 ;
        RECT 64.930 140.800 65.250 141.060 ;
        RECT 66.785 141.000 67.075 141.045 ;
        RECT 68.610 141.000 68.930 141.060 ;
        RECT 66.785 140.860 68.930 141.000 ;
        RECT 66.785 140.815 67.075 140.860 ;
        RECT 68.610 140.800 68.930 140.860 ;
        RECT 76.430 140.800 76.750 141.060 ;
        RECT 75.510 140.660 75.830 140.720 ;
        RECT 61.250 140.520 63.780 140.660 ;
        RECT 64.560 140.520 72.060 140.660 ;
        RECT 61.250 140.460 61.570 140.520 ;
        RECT 63.090 140.365 63.410 140.380 ;
        RECT 63.090 140.135 63.440 140.365 ;
        RECT 63.640 140.320 63.780 140.520 ;
        RECT 64.485 140.320 64.775 140.365 ;
        RECT 63.640 140.180 64.775 140.320 ;
        RECT 64.485 140.135 64.775 140.180 ;
        RECT 64.930 140.320 65.250 140.380 ;
        RECT 71.920 140.365 72.060 140.520 ;
        RECT 75.510 140.520 78.500 140.660 ;
        RECT 75.510 140.460 75.830 140.520 ;
        RECT 64.930 140.180 67.920 140.320 ;
        RECT 63.090 140.120 63.410 140.135 ;
        RECT 64.930 140.120 65.250 140.180 ;
        RECT 59.895 139.980 60.185 140.025 ;
        RECT 62.415 139.980 62.705 140.025 ;
        RECT 63.605 139.980 63.895 140.025 ;
        RECT 59.895 139.840 63.895 139.980 ;
        RECT 59.895 139.795 60.185 139.840 ;
        RECT 62.415 139.795 62.705 139.840 ;
        RECT 63.605 139.795 63.895 139.840 ;
        RECT 65.390 139.980 65.710 140.040 ;
        RECT 67.780 140.025 67.920 140.180 ;
        RECT 71.845 140.135 72.135 140.365 ;
        RECT 77.810 140.120 78.130 140.380 ;
        RECT 78.360 140.365 78.500 140.520 ;
        RECT 78.285 140.135 78.575 140.365 ;
        RECT 78.730 140.120 79.050 140.380 ;
        RECT 79.190 140.320 79.510 140.380 ;
        RECT 79.665 140.320 79.955 140.365 ;
        RECT 79.190 140.180 79.955 140.320 ;
        RECT 79.190 140.120 79.510 140.180 ;
        RECT 79.665 140.135 79.955 140.180 ;
        RECT 80.125 140.320 80.415 140.365 ;
        RECT 80.570 140.320 80.890 140.380 ;
        RECT 81.490 140.320 81.810 140.380 ;
        RECT 80.125 140.180 81.810 140.320 ;
        RECT 80.125 140.135 80.415 140.180 ;
        RECT 80.570 140.120 80.890 140.180 ;
        RECT 81.490 140.120 81.810 140.180 ;
        RECT 67.245 139.980 67.535 140.025 ;
        RECT 65.390 139.840 67.535 139.980 ;
        RECT 65.390 139.780 65.710 139.840 ;
        RECT 67.245 139.795 67.535 139.840 ;
        RECT 67.705 139.795 67.995 140.025 ;
        RECT 75.525 139.795 75.815 140.025 ;
        RECT 77.900 139.980 78.040 140.120 ;
        RECT 77.900 139.840 78.960 139.980 ;
        RECT 60.330 139.640 60.620 139.685 ;
        RECT 61.900 139.640 62.190 139.685 ;
        RECT 64.000 139.640 64.290 139.685 ;
        RECT 75.600 139.640 75.740 139.795 ;
        RECT 78.820 139.700 78.960 139.840 ;
        RECT 60.330 139.500 64.290 139.640 ;
        RECT 60.330 139.455 60.620 139.500 ;
        RECT 61.900 139.455 62.190 139.500 ;
        RECT 64.000 139.455 64.290 139.500 ;
        RECT 67.320 139.500 75.740 139.640 ;
        RECT 67.320 139.300 67.460 139.500 ;
        RECT 78.730 139.440 79.050 139.700 ;
        RECT 57.660 139.160 67.460 139.300 ;
        RECT 67.690 139.300 68.010 139.360 ;
        RECT 69.085 139.300 69.375 139.345 ;
        RECT 67.690 139.160 69.375 139.300 ;
        RECT 34.570 139.100 34.890 139.160 ;
        RECT 35.045 139.115 35.335 139.160 ;
        RECT 51.130 139.100 51.450 139.160 ;
        RECT 67.690 139.100 68.010 139.160 ;
        RECT 69.085 139.115 69.375 139.160 ;
        RECT 72.750 139.100 73.070 139.360 ;
        RECT 81.030 139.100 81.350 139.360 ;
        RECT 5.520 138.480 83.260 138.960 ;
        RECT 35.030 138.280 35.350 138.340 ;
        RECT 36.870 138.280 37.190 138.340 ;
        RECT 35.030 138.140 37.190 138.280 ;
        RECT 35.030 138.080 35.350 138.140 ;
        RECT 36.870 138.080 37.190 138.140 ;
        RECT 54.825 138.280 55.115 138.325 ;
        RECT 58.030 138.280 58.350 138.340 ;
        RECT 54.825 138.140 58.350 138.280 ;
        RECT 54.825 138.095 55.115 138.140 ;
        RECT 58.030 138.080 58.350 138.140 ;
        RECT 61.250 138.280 61.570 138.340 ;
        RECT 71.370 138.280 71.690 138.340 ;
        RECT 74.130 138.280 74.450 138.340 ;
        RECT 61.250 138.140 62.400 138.280 ;
        RECT 61.250 138.080 61.570 138.140 ;
        RECT 10.690 137.940 10.980 137.985 ;
        RECT 12.790 137.940 13.080 137.985 ;
        RECT 14.360 137.940 14.650 137.985 ;
        RECT 10.690 137.800 14.650 137.940 ;
        RECT 10.690 137.755 10.980 137.800 ;
        RECT 12.790 137.755 13.080 137.800 ;
        RECT 14.360 137.755 14.650 137.800 ;
        RECT 20.810 137.940 21.100 137.985 ;
        RECT 22.910 137.940 23.200 137.985 ;
        RECT 24.480 137.940 24.770 137.985 ;
        RECT 20.810 137.800 24.770 137.940 ;
        RECT 20.810 137.755 21.100 137.800 ;
        RECT 22.910 137.755 23.200 137.800 ;
        RECT 24.480 137.755 24.770 137.800 ;
        RECT 28.170 137.940 28.460 137.985 ;
        RECT 30.270 137.940 30.560 137.985 ;
        RECT 31.840 137.940 32.130 137.985 ;
        RECT 28.170 137.800 32.130 137.940 ;
        RECT 28.170 137.755 28.460 137.800 ;
        RECT 30.270 137.755 30.560 137.800 ;
        RECT 31.840 137.755 32.130 137.800 ;
        RECT 35.490 137.940 35.810 138.000 ;
        RECT 39.170 137.940 39.490 138.000 ;
        RECT 35.490 137.800 39.490 137.940 ;
        RECT 35.490 137.740 35.810 137.800 ;
        RECT 39.170 137.740 39.490 137.800 ;
        RECT 44.690 137.740 45.010 138.000 ;
        RECT 48.410 137.940 48.700 137.985 ;
        RECT 50.510 137.940 50.800 137.985 ;
        RECT 52.080 137.940 52.370 137.985 ;
        RECT 61.725 137.940 62.015 137.985 ;
        RECT 48.410 137.800 52.370 137.940 ;
        RECT 48.410 137.755 48.700 137.800 ;
        RECT 50.510 137.755 50.800 137.800 ;
        RECT 52.080 137.755 52.370 137.800 ;
        RECT 55.360 137.800 62.015 137.940 ;
        RECT 62.260 137.940 62.400 138.140 ;
        RECT 71.370 138.140 75.740 138.280 ;
        RECT 71.370 138.080 71.690 138.140 ;
        RECT 74.130 138.080 74.450 138.140 ;
        RECT 70.950 137.940 71.240 137.985 ;
        RECT 73.050 137.940 73.340 137.985 ;
        RECT 74.620 137.940 74.910 137.985 ;
        RECT 62.260 137.800 64.700 137.940 ;
        RECT 11.085 137.600 11.375 137.645 ;
        RECT 12.275 137.600 12.565 137.645 ;
        RECT 14.795 137.600 15.085 137.645 ;
        RECT 20.325 137.600 20.615 137.645 ;
        RECT 21.205 137.600 21.495 137.645 ;
        RECT 22.395 137.600 22.685 137.645 ;
        RECT 24.915 137.600 25.205 137.645 ;
        RECT 11.085 137.460 15.085 137.600 ;
        RECT 11.085 137.415 11.375 137.460 ;
        RECT 12.275 137.415 12.565 137.460 ;
        RECT 14.795 137.415 15.085 137.460 ;
        RECT 18.560 137.460 21.000 137.600 ;
        RECT 10.205 137.260 10.495 137.305 ;
        RECT 13.870 137.260 14.190 137.320 ;
        RECT 18.560 137.260 18.700 137.460 ;
        RECT 20.325 137.415 20.615 137.460 ;
        RECT 20.860 137.320 21.000 137.460 ;
        RECT 21.205 137.460 25.205 137.600 ;
        RECT 21.205 137.415 21.495 137.460 ;
        RECT 22.395 137.415 22.685 137.460 ;
        RECT 24.915 137.415 25.205 137.460 ;
        RECT 28.565 137.600 28.855 137.645 ;
        RECT 29.755 137.600 30.045 137.645 ;
        RECT 32.275 137.600 32.565 137.645 ;
        RECT 28.565 137.460 32.565 137.600 ;
        RECT 39.260 137.600 39.400 137.740 ;
        RECT 48.805 137.600 49.095 137.645 ;
        RECT 49.995 137.600 50.285 137.645 ;
        RECT 52.515 137.600 52.805 137.645 ;
        RECT 39.260 137.460 45.840 137.600 ;
        RECT 28.565 137.415 28.855 137.460 ;
        RECT 29.755 137.415 30.045 137.460 ;
        RECT 32.275 137.415 32.565 137.460 ;
        RECT 10.205 137.120 18.700 137.260 ;
        RECT 10.205 137.075 10.495 137.120 ;
        RECT 13.870 137.060 14.190 137.120 ;
        RECT 18.930 137.060 19.250 137.320 ;
        RECT 19.865 137.260 20.155 137.305 ;
        RECT 19.865 137.120 20.540 137.260 ;
        RECT 19.865 137.075 20.155 137.120 ;
        RECT 20.400 136.980 20.540 137.120 ;
        RECT 20.770 137.060 21.090 137.320 ;
        RECT 27.685 137.260 27.975 137.305 ;
        RECT 28.130 137.260 28.450 137.320 ;
        RECT 37.805 137.260 38.095 137.305 ;
        RECT 27.685 137.120 28.450 137.260 ;
        RECT 27.685 137.075 27.975 137.120 ;
        RECT 28.130 137.060 28.450 137.120 ;
        RECT 34.660 137.120 38.095 137.260 ;
        RECT 11.540 136.920 11.830 136.965 ;
        RECT 12.030 136.920 12.350 136.980 ;
        RECT 11.540 136.780 12.350 136.920 ;
        RECT 11.540 136.735 11.830 136.780 ;
        RECT 12.030 136.720 12.350 136.780 ;
        RECT 20.310 136.720 20.630 136.980 ;
        RECT 21.660 136.920 21.950 136.965 ;
        RECT 23.070 136.920 23.390 136.980 ;
        RECT 21.660 136.780 23.390 136.920 ;
        RECT 21.660 136.735 21.950 136.780 ;
        RECT 23.070 136.720 23.390 136.780 ;
        RECT 29.020 136.920 29.310 136.965 ;
        RECT 29.970 136.920 30.290 136.980 ;
        RECT 29.020 136.780 30.290 136.920 ;
        RECT 29.020 136.735 29.310 136.780 ;
        RECT 29.970 136.720 30.290 136.780 ;
        RECT 16.630 136.580 16.950 136.640 ;
        RECT 17.105 136.580 17.395 136.625 ;
        RECT 16.630 136.440 17.395 136.580 ;
        RECT 16.630 136.380 16.950 136.440 ;
        RECT 17.105 136.395 17.395 136.440 ;
        RECT 19.390 136.380 19.710 136.640 ;
        RECT 26.290 136.580 26.610 136.640 ;
        RECT 27.225 136.580 27.515 136.625 ;
        RECT 26.290 136.440 27.515 136.580 ;
        RECT 26.290 136.380 26.610 136.440 ;
        RECT 27.225 136.395 27.515 136.440 ;
        RECT 31.350 136.580 31.670 136.640 ;
        RECT 33.650 136.580 33.970 136.640 ;
        RECT 34.660 136.625 34.800 137.120 ;
        RECT 37.805 137.075 38.095 137.120 ;
        RECT 43.770 137.060 44.090 137.320 ;
        RECT 45.700 137.305 45.840 137.460 ;
        RECT 48.805 137.460 52.805 137.600 ;
        RECT 48.805 137.415 49.095 137.460 ;
        RECT 49.995 137.415 50.285 137.460 ;
        RECT 52.515 137.415 52.805 137.460 ;
        RECT 44.705 137.075 44.995 137.305 ;
        RECT 45.625 137.075 45.915 137.305 ;
        RECT 47.925 137.260 48.215 137.305 ;
        RECT 48.370 137.260 48.690 137.320 ;
        RECT 47.925 137.120 48.690 137.260 ;
        RECT 47.925 137.075 48.215 137.120 ;
        RECT 36.410 136.920 36.730 136.980 ;
        RECT 44.780 136.920 44.920 137.075 ;
        RECT 48.370 137.060 48.690 137.120 ;
        RECT 49.260 137.260 49.550 137.305 ;
        RECT 55.360 137.260 55.500 137.800 ;
        RECT 61.725 137.755 62.015 137.800 ;
        RECT 55.730 137.600 56.050 137.660 ;
        RECT 58.045 137.600 58.335 137.645 ;
        RECT 59.410 137.600 59.730 137.660 ;
        RECT 55.730 137.460 58.335 137.600 ;
        RECT 55.730 137.400 56.050 137.460 ;
        RECT 58.045 137.415 58.335 137.460 ;
        RECT 58.580 137.460 59.730 137.600 ;
        RECT 49.260 137.120 55.500 137.260 ;
        RECT 49.260 137.075 49.550 137.120 ;
        RECT 36.410 136.780 44.920 136.920 ;
        RECT 52.970 136.920 53.290 136.980 ;
        RECT 55.820 136.920 55.960 137.400 ;
        RECT 57.125 137.260 57.415 137.305 ;
        RECT 58.580 137.260 58.720 137.460 ;
        RECT 59.410 137.400 59.730 137.460 ;
        RECT 64.010 137.400 64.330 137.660 ;
        RECT 64.560 137.645 64.700 137.800 ;
        RECT 70.950 137.800 74.910 137.940 ;
        RECT 70.950 137.755 71.240 137.800 ;
        RECT 73.050 137.755 73.340 137.800 ;
        RECT 74.620 137.755 74.910 137.800 ;
        RECT 64.485 137.415 64.775 137.645 ;
        RECT 67.230 137.600 67.550 137.660 ;
        RECT 68.625 137.600 68.915 137.645 ;
        RECT 67.230 137.460 68.915 137.600 ;
        RECT 67.230 137.400 67.550 137.460 ;
        RECT 68.625 137.415 68.915 137.460 ;
        RECT 71.345 137.600 71.635 137.645 ;
        RECT 72.535 137.600 72.825 137.645 ;
        RECT 75.055 137.600 75.345 137.645 ;
        RECT 71.345 137.460 75.345 137.600 ;
        RECT 75.600 137.600 75.740 138.140 ;
        RECT 75.600 137.460 81.260 137.600 ;
        RECT 71.345 137.415 71.635 137.460 ;
        RECT 72.535 137.415 72.825 137.460 ;
        RECT 75.055 137.415 75.345 137.460 ;
        RECT 57.125 137.120 58.720 137.260 ;
        RECT 58.965 137.260 59.255 137.305 ;
        RECT 64.930 137.260 65.250 137.320 ;
        RECT 58.965 137.120 65.250 137.260 ;
        RECT 57.125 137.075 57.415 137.120 ;
        RECT 58.965 137.075 59.255 137.120 ;
        RECT 64.930 137.060 65.250 137.120 ;
        RECT 67.690 137.060 68.010 137.320 ;
        RECT 70.465 137.260 70.755 137.305 ;
        RECT 74.590 137.260 74.910 137.320 ;
        RECT 70.465 137.120 74.910 137.260 ;
        RECT 70.465 137.075 70.755 137.120 ;
        RECT 74.590 137.060 74.910 137.120 ;
        RECT 78.730 137.260 79.050 137.320 ;
        RECT 79.205 137.260 79.495 137.305 ;
        RECT 78.730 137.120 79.495 137.260 ;
        RECT 78.730 137.060 79.050 137.120 ;
        RECT 79.205 137.075 79.495 137.120 ;
        RECT 79.665 137.075 79.955 137.305 ;
        RECT 63.565 136.920 63.855 136.965 ;
        RECT 52.970 136.780 55.960 136.920 ;
        RECT 61.340 136.780 63.855 136.920 ;
        RECT 36.410 136.720 36.730 136.780 ;
        RECT 52.970 136.720 53.290 136.780 ;
        RECT 34.585 136.580 34.875 136.625 ;
        RECT 31.350 136.440 34.875 136.580 ;
        RECT 31.350 136.380 31.670 136.440 ;
        RECT 33.650 136.380 33.970 136.440 ;
        RECT 34.585 136.395 34.875 136.440 ;
        RECT 35.030 136.380 35.350 136.640 ;
        RECT 40.565 136.580 40.855 136.625 ;
        RECT 42.390 136.580 42.710 136.640 ;
        RECT 40.565 136.440 42.710 136.580 ;
        RECT 40.565 136.395 40.855 136.440 ;
        RECT 42.390 136.380 42.710 136.440 ;
        RECT 56.190 136.380 56.510 136.640 ;
        RECT 59.410 136.380 59.730 136.640 ;
        RECT 61.340 136.625 61.480 136.780 ;
        RECT 63.565 136.735 63.855 136.780 ;
        RECT 71.800 136.920 72.090 136.965 ;
        RECT 73.670 136.920 73.990 136.980 ;
        RECT 71.800 136.780 73.990 136.920 ;
        RECT 71.800 136.735 72.090 136.780 ;
        RECT 73.670 136.720 73.990 136.780 ;
        RECT 76.890 136.920 77.210 136.980 ;
        RECT 78.270 136.920 78.590 136.980 ;
        RECT 79.740 136.920 79.880 137.075 ;
        RECT 80.110 137.060 80.430 137.320 ;
        RECT 80.570 137.260 80.890 137.320 ;
        RECT 81.120 137.305 81.260 137.460 ;
        RECT 81.045 137.260 81.335 137.305 ;
        RECT 80.570 137.120 81.335 137.260 ;
        RECT 80.570 137.060 80.890 137.120 ;
        RECT 81.045 137.075 81.335 137.120 ;
        RECT 76.890 136.780 79.880 136.920 ;
        RECT 76.890 136.720 77.210 136.780 ;
        RECT 78.270 136.720 78.590 136.780 ;
        RECT 61.265 136.395 61.555 136.625 ;
        RECT 65.850 136.380 66.170 136.640 ;
        RECT 68.165 136.580 68.455 136.625 ;
        RECT 75.510 136.580 75.830 136.640 ;
        RECT 68.165 136.440 75.830 136.580 ;
        RECT 68.165 136.395 68.455 136.440 ;
        RECT 75.510 136.380 75.830 136.440 ;
        RECT 76.430 136.580 76.750 136.640 ;
        RECT 77.350 136.580 77.670 136.640 ;
        RECT 76.430 136.440 77.670 136.580 ;
        RECT 76.430 136.380 76.750 136.440 ;
        RECT 77.350 136.380 77.670 136.440 ;
        RECT 77.810 136.380 78.130 136.640 ;
        RECT 5.520 135.760 83.260 136.240 ;
        RECT 10.650 135.560 10.970 135.620 ;
        RECT 14.330 135.560 14.650 135.620 ;
        RECT 19.390 135.560 19.710 135.620 ;
        RECT 10.650 135.420 12.260 135.560 ;
        RECT 10.650 135.360 10.970 135.420 ;
        RECT 7.905 135.220 8.195 135.265 ;
        RECT 11.570 135.220 11.890 135.280 ;
        RECT 7.905 135.080 11.890 135.220 ;
        RECT 12.120 135.220 12.260 135.420 ;
        RECT 13.500 135.420 14.650 135.560 ;
        RECT 13.500 135.220 13.640 135.420 ;
        RECT 14.330 135.360 14.650 135.420 ;
        RECT 15.800 135.420 19.710 135.560 ;
        RECT 12.120 135.080 13.640 135.220 ;
        RECT 7.905 135.035 8.195 135.080 ;
        RECT 11.570 135.020 11.890 135.080 ;
        RECT 13.870 135.020 14.190 135.280 ;
        RECT 14.930 135.220 15.220 135.265 ;
        RECT 15.800 135.220 15.940 135.420 ;
        RECT 19.390 135.360 19.710 135.420 ;
        RECT 23.085 135.560 23.375 135.605 ;
        RECT 23.530 135.560 23.850 135.620 ;
        RECT 23.085 135.420 23.850 135.560 ;
        RECT 23.085 135.375 23.375 135.420 ;
        RECT 23.530 135.360 23.850 135.420 ;
        RECT 38.725 135.560 39.015 135.605 ;
        RECT 41.010 135.560 41.330 135.620 ;
        RECT 38.725 135.420 41.330 135.560 ;
        RECT 38.725 135.375 39.015 135.420 ;
        RECT 41.010 135.360 41.330 135.420 ;
        RECT 43.770 135.560 44.090 135.620 ;
        RECT 47.005 135.560 47.295 135.605 ;
        RECT 43.770 135.420 47.295 135.560 ;
        RECT 43.770 135.360 44.090 135.420 ;
        RECT 47.005 135.375 47.295 135.420 ;
        RECT 51.130 135.560 51.450 135.620 ;
        RECT 61.250 135.560 61.570 135.620 ;
        RECT 51.130 135.420 61.570 135.560 ;
        RECT 51.130 135.360 51.450 135.420 ;
        RECT 61.250 135.360 61.570 135.420 ;
        RECT 62.645 135.560 62.935 135.605 ;
        RECT 63.090 135.560 63.410 135.620 ;
        RECT 62.645 135.420 63.410 135.560 ;
        RECT 62.645 135.375 62.935 135.420 ;
        RECT 63.090 135.360 63.410 135.420 ;
        RECT 64.485 135.560 64.775 135.605 ;
        RECT 72.750 135.560 73.070 135.620 ;
        RECT 64.485 135.420 73.070 135.560 ;
        RECT 64.485 135.375 64.775 135.420 ;
        RECT 72.750 135.360 73.070 135.420 ;
        RECT 20.770 135.220 21.090 135.280 ;
        RECT 35.490 135.220 35.810 135.280 ;
        RECT 39.630 135.220 39.950 135.280 ;
        RECT 48.370 135.220 48.690 135.280 ;
        RECT 58.045 135.220 58.335 135.265 ;
        RECT 14.930 135.080 15.940 135.220 ;
        RECT 16.715 135.080 21.090 135.220 ;
        RECT 14.930 135.035 15.220 135.080 ;
        RECT 7.445 134.695 7.735 134.925 ;
        RECT 7.520 134.200 7.660 134.695 ;
        RECT 8.350 134.680 8.670 134.940 ;
        RECT 8.825 134.880 9.115 134.925 ;
        RECT 16.130 134.880 16.420 134.925 ;
        RECT 16.715 134.880 16.855 135.080 ;
        RECT 20.770 135.020 21.090 135.080 ;
        RECT 31.900 135.080 40.320 135.220 ;
        RECT 17.550 134.925 17.870 134.940 ;
        RECT 24.910 134.925 25.230 134.940 ;
        RECT 31.900 134.925 32.040 135.080 ;
        RECT 35.490 135.020 35.810 135.080 ;
        RECT 39.630 135.020 39.950 135.080 ;
        RECT 17.520 134.880 17.870 134.925 ;
        RECT 8.825 134.740 12.720 134.880 ;
        RECT 8.825 134.695 9.115 134.740 ;
        RECT 10.190 134.340 10.510 134.600 ;
        RECT 11.110 134.585 11.430 134.600 ;
        RECT 12.580 134.585 12.720 134.740 ;
        RECT 16.130 134.740 16.855 134.880 ;
        RECT 17.355 134.740 17.870 134.880 ;
        RECT 16.130 134.695 16.420 134.740 ;
        RECT 17.520 134.695 17.870 134.740 ;
        RECT 24.880 134.695 25.230 134.925 ;
        RECT 31.825 134.695 32.115 134.925 ;
        RECT 33.160 134.880 33.450 134.925 ;
        RECT 34.570 134.880 34.890 134.940 ;
        RECT 40.180 134.925 40.320 135.080 ;
        RECT 48.370 135.080 58.335 135.220 ;
        RECT 48.370 135.020 48.690 135.080 ;
        RECT 58.045 135.035 58.335 135.080 ;
        RECT 62.185 135.220 62.475 135.265 ;
        RECT 66.310 135.220 66.630 135.280 ;
        RECT 62.185 135.080 66.630 135.220 ;
        RECT 62.185 135.035 62.475 135.080 ;
        RECT 66.310 135.020 66.630 135.080 ;
        RECT 75.940 135.220 76.230 135.265 ;
        RECT 77.810 135.220 78.130 135.280 ;
        RECT 75.940 135.080 78.130 135.220 ;
        RECT 75.940 135.035 76.230 135.080 ;
        RECT 77.810 135.020 78.130 135.080 ;
        RECT 33.160 134.740 34.890 134.880 ;
        RECT 33.160 134.695 33.450 134.740 ;
        RECT 17.550 134.680 17.870 134.695 ;
        RECT 24.910 134.680 25.230 134.695 ;
        RECT 34.570 134.680 34.890 134.740 ;
        RECT 40.105 134.695 40.395 134.925 ;
        RECT 40.550 134.880 40.870 134.940 ;
        RECT 41.385 134.880 41.675 134.925 ;
        RECT 40.550 134.740 41.675 134.880 ;
        RECT 40.550 134.680 40.870 134.740 ;
        RECT 41.385 134.695 41.675 134.740 ;
        RECT 49.765 134.695 50.055 134.925 ;
        RECT 50.225 134.880 50.515 134.925 ;
        RECT 52.065 134.880 52.355 134.925 ;
        RECT 50.225 134.740 52.355 134.880 ;
        RECT 50.225 134.695 50.515 134.740 ;
        RECT 52.065 134.695 52.355 134.740 ;
        RECT 64.945 134.880 65.235 134.925 ;
        RECT 66.770 134.880 67.090 134.940 ;
        RECT 64.945 134.740 67.090 134.880 ;
        RECT 64.945 134.695 65.235 134.740 ;
        RECT 11.110 134.355 11.540 134.585 ;
        RECT 12.505 134.540 12.795 134.585 ;
        RECT 14.790 134.540 15.110 134.600 ;
        RECT 12.505 134.400 15.110 134.540 ;
        RECT 12.505 134.355 12.795 134.400 ;
        RECT 11.110 134.340 11.430 134.355 ;
        RECT 14.790 134.340 15.110 134.400 ;
        RECT 17.065 134.540 17.355 134.585 ;
        RECT 18.255 134.540 18.545 134.585 ;
        RECT 20.775 134.540 21.065 134.585 ;
        RECT 17.065 134.400 21.065 134.540 ;
        RECT 17.065 134.355 17.355 134.400 ;
        RECT 18.255 134.355 18.545 134.400 ;
        RECT 20.775 134.355 21.065 134.400 ;
        RECT 23.545 134.355 23.835 134.585 ;
        RECT 24.425 134.540 24.715 134.585 ;
        RECT 25.615 134.540 25.905 134.585 ;
        RECT 28.135 134.540 28.425 134.585 ;
        RECT 24.425 134.400 28.425 134.540 ;
        RECT 24.425 134.355 24.715 134.400 ;
        RECT 25.615 134.355 25.905 134.400 ;
        RECT 28.135 134.355 28.425 134.400 ;
        RECT 32.705 134.540 32.995 134.585 ;
        RECT 33.895 134.540 34.185 134.585 ;
        RECT 36.415 134.540 36.705 134.585 ;
        RECT 32.705 134.400 36.705 134.540 ;
        RECT 32.705 134.355 32.995 134.400 ;
        RECT 33.895 134.355 34.185 134.400 ;
        RECT 36.415 134.355 36.705 134.400 ;
        RECT 40.985 134.540 41.275 134.585 ;
        RECT 42.175 134.540 42.465 134.585 ;
        RECT 44.695 134.540 44.985 134.585 ;
        RECT 40.985 134.400 44.985 134.540 ;
        RECT 40.985 134.355 41.275 134.400 ;
        RECT 42.175 134.355 42.465 134.400 ;
        RECT 44.695 134.355 44.985 134.400 ;
        RECT 7.520 134.060 10.420 134.200 ;
        RECT 10.280 133.860 10.420 134.060 ;
        RECT 12.030 134.000 12.350 134.260 ;
        RECT 15.250 134.200 15.570 134.260 ;
        RECT 15.725 134.200 16.015 134.245 ;
        RECT 15.250 134.060 16.015 134.200 ;
        RECT 15.250 134.000 15.570 134.060 ;
        RECT 15.725 134.015 16.015 134.060 ;
        RECT 16.670 134.200 16.960 134.245 ;
        RECT 18.770 134.200 19.060 134.245 ;
        RECT 20.340 134.200 20.630 134.245 ;
        RECT 16.670 134.060 20.630 134.200 ;
        RECT 16.670 134.015 16.960 134.060 ;
        RECT 18.770 134.015 19.060 134.060 ;
        RECT 20.340 134.015 20.630 134.060 ;
        RECT 17.090 133.860 17.410 133.920 ;
        RECT 10.280 133.720 17.410 133.860 ;
        RECT 17.090 133.660 17.410 133.720 ;
        RECT 20.770 133.860 21.090 133.920 ;
        RECT 23.620 133.860 23.760 134.355 ;
        RECT 24.030 134.200 24.320 134.245 ;
        RECT 26.130 134.200 26.420 134.245 ;
        RECT 27.700 134.200 27.990 134.245 ;
        RECT 24.030 134.060 27.990 134.200 ;
        RECT 24.030 134.015 24.320 134.060 ;
        RECT 26.130 134.015 26.420 134.060 ;
        RECT 27.700 134.015 27.990 134.060 ;
        RECT 32.310 134.200 32.600 134.245 ;
        RECT 34.410 134.200 34.700 134.245 ;
        RECT 35.980 134.200 36.270 134.245 ;
        RECT 32.310 134.060 36.270 134.200 ;
        RECT 32.310 134.015 32.600 134.060 ;
        RECT 34.410 134.015 34.700 134.060 ;
        RECT 35.980 134.015 36.270 134.060 ;
        RECT 40.590 134.200 40.880 134.245 ;
        RECT 42.690 134.200 42.980 134.245 ;
        RECT 44.260 134.200 44.550 134.245 ;
        RECT 49.840 134.200 49.980 134.695 ;
        RECT 66.770 134.680 67.090 134.740 ;
        RECT 72.865 134.880 73.155 134.925 ;
        RECT 73.670 134.880 73.990 134.940 ;
        RECT 72.865 134.740 73.990 134.880 ;
        RECT 72.865 134.695 73.155 134.740 ;
        RECT 73.670 134.680 73.990 134.740 ;
        RECT 74.145 134.880 74.435 134.925 ;
        RECT 74.590 134.880 74.910 134.940 ;
        RECT 74.145 134.740 74.910 134.880 ;
        RECT 74.145 134.695 74.435 134.740 ;
        RECT 74.590 134.680 74.910 134.740 ;
        RECT 51.130 134.340 51.450 134.600 ;
        RECT 51.590 134.540 51.910 134.600 ;
        RECT 54.825 134.540 55.115 134.585 ;
        RECT 51.590 134.400 55.115 134.540 ;
        RECT 51.590 134.340 51.910 134.400 ;
        RECT 54.825 134.355 55.115 134.400 ;
        RECT 63.090 134.540 63.410 134.600 ;
        RECT 65.405 134.540 65.695 134.585 ;
        RECT 63.090 134.400 65.695 134.540 ;
        RECT 63.090 134.340 63.410 134.400 ;
        RECT 65.405 134.355 65.695 134.400 ;
        RECT 69.555 134.540 69.845 134.585 ;
        RECT 72.075 134.540 72.365 134.585 ;
        RECT 73.265 134.540 73.555 134.585 ;
        RECT 69.555 134.400 73.555 134.540 ;
        RECT 69.555 134.355 69.845 134.400 ;
        RECT 72.075 134.355 72.365 134.400 ;
        RECT 73.265 134.355 73.555 134.400 ;
        RECT 75.485 134.540 75.775 134.585 ;
        RECT 76.675 134.540 76.965 134.585 ;
        RECT 79.195 134.540 79.485 134.585 ;
        RECT 75.485 134.400 79.485 134.540 ;
        RECT 75.485 134.355 75.775 134.400 ;
        RECT 76.675 134.355 76.965 134.400 ;
        RECT 79.195 134.355 79.485 134.400 ;
        RECT 40.590 134.060 44.550 134.200 ;
        RECT 40.590 134.015 40.880 134.060 ;
        RECT 42.690 134.015 42.980 134.060 ;
        RECT 44.260 134.015 44.550 134.060 ;
        RECT 44.780 134.060 49.980 134.200 ;
        RECT 56.190 134.200 56.510 134.260 ;
        RECT 69.990 134.200 70.280 134.245 ;
        RECT 71.560 134.200 71.850 134.245 ;
        RECT 73.660 134.200 73.950 134.245 ;
        RECT 56.190 134.060 69.760 134.200 ;
        RECT 28.130 133.860 28.450 133.920 ;
        RECT 20.770 133.720 28.450 133.860 ;
        RECT 20.770 133.660 21.090 133.720 ;
        RECT 28.130 133.660 28.450 133.720 ;
        RECT 30.430 133.660 30.750 133.920 ;
        RECT 37.330 133.860 37.650 133.920 ;
        RECT 44.780 133.860 44.920 134.060 ;
        RECT 56.190 134.000 56.510 134.060 ;
        RECT 37.330 133.720 44.920 133.860 ;
        RECT 37.330 133.660 37.650 133.720 ;
        RECT 47.910 133.660 48.230 133.920 ;
        RECT 67.230 133.660 67.550 133.920 ;
        RECT 69.620 133.860 69.760 134.060 ;
        RECT 69.990 134.060 73.950 134.200 ;
        RECT 69.990 134.015 70.280 134.060 ;
        RECT 71.560 134.015 71.850 134.060 ;
        RECT 73.660 134.015 73.950 134.060 ;
        RECT 75.090 134.200 75.380 134.245 ;
        RECT 77.190 134.200 77.480 134.245 ;
        RECT 78.760 134.200 79.050 134.245 ;
        RECT 75.090 134.060 79.050 134.200 ;
        RECT 75.090 134.015 75.380 134.060 ;
        RECT 77.190 134.015 77.480 134.060 ;
        RECT 78.760 134.015 79.050 134.060 ;
        RECT 76.430 133.860 76.750 133.920 ;
        RECT 69.620 133.720 76.750 133.860 ;
        RECT 76.430 133.660 76.750 133.720 ;
        RECT 81.490 133.660 81.810 133.920 ;
        RECT 5.520 133.040 83.260 133.520 ;
        RECT 9.745 132.840 10.035 132.885 ;
        RECT 11.110 132.840 11.430 132.900 ;
        RECT 9.745 132.700 11.430 132.840 ;
        RECT 9.745 132.655 10.035 132.700 ;
        RECT 11.110 132.640 11.430 132.700 ;
        RECT 12.950 132.640 13.270 132.900 ;
        RECT 13.870 132.840 14.190 132.900 ;
        RECT 18.930 132.840 19.250 132.900 ;
        RECT 31.825 132.840 32.115 132.885 ;
        RECT 36.410 132.840 36.730 132.900 ;
        RECT 13.870 132.700 18.700 132.840 ;
        RECT 13.870 132.640 14.190 132.700 ;
        RECT 8.350 132.500 8.670 132.560 ;
        RECT 18.025 132.500 18.315 132.545 ;
        RECT 8.350 132.360 18.315 132.500 ;
        RECT 18.560 132.500 18.700 132.700 ;
        RECT 18.930 132.700 30.660 132.840 ;
        RECT 18.930 132.640 19.250 132.700 ;
        RECT 18.560 132.360 21.920 132.500 ;
        RECT 8.350 132.300 8.670 132.360 ;
        RECT 18.025 132.315 18.315 132.360 ;
        RECT 12.030 131.960 12.350 132.220 ;
        RECT 12.490 132.160 12.810 132.220 ;
        RECT 13.760 132.160 14.050 132.205 ;
        RECT 12.490 132.020 14.050 132.160 ;
        RECT 12.490 131.960 12.810 132.020 ;
        RECT 13.760 131.975 14.050 132.020 ;
        RECT 14.805 132.160 15.095 132.205 ;
        RECT 21.230 132.160 21.550 132.220 ;
        RECT 14.805 132.020 21.550 132.160 ;
        RECT 14.805 131.975 15.095 132.020 ;
        RECT 21.230 131.960 21.550 132.020 ;
        RECT 11.585 131.820 11.875 131.865 ;
        RECT 15.710 131.820 16.030 131.880 ;
        RECT 16.185 131.820 16.475 131.865 ;
        RECT 11.585 131.680 15.480 131.820 ;
        RECT 11.585 131.635 11.875 131.680 ;
        RECT 14.330 130.940 14.650 131.200 ;
        RECT 15.340 131.140 15.480 131.680 ;
        RECT 15.710 131.680 16.475 131.820 ;
        RECT 15.710 131.620 16.030 131.680 ;
        RECT 16.185 131.635 16.475 131.680 ;
        RECT 16.630 131.620 16.950 131.880 ;
        RECT 18.025 131.820 18.315 131.865 ;
        RECT 19.390 131.820 19.710 131.880 ;
        RECT 18.025 131.680 19.710 131.820 ;
        RECT 18.025 131.635 18.315 131.680 ;
        RECT 19.390 131.620 19.710 131.680 ;
        RECT 19.865 131.820 20.155 131.865 ;
        RECT 21.780 131.820 21.920 132.360 ;
        RECT 23.070 132.300 23.390 132.560 ;
        RECT 29.065 132.500 29.355 132.545 ;
        RECT 29.970 132.500 30.290 132.560 ;
        RECT 23.620 132.360 28.360 132.500 ;
        RECT 23.620 132.205 23.760 132.360 ;
        RECT 23.545 131.975 23.835 132.205 ;
        RECT 23.990 132.160 24.310 132.220 ;
        RECT 24.925 132.160 25.215 132.205 ;
        RECT 23.990 132.020 25.215 132.160 ;
        RECT 23.620 131.820 23.760 131.975 ;
        RECT 23.990 131.960 24.310 132.020 ;
        RECT 24.925 131.975 25.215 132.020 ;
        RECT 25.370 131.960 25.690 132.220 ;
        RECT 25.970 132.160 26.260 132.205 ;
        RECT 27.670 132.160 27.990 132.220 ;
        RECT 25.970 132.020 27.990 132.160 ;
        RECT 25.970 131.975 26.260 132.020 ;
        RECT 27.670 131.960 27.990 132.020 ;
        RECT 19.865 131.680 23.760 131.820 ;
        RECT 26.750 131.820 27.070 131.880 ;
        RECT 27.225 131.820 27.515 131.865 ;
        RECT 26.750 131.680 27.515 131.820 ;
        RECT 19.865 131.635 20.155 131.680 ;
        RECT 26.750 131.620 27.070 131.680 ;
        RECT 27.225 131.635 27.515 131.680 ;
        RECT 17.550 131.480 17.870 131.540 ;
        RECT 18.930 131.480 19.250 131.540 ;
        RECT 22.150 131.525 22.470 131.540 ;
        RECT 21.705 131.480 21.995 131.525 ;
        RECT 17.550 131.340 21.995 131.480 ;
        RECT 17.550 131.280 17.870 131.340 ;
        RECT 18.930 131.280 19.250 131.340 ;
        RECT 21.705 131.295 21.995 131.340 ;
        RECT 22.150 131.295 22.580 131.525 ;
        RECT 23.990 131.480 24.310 131.540 ;
        RECT 26.290 131.480 26.610 131.540 ;
        RECT 27.685 131.480 27.975 131.525 ;
        RECT 23.990 131.340 27.975 131.480 ;
        RECT 28.220 131.480 28.360 132.360 ;
        RECT 29.065 132.360 30.290 132.500 ;
        RECT 29.065 132.315 29.355 132.360 ;
        RECT 29.970 132.300 30.290 132.360 ;
        RECT 28.605 131.820 28.895 131.865 ;
        RECT 29.970 131.820 30.290 131.880 ;
        RECT 30.520 131.865 30.660 132.700 ;
        RECT 31.825 132.700 36.730 132.840 ;
        RECT 31.825 132.655 32.115 132.700 ;
        RECT 36.410 132.640 36.730 132.700 ;
        RECT 40.105 132.840 40.395 132.885 ;
        RECT 40.550 132.840 40.870 132.900 ;
        RECT 46.530 132.840 46.850 132.900 ;
        RECT 51.130 132.840 51.450 132.900 ;
        RECT 40.105 132.700 40.870 132.840 ;
        RECT 40.105 132.655 40.395 132.700 ;
        RECT 40.550 132.640 40.870 132.700 ;
        RECT 44.780 132.700 51.450 132.840 ;
        RECT 33.230 132.500 33.520 132.545 ;
        RECT 35.330 132.500 35.620 132.545 ;
        RECT 36.900 132.500 37.190 132.545 ;
        RECT 33.230 132.360 37.190 132.500 ;
        RECT 33.230 132.315 33.520 132.360 ;
        RECT 35.330 132.315 35.620 132.360 ;
        RECT 36.900 132.315 37.190 132.360 ;
        RECT 33.625 132.160 33.915 132.205 ;
        RECT 34.815 132.160 35.105 132.205 ;
        RECT 37.335 132.160 37.625 132.205 ;
        RECT 33.625 132.020 37.625 132.160 ;
        RECT 33.625 131.975 33.915 132.020 ;
        RECT 34.815 131.975 35.105 132.020 ;
        RECT 37.335 131.975 37.625 132.020 ;
        RECT 42.390 131.960 42.710 132.220 ;
        RECT 43.325 132.160 43.615 132.205 ;
        RECT 44.780 132.160 44.920 132.700 ;
        RECT 46.530 132.640 46.850 132.700 ;
        RECT 51.130 132.640 51.450 132.700 ;
        RECT 51.590 132.640 51.910 132.900 ;
        RECT 53.890 132.840 54.210 132.900 ;
        RECT 70.465 132.840 70.755 132.885 ;
        RECT 53.890 132.700 70.755 132.840 ;
        RECT 53.890 132.640 54.210 132.700 ;
        RECT 70.465 132.655 70.755 132.700 ;
        RECT 73.670 132.840 73.990 132.900 ;
        RECT 77.825 132.840 78.115 132.885 ;
        RECT 73.670 132.700 78.115 132.840 ;
        RECT 73.670 132.640 73.990 132.700 ;
        RECT 77.825 132.655 78.115 132.700 ;
        RECT 45.190 132.500 45.480 132.545 ;
        RECT 47.290 132.500 47.580 132.545 ;
        RECT 48.860 132.500 49.150 132.545 ;
        RECT 45.190 132.360 49.150 132.500 ;
        RECT 45.190 132.315 45.480 132.360 ;
        RECT 47.290 132.315 47.580 132.360 ;
        RECT 48.860 132.315 49.150 132.360 ;
        RECT 52.550 132.500 52.840 132.545 ;
        RECT 54.650 132.500 54.940 132.545 ;
        RECT 56.220 132.500 56.510 132.545 ;
        RECT 52.550 132.360 56.510 132.500 ;
        RECT 52.550 132.315 52.840 132.360 ;
        RECT 54.650 132.315 54.940 132.360 ;
        RECT 56.220 132.315 56.510 132.360 ;
        RECT 59.425 132.500 59.715 132.545 ;
        RECT 59.870 132.500 60.190 132.560 ;
        RECT 59.425 132.360 60.190 132.500 ;
        RECT 59.425 132.315 59.715 132.360 ;
        RECT 59.870 132.300 60.190 132.360 ;
        RECT 62.170 132.500 62.460 132.545 ;
        RECT 63.740 132.500 64.030 132.545 ;
        RECT 65.840 132.500 66.130 132.545 ;
        RECT 62.170 132.360 66.130 132.500 ;
        RECT 62.170 132.315 62.460 132.360 ;
        RECT 63.740 132.315 64.030 132.360 ;
        RECT 65.840 132.315 66.130 132.360 ;
        RECT 72.750 132.500 73.070 132.560 ;
        RECT 72.750 132.360 79.880 132.500 ;
        RECT 72.750 132.300 73.070 132.360 ;
        RECT 43.325 132.020 44.920 132.160 ;
        RECT 45.585 132.160 45.875 132.205 ;
        RECT 46.775 132.160 47.065 132.205 ;
        RECT 49.295 132.160 49.585 132.205 ;
        RECT 45.585 132.020 49.585 132.160 ;
        RECT 43.325 131.975 43.615 132.020 ;
        RECT 45.585 131.975 45.875 132.020 ;
        RECT 46.775 131.975 47.065 132.020 ;
        RECT 49.295 131.975 49.585 132.020 ;
        RECT 52.945 132.160 53.235 132.205 ;
        RECT 54.135 132.160 54.425 132.205 ;
        RECT 56.655 132.160 56.945 132.205 ;
        RECT 52.945 132.020 56.945 132.160 ;
        RECT 52.945 131.975 53.235 132.020 ;
        RECT 54.135 131.975 54.425 132.020 ;
        RECT 56.655 131.975 56.945 132.020 ;
        RECT 61.735 132.160 62.025 132.205 ;
        RECT 64.255 132.160 64.545 132.205 ;
        RECT 65.445 132.160 65.735 132.205 ;
        RECT 68.150 132.160 68.470 132.220 ;
        RECT 61.735 132.020 65.735 132.160 ;
        RECT 61.735 131.975 62.025 132.020 ;
        RECT 64.255 131.975 64.545 132.020 ;
        RECT 65.445 131.975 65.735 132.020 ;
        RECT 67.780 132.020 68.470 132.160 ;
        RECT 28.605 131.680 30.290 131.820 ;
        RECT 28.605 131.635 28.895 131.680 ;
        RECT 29.970 131.620 30.290 131.680 ;
        RECT 30.445 131.635 30.735 131.865 ;
        RECT 31.350 131.620 31.670 131.880 ;
        RECT 32.285 131.635 32.575 131.865 ;
        RECT 32.745 131.820 33.035 131.865 ;
        RECT 35.490 131.820 35.810 131.880 ;
        RECT 39.630 131.820 39.950 131.880 ;
        RECT 44.705 131.820 44.995 131.865 ;
        RECT 32.745 131.680 44.995 131.820 ;
        RECT 32.745 131.635 33.035 131.680 ;
        RECT 29.050 131.480 29.370 131.540 ;
        RECT 28.220 131.340 29.370 131.480 ;
        RECT 32.360 131.480 32.500 131.635 ;
        RECT 35.490 131.620 35.810 131.680 ;
        RECT 39.630 131.620 39.950 131.680 ;
        RECT 44.705 131.635 44.995 131.680 ;
        RECT 46.040 131.820 46.330 131.865 ;
        RECT 47.910 131.820 48.230 131.880 ;
        RECT 46.040 131.680 48.230 131.820 ;
        RECT 46.040 131.635 46.330 131.680 ;
        RECT 47.910 131.620 48.230 131.680 ;
        RECT 48.370 131.820 48.690 131.880 ;
        RECT 52.065 131.820 52.355 131.865 ;
        RECT 48.370 131.680 52.355 131.820 ;
        RECT 48.370 131.620 48.690 131.680 ;
        RECT 52.065 131.635 52.355 131.680 ;
        RECT 65.045 131.820 65.335 131.865 ;
        RECT 65.850 131.820 66.170 131.880 ;
        RECT 65.045 131.680 66.170 131.820 ;
        RECT 65.045 131.635 65.335 131.680 ;
        RECT 65.850 131.620 66.170 131.680 ;
        RECT 66.325 131.820 66.615 131.865 ;
        RECT 66.325 131.680 67.000 131.820 ;
        RECT 66.325 131.635 66.615 131.680 ;
        RECT 34.080 131.480 34.370 131.525 ;
        RECT 34.570 131.480 34.890 131.540 ;
        RECT 32.360 131.340 33.880 131.480 ;
        RECT 22.150 131.280 22.470 131.295 ;
        RECT 23.990 131.280 24.310 131.340 ;
        RECT 26.290 131.280 26.610 131.340 ;
        RECT 27.685 131.295 27.975 131.340 ;
        RECT 29.050 131.280 29.370 131.340 ;
        RECT 16.170 131.140 16.490 131.200 ;
        RECT 17.105 131.140 17.395 131.185 ;
        RECT 15.340 131.000 17.395 131.140 ;
        RECT 16.170 130.940 16.490 131.000 ;
        RECT 17.105 130.955 17.395 131.000 ;
        RECT 21.230 131.140 21.550 131.200 ;
        RECT 23.070 131.140 23.390 131.200 ;
        RECT 21.230 131.000 23.390 131.140 ;
        RECT 21.230 130.940 21.550 131.000 ;
        RECT 23.070 130.940 23.390 131.000 ;
        RECT 24.910 131.140 25.230 131.200 ;
        RECT 26.765 131.140 27.055 131.185 ;
        RECT 24.910 131.000 27.055 131.140 ;
        RECT 24.910 130.940 25.230 131.000 ;
        RECT 26.765 130.955 27.055 131.000 ;
        RECT 28.110 131.140 28.400 131.185 ;
        RECT 28.590 131.140 28.910 131.200 ;
        RECT 28.110 131.000 28.910 131.140 ;
        RECT 28.110 130.955 28.400 131.000 ;
        RECT 28.590 130.940 28.910 131.000 ;
        RECT 29.510 131.140 29.830 131.200 ;
        RECT 29.985 131.140 30.275 131.185 ;
        RECT 29.510 131.000 30.275 131.140 ;
        RECT 33.740 131.140 33.880 131.340 ;
        RECT 34.080 131.340 34.890 131.480 ;
        RECT 34.080 131.295 34.370 131.340 ;
        RECT 34.570 131.280 34.890 131.340 ;
        RECT 41.945 131.480 42.235 131.525 ;
        RECT 48.830 131.480 49.150 131.540 ;
        RECT 53.430 131.525 53.750 131.540 ;
        RECT 41.945 131.340 49.150 131.480 ;
        RECT 41.945 131.295 42.235 131.340 ;
        RECT 48.830 131.280 49.150 131.340 ;
        RECT 53.400 131.295 53.750 131.525 ;
        RECT 53.430 131.280 53.750 131.295 ;
        RECT 66.860 131.200 67.000 131.680 ;
        RECT 67.780 131.525 67.920 132.020 ;
        RECT 68.150 131.960 68.470 132.020 ;
        RECT 69.545 132.160 69.835 132.205 ;
        RECT 69.545 132.020 77.580 132.160 ;
        RECT 69.545 131.975 69.835 132.020 ;
        RECT 69.070 131.820 69.390 131.880 ;
        RECT 73.225 131.820 73.515 131.865 ;
        RECT 69.070 131.680 73.515 131.820 ;
        RECT 69.070 131.620 69.390 131.680 ;
        RECT 73.225 131.635 73.515 131.680 ;
        RECT 76.905 131.635 77.195 131.865 ;
        RECT 67.705 131.295 67.995 131.525 ;
        RECT 68.625 131.295 68.915 131.525 ;
        RECT 69.530 131.480 69.850 131.540 ;
        RECT 76.980 131.480 77.120 131.635 ;
        RECT 69.530 131.340 77.120 131.480 ;
        RECT 77.440 131.480 77.580 132.020 ;
        RECT 79.190 131.620 79.510 131.880 ;
        RECT 79.740 131.865 79.880 132.360 ;
        RECT 79.665 131.635 79.955 131.865 ;
        RECT 80.125 131.635 80.415 131.865 ;
        RECT 80.570 131.820 80.890 131.880 ;
        RECT 81.045 131.820 81.335 131.865 ;
        RECT 80.570 131.680 81.335 131.820 ;
        RECT 80.200 131.480 80.340 131.635 ;
        RECT 80.570 131.620 80.890 131.680 ;
        RECT 81.045 131.635 81.335 131.680 ;
        RECT 77.440 131.340 80.340 131.480 ;
        RECT 38.250 131.140 38.570 131.200 ;
        RECT 33.740 131.000 38.570 131.140 ;
        RECT 29.510 130.940 29.830 131.000 ;
        RECT 29.985 130.955 30.275 131.000 ;
        RECT 38.250 130.940 38.570 131.000 ;
        RECT 39.170 131.140 39.490 131.200 ;
        RECT 39.645 131.140 39.935 131.185 ;
        RECT 39.170 131.000 39.935 131.140 ;
        RECT 39.170 130.940 39.490 131.000 ;
        RECT 39.645 130.955 39.935 131.000 ;
        RECT 58.950 130.940 59.270 131.200 ;
        RECT 66.770 130.940 67.090 131.200 ;
        RECT 67.230 131.140 67.550 131.200 ;
        RECT 68.700 131.140 68.840 131.295 ;
        RECT 69.530 131.280 69.850 131.340 ;
        RECT 67.230 131.000 68.840 131.140 ;
        RECT 67.230 130.940 67.550 131.000 ;
        RECT 74.130 130.940 74.450 131.200 ;
        RECT 5.520 130.320 83.260 130.800 ;
        RECT 19.850 130.120 20.170 130.180 ;
        RECT 17.640 129.980 20.170 130.120 ;
        RECT 12.030 129.780 12.350 129.840 ;
        RECT 15.710 129.780 16.030 129.840 ;
        RECT 16.630 129.825 16.950 129.840 ;
        RECT 17.640 129.825 17.780 129.980 ;
        RECT 19.850 129.920 20.170 129.980 ;
        RECT 26.750 130.165 27.070 130.180 ;
        RECT 26.750 129.935 27.160 130.165 ;
        RECT 27.670 130.120 27.990 130.180 ;
        RECT 28.605 130.120 28.895 130.165 ;
        RECT 27.670 129.980 28.895 130.120 ;
        RECT 26.750 129.920 27.070 129.935 ;
        RECT 27.670 129.920 27.990 129.980 ;
        RECT 28.605 129.935 28.895 129.980 ;
        RECT 34.570 130.120 34.890 130.180 ;
        RECT 35.505 130.120 35.795 130.165 ;
        RECT 34.570 129.980 35.795 130.120 ;
        RECT 34.570 129.920 34.890 129.980 ;
        RECT 35.505 129.935 35.795 129.980 ;
        RECT 46.070 130.120 46.390 130.180 ;
        RECT 47.925 130.120 48.215 130.165 ;
        RECT 46.070 129.980 48.215 130.120 ;
        RECT 46.070 129.920 46.390 129.980 ;
        RECT 47.925 129.935 48.215 129.980 ;
        RECT 48.385 130.120 48.675 130.165 ;
        RECT 48.830 130.120 49.150 130.180 ;
        RECT 48.385 129.980 49.150 130.120 ;
        RECT 48.385 129.935 48.675 129.980 ;
        RECT 48.830 129.920 49.150 129.980 ;
        RECT 52.985 130.120 53.275 130.165 ;
        RECT 53.430 130.120 53.750 130.180 ;
        RECT 52.985 129.980 53.750 130.120 ;
        RECT 52.985 129.935 53.275 129.980 ;
        RECT 53.430 129.920 53.750 129.980 ;
        RECT 53.890 130.120 54.210 130.180 ;
        RECT 54.825 130.120 55.115 130.165 ;
        RECT 71.385 130.120 71.675 130.165 ;
        RECT 53.890 129.980 55.115 130.120 ;
        RECT 53.890 129.920 54.210 129.980 ;
        RECT 54.825 129.935 55.115 129.980 ;
        RECT 65.480 129.980 71.675 130.120 ;
        RECT 16.485 129.780 16.950 129.825 ;
        RECT 12.030 129.640 16.950 129.780 ;
        RECT 12.030 129.580 12.350 129.640 ;
        RECT 15.710 129.580 16.030 129.640 ;
        RECT 16.485 129.595 16.950 129.640 ;
        RECT 17.565 129.595 17.855 129.825 ;
        RECT 20.785 129.780 21.075 129.825 ;
        RECT 23.530 129.780 23.850 129.840 ;
        RECT 20.785 129.640 23.850 129.780 ;
        RECT 20.785 129.595 21.075 129.640 ;
        RECT 16.630 129.580 16.950 129.595 ;
        RECT 23.530 129.580 23.850 129.640 ;
        RECT 25.845 129.780 26.135 129.825 ;
        RECT 30.430 129.780 30.750 129.840 ;
        RECT 25.845 129.640 30.750 129.780 ;
        RECT 25.845 129.595 26.135 129.640 ;
        RECT 30.430 129.580 30.750 129.640 ;
        RECT 35.965 129.780 36.255 129.825 ;
        RECT 41.010 129.780 41.330 129.840 ;
        RECT 35.965 129.640 41.330 129.780 ;
        RECT 35.965 129.595 36.255 129.640 ;
        RECT 41.010 129.580 41.330 129.640 ;
        RECT 50.225 129.780 50.515 129.825 ;
        RECT 60.330 129.780 60.650 129.840 ;
        RECT 50.225 129.640 60.650 129.780 ;
        RECT 50.225 129.595 50.515 129.640 ;
        RECT 60.330 129.580 60.650 129.640 ;
        RECT 64.640 129.780 64.930 129.825 ;
        RECT 65.480 129.780 65.620 129.980 ;
        RECT 71.385 129.935 71.675 129.980 ;
        RECT 73.225 130.120 73.515 130.165 ;
        RECT 74.130 130.120 74.450 130.180 ;
        RECT 73.225 129.980 74.450 130.120 ;
        RECT 73.225 129.935 73.515 129.980 ;
        RECT 74.130 129.920 74.450 129.980 ;
        RECT 75.510 129.920 75.830 130.180 ;
        RECT 66.770 129.780 67.090 129.840 ;
        RECT 70.465 129.780 70.755 129.825 ;
        RECT 74.590 129.780 74.910 129.840 ;
        RECT 80.585 129.780 80.875 129.825 ;
        RECT 64.640 129.640 65.620 129.780 ;
        RECT 65.940 129.640 74.910 129.780 ;
        RECT 64.640 129.595 64.930 129.640 ;
        RECT 16.720 129.440 16.860 129.580 ;
        RECT 18.945 129.440 19.235 129.485 ;
        RECT 16.720 129.300 19.235 129.440 ;
        RECT 18.945 129.255 19.235 129.300 ;
        RECT 19.405 129.255 19.695 129.485 ;
        RECT 23.085 129.440 23.375 129.485 ;
        RECT 23.990 129.440 24.310 129.500 ;
        RECT 23.085 129.300 24.310 129.440 ;
        RECT 23.085 129.255 23.375 129.300 ;
        RECT 19.480 129.100 19.620 129.255 ;
        RECT 23.990 129.240 24.310 129.300 ;
        RECT 28.145 129.440 28.435 129.485 ;
        RECT 28.590 129.440 28.910 129.500 ;
        RECT 28.145 129.300 28.910 129.440 ;
        RECT 28.145 129.255 28.435 129.300 ;
        RECT 28.590 129.240 28.910 129.300 ;
        RECT 29.050 129.240 29.370 129.500 ;
        RECT 30.905 129.440 31.195 129.485 ;
        RECT 39.170 129.440 39.490 129.500 ;
        RECT 30.905 129.300 39.490 129.440 ;
        RECT 30.905 129.255 31.195 129.300 ;
        RECT 39.170 129.240 39.490 129.300 ;
        RECT 39.630 129.440 39.950 129.500 ;
        RECT 42.360 129.440 42.650 129.485 ;
        RECT 45.150 129.440 45.470 129.500 ;
        RECT 39.630 129.300 41.240 129.440 ;
        RECT 39.630 129.240 39.950 129.300 ;
        RECT 17.640 128.960 19.620 129.100 ;
        RECT 21.245 129.100 21.535 129.145 ;
        RECT 22.150 129.100 22.470 129.160 ;
        RECT 21.245 128.960 22.470 129.100 ;
        RECT 15.725 128.760 16.015 128.805 ;
        RECT 17.090 128.760 17.410 128.820 ;
        RECT 15.725 128.620 17.410 128.760 ;
        RECT 15.725 128.575 16.015 128.620 ;
        RECT 17.090 128.560 17.410 128.620 ;
        RECT 16.170 128.420 16.490 128.480 ;
        RECT 16.645 128.420 16.935 128.465 ;
        RECT 17.640 128.420 17.780 128.960 ;
        RECT 21.245 128.915 21.535 128.960 ;
        RECT 22.150 128.900 22.470 128.960 ;
        RECT 23.545 129.100 23.835 129.145 ;
        RECT 26.750 129.100 27.070 129.160 ;
        RECT 23.545 128.960 27.070 129.100 ;
        RECT 23.545 128.915 23.835 128.960 ;
        RECT 18.025 128.760 18.315 128.805 ;
        RECT 20.310 128.760 20.630 128.820 ;
        RECT 23.620 128.760 23.760 128.915 ;
        RECT 26.750 128.900 27.070 128.960 ;
        RECT 32.730 128.900 33.050 129.160 ;
        RECT 41.100 129.145 41.240 129.300 ;
        RECT 42.360 129.300 45.470 129.440 ;
        RECT 42.360 129.255 42.650 129.300 ;
        RECT 45.150 129.240 45.470 129.300 ;
        RECT 50.685 129.440 50.975 129.485 ;
        RECT 52.050 129.440 52.370 129.500 ;
        RECT 50.685 129.300 52.370 129.440 ;
        RECT 50.685 129.255 50.975 129.300 ;
        RECT 52.050 129.240 52.370 129.300 ;
        RECT 55.285 129.440 55.575 129.485 ;
        RECT 58.490 129.440 58.810 129.500 ;
        RECT 65.940 129.485 66.080 129.640 ;
        RECT 66.770 129.580 67.090 129.640 ;
        RECT 70.465 129.595 70.755 129.640 ;
        RECT 74.590 129.580 74.910 129.640 ;
        RECT 75.600 129.640 77.120 129.780 ;
        RECT 55.285 129.300 58.810 129.440 ;
        RECT 55.285 129.255 55.575 129.300 ;
        RECT 58.490 129.240 58.810 129.300 ;
        RECT 65.865 129.255 66.155 129.485 ;
        RECT 66.310 129.240 66.630 129.500 ;
        RECT 67.230 129.440 67.550 129.500 ;
        RECT 75.600 129.440 75.740 129.640 ;
        RECT 67.230 129.300 75.740 129.440 ;
        RECT 75.970 129.440 76.290 129.500 ;
        RECT 76.980 129.485 77.120 129.640 ;
        RECT 79.280 129.640 80.875 129.780 ;
        RECT 76.445 129.440 76.735 129.485 ;
        RECT 75.970 129.300 76.735 129.440 ;
        RECT 67.230 129.240 67.550 129.300 ;
        RECT 75.970 129.240 76.290 129.300 ;
        RECT 76.445 129.255 76.735 129.300 ;
        RECT 76.905 129.255 77.195 129.485 ;
        RECT 77.810 129.240 78.130 129.500 ;
        RECT 78.270 129.240 78.590 129.500 ;
        RECT 41.025 128.915 41.315 129.145 ;
        RECT 41.905 129.100 42.195 129.145 ;
        RECT 43.095 129.100 43.385 129.145 ;
        RECT 45.615 129.100 45.905 129.145 ;
        RECT 41.905 128.960 45.905 129.100 ;
        RECT 41.905 128.915 42.195 128.960 ;
        RECT 43.095 128.915 43.385 128.960 ;
        RECT 45.615 128.915 45.905 128.960 ;
        RECT 51.130 129.100 51.450 129.160 ;
        RECT 52.970 129.100 53.290 129.160 ;
        RECT 51.130 128.960 53.290 129.100 ;
        RECT 51.130 128.900 51.450 128.960 ;
        RECT 52.970 128.900 53.290 128.960 ;
        RECT 55.745 128.915 56.035 129.145 ;
        RECT 61.275 129.100 61.565 129.145 ;
        RECT 63.795 129.100 64.085 129.145 ;
        RECT 64.985 129.100 65.275 129.145 ;
        RECT 61.275 128.960 65.275 129.100 ;
        RECT 61.275 128.915 61.565 128.960 ;
        RECT 63.795 128.915 64.085 128.960 ;
        RECT 64.985 128.915 65.275 128.960 ;
        RECT 72.290 129.100 72.610 129.160 ;
        RECT 73.685 129.100 73.975 129.145 ;
        RECT 72.290 128.960 73.975 129.100 ;
        RECT 18.025 128.620 23.760 128.760 ;
        RECT 30.445 128.760 30.735 128.805 ;
        RECT 35.950 128.760 36.270 128.820 ;
        RECT 30.445 128.620 36.270 128.760 ;
        RECT 18.025 128.575 18.315 128.620 ;
        RECT 20.310 128.560 20.630 128.620 ;
        RECT 30.445 128.575 30.735 128.620 ;
        RECT 35.950 128.560 36.270 128.620 ;
        RECT 41.510 128.760 41.800 128.805 ;
        RECT 43.610 128.760 43.900 128.805 ;
        RECT 45.180 128.760 45.470 128.805 ;
        RECT 41.510 128.620 45.470 128.760 ;
        RECT 41.510 128.575 41.800 128.620 ;
        RECT 43.610 128.575 43.900 128.620 ;
        RECT 45.180 128.575 45.470 128.620 ;
        RECT 54.810 128.760 55.130 128.820 ;
        RECT 55.820 128.760 55.960 128.915 ;
        RECT 72.290 128.900 72.610 128.960 ;
        RECT 73.685 128.915 73.975 128.960 ;
        RECT 74.130 128.900 74.450 129.160 ;
        RECT 54.810 128.620 55.960 128.760 ;
        RECT 61.710 128.760 62.000 128.805 ;
        RECT 63.280 128.760 63.570 128.805 ;
        RECT 65.380 128.760 65.670 128.805 ;
        RECT 61.710 128.620 65.670 128.760 ;
        RECT 54.810 128.560 55.130 128.620 ;
        RECT 61.710 128.575 62.000 128.620 ;
        RECT 63.280 128.575 63.570 128.620 ;
        RECT 65.380 128.575 65.670 128.620 ;
        RECT 71.830 128.760 72.150 128.820 ;
        RECT 78.745 128.760 79.035 128.805 ;
        RECT 71.830 128.620 79.035 128.760 ;
        RECT 71.830 128.560 72.150 128.620 ;
        RECT 78.745 128.575 79.035 128.620 ;
        RECT 79.280 128.480 79.420 129.640 ;
        RECT 80.585 129.595 80.875 129.640 ;
        RECT 79.665 129.255 79.955 129.485 ;
        RECT 79.740 129.100 79.880 129.255 ;
        RECT 81.030 129.100 81.350 129.160 ;
        RECT 79.740 128.960 81.350 129.100 ;
        RECT 81.030 128.900 81.350 128.960 ;
        RECT 16.170 128.280 17.780 128.420 ;
        RECT 23.990 128.420 24.310 128.480 ;
        RECT 26.765 128.420 27.055 128.465 ;
        RECT 23.990 128.280 27.055 128.420 ;
        RECT 16.170 128.220 16.490 128.280 ;
        RECT 16.645 128.235 16.935 128.280 ;
        RECT 23.990 128.220 24.310 128.280 ;
        RECT 26.765 128.235 27.055 128.280 ;
        RECT 27.685 128.420 27.975 128.465 ;
        RECT 29.050 128.420 29.370 128.480 ;
        RECT 27.685 128.280 29.370 128.420 ;
        RECT 27.685 128.235 27.975 128.280 ;
        RECT 29.050 128.220 29.370 128.280 ;
        RECT 58.965 128.420 59.255 128.465 ;
        RECT 59.410 128.420 59.730 128.480 ;
        RECT 69.530 128.420 69.850 128.480 ;
        RECT 58.965 128.280 69.850 128.420 ;
        RECT 58.965 128.235 59.255 128.280 ;
        RECT 59.410 128.220 59.730 128.280 ;
        RECT 69.530 128.220 69.850 128.280 ;
        RECT 70.910 128.420 71.230 128.480 ;
        RECT 79.190 128.420 79.510 128.480 ;
        RECT 70.910 128.280 79.510 128.420 ;
        RECT 70.910 128.220 71.230 128.280 ;
        RECT 79.190 128.220 79.510 128.280 ;
        RECT 5.520 127.600 83.260 128.080 ;
        RECT 32.730 127.400 33.050 127.460 ;
        RECT 33.205 127.400 33.495 127.445 ;
        RECT 32.730 127.260 33.495 127.400 ;
        RECT 32.730 127.200 33.050 127.260 ;
        RECT 33.205 127.215 33.495 127.260 ;
        RECT 35.030 127.200 35.350 127.460 ;
        RECT 38.250 127.200 38.570 127.460 ;
        RECT 39.170 127.200 39.490 127.460 ;
        RECT 40.550 127.200 40.870 127.460 ;
        RECT 45.150 127.200 45.470 127.460 ;
        RECT 55.270 127.200 55.590 127.460 ;
        RECT 63.090 127.400 63.410 127.460 ;
        RECT 74.130 127.400 74.450 127.460 ;
        RECT 63.090 127.260 74.450 127.400 ;
        RECT 63.090 127.200 63.410 127.260 ;
        RECT 74.130 127.200 74.450 127.260 ;
        RECT 34.110 127.060 34.430 127.120 ;
        RECT 41.470 127.060 41.790 127.120 ;
        RECT 75.090 127.060 75.380 127.105 ;
        RECT 77.190 127.060 77.480 127.105 ;
        RECT 78.760 127.060 79.050 127.105 ;
        RECT 33.740 126.920 34.430 127.060 ;
        RECT 23.070 126.720 23.390 126.780 ;
        RECT 33.190 126.720 33.510 126.780 ;
        RECT 33.740 126.765 33.880 126.920 ;
        RECT 34.110 126.860 34.430 126.920 ;
        RECT 38.340 126.920 41.790 127.060 ;
        RECT 23.070 126.580 33.510 126.720 ;
        RECT 23.070 126.520 23.390 126.580 ;
        RECT 33.190 126.520 33.510 126.580 ;
        RECT 33.665 126.535 33.955 126.765 ;
        RECT 38.340 126.720 38.480 126.920 ;
        RECT 41.470 126.860 41.790 126.920 ;
        RECT 42.020 126.920 73.440 127.060 ;
        RECT 34.200 126.580 38.480 126.720 ;
        RECT 38.710 126.720 39.030 126.780 ;
        RECT 39.645 126.720 39.935 126.765 ;
        RECT 38.710 126.580 39.935 126.720 ;
        RECT 4.210 126.380 4.530 126.440 ;
        RECT 34.200 126.425 34.340 126.580 ;
        RECT 38.710 126.520 39.030 126.580 ;
        RECT 39.645 126.535 39.935 126.580 ;
        RECT 6.985 126.380 7.275 126.425 ;
        RECT 4.210 126.240 7.275 126.380 ;
        RECT 4.210 126.180 4.530 126.240 ;
        RECT 6.985 126.195 7.275 126.240 ;
        RECT 34.125 126.195 34.415 126.425 ;
        RECT 35.505 126.380 35.795 126.425 ;
        RECT 35.950 126.380 36.270 126.440 ;
        RECT 35.505 126.240 36.270 126.380 ;
        RECT 35.505 126.195 35.795 126.240 ;
        RECT 35.950 126.180 36.270 126.240 ;
        RECT 37.345 126.380 37.635 126.425 ;
        RECT 39.170 126.380 39.490 126.440 ;
        RECT 37.345 126.240 39.490 126.380 ;
        RECT 37.345 126.195 37.635 126.240 ;
        RECT 39.170 126.180 39.490 126.240 ;
        RECT 40.090 126.180 40.410 126.440 ;
        RECT 28.130 125.840 28.450 126.100 ;
        RECT 32.285 126.040 32.575 126.085 ;
        RECT 41.010 126.040 41.330 126.100 ;
        RECT 32.285 125.900 41.330 126.040 ;
        RECT 32.285 125.855 32.575 125.900 ;
        RECT 41.010 125.840 41.330 125.900 ;
        RECT 7.905 125.700 8.195 125.745 ;
        RECT 17.550 125.700 17.870 125.760 ;
        RECT 7.905 125.560 17.870 125.700 ;
        RECT 7.905 125.515 8.195 125.560 ;
        RECT 17.550 125.500 17.870 125.560 ;
        RECT 39.630 125.700 39.950 125.760 ;
        RECT 42.020 125.700 42.160 126.920 ;
        RECT 43.785 126.720 44.075 126.765 ;
        RECT 44.230 126.720 44.550 126.780 ;
        RECT 43.785 126.580 44.550 126.720 ;
        RECT 43.785 126.535 44.075 126.580 ;
        RECT 44.230 126.520 44.550 126.580 ;
        RECT 46.530 126.720 46.850 126.780 ;
        RECT 47.925 126.720 48.215 126.765 ;
        RECT 46.530 126.580 48.215 126.720 ;
        RECT 46.530 126.520 46.850 126.580 ;
        RECT 47.925 126.535 48.215 126.580 ;
        RECT 56.650 126.520 56.970 126.780 ;
        RECT 59.870 126.720 60.190 126.780 ;
        RECT 65.865 126.720 66.155 126.765 ;
        RECT 59.870 126.580 66.155 126.720 ;
        RECT 59.870 126.520 60.190 126.580 ;
        RECT 65.865 126.535 66.155 126.580 ;
        RECT 69.070 126.720 69.390 126.780 ;
        RECT 69.070 126.580 72.060 126.720 ;
        RECT 69.070 126.520 69.390 126.580 ;
        RECT 46.070 126.380 46.390 126.440 ;
        RECT 52.065 126.380 52.355 126.425 ;
        RECT 46.070 126.240 52.355 126.380 ;
        RECT 46.070 126.180 46.390 126.240 ;
        RECT 52.065 126.195 52.355 126.240 ;
        RECT 56.190 126.180 56.510 126.440 ;
        RECT 61.725 126.195 62.015 126.425 ;
        RECT 47.005 126.040 47.295 126.085 ;
        RECT 50.670 126.040 50.990 126.100 ;
        RECT 47.005 125.900 50.990 126.040 ;
        RECT 61.800 126.040 61.940 126.195 ;
        RECT 64.930 126.180 65.250 126.440 ;
        RECT 70.450 126.380 70.770 126.440 ;
        RECT 71.920 126.425 72.060 126.580 ;
        RECT 72.290 126.520 72.610 126.780 ;
        RECT 71.385 126.380 71.675 126.425 ;
        RECT 70.450 126.240 71.675 126.380 ;
        RECT 70.450 126.180 70.770 126.240 ;
        RECT 71.385 126.195 71.675 126.240 ;
        RECT 71.845 126.195 72.135 126.425 ;
        RECT 69.990 126.040 70.310 126.100 ;
        RECT 61.800 125.900 70.310 126.040 ;
        RECT 47.005 125.855 47.295 125.900 ;
        RECT 50.670 125.840 50.990 125.900 ;
        RECT 69.990 125.840 70.310 125.900 ;
        RECT 39.630 125.560 42.160 125.700 ;
        RECT 47.465 125.700 47.755 125.745 ;
        RECT 49.305 125.700 49.595 125.745 ;
        RECT 47.465 125.560 49.595 125.700 ;
        RECT 39.630 125.500 39.950 125.560 ;
        RECT 47.465 125.515 47.755 125.560 ;
        RECT 49.305 125.515 49.595 125.560 ;
        RECT 59.885 125.700 60.175 125.745 ;
        RECT 60.330 125.700 60.650 125.760 ;
        RECT 59.885 125.560 60.650 125.700 ;
        RECT 59.885 125.515 60.175 125.560 ;
        RECT 60.330 125.500 60.650 125.560 ;
        RECT 60.790 125.500 61.110 125.760 ;
        RECT 61.250 125.700 61.570 125.760 ;
        RECT 62.185 125.700 62.475 125.745 ;
        RECT 61.250 125.560 62.475 125.700 ;
        RECT 61.250 125.500 61.570 125.560 ;
        RECT 62.185 125.515 62.475 125.560 ;
        RECT 66.770 125.700 67.090 125.760 ;
        RECT 69.085 125.700 69.375 125.745 ;
        RECT 66.770 125.560 69.375 125.700 ;
        RECT 66.770 125.500 67.090 125.560 ;
        RECT 69.085 125.515 69.375 125.560 ;
        RECT 70.465 125.700 70.755 125.745 ;
        RECT 72.380 125.700 72.520 126.520 ;
        RECT 73.300 126.425 73.440 126.920 ;
        RECT 75.090 126.920 79.050 127.060 ;
        RECT 75.090 126.875 75.380 126.920 ;
        RECT 77.190 126.875 77.480 126.920 ;
        RECT 78.760 126.875 79.050 126.920 ;
        RECT 74.590 126.520 74.910 126.780 ;
        RECT 75.485 126.720 75.775 126.765 ;
        RECT 76.675 126.720 76.965 126.765 ;
        RECT 79.195 126.720 79.485 126.765 ;
        RECT 75.485 126.580 79.485 126.720 ;
        RECT 75.485 126.535 75.775 126.580 ;
        RECT 76.675 126.535 76.965 126.580 ;
        RECT 79.195 126.535 79.485 126.580 ;
        RECT 72.765 126.195 73.055 126.425 ;
        RECT 73.225 126.195 73.515 126.425 ;
        RECT 70.465 125.560 72.520 125.700 ;
        RECT 72.840 125.700 72.980 126.195 ;
        RECT 75.970 126.085 76.290 126.100 ;
        RECT 75.940 125.855 76.290 126.085 ;
        RECT 75.970 125.840 76.290 125.855 ;
        RECT 77.810 125.700 78.130 125.760 ;
        RECT 72.840 125.560 78.130 125.700 ;
        RECT 70.465 125.515 70.755 125.560 ;
        RECT 77.810 125.500 78.130 125.560 ;
        RECT 81.030 125.700 81.350 125.760 ;
        RECT 81.505 125.700 81.795 125.745 ;
        RECT 81.030 125.560 81.795 125.700 ;
        RECT 81.030 125.500 81.350 125.560 ;
        RECT 81.505 125.515 81.795 125.560 ;
        RECT 5.520 124.880 83.260 125.360 ;
        RECT 10.190 124.680 10.510 124.740 ;
        RECT 23.070 124.680 23.390 124.740 ;
        RECT 10.190 124.540 23.390 124.680 ;
        RECT 10.190 124.480 10.510 124.540 ;
        RECT 23.070 124.480 23.390 124.540 ;
        RECT 38.250 124.680 38.570 124.740 ;
        RECT 40.550 124.680 40.870 124.740 ;
        RECT 43.785 124.680 44.075 124.725 ;
        RECT 38.250 124.540 40.320 124.680 ;
        RECT 38.250 124.480 38.570 124.540 ;
        RECT 18.010 124.340 18.330 124.400 ;
        RECT 23.530 124.340 23.850 124.400 ;
        RECT 39.170 124.340 39.490 124.400 ;
        RECT 18.010 124.200 20.080 124.340 ;
        RECT 18.010 124.140 18.330 124.200 ;
        RECT 19.940 124.060 20.080 124.200 ;
        RECT 20.860 124.200 23.850 124.340 ;
        RECT 9.745 124.000 10.035 124.045 ;
        RECT 14.330 124.000 14.650 124.060 ;
        RECT 17.090 124.000 17.410 124.060 ;
        RECT 9.745 123.860 17.410 124.000 ;
        RECT 9.745 123.815 10.035 123.860 ;
        RECT 14.330 123.800 14.650 123.860 ;
        RECT 17.090 123.800 17.410 123.860 ;
        RECT 17.550 123.800 17.870 124.060 ;
        RECT 19.850 123.800 20.170 124.060 ;
        RECT 20.860 124.045 21.000 124.200 ;
        RECT 23.530 124.140 23.850 124.200 ;
        RECT 35.120 124.200 39.490 124.340 ;
        RECT 40.180 124.340 40.320 124.540 ;
        RECT 40.550 124.540 44.075 124.680 ;
        RECT 40.550 124.480 40.870 124.540 ;
        RECT 43.785 124.495 44.075 124.540 ;
        RECT 46.530 124.480 46.850 124.740 ;
        RECT 56.650 124.480 56.970 124.740 ;
        RECT 64.485 124.680 64.775 124.725 ;
        RECT 64.930 124.680 65.250 124.740 ;
        RECT 64.485 124.540 65.250 124.680 ;
        RECT 64.485 124.495 64.775 124.540 ;
        RECT 64.930 124.480 65.250 124.540 ;
        RECT 66.770 124.480 67.090 124.740 ;
        RECT 67.690 124.680 68.010 124.740 ;
        RECT 78.730 124.680 79.050 124.740 ;
        RECT 67.690 124.540 79.050 124.680 ;
        RECT 67.690 124.480 68.010 124.540 ;
        RECT 78.730 124.480 79.050 124.540 ;
        RECT 40.180 124.200 41.700 124.340 ;
        RECT 20.785 123.815 21.075 124.045 ;
        RECT 23.085 124.000 23.375 124.045 ;
        RECT 21.320 123.860 23.375 124.000 ;
        RECT 9.270 123.705 9.590 123.720 ;
        RECT 9.160 123.475 9.590 123.705 ;
        RECT 11.585 123.660 11.875 123.705 ;
        RECT 12.950 123.660 13.270 123.720 ;
        RECT 11.585 123.520 13.270 123.660 ;
        RECT 11.585 123.475 11.875 123.520 ;
        RECT 9.270 123.460 9.590 123.475 ;
        RECT 12.950 123.460 13.270 123.520 ;
        RECT 19.390 123.460 19.710 123.720 ;
        RECT 18.930 123.320 19.250 123.380 ;
        RECT 21.320 123.320 21.460 123.860 ;
        RECT 23.085 123.815 23.375 123.860 ;
        RECT 26.305 123.815 26.595 124.045 ;
        RECT 27.225 123.815 27.515 124.045 ;
        RECT 24.005 123.660 24.295 123.705 ;
        RECT 24.450 123.660 24.770 123.720 ;
        RECT 24.005 123.520 24.770 123.660 ;
        RECT 24.005 123.475 24.295 123.520 ;
        RECT 24.450 123.460 24.770 123.520 ;
        RECT 18.930 123.180 21.460 123.320 ;
        RECT 21.705 123.320 21.995 123.365 ;
        RECT 23.070 123.320 23.390 123.380 ;
        RECT 21.705 123.180 23.390 123.320 ;
        RECT 26.380 123.320 26.520 123.815 ;
        RECT 27.300 123.660 27.440 123.815 ;
        RECT 28.130 123.800 28.450 124.060 ;
        RECT 29.050 124.000 29.370 124.060 ;
        RECT 31.825 124.000 32.115 124.045 ;
        RECT 29.050 123.860 32.115 124.000 ;
        RECT 29.050 123.800 29.370 123.860 ;
        RECT 31.825 123.815 32.115 123.860 ;
        RECT 32.745 123.815 33.035 124.045 ;
        RECT 34.125 124.000 34.415 124.045 ;
        RECT 35.120 124.000 35.260 124.200 ;
        RECT 39.170 124.140 39.490 124.200 ;
        RECT 35.490 124.045 35.810 124.060 ;
        RECT 34.125 123.860 35.260 124.000 ;
        RECT 34.125 123.815 34.415 123.860 ;
        RECT 35.460 123.815 35.810 124.045 ;
        RECT 41.560 124.000 41.700 124.200 ;
        RECT 43.310 124.140 43.630 124.400 ;
        RECT 75.050 124.340 75.370 124.400 ;
        RECT 81.030 124.340 81.350 124.400 ;
        RECT 72.380 124.200 75.370 124.340 ;
        RECT 46.085 124.000 46.375 124.045 ;
        RECT 41.560 123.860 46.375 124.000 ;
        RECT 46.085 123.815 46.375 123.860 ;
        RECT 48.370 124.000 48.690 124.060 ;
        RECT 49.765 124.000 50.055 124.045 ;
        RECT 48.370 123.860 50.055 124.000 ;
        RECT 32.285 123.660 32.575 123.705 ;
        RECT 27.300 123.520 32.575 123.660 ;
        RECT 32.285 123.475 32.575 123.520 ;
        RECT 29.050 123.320 29.370 123.380 ;
        RECT 30.890 123.320 31.210 123.380 ;
        RECT 26.380 123.180 31.210 123.320 ;
        RECT 18.930 123.120 19.250 123.180 ;
        RECT 21.705 123.135 21.995 123.180 ;
        RECT 23.070 123.120 23.390 123.180 ;
        RECT 29.050 123.120 29.370 123.180 ;
        RECT 30.890 123.120 31.210 123.180 ;
        RECT 31.350 123.320 31.670 123.380 ;
        RECT 32.820 123.320 32.960 123.815 ;
        RECT 35.490 123.800 35.810 123.815 ;
        RECT 48.370 123.800 48.690 123.860 ;
        RECT 49.765 123.815 50.055 123.860 ;
        RECT 51.100 124.000 51.390 124.045 ;
        RECT 56.190 124.000 56.510 124.060 ;
        RECT 51.100 123.860 56.510 124.000 ;
        RECT 51.100 123.815 51.390 123.860 ;
        RECT 56.190 123.800 56.510 123.860 ;
        RECT 58.030 124.000 58.350 124.060 ;
        RECT 58.865 124.000 59.155 124.045 ;
        RECT 58.030 123.860 59.155 124.000 ;
        RECT 58.030 123.800 58.350 123.860 ;
        RECT 58.865 123.815 59.155 123.860 ;
        RECT 61.710 124.000 62.030 124.060 ;
        RECT 67.245 124.000 67.535 124.045 ;
        RECT 68.610 124.000 68.930 124.060 ;
        RECT 61.710 123.860 62.860 124.000 ;
        RECT 61.710 123.800 62.030 123.860 ;
        RECT 35.005 123.660 35.295 123.705 ;
        RECT 36.195 123.660 36.485 123.705 ;
        RECT 38.715 123.660 39.005 123.705 ;
        RECT 35.005 123.520 39.005 123.660 ;
        RECT 35.005 123.475 35.295 123.520 ;
        RECT 36.195 123.475 36.485 123.520 ;
        RECT 38.715 123.475 39.005 123.520 ;
        RECT 41.470 123.660 41.790 123.720 ;
        RECT 44.705 123.660 44.995 123.705 ;
        RECT 46.530 123.660 46.850 123.720 ;
        RECT 41.470 123.520 46.850 123.660 ;
        RECT 41.470 123.460 41.790 123.520 ;
        RECT 44.705 123.475 44.995 123.520 ;
        RECT 46.530 123.460 46.850 123.520 ;
        RECT 50.645 123.660 50.935 123.705 ;
        RECT 51.835 123.660 52.125 123.705 ;
        RECT 54.355 123.660 54.645 123.705 ;
        RECT 50.645 123.520 54.645 123.660 ;
        RECT 50.645 123.475 50.935 123.520 ;
        RECT 51.835 123.475 52.125 123.520 ;
        RECT 54.355 123.475 54.645 123.520 ;
        RECT 57.570 123.460 57.890 123.720 ;
        RECT 58.465 123.660 58.755 123.705 ;
        RECT 59.655 123.660 59.945 123.705 ;
        RECT 62.175 123.660 62.465 123.705 ;
        RECT 58.465 123.520 62.465 123.660 ;
        RECT 58.465 123.475 58.755 123.520 ;
        RECT 59.655 123.475 59.945 123.520 ;
        RECT 62.175 123.475 62.465 123.520 ;
        RECT 31.350 123.180 32.960 123.320 ;
        RECT 34.610 123.320 34.900 123.365 ;
        RECT 36.710 123.320 37.000 123.365 ;
        RECT 38.280 123.320 38.570 123.365 ;
        RECT 34.610 123.180 38.570 123.320 ;
        RECT 31.350 123.120 31.670 123.180 ;
        RECT 34.610 123.135 34.900 123.180 ;
        RECT 36.710 123.135 37.000 123.180 ;
        RECT 38.280 123.135 38.570 123.180 ;
        RECT 50.250 123.320 50.540 123.365 ;
        RECT 52.350 123.320 52.640 123.365 ;
        RECT 53.920 123.320 54.210 123.365 ;
        RECT 50.250 123.180 54.210 123.320 ;
        RECT 50.250 123.135 50.540 123.180 ;
        RECT 52.350 123.135 52.640 123.180 ;
        RECT 53.920 123.135 54.210 123.180 ;
        RECT 58.070 123.320 58.360 123.365 ;
        RECT 60.170 123.320 60.460 123.365 ;
        RECT 61.740 123.320 62.030 123.365 ;
        RECT 58.070 123.180 62.030 123.320 ;
        RECT 62.720 123.320 62.860 123.860 ;
        RECT 67.245 123.860 68.930 124.000 ;
        RECT 67.245 123.815 67.535 123.860 ;
        RECT 68.610 123.800 68.930 123.860 ;
        RECT 70.465 123.815 70.755 124.045 ;
        RECT 70.925 124.000 71.215 124.045 ;
        RECT 71.370 124.000 71.690 124.060 ;
        RECT 70.925 123.860 71.690 124.000 ;
        RECT 70.925 123.815 71.215 123.860 ;
        RECT 63.090 123.660 63.410 123.720 ;
        RECT 67.705 123.660 67.995 123.705 ;
        RECT 63.090 123.520 67.995 123.660 ;
        RECT 70.540 123.660 70.680 123.815 ;
        RECT 71.370 123.800 71.690 123.860 ;
        RECT 71.830 123.800 72.150 124.060 ;
        RECT 72.380 124.045 72.520 124.200 ;
        RECT 75.050 124.140 75.370 124.200 ;
        RECT 75.600 124.200 81.350 124.340 ;
        RECT 72.305 123.815 72.595 124.045 ;
        RECT 72.750 123.800 73.070 124.060 ;
        RECT 74.590 123.800 74.910 124.060 ;
        RECT 75.600 124.000 75.740 124.200 ;
        RECT 81.030 124.140 81.350 124.200 ;
        RECT 75.140 123.860 75.740 124.000 ;
        RECT 75.940 124.000 76.230 124.045 ;
        RECT 77.350 124.000 77.670 124.060 ;
        RECT 75.940 123.860 77.670 124.000 ;
        RECT 75.140 123.660 75.280 123.860 ;
        RECT 75.940 123.815 76.230 123.860 ;
        RECT 77.350 123.800 77.670 123.860 ;
        RECT 70.540 123.520 75.280 123.660 ;
        RECT 75.485 123.660 75.775 123.705 ;
        RECT 76.675 123.660 76.965 123.705 ;
        RECT 79.195 123.660 79.485 123.705 ;
        RECT 75.485 123.520 79.485 123.660 ;
        RECT 63.090 123.460 63.410 123.520 ;
        RECT 67.705 123.475 67.995 123.520 ;
        RECT 75.485 123.475 75.775 123.520 ;
        RECT 76.675 123.475 76.965 123.520 ;
        RECT 79.195 123.475 79.485 123.520 ;
        RECT 62.720 123.180 69.300 123.320 ;
        RECT 58.070 123.135 58.360 123.180 ;
        RECT 60.170 123.135 60.460 123.180 ;
        RECT 61.740 123.135 62.030 123.180 ;
        RECT 8.365 122.980 8.655 123.025 ;
        RECT 8.810 122.980 9.130 123.040 ;
        RECT 8.365 122.840 9.130 122.980 ;
        RECT 8.365 122.795 8.655 122.840 ;
        RECT 8.810 122.780 9.130 122.840 ;
        RECT 17.090 122.980 17.410 123.040 ;
        RECT 18.485 122.980 18.775 123.025 ;
        RECT 20.310 122.980 20.630 123.040 ;
        RECT 17.090 122.840 20.630 122.980 ;
        RECT 17.090 122.780 17.410 122.840 ;
        RECT 18.485 122.795 18.775 122.840 ;
        RECT 20.310 122.780 20.630 122.840 ;
        RECT 22.165 122.980 22.455 123.025 ;
        RECT 23.530 122.980 23.850 123.040 ;
        RECT 22.165 122.840 23.850 122.980 ;
        RECT 22.165 122.795 22.455 122.840 ;
        RECT 23.530 122.780 23.850 122.840 ;
        RECT 27.210 122.780 27.530 123.040 ;
        RECT 38.710 122.980 39.030 123.040 ;
        RECT 41.025 122.980 41.315 123.025 ;
        RECT 38.710 122.840 41.315 122.980 ;
        RECT 38.710 122.780 39.030 122.840 ;
        RECT 41.025 122.795 41.315 122.840 ;
        RECT 41.485 122.980 41.775 123.025 ;
        RECT 42.390 122.980 42.710 123.040 ;
        RECT 41.485 122.840 42.710 122.980 ;
        RECT 41.485 122.795 41.775 122.840 ;
        RECT 42.390 122.780 42.710 122.840 ;
        RECT 57.110 122.980 57.430 123.040 ;
        RECT 64.010 122.980 64.330 123.040 ;
        RECT 57.110 122.840 64.330 122.980 ;
        RECT 57.110 122.780 57.430 122.840 ;
        RECT 64.010 122.780 64.330 122.840 ;
        RECT 64.930 122.780 65.250 123.040 ;
        RECT 69.160 122.980 69.300 123.180 ;
        RECT 69.530 123.120 69.850 123.380 ;
        RECT 70.450 123.320 70.770 123.380 ;
        RECT 71.830 123.320 72.150 123.380 ;
        RECT 70.450 123.180 72.150 123.320 ;
        RECT 70.450 123.120 70.770 123.180 ;
        RECT 71.830 123.120 72.150 123.180 ;
        RECT 73.670 123.320 73.990 123.380 ;
        RECT 74.590 123.320 74.910 123.380 ;
        RECT 73.670 123.180 74.910 123.320 ;
        RECT 73.670 123.120 73.990 123.180 ;
        RECT 74.590 123.120 74.910 123.180 ;
        RECT 75.090 123.320 75.380 123.365 ;
        RECT 77.190 123.320 77.480 123.365 ;
        RECT 78.760 123.320 79.050 123.365 ;
        RECT 75.090 123.180 79.050 123.320 ;
        RECT 75.090 123.135 75.380 123.180 ;
        RECT 77.190 123.135 77.480 123.180 ;
        RECT 78.760 123.135 79.050 123.180 ;
        RECT 73.210 122.980 73.530 123.040 ;
        RECT 69.160 122.840 73.530 122.980 ;
        RECT 73.210 122.780 73.530 122.840 ;
        RECT 74.145 122.980 74.435 123.025 ;
        RECT 75.970 122.980 76.290 123.040 ;
        RECT 74.145 122.840 76.290 122.980 ;
        RECT 74.145 122.795 74.435 122.840 ;
        RECT 75.970 122.780 76.290 122.840 ;
        RECT 76.430 122.980 76.750 123.040 ;
        RECT 78.270 122.980 78.590 123.040 ;
        RECT 76.430 122.840 78.590 122.980 ;
        RECT 76.430 122.780 76.750 122.840 ;
        RECT 78.270 122.780 78.590 122.840 ;
        RECT 79.190 122.980 79.510 123.040 ;
        RECT 81.505 122.980 81.795 123.025 ;
        RECT 79.190 122.840 81.795 122.980 ;
        RECT 79.190 122.780 79.510 122.840 ;
        RECT 81.505 122.795 81.795 122.840 ;
        RECT 5.520 122.160 83.260 122.640 ;
        RECT 9.270 121.960 9.590 122.020 ;
        RECT 14.805 121.960 15.095 122.005 ;
        RECT 9.270 121.820 15.095 121.960 ;
        RECT 9.270 121.760 9.590 121.820 ;
        RECT 14.805 121.775 15.095 121.820 ;
        RECT 21.230 121.960 21.550 122.020 ;
        RECT 24.450 121.960 24.770 122.020 ;
        RECT 21.230 121.820 24.770 121.960 ;
        RECT 21.230 121.760 21.550 121.820 ;
        RECT 24.450 121.760 24.770 121.820 ;
        RECT 26.750 121.960 27.070 122.020 ;
        RECT 30.890 121.960 31.210 122.020 ;
        RECT 33.205 121.960 33.495 122.005 ;
        RECT 26.750 121.820 30.660 121.960 ;
        RECT 26.750 121.760 27.070 121.820 ;
        RECT 7.930 121.620 8.220 121.665 ;
        RECT 10.030 121.620 10.320 121.665 ;
        RECT 11.600 121.620 11.890 121.665 ;
        RECT 7.930 121.480 11.890 121.620 ;
        RECT 7.930 121.435 8.220 121.480 ;
        RECT 10.030 121.435 10.320 121.480 ;
        RECT 11.600 121.435 11.890 121.480 ;
        RECT 19.405 121.620 19.695 121.665 ;
        RECT 19.850 121.620 20.170 121.680 ;
        RECT 19.405 121.480 20.170 121.620 ;
        RECT 24.540 121.620 24.680 121.760 ;
        RECT 30.520 121.620 30.660 121.820 ;
        RECT 30.890 121.820 33.495 121.960 ;
        RECT 30.890 121.760 31.210 121.820 ;
        RECT 33.205 121.775 33.495 121.820 ;
        RECT 35.490 121.960 35.810 122.020 ;
        RECT 35.965 121.960 36.255 122.005 ;
        RECT 35.490 121.820 36.255 121.960 ;
        RECT 35.490 121.760 35.810 121.820 ;
        RECT 35.965 121.775 36.255 121.820 ;
        RECT 36.885 121.960 37.175 122.005 ;
        RECT 44.230 121.960 44.550 122.020 ;
        RECT 36.885 121.820 44.550 121.960 ;
        RECT 36.885 121.775 37.175 121.820 ;
        RECT 44.230 121.760 44.550 121.820 ;
        RECT 50.670 121.760 50.990 122.020 ;
        RECT 51.130 121.960 51.450 122.020 ;
        RECT 53.430 121.960 53.750 122.020 ;
        RECT 61.250 121.960 61.570 122.020 ;
        RECT 51.130 121.820 53.750 121.960 ;
        RECT 51.130 121.760 51.450 121.820 ;
        RECT 53.430 121.760 53.750 121.820 ;
        RECT 54.900 121.820 61.570 121.960 ;
        RECT 39.630 121.620 39.920 121.665 ;
        RECT 41.200 121.620 41.490 121.665 ;
        RECT 43.300 121.620 43.590 121.665 ;
        RECT 54.900 121.620 55.040 121.820 ;
        RECT 61.250 121.760 61.570 121.820 ;
        RECT 65.850 121.960 66.170 122.020 ;
        RECT 71.370 121.960 71.690 122.020 ;
        RECT 74.590 121.960 74.910 122.020 ;
        RECT 65.850 121.820 67.000 121.960 ;
        RECT 65.850 121.760 66.170 121.820 ;
        RECT 24.540 121.480 30.200 121.620 ;
        RECT 30.520 121.480 32.500 121.620 ;
        RECT 19.405 121.435 19.695 121.480 ;
        RECT 19.850 121.420 20.170 121.480 ;
        RECT 8.325 121.280 8.615 121.325 ;
        RECT 9.515 121.280 9.805 121.325 ;
        RECT 12.035 121.280 12.325 121.325 ;
        RECT 15.250 121.280 15.570 121.340 ;
        RECT 23.085 121.280 23.375 121.325 ;
        RECT 8.325 121.140 12.325 121.280 ;
        RECT 8.325 121.095 8.615 121.140 ;
        RECT 9.515 121.095 9.805 121.140 ;
        RECT 12.035 121.095 12.325 121.140 ;
        RECT 14.420 121.140 23.375 121.280 ;
        RECT 6.970 120.940 7.290 121.000 ;
        RECT 8.810 120.985 9.130 121.000 ;
        RECT 7.445 120.940 7.735 120.985 ;
        RECT 8.780 120.940 9.130 120.985 ;
        RECT 6.970 120.800 7.735 120.940 ;
        RECT 8.615 120.800 9.130 120.940 ;
        RECT 6.970 120.740 7.290 120.800 ;
        RECT 7.445 120.755 7.735 120.800 ;
        RECT 8.780 120.755 9.130 120.800 ;
        RECT 8.810 120.740 9.130 120.755 ;
        RECT 10.190 120.940 10.510 121.000 ;
        RECT 14.420 120.940 14.560 121.140 ;
        RECT 15.250 121.080 15.570 121.140 ;
        RECT 23.085 121.095 23.375 121.140 ;
        RECT 10.190 120.800 14.560 120.940 ;
        RECT 10.190 120.740 10.510 120.800 ;
        RECT 14.790 120.740 15.110 121.000 ;
        RECT 15.710 120.740 16.030 121.000 ;
        RECT 17.090 120.985 17.410 121.000 ;
        RECT 17.090 120.755 17.545 120.985 ;
        RECT 17.090 120.740 17.410 120.755 ;
        RECT 18.010 120.740 18.330 121.000 ;
        RECT 18.945 120.755 19.235 120.985 ;
        RECT 19.865 120.755 20.155 120.985 ;
        RECT 20.310 120.940 20.630 121.000 ;
        RECT 20.785 120.940 21.075 120.985 ;
        RECT 20.310 120.800 21.075 120.940 ;
        RECT 23.160 120.940 23.300 121.095 ;
        RECT 24.910 121.080 25.230 121.340 ;
        RECT 25.510 121.280 25.800 121.325 ;
        RECT 27.210 121.280 27.530 121.340 ;
        RECT 25.510 121.140 27.530 121.280 ;
        RECT 25.510 121.095 25.800 121.140 ;
        RECT 27.210 121.080 27.530 121.140 ;
        RECT 28.145 121.280 28.435 121.325 ;
        RECT 29.510 121.280 29.830 121.340 ;
        RECT 28.145 121.140 29.830 121.280 ;
        RECT 28.145 121.095 28.435 121.140 ;
        RECT 26.765 120.940 27.055 120.985 ;
        RECT 28.220 120.940 28.360 121.095 ;
        RECT 29.510 121.080 29.830 121.140 ;
        RECT 23.160 120.800 27.055 120.940 ;
        RECT 12.950 120.600 13.270 120.660 ;
        RECT 15.800 120.600 15.940 120.740 ;
        RECT 12.950 120.460 15.940 120.600 ;
        RECT 16.185 120.600 16.475 120.645 ;
        RECT 16.630 120.600 16.950 120.660 ;
        RECT 19.020 120.600 19.160 120.755 ;
        RECT 16.185 120.460 19.160 120.600 ;
        RECT 12.950 120.400 13.270 120.460 ;
        RECT 16.185 120.415 16.475 120.460 ;
        RECT 16.630 120.400 16.950 120.460 ;
        RECT 14.345 120.260 14.635 120.305 ;
        RECT 15.250 120.260 15.570 120.320 ;
        RECT 14.345 120.120 15.570 120.260 ;
        RECT 14.345 120.075 14.635 120.120 ;
        RECT 15.250 120.060 15.570 120.120 ;
        RECT 15.710 120.260 16.030 120.320 ;
        RECT 19.940 120.260 20.080 120.755 ;
        RECT 20.310 120.740 20.630 120.800 ;
        RECT 20.785 120.755 21.075 120.800 ;
        RECT 26.765 120.755 27.055 120.800 ;
        RECT 27.300 120.800 28.360 120.940 ;
        RECT 30.060 120.940 30.200 121.480 ;
        RECT 32.360 120.985 32.500 121.480 ;
        RECT 39.630 121.480 43.590 121.620 ;
        RECT 39.630 121.435 39.920 121.480 ;
        RECT 41.200 121.435 41.490 121.480 ;
        RECT 43.300 121.435 43.590 121.480 ;
        RECT 48.920 121.480 55.040 121.620 ;
        RECT 55.270 121.620 55.590 121.680 ;
        RECT 59.870 121.620 60.190 121.680 ;
        RECT 55.270 121.480 60.190 121.620 ;
        RECT 35.045 121.280 35.335 121.325 ;
        RECT 36.870 121.280 37.190 121.340 ;
        RECT 35.045 121.140 37.190 121.280 ;
        RECT 35.045 121.095 35.335 121.140 ;
        RECT 36.870 121.080 37.190 121.140 ;
        RECT 39.195 121.280 39.485 121.325 ;
        RECT 41.715 121.280 42.005 121.325 ;
        RECT 42.905 121.280 43.195 121.325 ;
        RECT 39.195 121.140 43.195 121.280 ;
        RECT 39.195 121.095 39.485 121.140 ;
        RECT 41.715 121.095 42.005 121.140 ;
        RECT 42.905 121.095 43.195 121.140 ;
        RECT 31.825 120.940 32.115 120.985 ;
        RECT 30.060 120.800 32.115 120.940 ;
        RECT 24.465 120.600 24.755 120.645 ;
        RECT 25.830 120.600 26.150 120.660 ;
        RECT 27.300 120.600 27.440 120.800 ;
        RECT 31.825 120.755 32.115 120.800 ;
        RECT 32.285 120.755 32.575 120.985 ;
        RECT 34.585 120.940 34.875 120.985 ;
        RECT 37.790 120.940 38.110 121.000 ;
        RECT 34.585 120.800 38.110 120.940 ;
        RECT 34.585 120.755 34.875 120.800 ;
        RECT 37.790 120.740 38.110 120.800 ;
        RECT 42.390 120.985 42.710 121.000 ;
        RECT 42.390 120.940 42.740 120.985 ;
        RECT 43.785 120.940 44.075 120.985 ;
        RECT 46.070 120.940 46.390 121.000 ;
        RECT 48.920 120.985 49.060 121.480 ;
        RECT 55.270 121.420 55.590 121.480 ;
        RECT 59.870 121.420 60.190 121.480 ;
        RECT 62.630 121.620 62.920 121.665 ;
        RECT 64.200 121.620 64.490 121.665 ;
        RECT 66.300 121.620 66.590 121.665 ;
        RECT 62.630 121.480 66.590 121.620 ;
        RECT 62.630 121.435 62.920 121.480 ;
        RECT 64.200 121.435 64.490 121.480 ;
        RECT 66.300 121.435 66.590 121.480 ;
        RECT 52.970 121.080 53.290 121.340 ;
        RECT 53.430 121.080 53.750 121.340 ;
        RECT 57.110 121.280 57.430 121.340 ;
        RECT 60.790 121.280 61.110 121.340 ;
        RECT 66.860 121.325 67.000 121.820 ;
        RECT 71.370 121.820 74.910 121.960 ;
        RECT 71.370 121.760 71.690 121.820 ;
        RECT 74.590 121.760 74.910 121.820 ;
        RECT 77.350 121.760 77.670 122.020 ;
        RECT 77.810 121.760 78.130 122.020 ;
        RECT 68.150 121.620 68.470 121.680 ;
        RECT 69.990 121.620 70.310 121.680 ;
        RECT 68.150 121.480 70.310 121.620 ;
        RECT 68.150 121.420 68.470 121.480 ;
        RECT 69.990 121.420 70.310 121.480 ;
        RECT 72.750 121.420 73.070 121.680 ;
        RECT 75.510 121.620 75.830 121.680 ;
        RECT 75.510 121.480 78.960 121.620 ;
        RECT 75.510 121.420 75.830 121.480 ;
        RECT 56.280 121.140 57.430 121.280 ;
        RECT 42.390 120.800 42.905 120.940 ;
        RECT 43.785 120.800 46.390 120.940 ;
        RECT 42.390 120.755 42.740 120.800 ;
        RECT 43.785 120.755 44.075 120.800 ;
        RECT 42.390 120.740 42.710 120.755 ;
        RECT 46.070 120.740 46.390 120.800 ;
        RECT 48.845 120.755 49.135 120.985 ;
        RECT 49.290 120.740 49.610 121.000 ;
        RECT 56.280 120.985 56.420 121.140 ;
        RECT 57.110 121.080 57.430 121.140 ;
        RECT 57.660 121.140 61.110 121.280 ;
        RECT 50.225 120.940 50.515 120.985 ;
        RECT 56.205 120.940 56.495 120.985 ;
        RECT 50.225 120.800 56.495 120.940 ;
        RECT 50.225 120.755 50.515 120.800 ;
        RECT 56.205 120.755 56.495 120.800 ;
        RECT 56.650 120.740 56.970 121.000 ;
        RECT 57.660 120.985 57.800 121.140 ;
        RECT 60.790 121.080 61.110 121.140 ;
        RECT 62.195 121.280 62.485 121.325 ;
        RECT 64.715 121.280 65.005 121.325 ;
        RECT 65.905 121.280 66.195 121.325 ;
        RECT 62.195 121.140 66.195 121.280 ;
        RECT 62.195 121.095 62.485 121.140 ;
        RECT 64.715 121.095 65.005 121.140 ;
        RECT 65.905 121.095 66.195 121.140 ;
        RECT 66.785 121.095 67.075 121.325 ;
        RECT 69.070 121.280 69.390 121.340 ;
        RECT 68.700 121.140 69.390 121.280 ;
        RECT 57.585 120.755 57.875 120.985 ;
        RECT 58.045 120.940 58.335 120.985 ;
        RECT 58.490 120.940 58.810 121.000 ;
        RECT 58.045 120.800 58.810 120.940 ;
        RECT 58.045 120.755 58.335 120.800 ;
        RECT 58.490 120.740 58.810 120.800 ;
        RECT 58.965 120.940 59.255 120.985 ;
        RECT 61.250 120.940 61.570 121.000 ;
        RECT 58.965 120.800 61.570 120.940 ;
        RECT 58.965 120.755 59.255 120.800 ;
        RECT 61.250 120.740 61.570 120.800 ;
        RECT 67.705 120.940 67.995 120.985 ;
        RECT 68.150 120.940 68.470 121.000 ;
        RECT 68.700 120.985 68.840 121.140 ;
        RECT 69.070 121.080 69.390 121.140 ;
        RECT 69.530 121.280 69.850 121.340 ;
        RECT 72.840 121.280 72.980 121.420 ;
        RECT 69.530 121.140 76.200 121.280 ;
        RECT 69.530 121.080 69.850 121.140 ;
        RECT 71.920 120.985 72.060 121.140 ;
        RECT 67.705 120.800 68.470 120.940 ;
        RECT 67.705 120.755 67.995 120.800 ;
        RECT 68.150 120.740 68.470 120.800 ;
        RECT 68.625 120.755 68.915 120.985 ;
        RECT 71.845 120.755 72.135 120.985 ;
        RECT 72.290 120.740 72.610 121.000 ;
        RECT 72.765 120.740 73.055 120.970 ;
        RECT 73.685 120.940 73.975 120.985 ;
        RECT 74.145 120.940 74.435 120.985 ;
        RECT 74.590 120.940 74.910 121.000 ;
        RECT 73.685 120.800 74.910 120.940 ;
        RECT 73.685 120.755 73.975 120.800 ;
        RECT 74.145 120.755 74.435 120.800 ;
        RECT 74.590 120.740 74.910 120.800 ;
        RECT 75.050 120.740 75.370 121.000 ;
        RECT 76.060 120.985 76.200 121.140 ;
        RECT 75.525 120.755 75.815 120.985 ;
        RECT 75.985 120.755 76.275 120.985 ;
        RECT 77.810 120.940 78.130 121.000 ;
        RECT 78.820 120.985 78.960 121.480 ;
        RECT 78.745 120.940 79.035 120.985 ;
        RECT 77.810 120.800 79.035 120.940 ;
        RECT 24.465 120.460 27.440 120.600 ;
        RECT 27.670 120.600 27.990 120.660 ;
        RECT 29.190 120.600 29.480 120.645 ;
        RECT 27.670 120.460 29.480 120.600 ;
        RECT 24.465 120.415 24.755 120.460 ;
        RECT 25.830 120.400 26.150 120.460 ;
        RECT 27.670 120.400 27.990 120.460 ;
        RECT 29.190 120.415 29.480 120.460 ;
        RECT 30.430 120.400 30.750 120.660 ;
        RECT 49.765 120.600 50.055 120.645 ;
        RECT 62.630 120.600 62.950 120.660 ;
        RECT 49.765 120.460 62.950 120.600 ;
        RECT 49.765 120.415 50.055 120.460 ;
        RECT 62.630 120.400 62.950 120.460 ;
        RECT 64.930 120.600 65.250 120.660 ;
        RECT 65.450 120.600 65.740 120.645 ;
        RECT 64.930 120.460 65.740 120.600 ;
        RECT 64.930 120.400 65.250 120.460 ;
        RECT 65.450 120.415 65.740 120.460 ;
        RECT 69.545 120.600 69.835 120.645 ;
        RECT 72.840 120.600 72.980 120.740 ;
        RECT 69.545 120.460 72.980 120.600 ;
        RECT 75.600 120.600 75.740 120.755 ;
        RECT 77.810 120.740 78.130 120.800 ;
        RECT 78.745 120.755 79.035 120.800 ;
        RECT 80.585 120.940 80.875 120.985 ;
        RECT 81.030 120.940 81.350 121.000 ;
        RECT 80.585 120.800 81.350 120.940 ;
        RECT 80.585 120.755 80.875 120.800 ;
        RECT 81.030 120.740 81.350 120.800 ;
        RECT 76.890 120.600 77.210 120.660 ;
        RECT 75.600 120.460 77.210 120.600 ;
        RECT 69.545 120.415 69.835 120.460 ;
        RECT 76.890 120.400 77.210 120.460 ;
        RECT 79.190 120.400 79.510 120.660 ;
        RECT 79.650 120.600 79.970 120.660 ;
        RECT 81.950 120.600 82.270 120.660 ;
        RECT 79.650 120.460 82.270 120.600 ;
        RECT 79.650 120.400 79.970 120.460 ;
        RECT 81.950 120.400 82.270 120.460 ;
        RECT 15.710 120.120 20.080 120.260 ;
        RECT 20.310 120.260 20.630 120.320 ;
        RECT 21.245 120.260 21.535 120.305 ;
        RECT 20.310 120.120 21.535 120.260 ;
        RECT 15.710 120.060 16.030 120.120 ;
        RECT 20.310 120.060 20.630 120.120 ;
        RECT 21.245 120.075 21.535 120.120 ;
        RECT 26.305 120.260 26.595 120.305 ;
        RECT 26.750 120.260 27.070 120.320 ;
        RECT 26.305 120.120 27.070 120.260 ;
        RECT 26.305 120.075 26.595 120.120 ;
        RECT 26.750 120.060 27.070 120.120 ;
        RECT 27.210 120.260 27.530 120.320 ;
        RECT 28.605 120.260 28.895 120.305 ;
        RECT 27.210 120.120 28.895 120.260 ;
        RECT 27.210 120.060 27.530 120.120 ;
        RECT 28.605 120.075 28.895 120.120 ;
        RECT 29.985 120.260 30.275 120.305 ;
        RECT 30.890 120.260 31.210 120.320 ;
        RECT 29.985 120.120 31.210 120.260 ;
        RECT 29.985 120.075 30.275 120.120 ;
        RECT 30.890 120.060 31.210 120.120 ;
        RECT 31.350 120.060 31.670 120.320 ;
        RECT 48.370 120.060 48.690 120.320 ;
        RECT 52.525 120.260 52.815 120.305 ;
        RECT 54.810 120.260 55.130 120.320 ;
        RECT 52.525 120.120 55.130 120.260 ;
        RECT 52.525 120.075 52.815 120.120 ;
        RECT 54.810 120.060 55.130 120.120 ;
        RECT 55.285 120.260 55.575 120.305 ;
        RECT 55.730 120.260 56.050 120.320 ;
        RECT 56.650 120.260 56.970 120.320 ;
        RECT 55.285 120.120 56.970 120.260 ;
        RECT 55.285 120.075 55.575 120.120 ;
        RECT 55.730 120.060 56.050 120.120 ;
        RECT 56.650 120.060 56.970 120.120 ;
        RECT 57.110 120.060 57.430 120.320 ;
        RECT 58.490 120.060 58.810 120.320 ;
        RECT 70.450 120.060 70.770 120.320 ;
        RECT 70.910 120.260 71.230 120.320 ;
        RECT 79.280 120.260 79.420 120.400 ;
        RECT 70.910 120.120 79.420 120.260 ;
        RECT 70.910 120.060 71.230 120.120 ;
        RECT 5.520 119.440 83.260 119.920 ;
        RECT 14.790 119.040 15.110 119.300 ;
        RECT 52.970 119.040 53.290 119.300 ;
        RECT 64.010 119.240 64.330 119.300 ;
        RECT 64.930 119.240 65.250 119.300 ;
        RECT 57.660 119.100 61.020 119.240 ;
        RECT 57.660 118.960 57.800 119.100 ;
        RECT 28.130 118.900 28.450 118.960 ;
        RECT 7.060 118.760 28.450 118.900 ;
        RECT 7.060 118.620 7.200 118.760 ;
        RECT 6.970 118.360 7.290 118.620 ;
        RECT 8.350 118.605 8.670 118.620 ;
        RECT 8.320 118.375 8.670 118.605 ;
        RECT 8.350 118.360 8.670 118.375 ;
        RECT 14.330 118.360 14.650 118.620 ;
        RECT 15.250 118.360 15.570 118.620 ;
        RECT 15.710 118.360 16.030 118.620 ;
        RECT 16.630 118.360 16.950 118.620 ;
        RECT 17.090 118.360 17.410 118.620 ;
        RECT 17.565 118.375 17.855 118.605 ;
        RECT 18.470 118.560 18.790 118.620 ;
        RECT 20.785 118.560 21.075 118.605 ;
        RECT 18.470 118.420 21.075 118.560 ;
        RECT 7.865 118.220 8.155 118.265 ;
        RECT 9.055 118.220 9.345 118.265 ;
        RECT 11.575 118.220 11.865 118.265 ;
        RECT 7.865 118.080 11.865 118.220 ;
        RECT 15.340 118.220 15.480 118.360 ;
        RECT 17.640 118.220 17.780 118.375 ;
        RECT 18.470 118.360 18.790 118.420 ;
        RECT 20.785 118.375 21.075 118.420 ;
        RECT 21.230 118.360 21.550 118.620 ;
        RECT 24.080 118.605 24.220 118.760 ;
        RECT 28.130 118.700 28.450 118.760 ;
        RECT 46.070 118.900 46.390 118.960 ;
        RECT 57.570 118.900 57.890 118.960 ;
        RECT 46.070 118.760 57.890 118.900 ;
        RECT 46.070 118.700 46.390 118.760 ;
        RECT 57.570 118.700 57.890 118.760 ;
        RECT 58.965 118.900 59.255 118.945 ;
        RECT 59.870 118.900 60.190 118.960 ;
        RECT 58.965 118.760 60.190 118.900 ;
        RECT 58.965 118.715 59.255 118.760 ;
        RECT 59.870 118.700 60.190 118.760 ;
        RECT 22.625 118.375 22.915 118.605 ;
        RECT 24.005 118.375 24.295 118.605 ;
        RECT 25.340 118.560 25.630 118.605 ;
        RECT 26.750 118.560 27.070 118.620 ;
        RECT 25.340 118.420 27.070 118.560 ;
        RECT 25.340 118.375 25.630 118.420 ;
        RECT 15.340 118.080 17.780 118.220 ;
        RECT 18.010 118.220 18.330 118.280 ;
        RECT 20.310 118.220 20.630 118.280 ;
        RECT 22.700 118.220 22.840 118.375 ;
        RECT 26.750 118.360 27.070 118.420 ;
        RECT 47.420 118.560 47.710 118.605 ;
        RECT 52.510 118.560 52.830 118.620 ;
        RECT 47.420 118.420 52.830 118.560 ;
        RECT 47.420 118.375 47.710 118.420 ;
        RECT 52.510 118.360 52.830 118.420 ;
        RECT 52.970 118.560 53.290 118.620 ;
        RECT 53.445 118.560 53.735 118.605 ;
        RECT 52.970 118.420 53.735 118.560 ;
        RECT 52.970 118.360 53.290 118.420 ;
        RECT 53.445 118.375 53.735 118.420 ;
        RECT 57.110 118.560 57.430 118.620 ;
        RECT 58.505 118.560 58.795 118.605 ;
        RECT 57.110 118.420 58.795 118.560 ;
        RECT 57.110 118.360 57.430 118.420 ;
        RECT 58.505 118.375 58.795 118.420 ;
        RECT 18.010 118.080 22.840 118.220 ;
        RECT 24.885 118.220 25.175 118.265 ;
        RECT 26.075 118.220 26.365 118.265 ;
        RECT 28.595 118.220 28.885 118.265 ;
        RECT 24.885 118.080 28.885 118.220 ;
        RECT 7.865 118.035 8.155 118.080 ;
        RECT 9.055 118.035 9.345 118.080 ;
        RECT 11.575 118.035 11.865 118.080 ;
        RECT 18.010 118.020 18.330 118.080 ;
        RECT 20.310 118.020 20.630 118.080 ;
        RECT 24.885 118.035 25.175 118.080 ;
        RECT 26.075 118.035 26.365 118.080 ;
        RECT 28.595 118.035 28.885 118.080 ;
        RECT 46.070 118.020 46.390 118.280 ;
        RECT 46.965 118.220 47.255 118.265 ;
        RECT 48.155 118.220 48.445 118.265 ;
        RECT 50.675 118.220 50.965 118.265 ;
        RECT 46.965 118.080 50.965 118.220 ;
        RECT 46.965 118.035 47.255 118.080 ;
        RECT 48.155 118.035 48.445 118.080 ;
        RECT 50.675 118.035 50.965 118.080 ;
        RECT 54.810 118.220 55.130 118.280 ;
        RECT 56.665 118.220 56.955 118.265 ;
        RECT 54.810 118.080 56.955 118.220 ;
        RECT 54.810 118.020 55.130 118.080 ;
        RECT 56.665 118.035 56.955 118.080 ;
        RECT 7.470 117.880 7.760 117.925 ;
        RECT 9.570 117.880 9.860 117.925 ;
        RECT 11.140 117.880 11.430 117.925 ;
        RECT 7.470 117.740 11.430 117.880 ;
        RECT 7.470 117.695 7.760 117.740 ;
        RECT 9.570 117.695 9.860 117.740 ;
        RECT 11.140 117.695 11.430 117.740 ;
        RECT 22.165 117.880 22.455 117.925 ;
        RECT 23.990 117.880 24.310 117.940 ;
        RECT 22.165 117.740 24.310 117.880 ;
        RECT 22.165 117.695 22.455 117.740 ;
        RECT 23.990 117.680 24.310 117.740 ;
        RECT 24.490 117.880 24.780 117.925 ;
        RECT 26.590 117.880 26.880 117.925 ;
        RECT 28.160 117.880 28.450 117.925 ;
        RECT 24.490 117.740 28.450 117.880 ;
        RECT 24.490 117.695 24.780 117.740 ;
        RECT 26.590 117.695 26.880 117.740 ;
        RECT 28.160 117.695 28.450 117.740 ;
        RECT 46.570 117.880 46.860 117.925 ;
        RECT 48.670 117.880 48.960 117.925 ;
        RECT 50.240 117.880 50.530 117.925 ;
        RECT 46.570 117.740 50.530 117.880 ;
        RECT 46.570 117.695 46.860 117.740 ;
        RECT 48.670 117.695 48.960 117.740 ;
        RECT 50.240 117.695 50.530 117.740 ;
        RECT 56.190 117.880 56.510 117.940 ;
        RECT 56.190 117.740 56.880 117.880 ;
        RECT 56.190 117.680 56.510 117.740 ;
        RECT 13.885 117.540 14.175 117.585 ;
        RECT 14.790 117.540 15.110 117.600 ;
        RECT 13.885 117.400 15.110 117.540 ;
        RECT 13.885 117.355 14.175 117.400 ;
        RECT 14.790 117.340 15.110 117.400 ;
        RECT 18.930 117.340 19.250 117.600 ;
        RECT 19.865 117.540 20.155 117.585 ;
        RECT 20.310 117.540 20.630 117.600 ;
        RECT 19.865 117.400 20.630 117.540 ;
        RECT 19.865 117.355 20.155 117.400 ;
        RECT 20.310 117.340 20.630 117.400 ;
        RECT 29.510 117.540 29.830 117.600 ;
        RECT 30.905 117.540 31.195 117.585 ;
        RECT 31.350 117.540 31.670 117.600 ;
        RECT 29.510 117.400 31.670 117.540 ;
        RECT 29.510 117.340 29.830 117.400 ;
        RECT 30.905 117.355 31.195 117.400 ;
        RECT 31.350 117.340 31.670 117.400 ;
        RECT 49.290 117.540 49.610 117.600 ;
        RECT 55.270 117.540 55.590 117.600 ;
        RECT 49.290 117.400 55.590 117.540 ;
        RECT 56.740 117.540 56.880 117.740 ;
        RECT 57.585 117.695 57.875 117.925 ;
        RECT 58.580 117.880 58.720 118.375 ;
        RECT 59.410 118.360 59.730 118.620 ;
        RECT 60.330 118.360 60.650 118.620 ;
        RECT 60.880 118.220 61.020 119.100 ;
        RECT 64.010 119.100 65.250 119.240 ;
        RECT 64.010 119.040 64.330 119.100 ;
        RECT 64.930 119.040 65.250 119.100 ;
        RECT 65.390 119.040 65.710 119.300 ;
        RECT 69.070 119.240 69.390 119.300 ;
        RECT 72.765 119.240 73.055 119.285 ;
        RECT 66.860 119.100 73.055 119.240 ;
        RECT 66.860 118.900 67.000 119.100 ;
        RECT 69.070 119.040 69.390 119.100 ;
        RECT 72.765 119.055 73.055 119.100 ;
        RECT 75.050 119.040 75.370 119.300 ;
        RECT 76.520 119.100 80.800 119.240 ;
        RECT 62.260 118.760 67.000 118.900 ;
        RECT 67.200 118.900 67.490 118.945 ;
        RECT 70.450 118.900 70.770 118.960 ;
        RECT 67.200 118.760 70.770 118.900 ;
        RECT 62.260 118.605 62.400 118.760 ;
        RECT 67.200 118.715 67.490 118.760 ;
        RECT 70.450 118.700 70.770 118.760 ;
        RECT 70.910 118.900 71.230 118.960 ;
        RECT 74.145 118.900 74.435 118.945 ;
        RECT 76.520 118.900 76.660 119.100 ;
        RECT 80.660 118.945 80.800 119.100 ;
        RECT 79.665 118.900 79.955 118.945 ;
        RECT 70.910 118.760 74.435 118.900 ;
        RECT 70.910 118.700 71.230 118.760 ;
        RECT 74.145 118.715 74.435 118.760 ;
        RECT 75.140 118.760 76.660 118.900 ;
        RECT 76.980 118.760 79.955 118.900 ;
        RECT 62.185 118.375 62.475 118.605 ;
        RECT 62.630 118.360 62.950 118.620 ;
        RECT 63.550 118.360 63.870 118.620 ;
        RECT 64.010 118.360 64.330 118.620 ;
        RECT 64.485 118.560 64.775 118.605 ;
        RECT 65.390 118.560 65.710 118.620 ;
        RECT 64.485 118.420 65.710 118.560 ;
        RECT 64.485 118.375 64.775 118.420 ;
        RECT 65.390 118.360 65.710 118.420 ;
        RECT 73.225 118.560 73.515 118.605 ;
        RECT 75.140 118.560 75.280 118.760 ;
        RECT 76.980 118.620 77.120 118.760 ;
        RECT 79.665 118.715 79.955 118.760 ;
        RECT 80.585 118.900 80.875 118.945 ;
        RECT 82.410 118.900 82.730 118.960 ;
        RECT 80.585 118.760 82.730 118.900 ;
        RECT 80.585 118.715 80.875 118.760 ;
        RECT 82.410 118.700 82.730 118.760 ;
        RECT 73.225 118.420 75.280 118.560 ;
        RECT 73.225 118.375 73.515 118.420 ;
        RECT 75.510 118.360 75.830 118.620 ;
        RECT 76.445 118.375 76.735 118.605 ;
        RECT 65.850 118.220 66.170 118.280 ;
        RECT 60.880 118.080 66.170 118.220 ;
        RECT 65.850 118.020 66.170 118.080 ;
        RECT 66.745 118.220 67.035 118.265 ;
        RECT 67.935 118.220 68.225 118.265 ;
        RECT 70.455 118.220 70.745 118.265 ;
        RECT 75.970 118.220 76.290 118.280 ;
        RECT 66.745 118.080 70.745 118.220 ;
        RECT 66.745 118.035 67.035 118.080 ;
        RECT 67.935 118.035 68.225 118.080 ;
        RECT 70.455 118.035 70.745 118.080 ;
        RECT 71.000 118.080 76.290 118.220 ;
        RECT 76.520 118.220 76.660 118.375 ;
        RECT 76.890 118.360 77.210 118.620 ;
        RECT 77.365 118.560 77.655 118.605 ;
        RECT 77.810 118.560 78.130 118.620 ;
        RECT 77.365 118.420 80.800 118.560 ;
        RECT 77.365 118.375 77.655 118.420 ;
        RECT 77.810 118.360 78.130 118.420 ;
        RECT 80.660 118.280 80.800 118.420 ;
        RECT 78.270 118.220 78.590 118.280 ;
        RECT 79.650 118.220 79.970 118.280 ;
        RECT 76.520 118.080 79.970 118.220 ;
        RECT 60.330 117.880 60.650 117.940 ;
        RECT 58.580 117.740 60.650 117.880 ;
        RECT 57.660 117.540 57.800 117.695 ;
        RECT 60.330 117.680 60.650 117.740 ;
        RECT 66.350 117.880 66.640 117.925 ;
        RECT 68.450 117.880 68.740 117.925 ;
        RECT 70.020 117.880 70.310 117.925 ;
        RECT 66.350 117.740 70.310 117.880 ;
        RECT 66.350 117.695 66.640 117.740 ;
        RECT 68.450 117.695 68.740 117.740 ;
        RECT 70.020 117.695 70.310 117.740 ;
        RECT 56.740 117.400 57.800 117.540 ;
        RECT 61.265 117.540 61.555 117.585 ;
        RECT 71.000 117.540 71.140 118.080 ;
        RECT 75.970 118.020 76.290 118.080 ;
        RECT 78.270 118.020 78.590 118.080 ;
        RECT 79.650 118.020 79.970 118.080 ;
        RECT 80.570 118.020 80.890 118.280 ;
        RECT 71.370 117.880 71.690 117.940 ;
        RECT 78.745 117.880 79.035 117.925 ;
        RECT 71.370 117.740 79.035 117.880 ;
        RECT 71.370 117.680 71.690 117.740 ;
        RECT 78.745 117.695 79.035 117.740 ;
        RECT 61.265 117.400 71.140 117.540 ;
        RECT 76.430 117.540 76.750 117.600 ;
        RECT 78.285 117.540 78.575 117.585 ;
        RECT 76.430 117.400 78.575 117.540 ;
        RECT 49.290 117.340 49.610 117.400 ;
        RECT 55.270 117.340 55.590 117.400 ;
        RECT 61.265 117.355 61.555 117.400 ;
        RECT 76.430 117.340 76.750 117.400 ;
        RECT 78.285 117.355 78.575 117.400 ;
        RECT 5.520 116.720 83.260 117.200 ;
        RECT 7.905 116.520 8.195 116.565 ;
        RECT 8.350 116.520 8.670 116.580 ;
        RECT 7.905 116.380 8.670 116.520 ;
        RECT 7.905 116.335 8.195 116.380 ;
        RECT 8.350 116.320 8.670 116.380 ;
        RECT 12.950 116.320 13.270 116.580 ;
        RECT 14.790 116.520 15.110 116.580 ;
        RECT 16.185 116.520 16.475 116.565 ;
        RECT 14.790 116.380 16.475 116.520 ;
        RECT 14.790 116.320 15.110 116.380 ;
        RECT 16.185 116.335 16.475 116.380 ;
        RECT 40.090 116.320 40.410 116.580 ;
        RECT 43.310 116.520 43.630 116.580 ;
        RECT 45.625 116.520 45.915 116.565 ;
        RECT 51.130 116.520 51.450 116.580 ;
        RECT 43.310 116.380 45.915 116.520 ;
        RECT 43.310 116.320 43.630 116.380 ;
        RECT 45.625 116.335 45.915 116.380 ;
        RECT 48.460 116.380 51.450 116.520 ;
        RECT 13.410 116.180 13.730 116.240 ;
        RECT 9.820 116.040 13.730 116.180 ;
        RECT 9.820 115.885 9.960 116.040 ;
        RECT 13.410 115.980 13.730 116.040 ;
        RECT 15.250 116.180 15.570 116.240 ;
        RECT 15.725 116.180 16.015 116.225 ;
        RECT 28.130 116.180 28.420 116.225 ;
        RECT 29.700 116.180 29.990 116.225 ;
        RECT 31.800 116.180 32.090 116.225 ;
        RECT 15.250 116.040 16.860 116.180 ;
        RECT 15.250 115.980 15.570 116.040 ;
        RECT 15.725 115.995 16.015 116.040 ;
        RECT 16.720 115.900 16.860 116.040 ;
        RECT 28.130 116.040 32.090 116.180 ;
        RECT 28.130 115.995 28.420 116.040 ;
        RECT 29.700 115.995 29.990 116.040 ;
        RECT 31.800 115.995 32.090 116.040 ;
        RECT 35.490 116.180 35.780 116.225 ;
        RECT 37.060 116.180 37.350 116.225 ;
        RECT 39.160 116.180 39.450 116.225 ;
        RECT 35.490 116.040 39.450 116.180 ;
        RECT 35.490 115.995 35.780 116.040 ;
        RECT 37.060 115.995 37.350 116.040 ;
        RECT 39.160 115.995 39.450 116.040 ;
        RECT 9.745 115.655 10.035 115.885 ;
        RECT 10.190 115.840 10.510 115.900 ;
        RECT 11.125 115.840 11.415 115.885 ;
        RECT 10.190 115.700 11.415 115.840 ;
        RECT 10.190 115.640 10.510 115.700 ;
        RECT 11.125 115.655 11.415 115.700 ;
        RECT 16.630 115.640 16.950 115.900 ;
        RECT 27.695 115.840 27.985 115.885 ;
        RECT 30.215 115.840 30.505 115.885 ;
        RECT 31.405 115.840 31.695 115.885 ;
        RECT 27.695 115.700 31.695 115.840 ;
        RECT 27.695 115.655 27.985 115.700 ;
        RECT 30.215 115.655 30.505 115.700 ;
        RECT 31.405 115.655 31.695 115.700 ;
        RECT 35.055 115.840 35.345 115.885 ;
        RECT 37.575 115.840 37.865 115.885 ;
        RECT 38.765 115.840 39.055 115.885 ;
        RECT 35.055 115.700 39.055 115.840 ;
        RECT 35.055 115.655 35.345 115.700 ;
        RECT 37.575 115.655 37.865 115.700 ;
        RECT 38.765 115.655 39.055 115.700 ;
        RECT 39.645 115.840 39.935 115.885 ;
        RECT 41.470 115.840 41.790 115.900 ;
        RECT 39.645 115.700 41.790 115.840 ;
        RECT 39.645 115.655 39.935 115.700 ;
        RECT 41.470 115.640 41.790 115.700 ;
        RECT 47.450 115.840 47.770 115.900 ;
        RECT 48.460 115.885 48.600 116.380 ;
        RECT 51.130 116.320 51.450 116.380 ;
        RECT 52.510 116.520 52.830 116.580 ;
        RECT 53.445 116.520 53.735 116.565 ;
        RECT 52.510 116.380 53.735 116.520 ;
        RECT 52.510 116.320 52.830 116.380 ;
        RECT 53.445 116.335 53.735 116.380 ;
        RECT 55.270 116.520 55.590 116.580 ;
        RECT 55.745 116.520 56.035 116.565 ;
        RECT 55.270 116.380 56.035 116.520 ;
        RECT 55.270 116.320 55.590 116.380 ;
        RECT 55.745 116.335 56.035 116.380 ;
        RECT 56.190 116.520 56.510 116.580 ;
        RECT 57.125 116.520 57.415 116.565 ;
        RECT 56.190 116.380 57.415 116.520 ;
        RECT 56.190 116.320 56.510 116.380 ;
        RECT 57.125 116.335 57.415 116.380 ;
        RECT 57.585 116.520 57.875 116.565 ;
        RECT 58.030 116.520 58.350 116.580 ;
        RECT 57.585 116.380 58.350 116.520 ;
        RECT 57.585 116.335 57.875 116.380 ;
        RECT 58.030 116.320 58.350 116.380 ;
        RECT 58.965 116.520 59.255 116.565 ;
        RECT 59.410 116.520 59.730 116.580 ;
        RECT 58.965 116.380 59.730 116.520 ;
        RECT 58.965 116.335 59.255 116.380 ;
        RECT 59.410 116.320 59.730 116.380 ;
        RECT 60.330 116.320 60.650 116.580 ;
        RECT 67.230 116.520 67.550 116.580 ;
        RECT 68.150 116.520 68.470 116.580 ;
        RECT 77.350 116.520 77.670 116.580 ;
        RECT 67.230 116.380 68.470 116.520 ;
        RECT 67.230 116.320 67.550 116.380 ;
        RECT 68.150 116.320 68.470 116.380 ;
        RECT 71.920 116.380 77.670 116.520 ;
        RECT 60.420 116.180 60.560 116.320 ;
        RECT 69.530 116.180 69.850 116.240 ;
        RECT 59.500 116.040 60.560 116.180 ;
        RECT 61.800 116.040 69.850 116.180 ;
        RECT 48.385 115.840 48.675 115.885 ;
        RECT 47.450 115.700 48.675 115.840 ;
        RECT 47.450 115.640 47.770 115.700 ;
        RECT 48.385 115.655 48.675 115.700 ;
        RECT 50.670 115.840 50.990 115.900 ;
        RECT 50.670 115.700 55.500 115.840 ;
        RECT 50.670 115.640 50.990 115.700 ;
        RECT 9.285 115.500 9.575 115.545 ;
        RECT 10.650 115.500 10.970 115.560 ;
        RECT 9.285 115.360 10.970 115.500 ;
        RECT 9.285 115.315 9.575 115.360 ;
        RECT 10.650 115.300 10.970 115.360 ;
        RECT 11.570 115.300 11.890 115.560 ;
        RECT 12.505 115.500 12.795 115.545 ;
        RECT 14.330 115.500 14.650 115.560 ;
        RECT 12.505 115.360 14.650 115.500 ;
        RECT 12.505 115.315 12.795 115.360 ;
        RECT 14.330 115.300 14.650 115.360 ;
        RECT 14.790 115.300 15.110 115.560 ;
        RECT 16.170 115.300 16.490 115.560 ;
        RECT 18.930 115.300 19.250 115.560 ;
        RECT 19.865 115.315 20.155 115.545 ;
        RECT 20.325 115.315 20.615 115.545 ;
        RECT 20.770 115.500 21.090 115.560 ;
        RECT 30.890 115.545 31.210 115.560 ;
        RECT 23.545 115.500 23.835 115.545 ;
        RECT 20.770 115.360 23.835 115.500 ;
        RECT 8.700 115.160 8.990 115.205 ;
        RECT 12.045 115.160 12.335 115.205 ;
        RECT 15.250 115.160 15.570 115.220 ;
        RECT 19.940 115.160 20.080 115.315 ;
        RECT 8.700 115.020 12.335 115.160 ;
        RECT 8.700 114.975 8.990 115.020 ;
        RECT 12.045 114.975 12.335 115.020 ;
        RECT 14.420 115.020 15.570 115.160 ;
        RECT 12.490 114.820 12.810 114.880 ;
        RECT 14.420 114.865 14.560 115.020 ;
        RECT 15.250 114.960 15.570 115.020 ;
        RECT 18.100 115.020 20.080 115.160 ;
        RECT 20.400 115.160 20.540 115.315 ;
        RECT 20.770 115.300 21.090 115.360 ;
        RECT 23.545 115.315 23.835 115.360 ;
        RECT 30.890 115.500 31.240 115.545 ;
        RECT 31.810 115.500 32.130 115.560 ;
        RECT 32.285 115.500 32.575 115.545 ;
        RECT 30.890 115.360 31.405 115.500 ;
        RECT 31.810 115.360 32.575 115.500 ;
        RECT 30.890 115.315 31.240 115.360 ;
        RECT 30.890 115.300 31.210 115.315 ;
        RECT 31.810 115.300 32.130 115.360 ;
        RECT 32.285 115.315 32.575 115.360 ;
        RECT 40.105 115.315 40.395 115.545 ;
        RECT 41.025 115.500 41.315 115.545 ;
        RECT 42.850 115.500 43.170 115.560 ;
        RECT 41.025 115.360 43.170 115.500 ;
        RECT 41.025 115.315 41.315 115.360 ;
        RECT 21.230 115.160 21.550 115.220 ;
        RECT 22.625 115.160 22.915 115.205 ;
        RECT 38.420 115.160 38.710 115.205 ;
        RECT 40.180 115.160 40.320 115.315 ;
        RECT 42.850 115.300 43.170 115.360 ;
        RECT 47.925 115.500 48.215 115.545 ;
        RECT 48.830 115.500 49.150 115.560 ;
        RECT 49.765 115.500 50.055 115.545 ;
        RECT 47.925 115.360 50.055 115.500 ;
        RECT 47.925 115.315 48.215 115.360 ;
        RECT 48.830 115.300 49.150 115.360 ;
        RECT 49.765 115.315 50.055 115.360 ;
        RECT 53.430 115.500 53.750 115.560 ;
        RECT 54.365 115.500 54.655 115.545 ;
        RECT 53.430 115.360 54.655 115.500 ;
        RECT 53.430 115.300 53.750 115.360 ;
        RECT 54.365 115.315 54.655 115.360 ;
        RECT 54.810 115.300 55.130 115.560 ;
        RECT 55.360 115.500 55.500 115.700 ;
        RECT 58.030 115.680 58.350 115.940 ;
        RECT 58.505 115.880 58.795 115.885 ;
        RECT 58.950 115.880 59.270 115.900 ;
        RECT 59.500 115.885 59.640 116.040 ;
        RECT 58.505 115.740 59.270 115.880 ;
        RECT 58.505 115.655 58.795 115.740 ;
        RECT 58.950 115.640 59.270 115.740 ;
        RECT 59.425 115.655 59.715 115.885 ;
        RECT 60.330 115.840 60.650 115.900 ;
        RECT 61.800 115.840 61.940 116.040 ;
        RECT 69.530 115.980 69.850 116.040 ;
        RECT 60.330 115.700 61.940 115.840 ;
        RECT 60.330 115.640 60.650 115.700 ;
        RECT 56.190 115.500 56.510 115.560 ;
        RECT 55.360 115.360 56.510 115.500 ;
        RECT 56.190 115.300 56.510 115.360 ;
        RECT 56.650 115.300 56.970 115.560 ;
        RECT 59.870 115.300 60.190 115.560 ;
        RECT 61.250 115.300 61.570 115.560 ;
        RECT 61.800 115.545 61.940 115.700 ;
        RECT 62.170 115.840 62.490 115.900 ;
        RECT 63.565 115.840 63.855 115.885 ;
        RECT 62.170 115.700 63.855 115.840 ;
        RECT 62.170 115.640 62.490 115.700 ;
        RECT 63.565 115.655 63.855 115.700 ;
        RECT 64.930 115.840 65.250 115.900 ;
        RECT 67.230 115.840 67.550 115.900 ;
        RECT 64.930 115.700 67.550 115.840 ;
        RECT 64.930 115.640 65.250 115.700 ;
        RECT 67.230 115.640 67.550 115.700 ;
        RECT 61.725 115.315 62.015 115.545 ;
        RECT 63.105 115.500 63.395 115.545 ;
        RECT 64.010 115.500 64.330 115.560 ;
        RECT 63.105 115.360 64.330 115.500 ;
        RECT 63.105 115.315 63.395 115.360 ;
        RECT 64.010 115.300 64.330 115.360 ;
        RECT 70.450 115.300 70.770 115.560 ;
        RECT 71.370 115.300 71.690 115.560 ;
        RECT 71.920 115.545 72.060 116.380 ;
        RECT 77.350 116.320 77.670 116.380 ;
        RECT 74.630 116.180 74.920 116.225 ;
        RECT 76.730 116.180 77.020 116.225 ;
        RECT 78.300 116.180 78.590 116.225 ;
        RECT 74.630 116.040 78.590 116.180 ;
        RECT 74.630 115.995 74.920 116.040 ;
        RECT 76.730 115.995 77.020 116.040 ;
        RECT 78.300 115.995 78.590 116.040 ;
        RECT 75.025 115.840 75.315 115.885 ;
        RECT 76.215 115.840 76.505 115.885 ;
        RECT 78.735 115.840 79.025 115.885 ;
        RECT 75.025 115.700 79.025 115.840 ;
        RECT 75.025 115.655 75.315 115.700 ;
        RECT 76.215 115.655 76.505 115.700 ;
        RECT 78.735 115.655 79.025 115.700 ;
        RECT 71.845 115.315 72.135 115.545 ;
        RECT 72.290 115.300 72.610 115.560 ;
        RECT 74.145 115.500 74.435 115.545 ;
        RECT 72.840 115.360 74.435 115.500 ;
        RECT 41.930 115.160 42.250 115.220 ;
        RECT 60.790 115.160 61.110 115.220 ;
        RECT 20.400 115.020 23.760 115.160 ;
        RECT 18.100 114.865 18.240 115.020 ;
        RECT 21.230 114.960 21.550 115.020 ;
        RECT 22.625 114.975 22.915 115.020 ;
        RECT 23.620 114.880 23.760 115.020 ;
        RECT 38.420 115.020 39.860 115.160 ;
        RECT 40.180 115.020 42.250 115.160 ;
        RECT 38.420 114.975 38.710 115.020 ;
        RECT 13.885 114.820 14.175 114.865 ;
        RECT 12.490 114.680 14.175 114.820 ;
        RECT 12.490 114.620 12.810 114.680 ;
        RECT 13.885 114.635 14.175 114.680 ;
        RECT 14.345 114.635 14.635 114.865 ;
        RECT 18.025 114.635 18.315 114.865 ;
        RECT 22.165 114.820 22.455 114.865 ;
        RECT 23.070 114.820 23.390 114.880 ;
        RECT 22.165 114.680 23.390 114.820 ;
        RECT 22.165 114.635 22.455 114.680 ;
        RECT 23.070 114.620 23.390 114.680 ;
        RECT 23.530 114.620 23.850 114.880 ;
        RECT 23.990 114.820 24.310 114.880 ;
        RECT 24.465 114.820 24.755 114.865 ;
        RECT 23.990 114.680 24.755 114.820 ;
        RECT 23.990 114.620 24.310 114.680 ;
        RECT 24.465 114.635 24.755 114.680 ;
        RECT 25.385 114.820 25.675 114.865 ;
        RECT 26.750 114.820 27.070 114.880 ;
        RECT 25.385 114.680 27.070 114.820 ;
        RECT 25.385 114.635 25.675 114.680 ;
        RECT 26.750 114.620 27.070 114.680 ;
        RECT 32.745 114.820 33.035 114.865 ;
        RECT 34.570 114.820 34.890 114.880 ;
        RECT 32.745 114.680 34.890 114.820 ;
        RECT 39.720 114.820 39.860 115.020 ;
        RECT 41.930 114.960 42.250 115.020 ;
        RECT 47.080 115.020 61.110 115.160 ;
        RECT 47.080 114.820 47.220 115.020 ;
        RECT 60.790 114.960 61.110 115.020 ;
        RECT 62.185 115.160 62.475 115.205 ;
        RECT 63.550 115.160 63.870 115.220 ;
        RECT 62.185 115.020 63.870 115.160 ;
        RECT 62.185 114.975 62.475 115.020 ;
        RECT 63.550 114.960 63.870 115.020 ;
        RECT 67.245 115.160 67.535 115.205 ;
        RECT 69.530 115.160 69.850 115.220 ;
        RECT 72.840 115.160 72.980 115.360 ;
        RECT 74.145 115.315 74.435 115.360 ;
        RECT 67.245 115.020 72.980 115.160 ;
        RECT 73.685 115.160 73.975 115.205 ;
        RECT 75.370 115.160 75.660 115.205 ;
        RECT 73.685 115.020 75.660 115.160 ;
        RECT 67.245 114.975 67.535 115.020 ;
        RECT 69.530 114.960 69.850 115.020 ;
        RECT 73.685 114.975 73.975 115.020 ;
        RECT 75.370 114.975 75.660 115.020 ;
        RECT 39.720 114.680 47.220 114.820 ;
        RECT 32.745 114.635 33.035 114.680 ;
        RECT 34.570 114.620 34.890 114.680 ;
        RECT 47.450 114.620 47.770 114.880 ;
        RECT 52.970 114.620 53.290 114.880 ;
        RECT 55.730 114.820 56.050 114.880 ;
        RECT 59.870 114.820 60.190 114.880 ;
        RECT 55.730 114.680 60.190 114.820 ;
        RECT 55.730 114.620 56.050 114.680 ;
        RECT 59.870 114.620 60.190 114.680 ;
        RECT 60.345 114.820 60.635 114.865 ;
        RECT 65.850 114.820 66.170 114.880 ;
        RECT 60.345 114.680 66.170 114.820 ;
        RECT 60.345 114.635 60.635 114.680 ;
        RECT 65.850 114.620 66.170 114.680 ;
        RECT 66.770 114.620 67.090 114.880 ;
        RECT 70.450 114.820 70.770 114.880 ;
        RECT 74.130 114.820 74.450 114.880 ;
        RECT 70.450 114.680 74.450 114.820 ;
        RECT 70.450 114.620 70.770 114.680 ;
        RECT 74.130 114.620 74.450 114.680 ;
        RECT 76.890 114.820 77.210 114.880 ;
        RECT 81.045 114.820 81.335 114.865 ;
        RECT 76.890 114.680 81.335 114.820 ;
        RECT 76.890 114.620 77.210 114.680 ;
        RECT 81.045 114.635 81.335 114.680 ;
        RECT 5.520 114.000 83.260 114.480 ;
        RECT 11.110 113.800 11.430 113.860 ;
        RECT 12.490 113.845 12.810 113.860 ;
        RECT 12.490 113.800 12.875 113.845 ;
        RECT 9.820 113.660 12.875 113.800 ;
        RECT 9.820 113.165 9.960 113.660 ;
        RECT 11.110 113.600 11.430 113.660 ;
        RECT 12.490 113.615 12.875 113.660 ;
        RECT 13.425 113.800 13.715 113.845 ;
        RECT 14.330 113.800 14.650 113.860 ;
        RECT 13.425 113.660 14.650 113.800 ;
        RECT 13.425 113.615 13.715 113.660 ;
        RECT 12.490 113.600 12.810 113.615 ;
        RECT 14.330 113.600 14.650 113.660 ;
        RECT 17.550 113.800 17.870 113.860 ;
        RECT 18.930 113.800 19.250 113.860 ;
        RECT 17.550 113.660 32.960 113.800 ;
        RECT 17.550 113.600 17.870 113.660 ;
        RECT 18.930 113.600 19.250 113.660 ;
        RECT 11.585 113.275 11.875 113.505 ;
        RECT 27.210 113.460 27.530 113.520 ;
        RECT 32.820 113.505 32.960 113.660 ;
        RECT 48.830 113.600 49.150 113.860 ;
        RECT 55.745 113.800 56.035 113.845 ;
        RECT 54.440 113.660 56.035 113.800 ;
        RECT 31.825 113.460 32.115 113.505 ;
        RECT 27.210 113.320 32.115 113.460 ;
        RECT 9.745 112.935 10.035 113.165 ;
        RECT 10.205 112.935 10.495 113.165 ;
        RECT 11.125 113.120 11.415 113.165 ;
        RECT 11.660 113.120 11.800 113.275 ;
        RECT 27.210 113.260 27.530 113.320 ;
        RECT 31.825 113.275 32.115 113.320 ;
        RECT 32.745 113.275 33.035 113.505 ;
        RECT 41.470 113.460 41.790 113.520 ;
        RECT 34.660 113.320 41.790 113.460 ;
        RECT 15.250 113.120 15.570 113.180 ;
        RECT 11.125 112.980 15.570 113.120 ;
        RECT 11.125 112.935 11.415 112.980 ;
        RECT 10.280 112.100 10.420 112.935 ;
        RECT 15.250 112.920 15.570 112.980 ;
        RECT 19.405 113.120 19.695 113.165 ;
        RECT 20.310 113.120 20.630 113.180 ;
        RECT 19.405 112.980 20.630 113.120 ;
        RECT 19.405 112.935 19.695 112.980 ;
        RECT 20.310 112.920 20.630 112.980 ;
        RECT 21.245 113.120 21.535 113.165 ;
        RECT 22.150 113.120 22.470 113.180 ;
        RECT 21.245 112.980 22.470 113.120 ;
        RECT 21.245 112.935 21.535 112.980 ;
        RECT 22.150 112.920 22.470 112.980 ;
        RECT 22.625 112.935 22.915 113.165 ;
        RECT 12.030 112.780 12.350 112.840 ;
        RECT 15.725 112.780 16.015 112.825 ;
        RECT 16.170 112.780 16.490 112.840 ;
        RECT 22.700 112.780 22.840 112.935 ;
        RECT 23.530 112.920 23.850 113.180 ;
        RECT 25.845 112.935 26.135 113.165 ;
        RECT 29.050 113.120 29.370 113.180 ;
        RECT 26.380 112.980 29.370 113.120 ;
        RECT 24.910 112.780 25.230 112.840 ;
        RECT 12.030 112.640 16.490 112.780 ;
        RECT 12.030 112.580 12.350 112.640 ;
        RECT 15.725 112.595 16.015 112.640 ;
        RECT 16.170 112.580 16.490 112.640 ;
        RECT 17.180 112.640 25.230 112.780 ;
        RECT 11.125 112.440 11.415 112.485 ;
        RECT 11.570 112.440 11.890 112.500 ;
        RECT 17.180 112.485 17.320 112.640 ;
        RECT 24.910 112.580 25.230 112.640 ;
        RECT 11.125 112.300 11.890 112.440 ;
        RECT 11.125 112.255 11.415 112.300 ;
        RECT 11.570 112.240 11.890 112.300 ;
        RECT 17.105 112.255 17.395 112.485 ;
        RECT 21.230 112.440 21.550 112.500 ;
        RECT 20.400 112.300 21.550 112.440 ;
        RECT 12.505 112.100 12.795 112.145 ;
        RECT 15.710 112.100 16.030 112.160 ;
        RECT 20.400 112.145 20.540 112.300 ;
        RECT 21.230 112.240 21.550 112.300 ;
        RECT 22.165 112.440 22.455 112.485 ;
        RECT 23.530 112.440 23.850 112.500 ;
        RECT 25.370 112.440 25.690 112.500 ;
        RECT 22.165 112.300 23.850 112.440 ;
        RECT 22.165 112.255 22.455 112.300 ;
        RECT 23.530 112.240 23.850 112.300 ;
        RECT 24.080 112.300 25.690 112.440 ;
        RECT 25.920 112.440 26.060 112.935 ;
        RECT 26.380 112.825 26.520 112.980 ;
        RECT 29.050 112.920 29.370 112.980 ;
        RECT 29.525 113.120 29.815 113.165 ;
        RECT 32.270 113.120 32.590 113.180 ;
        RECT 34.660 113.165 34.800 113.320 ;
        RECT 41.470 113.260 41.790 113.320 ;
        RECT 43.280 113.460 43.570 113.505 ;
        RECT 54.440 113.460 54.580 113.660 ;
        RECT 55.745 113.615 56.035 113.660 ;
        RECT 60.790 113.800 61.110 113.860 ;
        RECT 75.510 113.800 75.830 113.860 ;
        RECT 76.445 113.800 76.735 113.845 ;
        RECT 60.790 113.660 69.760 113.800 ;
        RECT 60.790 113.600 61.110 113.660 ;
        RECT 43.280 113.320 54.580 113.460 ;
        RECT 55.270 113.460 55.590 113.520 ;
        RECT 68.625 113.460 68.915 113.505 ;
        RECT 55.270 113.320 68.915 113.460 ;
        RECT 43.280 113.275 43.570 113.320 ;
        RECT 55.270 113.260 55.590 113.320 ;
        RECT 68.625 113.275 68.915 113.320 ;
        RECT 29.525 112.980 32.590 113.120 ;
        RECT 29.525 112.935 29.815 112.980 ;
        RECT 32.270 112.920 32.590 112.980 ;
        RECT 34.585 112.935 34.875 113.165 ;
        RECT 35.920 113.120 36.210 113.165 ;
        RECT 42.390 113.120 42.710 113.180 ;
        RECT 35.920 112.980 42.710 113.120 ;
        RECT 35.920 112.935 36.210 112.980 ;
        RECT 42.390 112.920 42.710 112.980 ;
        RECT 52.050 112.920 52.370 113.180 ;
        RECT 52.970 112.920 53.290 113.180 ;
        RECT 53.890 112.920 54.210 113.180 ;
        RECT 54.365 112.935 54.655 113.165 ;
        RECT 26.305 112.595 26.595 112.825 ;
        RECT 27.670 112.580 27.990 112.840 ;
        RECT 29.985 112.595 30.275 112.825 ;
        RECT 30.445 112.780 30.735 112.825 ;
        RECT 31.350 112.780 31.670 112.840 ;
        RECT 30.445 112.640 31.670 112.780 ;
        RECT 30.445 112.595 30.735 112.640 ;
        RECT 26.750 112.440 27.070 112.500 ;
        RECT 30.060 112.440 30.200 112.595 ;
        RECT 31.350 112.580 31.670 112.640 ;
        RECT 35.465 112.780 35.755 112.825 ;
        RECT 36.655 112.780 36.945 112.825 ;
        RECT 39.175 112.780 39.465 112.825 ;
        RECT 35.465 112.640 39.465 112.780 ;
        RECT 35.465 112.595 35.755 112.640 ;
        RECT 36.655 112.595 36.945 112.640 ;
        RECT 39.175 112.595 39.465 112.640 ;
        RECT 41.470 112.780 41.790 112.840 ;
        RECT 41.945 112.780 42.235 112.825 ;
        RECT 41.470 112.640 42.235 112.780 ;
        RECT 41.470 112.580 41.790 112.640 ;
        RECT 41.945 112.595 42.235 112.640 ;
        RECT 42.825 112.780 43.115 112.825 ;
        RECT 44.015 112.780 44.305 112.825 ;
        RECT 46.535 112.780 46.825 112.825 ;
        RECT 52.140 112.780 52.280 112.920 ;
        RECT 42.825 112.640 46.825 112.780 ;
        RECT 42.825 112.595 43.115 112.640 ;
        RECT 44.015 112.595 44.305 112.640 ;
        RECT 46.535 112.595 46.825 112.640 ;
        RECT 47.080 112.640 52.280 112.780 ;
        RECT 52.510 112.780 52.830 112.840 ;
        RECT 54.440 112.780 54.580 112.935 ;
        RECT 54.810 112.920 55.130 113.180 ;
        RECT 57.570 112.920 57.890 113.180 ;
        RECT 64.930 113.120 65.250 113.180 ;
        RECT 66.370 113.120 66.660 113.165 ;
        RECT 64.930 112.980 66.660 113.120 ;
        RECT 64.930 112.920 65.250 112.980 ;
        RECT 66.370 112.935 66.660 112.980 ;
        RECT 67.705 112.935 67.995 113.165 ;
        RECT 68.165 112.935 68.455 113.165 ;
        RECT 69.085 113.120 69.375 113.165 ;
        RECT 69.620 113.120 69.760 113.660 ;
        RECT 75.510 113.660 76.735 113.800 ;
        RECT 75.510 113.600 75.830 113.660 ;
        RECT 76.445 113.615 76.735 113.660 ;
        RECT 80.110 113.800 80.430 113.860 ;
        RECT 81.045 113.800 81.335 113.845 ;
        RECT 80.110 113.660 81.335 113.800 ;
        RECT 76.520 113.460 76.660 113.615 ;
        RECT 80.110 113.600 80.430 113.660 ;
        RECT 81.045 113.615 81.335 113.660 ;
        RECT 77.825 113.460 78.115 113.505 ;
        RECT 76.520 113.320 78.115 113.460 ;
        RECT 77.825 113.275 78.115 113.320 ;
        RECT 78.730 113.260 79.050 113.520 ;
        RECT 79.205 113.460 79.495 113.505 ;
        RECT 82.410 113.460 82.730 113.520 ;
        RECT 79.205 113.320 82.730 113.460 ;
        RECT 79.205 113.275 79.495 113.320 ;
        RECT 82.410 113.260 82.730 113.320 ;
        RECT 69.085 112.980 69.760 113.120 ;
        RECT 70.880 113.120 71.170 113.165 ;
        RECT 72.750 113.120 73.070 113.180 ;
        RECT 70.880 112.980 73.070 113.120 ;
        RECT 69.085 112.935 69.375 112.980 ;
        RECT 70.880 112.935 71.170 112.980 ;
        RECT 52.510 112.640 54.580 112.780 ;
        RECT 63.115 112.780 63.405 112.825 ;
        RECT 65.635 112.780 65.925 112.825 ;
        RECT 66.825 112.780 67.115 112.825 ;
        RECT 63.115 112.640 67.115 112.780 ;
        RECT 30.890 112.440 31.210 112.500 ;
        RECT 25.920 112.300 31.210 112.440 ;
        RECT 10.280 111.960 16.030 112.100 ;
        RECT 12.505 111.915 12.795 111.960 ;
        RECT 15.710 111.900 16.030 111.960 ;
        RECT 20.325 111.915 20.615 112.145 ;
        RECT 23.085 112.100 23.375 112.145 ;
        RECT 24.080 112.100 24.220 112.300 ;
        RECT 25.370 112.240 25.690 112.300 ;
        RECT 26.750 112.240 27.070 112.300 ;
        RECT 30.890 112.240 31.210 112.300 ;
        RECT 35.070 112.440 35.360 112.485 ;
        RECT 37.170 112.440 37.460 112.485 ;
        RECT 38.740 112.440 39.030 112.485 ;
        RECT 35.070 112.300 39.030 112.440 ;
        RECT 35.070 112.255 35.360 112.300 ;
        RECT 37.170 112.255 37.460 112.300 ;
        RECT 38.740 112.255 39.030 112.300 ;
        RECT 42.430 112.440 42.720 112.485 ;
        RECT 44.530 112.440 44.820 112.485 ;
        RECT 46.100 112.440 46.390 112.485 ;
        RECT 42.430 112.300 46.390 112.440 ;
        RECT 42.430 112.255 42.720 112.300 ;
        RECT 44.530 112.255 44.820 112.300 ;
        RECT 46.100 112.255 46.390 112.300 ;
        RECT 23.085 111.960 24.220 112.100 ;
        RECT 23.085 111.915 23.375 111.960 ;
        RECT 24.450 111.900 24.770 112.160 ;
        RECT 28.130 111.900 28.450 112.160 ;
        RECT 41.485 112.100 41.775 112.145 ;
        RECT 47.080 112.100 47.220 112.640 ;
        RECT 52.510 112.580 52.830 112.640 ;
        RECT 63.115 112.595 63.405 112.640 ;
        RECT 65.635 112.595 65.925 112.640 ;
        RECT 66.825 112.595 67.115 112.640 ;
        RECT 47.450 112.440 47.770 112.500 ;
        RECT 60.805 112.440 61.095 112.485 ;
        RECT 62.170 112.440 62.490 112.500 ;
        RECT 47.450 112.300 62.490 112.440 ;
        RECT 47.450 112.240 47.770 112.300 ;
        RECT 60.805 112.255 61.095 112.300 ;
        RECT 62.170 112.240 62.490 112.300 ;
        RECT 63.550 112.440 63.840 112.485 ;
        RECT 65.120 112.440 65.410 112.485 ;
        RECT 67.220 112.440 67.510 112.485 ;
        RECT 63.550 112.300 67.510 112.440 ;
        RECT 63.550 112.255 63.840 112.300 ;
        RECT 65.120 112.255 65.410 112.300 ;
        RECT 67.220 112.255 67.510 112.300 ;
        RECT 41.485 111.960 47.220 112.100 ;
        RECT 41.485 111.915 41.775 111.960 ;
        RECT 49.290 111.900 49.610 112.160 ;
        RECT 50.210 112.100 50.530 112.160 ;
        RECT 58.950 112.100 59.270 112.160 ;
        RECT 50.210 111.960 59.270 112.100 ;
        RECT 67.780 112.100 67.920 112.935 ;
        RECT 68.240 112.780 68.380 112.935 ;
        RECT 72.750 112.920 73.070 112.980 ;
        RECT 80.125 113.120 80.415 113.165 ;
        RECT 81.490 113.120 81.810 113.180 ;
        RECT 80.125 112.980 81.810 113.120 ;
        RECT 80.125 112.935 80.415 112.980 ;
        RECT 81.490 112.920 81.810 112.980 ;
        RECT 68.240 112.640 69.300 112.780 ;
        RECT 69.160 112.500 69.300 112.640 ;
        RECT 69.530 112.580 69.850 112.840 ;
        RECT 70.425 112.780 70.715 112.825 ;
        RECT 71.615 112.780 71.905 112.825 ;
        RECT 74.135 112.780 74.425 112.825 ;
        RECT 70.425 112.640 74.425 112.780 ;
        RECT 70.425 112.595 70.715 112.640 ;
        RECT 71.615 112.595 71.905 112.640 ;
        RECT 74.135 112.595 74.425 112.640 ;
        RECT 69.070 112.240 69.390 112.500 ;
        RECT 69.620 112.100 69.760 112.580 ;
        RECT 70.030 112.440 70.320 112.485 ;
        RECT 72.130 112.440 72.420 112.485 ;
        RECT 73.700 112.440 73.990 112.485 ;
        RECT 70.030 112.300 73.990 112.440 ;
        RECT 70.030 112.255 70.320 112.300 ;
        RECT 72.130 112.255 72.420 112.300 ;
        RECT 73.700 112.255 73.990 112.300 ;
        RECT 75.050 112.440 75.370 112.500 ;
        RECT 76.905 112.440 77.195 112.485 ;
        RECT 75.050 112.300 77.195 112.440 ;
        RECT 75.050 112.240 75.370 112.300 ;
        RECT 76.905 112.255 77.195 112.300 ;
        RECT 70.450 112.100 70.770 112.160 ;
        RECT 67.780 111.960 70.770 112.100 ;
        RECT 50.210 111.900 50.530 111.960 ;
        RECT 58.950 111.900 59.270 111.960 ;
        RECT 70.450 111.900 70.770 111.960 ;
        RECT 5.520 111.280 83.260 111.760 ;
        RECT 16.630 110.880 16.950 111.140 ;
        RECT 22.150 111.080 22.470 111.140 ;
        RECT 24.910 111.080 25.230 111.140 ;
        RECT 22.150 110.940 25.230 111.080 ;
        RECT 22.150 110.880 22.470 110.940 ;
        RECT 24.910 110.880 25.230 110.940 ;
        RECT 41.485 111.080 41.775 111.125 ;
        RECT 41.930 111.080 42.250 111.140 ;
        RECT 41.485 110.940 42.250 111.080 ;
        RECT 41.485 110.895 41.775 110.940 ;
        RECT 41.930 110.880 42.250 110.940 ;
        RECT 42.390 111.080 42.710 111.140 ;
        RECT 44.705 111.080 44.995 111.125 ;
        RECT 42.390 110.940 44.995 111.080 ;
        RECT 42.390 110.880 42.710 110.940 ;
        RECT 44.705 110.895 44.995 110.940 ;
        RECT 51.605 111.080 51.895 111.125 ;
        RECT 53.890 111.080 54.210 111.140 ;
        RECT 51.605 110.940 54.210 111.080 ;
        RECT 51.605 110.895 51.895 110.940 ;
        RECT 53.890 110.880 54.210 110.940 ;
        RECT 58.030 111.080 58.350 111.140 ;
        RECT 59.885 111.080 60.175 111.125 ;
        RECT 58.030 110.940 60.175 111.080 ;
        RECT 58.030 110.880 58.350 110.940 ;
        RECT 59.885 110.895 60.175 110.940 ;
        RECT 67.230 111.080 67.550 111.140 ;
        RECT 67.705 111.080 67.995 111.125 ;
        RECT 67.230 110.940 67.995 111.080 ;
        RECT 67.230 110.880 67.550 110.940 ;
        RECT 67.705 110.895 67.995 110.940 ;
        RECT 68.150 110.880 68.470 111.140 ;
        RECT 71.830 111.080 72.150 111.140 ;
        RECT 74.590 111.080 74.910 111.140 ;
        RECT 71.830 110.940 74.910 111.080 ;
        RECT 71.830 110.880 72.150 110.940 ;
        RECT 74.590 110.880 74.910 110.940 ;
        RECT 16.720 110.740 16.860 110.880 ;
        RECT 16.260 110.600 16.860 110.740 ;
        RECT 18.025 110.740 18.315 110.785 ;
        RECT 21.690 110.740 22.010 110.800 ;
        RECT 25.370 110.740 25.690 110.800 ;
        RECT 18.025 110.600 25.690 110.740 ;
        RECT 16.260 110.105 16.400 110.600 ;
        RECT 18.025 110.555 18.315 110.600 ;
        RECT 21.690 110.540 22.010 110.600 ;
        RECT 25.370 110.540 25.690 110.600 ;
        RECT 31.810 110.740 32.130 110.800 ;
        RECT 35.070 110.740 35.360 110.785 ;
        RECT 37.170 110.740 37.460 110.785 ;
        RECT 38.740 110.740 39.030 110.785 ;
        RECT 31.810 110.600 34.800 110.740 ;
        RECT 31.810 110.540 32.130 110.600 ;
        RECT 16.630 110.200 16.950 110.460 ;
        RECT 23.070 110.400 23.390 110.460 ;
        RECT 21.780 110.260 23.390 110.400 ;
        RECT 16.185 109.875 16.475 110.105 ;
        RECT 19.850 109.860 20.170 110.120 ;
        RECT 20.605 110.060 20.895 110.105 ;
        RECT 21.780 110.060 21.920 110.260 ;
        RECT 23.070 110.200 23.390 110.260 ;
        RECT 29.050 110.400 29.370 110.460 ;
        RECT 34.660 110.445 34.800 110.600 ;
        RECT 35.070 110.600 39.030 110.740 ;
        RECT 35.070 110.555 35.360 110.600 ;
        RECT 37.170 110.555 37.460 110.600 ;
        RECT 38.740 110.555 39.030 110.600 ;
        RECT 52.970 110.740 53.290 110.800 ;
        RECT 59.410 110.740 59.730 110.800 ;
        RECT 64.930 110.740 65.250 110.800 ;
        RECT 68.240 110.740 68.380 110.880 ;
        RECT 52.970 110.600 61.940 110.740 ;
        RECT 52.970 110.540 53.290 110.600 ;
        RECT 59.410 110.540 59.730 110.600 ;
        RECT 29.050 110.260 33.420 110.400 ;
        RECT 29.050 110.200 29.370 110.260 ;
        RECT 20.605 109.920 21.920 110.060 ;
        RECT 22.395 110.060 22.685 110.105 ;
        RECT 23.990 110.060 24.310 110.120 ;
        RECT 22.395 109.920 24.310 110.060 ;
        RECT 20.605 109.875 20.895 109.920 ;
        RECT 22.395 109.875 22.685 109.920 ;
        RECT 23.990 109.860 24.310 109.920 ;
        RECT 27.210 110.060 27.530 110.120 ;
        RECT 31.810 110.060 32.130 110.120 ;
        RECT 33.280 110.105 33.420 110.260 ;
        RECT 34.585 110.215 34.875 110.445 ;
        RECT 35.465 110.400 35.755 110.445 ;
        RECT 36.655 110.400 36.945 110.445 ;
        RECT 39.175 110.400 39.465 110.445 ;
        RECT 35.465 110.260 39.465 110.400 ;
        RECT 35.465 110.215 35.755 110.260 ;
        RECT 36.655 110.215 36.945 110.260 ;
        RECT 39.175 110.215 39.465 110.260 ;
        RECT 46.990 110.400 47.310 110.460 ;
        RECT 47.465 110.400 47.755 110.445 ;
        RECT 46.990 110.260 47.755 110.400 ;
        RECT 46.990 110.200 47.310 110.260 ;
        RECT 47.465 110.215 47.755 110.260 ;
        RECT 52.050 110.400 52.370 110.460 ;
        RECT 52.525 110.400 52.815 110.445 ;
        RECT 60.330 110.400 60.650 110.460 ;
        RECT 61.800 110.445 61.940 110.600 ;
        RECT 64.560 110.600 68.380 110.740 ;
        RECT 52.050 110.260 52.815 110.400 ;
        RECT 52.050 110.200 52.370 110.260 ;
        RECT 52.525 110.215 52.815 110.260 ;
        RECT 53.520 110.260 60.650 110.400 ;
        RECT 27.210 109.920 32.130 110.060 ;
        RECT 27.210 109.860 27.530 109.920 ;
        RECT 31.810 109.860 32.130 109.920 ;
        RECT 33.205 109.875 33.495 110.105 ;
        RECT 34.110 110.060 34.430 110.120 ;
        RECT 46.530 110.060 46.850 110.120 ;
        RECT 48.845 110.060 49.135 110.105 ;
        RECT 34.110 109.920 38.940 110.060 ;
        RECT 34.110 109.860 34.430 109.920 ;
        RECT 19.390 109.720 19.710 109.780 ;
        RECT 21.245 109.720 21.535 109.765 ;
        RECT 19.390 109.580 21.535 109.720 ;
        RECT 19.390 109.520 19.710 109.580 ;
        RECT 21.245 109.535 21.535 109.580 ;
        RECT 21.705 109.720 21.995 109.765 ;
        RECT 23.530 109.720 23.850 109.780 ;
        RECT 21.705 109.580 23.850 109.720 ;
        RECT 21.705 109.535 21.995 109.580 ;
        RECT 23.530 109.520 23.850 109.580 ;
        RECT 28.145 109.720 28.435 109.765 ;
        RECT 35.030 109.720 35.350 109.780 ;
        RECT 28.145 109.580 35.350 109.720 ;
        RECT 28.145 109.535 28.435 109.580 ;
        RECT 35.030 109.520 35.350 109.580 ;
        RECT 35.920 109.720 36.210 109.765 ;
        RECT 37.790 109.720 38.110 109.780 ;
        RECT 35.920 109.580 38.110 109.720 ;
        RECT 38.800 109.720 38.940 109.920 ;
        RECT 46.530 109.920 49.135 110.060 ;
        RECT 46.530 109.860 46.850 109.920 ;
        RECT 48.845 109.875 49.135 109.920 ;
        RECT 49.305 109.875 49.595 110.105 ;
        RECT 49.750 110.060 50.070 110.120 ;
        RECT 50.225 110.060 50.515 110.105 ;
        RECT 49.750 109.920 50.515 110.060 ;
        RECT 39.170 109.720 39.490 109.780 ;
        RECT 38.800 109.580 39.490 109.720 ;
        RECT 35.920 109.535 36.210 109.580 ;
        RECT 37.790 109.520 38.110 109.580 ;
        RECT 39.170 109.520 39.490 109.580 ;
        RECT 47.450 109.720 47.770 109.780 ;
        RECT 49.380 109.720 49.520 109.875 ;
        RECT 49.750 109.860 50.070 109.920 ;
        RECT 50.225 109.875 50.515 109.920 ;
        RECT 50.685 110.060 50.975 110.105 ;
        RECT 51.590 110.060 51.910 110.120 ;
        RECT 53.520 110.105 53.660 110.260 ;
        RECT 60.330 110.200 60.650 110.260 ;
        RECT 61.725 110.215 62.015 110.445 ;
        RECT 62.170 110.200 62.490 110.460 ;
        RECT 64.560 110.445 64.700 110.600 ;
        RECT 64.930 110.540 65.250 110.600 ;
        RECT 64.485 110.215 64.775 110.445 ;
        RECT 65.405 110.400 65.695 110.445 ;
        RECT 70.910 110.400 71.230 110.460 ;
        RECT 65.405 110.260 71.230 110.400 ;
        RECT 65.405 110.215 65.695 110.260 ;
        RECT 70.910 110.200 71.230 110.260 ;
        RECT 71.370 110.400 71.690 110.460 ;
        RECT 73.670 110.400 73.990 110.460 ;
        RECT 71.370 110.260 73.990 110.400 ;
        RECT 71.370 110.200 71.690 110.260 ;
        RECT 73.670 110.200 73.990 110.260 ;
        RECT 50.685 109.920 51.910 110.060 ;
        RECT 50.685 109.875 50.975 109.920 ;
        RECT 51.590 109.860 51.910 109.920 ;
        RECT 53.445 109.875 53.735 110.105 ;
        RECT 58.490 110.060 58.810 110.120 ;
        RECT 60.805 110.060 61.095 110.105 ;
        RECT 58.490 109.920 61.095 110.060 ;
        RECT 58.490 109.860 58.810 109.920 ;
        RECT 60.805 109.875 61.095 109.920 ;
        RECT 61.250 109.860 61.570 110.120 ;
        RECT 65.865 110.060 66.155 110.105 ;
        RECT 66.770 110.060 67.090 110.120 ;
        RECT 65.865 109.920 67.090 110.060 ;
        RECT 65.865 109.875 66.155 109.920 ;
        RECT 66.770 109.860 67.090 109.920 ;
        RECT 69.545 110.060 69.835 110.105 ;
        RECT 75.510 110.060 75.830 110.120 ;
        RECT 69.545 109.920 75.830 110.060 ;
        RECT 69.545 109.875 69.835 109.920 ;
        RECT 75.510 109.860 75.830 109.920 ;
        RECT 76.890 109.860 77.210 110.120 ;
        RECT 78.285 110.060 78.575 110.105 ;
        RECT 79.650 110.060 79.970 110.120 ;
        RECT 78.285 109.920 79.970 110.060 ;
        RECT 78.285 109.875 78.575 109.920 ;
        RECT 79.650 109.860 79.970 109.920 ;
        RECT 80.110 109.860 80.430 110.120 ;
        RECT 47.450 109.580 49.520 109.720 ;
        RECT 51.130 109.720 51.450 109.780 ;
        RECT 54.825 109.720 55.115 109.765 ;
        RECT 51.130 109.580 55.115 109.720 ;
        RECT 47.450 109.520 47.770 109.580 ;
        RECT 51.130 109.520 51.450 109.580 ;
        RECT 54.825 109.535 55.115 109.580 ;
        RECT 57.570 109.720 57.890 109.780 ;
        RECT 58.965 109.720 59.255 109.765 ;
        RECT 59.870 109.720 60.190 109.780 ;
        RECT 66.310 109.720 66.630 109.780 ;
        RECT 70.465 109.720 70.755 109.765 ;
        RECT 57.570 109.580 60.190 109.720 ;
        RECT 23.070 109.180 23.390 109.440 ;
        RECT 33.650 109.180 33.970 109.440 ;
        RECT 45.610 109.380 45.930 109.440 ;
        RECT 46.545 109.380 46.835 109.425 ;
        RECT 45.610 109.240 46.835 109.380 ;
        RECT 45.610 109.180 45.930 109.240 ;
        RECT 46.545 109.195 46.835 109.240 ;
        RECT 47.005 109.380 47.295 109.425 ;
        RECT 49.290 109.380 49.610 109.440 ;
        RECT 47.005 109.240 49.610 109.380 ;
        RECT 47.005 109.195 47.295 109.240 ;
        RECT 49.290 109.180 49.610 109.240 ;
        RECT 53.890 109.380 54.210 109.440 ;
        RECT 54.365 109.380 54.655 109.425 ;
        RECT 53.890 109.240 54.655 109.380 ;
        RECT 54.900 109.380 55.040 109.535 ;
        RECT 57.570 109.520 57.890 109.580 ;
        RECT 58.965 109.535 59.255 109.580 ;
        RECT 59.870 109.520 60.190 109.580 ;
        RECT 62.030 109.580 70.755 109.720 ;
        RECT 62.030 109.380 62.170 109.580 ;
        RECT 66.310 109.520 66.630 109.580 ;
        RECT 70.465 109.535 70.755 109.580 ;
        RECT 72.290 109.720 72.610 109.780 ;
        RECT 74.145 109.720 74.435 109.765 ;
        RECT 76.430 109.720 76.750 109.780 ;
        RECT 72.290 109.580 74.435 109.720 ;
        RECT 72.290 109.520 72.610 109.580 ;
        RECT 74.145 109.535 74.435 109.580 ;
        RECT 74.680 109.580 76.750 109.720 ;
        RECT 54.900 109.240 62.170 109.380 ;
        RECT 68.625 109.380 68.915 109.425 ;
        RECT 74.680 109.380 74.820 109.580 ;
        RECT 76.430 109.520 76.750 109.580 ;
        RECT 68.625 109.240 74.820 109.380 ;
        RECT 53.890 109.180 54.210 109.240 ;
        RECT 54.365 109.195 54.655 109.240 ;
        RECT 68.625 109.195 68.915 109.240 ;
        RECT 75.970 109.180 76.290 109.440 ;
        RECT 79.190 109.180 79.510 109.440 ;
        RECT 81.030 109.180 81.350 109.440 ;
        RECT 5.520 108.560 83.260 109.040 ;
        RECT 18.010 108.360 18.330 108.420 ;
        RECT 14.880 108.220 18.330 108.360 ;
        RECT 4.210 107.680 4.530 107.740 ;
        RECT 6.985 107.680 7.275 107.725 ;
        RECT 4.210 107.540 7.275 107.680 ;
        RECT 4.210 107.480 4.530 107.540 ;
        RECT 6.985 107.495 7.275 107.540 ;
        RECT 14.345 107.680 14.635 107.725 ;
        RECT 14.880 107.680 15.020 108.220 ;
        RECT 18.010 108.160 18.330 108.220 ;
        RECT 19.390 108.160 19.710 108.420 ;
        RECT 26.290 108.160 26.610 108.420 ;
        RECT 26.750 108.160 27.070 108.420 ;
        RECT 37.790 108.160 38.110 108.420 ;
        RECT 54.350 108.160 54.670 108.420 ;
        RECT 60.330 108.360 60.650 108.420 ;
        RECT 61.710 108.360 62.030 108.420 ;
        RECT 60.330 108.220 62.030 108.360 ;
        RECT 60.330 108.160 60.650 108.220 ;
        RECT 61.710 108.160 62.030 108.220 ;
        RECT 70.450 108.360 70.770 108.420 ;
        RECT 72.290 108.360 72.610 108.420 ;
        RECT 70.450 108.220 72.610 108.360 ;
        RECT 70.450 108.160 70.770 108.220 ;
        RECT 72.290 108.160 72.610 108.220 ;
        RECT 72.750 108.160 73.070 108.420 ;
        RECT 77.365 108.360 77.655 108.405 ;
        RECT 80.110 108.360 80.430 108.420 ;
        RECT 77.365 108.220 80.430 108.360 ;
        RECT 77.365 108.175 77.655 108.220 ;
        RECT 80.110 108.160 80.430 108.220 ;
        RECT 17.565 108.020 17.855 108.065 ;
        RECT 15.800 107.880 17.855 108.020 ;
        RECT 15.800 107.740 15.940 107.880 ;
        RECT 17.565 107.835 17.855 107.880 ;
        RECT 23.545 108.020 23.835 108.065 ;
        RECT 24.910 108.020 25.230 108.080 ;
        RECT 23.545 107.880 25.230 108.020 ;
        RECT 23.545 107.835 23.835 107.880 ;
        RECT 24.910 107.820 25.230 107.880 ;
        RECT 27.350 108.020 27.640 108.065 ;
        RECT 28.130 108.020 28.450 108.080 ;
        RECT 27.350 107.880 28.450 108.020 ;
        RECT 27.350 107.835 27.640 107.880 ;
        RECT 28.130 107.820 28.450 107.880 ;
        RECT 29.050 108.020 29.370 108.080 ;
        RECT 30.445 108.020 30.735 108.065 ;
        RECT 30.890 108.020 31.210 108.080 ;
        RECT 34.110 108.020 34.430 108.080 ;
        RECT 29.050 107.880 34.430 108.020 ;
        RECT 29.050 107.820 29.370 107.880 ;
        RECT 30.445 107.835 30.735 107.880 ;
        RECT 30.890 107.820 31.210 107.880 ;
        RECT 34.110 107.820 34.430 107.880 ;
        RECT 35.030 108.020 35.350 108.080 ;
        RECT 41.010 108.020 41.330 108.080 ;
        RECT 51.130 108.020 51.450 108.080 ;
        RECT 35.030 107.880 51.450 108.020 ;
        RECT 35.030 107.820 35.350 107.880 ;
        RECT 41.010 107.820 41.330 107.880 ;
        RECT 51.130 107.820 51.450 107.880 ;
        RECT 52.050 108.020 52.370 108.080 ;
        RECT 56.190 108.020 56.510 108.080 ;
        RECT 61.250 108.020 61.570 108.080 ;
        RECT 52.050 107.880 56.510 108.020 ;
        RECT 52.050 107.820 52.370 107.880 ;
        RECT 56.190 107.820 56.510 107.880 ;
        RECT 59.500 107.880 61.570 108.020 ;
        RECT 14.345 107.540 15.020 107.680 ;
        RECT 15.265 107.680 15.555 107.725 ;
        RECT 15.710 107.680 16.030 107.740 ;
        RECT 15.265 107.540 16.030 107.680 ;
        RECT 14.345 107.495 14.635 107.540 ;
        RECT 15.265 107.495 15.555 107.540 ;
        RECT 15.710 107.480 16.030 107.540 ;
        RECT 16.185 107.495 16.475 107.725 ;
        RECT 16.630 107.680 16.950 107.740 ;
        RECT 17.105 107.680 17.395 107.725 ;
        RECT 16.630 107.540 17.395 107.680 ;
        RECT 14.805 107.340 15.095 107.385 ;
        RECT 16.260 107.340 16.400 107.495 ;
        RECT 16.630 107.480 16.950 107.540 ;
        RECT 17.105 107.495 17.395 107.540 ;
        RECT 18.025 107.495 18.315 107.725 ;
        RECT 19.390 107.680 19.710 107.740 ;
        RECT 20.325 107.680 20.615 107.725 ;
        RECT 19.390 107.540 20.615 107.680 ;
        RECT 14.805 107.200 16.400 107.340 ;
        RECT 18.100 107.340 18.240 107.495 ;
        RECT 19.390 107.480 19.710 107.540 ;
        RECT 20.325 107.495 20.615 107.540 ;
        RECT 20.785 107.495 21.075 107.725 ;
        RECT 20.860 107.340 21.000 107.495 ;
        RECT 21.690 107.480 22.010 107.740 ;
        RECT 22.150 107.480 22.470 107.740 ;
        RECT 24.450 107.680 24.770 107.740 ;
        RECT 24.450 107.540 26.060 107.680 ;
        RECT 24.450 107.480 24.770 107.540 ;
        RECT 24.540 107.340 24.680 107.480 ;
        RECT 18.100 107.200 24.680 107.340 ;
        RECT 24.925 107.340 25.215 107.385 ;
        RECT 25.370 107.340 25.690 107.400 ;
        RECT 24.925 107.200 25.690 107.340 ;
        RECT 25.920 107.340 26.060 107.540 ;
        RECT 29.510 107.480 29.830 107.740 ;
        RECT 32.745 107.680 33.035 107.725 ;
        RECT 33.190 107.680 33.510 107.740 ;
        RECT 30.060 107.540 31.580 107.680 ;
        RECT 30.060 107.340 30.200 107.540 ;
        RECT 30.890 107.445 31.180 107.540 ;
        RECT 25.920 107.200 30.200 107.340 ;
        RECT 31.440 107.340 31.580 107.540 ;
        RECT 32.745 107.540 33.510 107.680 ;
        RECT 32.745 107.495 33.035 107.540 ;
        RECT 33.190 107.480 33.510 107.540 ;
        RECT 34.570 107.480 34.890 107.740 ;
        RECT 38.265 107.495 38.555 107.725 ;
        RECT 38.340 107.340 38.480 107.495 ;
        RECT 39.170 107.480 39.490 107.740 ;
        RECT 46.070 107.680 46.390 107.740 ;
        RECT 48.830 107.725 49.150 107.740 ;
        RECT 47.465 107.680 47.755 107.725 ;
        RECT 46.070 107.540 47.755 107.680 ;
        RECT 46.070 107.480 46.390 107.540 ;
        RECT 47.465 107.495 47.755 107.540 ;
        RECT 48.800 107.495 49.150 107.725 ;
        RECT 48.830 107.480 49.150 107.495 ;
        RECT 53.890 107.680 54.210 107.740 ;
        RECT 54.825 107.680 55.115 107.725 ;
        RECT 57.110 107.680 57.430 107.740 ;
        RECT 53.890 107.540 57.430 107.680 ;
        RECT 53.890 107.480 54.210 107.540 ;
        RECT 54.825 107.495 55.115 107.540 ;
        RECT 57.110 107.480 57.430 107.540 ;
        RECT 57.570 107.480 57.890 107.740 ;
        RECT 58.490 107.480 58.810 107.740 ;
        RECT 59.500 107.400 59.640 107.880 ;
        RECT 61.250 107.820 61.570 107.880 ;
        RECT 71.830 107.820 72.150 108.080 ;
        RECT 73.670 108.020 73.990 108.080 ;
        RECT 77.810 108.020 78.130 108.080 ;
        RECT 73.670 107.880 78.130 108.020 ;
        RECT 73.670 107.820 73.990 107.880 ;
        RECT 60.345 107.680 60.635 107.725 ;
        RECT 61.710 107.680 62.030 107.790 ;
        RECT 63.090 107.725 63.410 107.740 ;
        RECT 60.345 107.540 62.030 107.680 ;
        RECT 60.345 107.495 60.635 107.540 ;
        RECT 61.710 107.530 62.030 107.540 ;
        RECT 63.060 107.495 63.410 107.725 ;
        RECT 71.920 107.680 72.060 107.820 ;
        RECT 74.145 107.680 74.435 107.725 ;
        RECT 71.920 107.540 74.435 107.680 ;
        RECT 74.145 107.495 74.435 107.540 ;
        RECT 63.090 107.480 63.410 107.495 ;
        RECT 74.590 107.480 74.910 107.740 ;
        RECT 75.050 107.480 75.370 107.740 ;
        RECT 76.060 107.725 76.200 107.880 ;
        RECT 77.810 107.820 78.130 107.880 ;
        RECT 75.985 107.495 76.275 107.725 ;
        RECT 76.445 107.495 76.735 107.725 ;
        RECT 78.745 107.680 79.035 107.725 ;
        RECT 79.190 107.680 79.510 107.740 ;
        RECT 78.745 107.540 79.510 107.680 ;
        RECT 78.745 107.495 79.035 107.540 ;
        RECT 31.440 107.200 38.480 107.340 ;
        RECT 14.805 107.155 15.095 107.200 ;
        RECT 24.925 107.155 25.215 107.200 ;
        RECT 25.370 107.140 25.690 107.200 ;
        RECT 44.690 107.140 45.010 107.400 ;
        RECT 48.345 107.340 48.635 107.385 ;
        RECT 49.535 107.340 49.825 107.385 ;
        RECT 52.055 107.340 52.345 107.385 ;
        RECT 48.345 107.200 52.345 107.340 ;
        RECT 48.345 107.155 48.635 107.200 ;
        RECT 49.535 107.155 49.825 107.200 ;
        RECT 52.055 107.155 52.345 107.200 ;
        RECT 55.285 107.340 55.575 107.385 ;
        RECT 55.730 107.340 56.050 107.400 ;
        RECT 55.285 107.200 56.050 107.340 ;
        RECT 55.285 107.155 55.575 107.200 ;
        RECT 55.730 107.140 56.050 107.200 ;
        RECT 56.650 107.140 56.970 107.400 ;
        RECT 58.965 107.155 59.255 107.385 ;
        RECT 26.290 107.000 26.610 107.060 ;
        RECT 31.825 107.000 32.115 107.045 ;
        RECT 26.290 106.860 32.115 107.000 ;
        RECT 26.290 106.800 26.610 106.860 ;
        RECT 31.825 106.815 32.115 106.860 ;
        RECT 47.950 107.000 48.240 107.045 ;
        RECT 50.050 107.000 50.340 107.045 ;
        RECT 51.620 107.000 51.910 107.045 ;
        RECT 56.740 107.000 56.880 107.140 ;
        RECT 59.040 107.000 59.180 107.155 ;
        RECT 59.410 107.140 59.730 107.400 ;
        RECT 59.870 107.340 60.190 107.400 ;
        RECT 61.725 107.340 62.015 107.385 ;
        RECT 59.870 107.200 62.015 107.340 ;
        RECT 59.870 107.140 60.190 107.200 ;
        RECT 61.725 107.155 62.015 107.200 ;
        RECT 62.605 107.340 62.895 107.385 ;
        RECT 63.795 107.340 64.085 107.385 ;
        RECT 66.315 107.340 66.605 107.385 ;
        RECT 62.605 107.200 66.605 107.340 ;
        RECT 62.605 107.155 62.895 107.200 ;
        RECT 63.795 107.155 64.085 107.200 ;
        RECT 66.315 107.155 66.605 107.200 ;
        RECT 71.845 107.340 72.135 107.385 ;
        RECT 76.520 107.340 76.660 107.495 ;
        RECT 79.190 107.480 79.510 107.540 ;
        RECT 79.665 107.495 79.955 107.725 ;
        RECT 79.740 107.340 79.880 107.495 ;
        RECT 80.110 107.480 80.430 107.740 ;
        RECT 82.410 107.340 82.730 107.400 ;
        RECT 71.845 107.200 76.660 107.340 ;
        RECT 79.280 107.200 82.730 107.340 ;
        RECT 71.845 107.155 72.135 107.200 ;
        RECT 47.950 106.860 51.910 107.000 ;
        RECT 47.950 106.815 48.240 106.860 ;
        RECT 50.050 106.815 50.340 106.860 ;
        RECT 51.620 106.815 51.910 106.860 ;
        RECT 54.900 106.860 59.180 107.000 ;
        RECT 62.210 107.000 62.500 107.045 ;
        RECT 64.310 107.000 64.600 107.045 ;
        RECT 65.880 107.000 66.170 107.045 ;
        RECT 62.210 106.860 66.170 107.000 ;
        RECT 7.905 106.660 8.195 106.705 ;
        RECT 17.090 106.660 17.410 106.720 ;
        RECT 7.905 106.520 17.410 106.660 ;
        RECT 7.905 106.475 8.195 106.520 ;
        RECT 17.090 106.460 17.410 106.520 ;
        RECT 18.945 106.660 19.235 106.705 ;
        RECT 19.390 106.660 19.710 106.720 ;
        RECT 18.945 106.520 19.710 106.660 ;
        RECT 18.945 106.475 19.235 106.520 ;
        RECT 19.390 106.460 19.710 106.520 ;
        RECT 22.625 106.660 22.915 106.705 ;
        RECT 23.530 106.660 23.850 106.720 ;
        RECT 22.625 106.520 23.850 106.660 ;
        RECT 22.625 106.475 22.915 106.520 ;
        RECT 23.530 106.460 23.850 106.520 ;
        RECT 28.130 106.460 28.450 106.720 ;
        RECT 28.605 106.660 28.895 106.705 ;
        RECT 29.050 106.660 29.370 106.720 ;
        RECT 28.605 106.520 29.370 106.660 ;
        RECT 28.605 106.475 28.895 106.520 ;
        RECT 29.050 106.460 29.370 106.520 ;
        RECT 32.730 106.660 33.050 106.720 ;
        RECT 38.265 106.660 38.555 106.705 ;
        RECT 32.730 106.520 38.555 106.660 ;
        RECT 32.730 106.460 33.050 106.520 ;
        RECT 38.265 106.475 38.555 106.520 ;
        RECT 43.310 106.660 43.630 106.720 ;
        RECT 47.450 106.660 47.770 106.720 ;
        RECT 54.900 106.705 55.040 106.860 ;
        RECT 62.210 106.815 62.500 106.860 ;
        RECT 64.310 106.815 64.600 106.860 ;
        RECT 65.880 106.815 66.170 106.860 ;
        RECT 68.625 107.000 68.915 107.045 ;
        RECT 71.920 107.000 72.060 107.155 ;
        RECT 79.280 107.060 79.420 107.200 ;
        RECT 82.410 107.140 82.730 107.200 ;
        RECT 68.625 106.860 72.060 107.000 ;
        RECT 76.890 107.000 77.210 107.060 ;
        RECT 77.825 107.000 78.115 107.045 ;
        RECT 76.890 106.860 78.115 107.000 ;
        RECT 68.625 106.815 68.915 106.860 ;
        RECT 76.890 106.800 77.210 106.860 ;
        RECT 77.825 106.815 78.115 106.860 ;
        RECT 79.190 106.800 79.510 107.060 ;
        RECT 54.825 106.660 55.115 106.705 ;
        RECT 43.310 106.520 55.115 106.660 ;
        RECT 43.310 106.460 43.630 106.520 ;
        RECT 47.450 106.460 47.770 106.520 ;
        RECT 54.825 106.475 55.115 106.520 ;
        RECT 56.665 106.660 56.955 106.705 ;
        RECT 59.410 106.660 59.730 106.720 ;
        RECT 56.665 106.520 59.730 106.660 ;
        RECT 56.665 106.475 56.955 106.520 ;
        RECT 59.410 106.460 59.730 106.520 ;
        RECT 61.265 106.660 61.555 106.705 ;
        RECT 66.310 106.660 66.630 106.720 ;
        RECT 61.265 106.520 66.630 106.660 ;
        RECT 61.265 106.475 61.555 106.520 ;
        RECT 66.310 106.460 66.630 106.520 ;
        RECT 69.070 106.460 69.390 106.720 ;
        RECT 71.370 106.660 71.690 106.720 ;
        RECT 74.590 106.660 74.910 106.720 ;
        RECT 71.370 106.520 74.910 106.660 ;
        RECT 71.370 106.460 71.690 106.520 ;
        RECT 74.590 106.460 74.910 106.520 ;
        RECT 81.045 106.660 81.335 106.705 ;
        RECT 81.490 106.660 81.810 106.720 ;
        RECT 81.045 106.520 81.810 106.660 ;
        RECT 81.045 106.475 81.335 106.520 ;
        RECT 81.490 106.460 81.810 106.520 ;
        RECT 5.520 105.840 83.260 106.320 ;
        RECT 16.630 105.440 16.950 105.700 ;
        RECT 18.930 105.440 19.250 105.700 ;
        RECT 30.905 105.640 31.195 105.685 ;
        RECT 36.410 105.640 36.730 105.700 ;
        RECT 21.320 105.500 25.140 105.640 ;
        RECT 10.190 105.300 10.510 105.360 ;
        RECT 11.125 105.300 11.415 105.345 ;
        RECT 10.190 105.160 15.480 105.300 ;
        RECT 10.190 105.100 10.510 105.160 ;
        RECT 11.125 105.115 11.415 105.160 ;
        RECT 8.365 104.960 8.655 105.005 ;
        RECT 10.650 104.960 10.970 105.020 ;
        RECT 13.425 104.960 13.715 105.005 ;
        RECT 8.365 104.820 13.715 104.960 ;
        RECT 8.365 104.775 8.655 104.820 ;
        RECT 10.650 104.760 10.970 104.820 ;
        RECT 13.425 104.775 13.715 104.820 ;
        RECT 13.870 104.760 14.190 105.020 ;
        RECT 15.340 105.005 15.480 105.160 ;
        RECT 15.265 104.960 15.555 105.005 ;
        RECT 15.265 104.820 17.780 104.960 ;
        RECT 15.265 104.775 15.555 104.820 ;
        RECT 8.825 104.620 9.115 104.665 ;
        RECT 12.030 104.620 12.350 104.680 ;
        RECT 8.825 104.480 12.350 104.620 ;
        RECT 8.825 104.435 9.115 104.480 ;
        RECT 12.030 104.420 12.350 104.480 ;
        RECT 12.840 104.435 13.130 104.665 ;
        RECT 14.330 104.620 14.650 104.680 ;
        RECT 15.725 104.620 16.015 104.665 ;
        RECT 14.330 104.480 16.015 104.620 ;
        RECT 11.110 104.080 11.430 104.340 ;
        RECT 12.915 104.280 13.055 104.435 ;
        RECT 14.330 104.420 14.650 104.480 ;
        RECT 15.725 104.435 16.015 104.480 ;
        RECT 16.495 104.620 16.785 104.665 ;
        RECT 17.090 104.620 17.410 104.680 ;
        RECT 16.495 104.480 17.410 104.620 ;
        RECT 16.495 104.435 16.785 104.480 ;
        RECT 17.090 104.420 17.410 104.480 ;
        RECT 14.790 104.280 15.110 104.340 ;
        RECT 12.915 104.140 15.110 104.280 ;
        RECT 17.640 104.280 17.780 104.820 ;
        RECT 19.850 104.620 20.140 104.665 ;
        RECT 21.320 104.620 21.460 105.500 ;
        RECT 25.000 105.360 25.140 105.500 ;
        RECT 30.905 105.500 36.730 105.640 ;
        RECT 30.905 105.455 31.195 105.500 ;
        RECT 36.410 105.440 36.730 105.500 ;
        RECT 41.485 105.640 41.775 105.685 ;
        RECT 42.390 105.640 42.710 105.700 ;
        RECT 41.485 105.500 42.710 105.640 ;
        RECT 41.485 105.455 41.775 105.500 ;
        RECT 42.390 105.440 42.710 105.500 ;
        RECT 48.830 105.440 49.150 105.700 ;
        RECT 53.905 105.640 54.195 105.685 ;
        RECT 58.490 105.640 58.810 105.700 ;
        RECT 53.905 105.500 58.810 105.640 ;
        RECT 53.905 105.455 54.195 105.500 ;
        RECT 58.490 105.440 58.810 105.500 ;
        RECT 61.710 105.440 62.030 105.700 ;
        RECT 63.090 105.640 63.410 105.700 ;
        RECT 63.565 105.640 63.855 105.685 ;
        RECT 63.090 105.500 63.855 105.640 ;
        RECT 63.090 105.440 63.410 105.500 ;
        RECT 63.565 105.455 63.855 105.500 ;
        RECT 68.610 105.640 68.930 105.700 ;
        RECT 75.510 105.640 75.830 105.700 ;
        RECT 68.610 105.500 75.830 105.640 ;
        RECT 68.610 105.440 68.930 105.500 ;
        RECT 75.510 105.440 75.830 105.500 ;
        RECT 23.990 105.300 24.310 105.360 ;
        RECT 22.240 105.160 24.310 105.300 ;
        RECT 22.240 105.005 22.380 105.160 ;
        RECT 23.990 105.100 24.310 105.160 ;
        RECT 24.910 105.300 25.230 105.360 ;
        RECT 31.350 105.300 31.670 105.360 ;
        RECT 24.910 105.160 31.670 105.300 ;
        RECT 24.910 105.100 25.230 105.160 ;
        RECT 31.350 105.100 31.670 105.160 ;
        RECT 31.810 105.300 32.130 105.360 ;
        RECT 35.070 105.300 35.360 105.345 ;
        RECT 37.170 105.300 37.460 105.345 ;
        RECT 38.740 105.300 39.030 105.345 ;
        RECT 31.810 105.160 34.800 105.300 ;
        RECT 31.810 105.100 32.130 105.160 ;
        RECT 22.165 104.775 22.455 105.005 ;
        RECT 25.370 104.960 25.690 105.020 ;
        RECT 27.685 104.960 27.975 105.005 ;
        RECT 23.160 104.820 27.975 104.960 ;
        RECT 19.850 104.480 21.460 104.620 ;
        RECT 19.850 104.435 20.140 104.480 ;
        RECT 21.690 104.420 22.010 104.680 ;
        RECT 22.610 104.420 22.930 104.680 ;
        RECT 23.160 104.280 23.300 104.820 ;
        RECT 25.370 104.760 25.690 104.820 ;
        RECT 27.685 104.775 27.975 104.820 ;
        RECT 33.650 104.760 33.970 105.020 ;
        RECT 34.660 105.005 34.800 105.160 ;
        RECT 35.070 105.160 39.030 105.300 ;
        RECT 35.070 105.115 35.360 105.160 ;
        RECT 37.170 105.115 37.460 105.160 ;
        RECT 38.740 105.115 39.030 105.160 ;
        RECT 50.670 105.100 50.990 105.360 ;
        RECT 51.590 105.300 51.910 105.360 ;
        RECT 54.350 105.300 54.670 105.360 ;
        RECT 58.030 105.300 58.350 105.360 ;
        RECT 62.645 105.300 62.935 105.345 ;
        RECT 64.010 105.300 64.330 105.360 ;
        RECT 51.590 105.160 53.660 105.300 ;
        RECT 51.590 105.100 51.910 105.160 ;
        RECT 34.585 104.775 34.875 105.005 ;
        RECT 35.465 104.960 35.755 105.005 ;
        RECT 36.655 104.960 36.945 105.005 ;
        RECT 39.175 104.960 39.465 105.005 ;
        RECT 35.465 104.820 39.465 104.960 ;
        RECT 35.465 104.775 35.755 104.820 ;
        RECT 36.655 104.775 36.945 104.820 ;
        RECT 39.175 104.775 39.465 104.820 ;
        RECT 46.530 104.960 46.850 105.020 ;
        RECT 50.225 104.960 50.515 105.005 ;
        RECT 46.530 104.820 52.280 104.960 ;
        RECT 46.530 104.760 46.850 104.820 ;
        RECT 50.225 104.775 50.515 104.820 ;
        RECT 24.005 104.620 24.295 104.665 ;
        RECT 24.450 104.620 24.770 104.680 ;
        RECT 24.005 104.480 24.770 104.620 ;
        RECT 24.005 104.435 24.295 104.480 ;
        RECT 17.640 104.140 23.300 104.280 ;
        RECT 14.790 104.080 15.110 104.140 ;
        RECT 24.080 104.000 24.220 104.435 ;
        RECT 24.450 104.420 24.770 104.480 ;
        RECT 26.290 104.620 26.610 104.680 ;
        RECT 29.065 104.620 29.355 104.665 ;
        RECT 26.290 104.480 29.355 104.620 ;
        RECT 26.290 104.420 26.610 104.480 ;
        RECT 29.065 104.435 29.355 104.480 ;
        RECT 32.270 104.620 32.590 104.680 ;
        RECT 33.205 104.620 33.495 104.665 ;
        RECT 32.270 104.480 33.495 104.620 ;
        RECT 32.270 104.420 32.590 104.480 ;
        RECT 33.205 104.435 33.495 104.480 ;
        RECT 41.470 104.620 41.790 104.680 ;
        RECT 44.690 104.620 45.010 104.680 ;
        RECT 41.470 104.480 45.010 104.620 ;
        RECT 41.470 104.420 41.790 104.480 ;
        RECT 44.690 104.420 45.010 104.480 ;
        RECT 49.750 104.420 50.070 104.680 ;
        RECT 51.145 104.620 51.435 104.665 ;
        RECT 51.590 104.620 51.910 104.680 ;
        RECT 52.140 104.665 52.280 104.820 ;
        RECT 51.145 104.480 51.910 104.620 ;
        RECT 51.145 104.435 51.435 104.480 ;
        RECT 51.590 104.420 51.910 104.480 ;
        RECT 52.065 104.435 52.355 104.665 ;
        RECT 52.970 104.420 53.290 104.680 ;
        RECT 53.520 104.665 53.660 105.160 ;
        RECT 54.350 105.160 55.040 105.300 ;
        RECT 54.350 105.100 54.670 105.160 ;
        RECT 54.900 105.005 55.040 105.160 ;
        RECT 58.030 105.160 62.400 105.300 ;
        RECT 58.030 105.100 58.350 105.160 ;
        RECT 54.825 104.775 55.115 105.005 ;
        RECT 53.445 104.620 53.735 104.665 ;
        RECT 53.890 104.620 54.210 104.680 ;
        RECT 53.445 104.480 54.210 104.620 ;
        RECT 53.445 104.435 53.735 104.480 ;
        RECT 53.890 104.420 54.210 104.480 ;
        RECT 54.365 104.620 54.655 104.665 ;
        RECT 58.120 104.620 58.260 105.100 ;
        RECT 60.790 104.960 61.110 105.020 ;
        RECT 59.960 104.820 61.110 104.960 ;
        RECT 54.365 104.480 58.260 104.620 ;
        RECT 54.365 104.435 54.655 104.480 ;
        RECT 58.490 104.420 58.810 104.680 ;
        RECT 59.410 104.420 59.730 104.680 ;
        RECT 59.960 104.665 60.100 104.820 ;
        RECT 60.790 104.760 61.110 104.820 ;
        RECT 59.885 104.435 60.175 104.665 ;
        RECT 60.345 104.620 60.635 104.665 ;
        RECT 61.250 104.620 61.570 104.680 ;
        RECT 62.260 104.665 62.400 105.160 ;
        RECT 62.645 105.160 64.330 105.300 ;
        RECT 62.645 105.115 62.935 105.160 ;
        RECT 64.010 105.100 64.330 105.160 ;
        RECT 64.930 105.300 65.250 105.360 ;
        RECT 71.830 105.300 72.150 105.360 ;
        RECT 64.930 105.160 72.150 105.300 ;
        RECT 64.930 105.100 65.250 105.160 ;
        RECT 71.830 105.100 72.150 105.160 ;
        RECT 75.090 105.300 75.380 105.345 ;
        RECT 77.190 105.300 77.480 105.345 ;
        RECT 78.760 105.300 79.050 105.345 ;
        RECT 75.090 105.160 79.050 105.300 ;
        RECT 75.090 105.115 75.380 105.160 ;
        RECT 77.190 105.115 77.480 105.160 ;
        RECT 78.760 105.115 79.050 105.160 ;
        RECT 65.850 104.760 66.170 105.020 ;
        RECT 66.310 104.760 66.630 105.020 ;
        RECT 75.485 104.960 75.775 105.005 ;
        RECT 76.675 104.960 76.965 105.005 ;
        RECT 79.195 104.960 79.485 105.005 ;
        RECT 75.485 104.820 79.485 104.960 ;
        RECT 75.485 104.775 75.775 104.820 ;
        RECT 76.675 104.775 76.965 104.820 ;
        RECT 79.195 104.775 79.485 104.820 ;
        RECT 60.345 104.480 61.570 104.620 ;
        RECT 60.345 104.435 60.635 104.480 ;
        RECT 61.250 104.420 61.570 104.480 ;
        RECT 62.185 104.435 62.475 104.665 ;
        RECT 63.090 104.620 63.410 104.680 ;
        RECT 64.470 104.620 64.790 104.680 ;
        RECT 63.090 104.480 64.790 104.620 ;
        RECT 63.090 104.420 63.410 104.480 ;
        RECT 64.470 104.420 64.790 104.480 ;
        RECT 65.405 104.620 65.695 104.665 ;
        RECT 69.070 104.620 69.390 104.680 ;
        RECT 65.405 104.480 69.390 104.620 ;
        RECT 65.405 104.435 65.695 104.480 ;
        RECT 69.070 104.420 69.390 104.480 ;
        RECT 70.910 104.620 71.230 104.680 ;
        RECT 72.290 104.620 72.610 104.680 ;
        RECT 74.605 104.620 74.895 104.665 ;
        RECT 70.910 104.480 74.895 104.620 ;
        RECT 70.910 104.420 71.230 104.480 ;
        RECT 72.290 104.420 72.610 104.480 ;
        RECT 74.605 104.435 74.895 104.480 ;
        RECT 26.750 104.280 27.070 104.340 ;
        RECT 29.525 104.280 29.815 104.325 ;
        RECT 26.750 104.140 29.815 104.280 ;
        RECT 26.750 104.080 27.070 104.140 ;
        RECT 29.525 104.095 29.815 104.140 ;
        RECT 30.110 104.280 30.400 104.325 ;
        RECT 35.920 104.280 36.210 104.325 ;
        RECT 44.230 104.280 44.550 104.340 ;
        RECT 30.110 104.140 31.580 104.280 ;
        RECT 30.110 104.095 30.400 104.140 ;
        RECT 7.430 103.740 7.750 104.000 ;
        RECT 12.030 103.740 12.350 104.000 ;
        RECT 19.865 103.940 20.155 103.985 ;
        RECT 23.990 103.940 24.310 104.000 ;
        RECT 31.440 103.985 31.580 104.140 ;
        RECT 35.920 104.140 44.550 104.280 ;
        RECT 35.920 104.095 36.210 104.140 ;
        RECT 44.230 104.080 44.550 104.140 ;
        RECT 52.525 104.280 52.815 104.325 ;
        RECT 54.810 104.280 55.130 104.340 ;
        RECT 69.990 104.280 70.310 104.340 ;
        RECT 52.525 104.140 62.400 104.280 ;
        RECT 52.525 104.095 52.815 104.140 ;
        RECT 54.810 104.080 55.130 104.140 ;
        RECT 62.260 104.000 62.400 104.140 ;
        RECT 69.990 104.140 71.600 104.280 ;
        RECT 69.990 104.080 70.310 104.140 ;
        RECT 19.865 103.800 24.310 103.940 ;
        RECT 19.865 103.755 20.155 103.800 ;
        RECT 23.990 103.740 24.310 103.800 ;
        RECT 31.365 103.755 31.655 103.985 ;
        RECT 55.270 103.940 55.590 104.000 ;
        RECT 58.045 103.940 58.335 103.985 ;
        RECT 55.270 103.800 58.335 103.940 ;
        RECT 55.270 103.740 55.590 103.800 ;
        RECT 58.045 103.755 58.335 103.800 ;
        RECT 62.170 103.740 62.490 104.000 ;
        RECT 64.470 103.940 64.790 104.000 ;
        RECT 70.925 103.940 71.215 103.985 ;
        RECT 64.470 103.800 71.215 103.940 ;
        RECT 71.460 103.940 71.600 104.140 ;
        RECT 71.830 104.080 72.150 104.340 ;
        RECT 72.765 104.095 73.055 104.325 ;
        RECT 75.050 104.280 75.370 104.340 ;
        RECT 75.830 104.280 76.120 104.325 ;
        RECT 75.050 104.140 76.120 104.280 ;
        RECT 72.840 103.940 72.980 104.095 ;
        RECT 75.050 104.080 75.370 104.140 ;
        RECT 75.830 104.095 76.120 104.140 ;
        RECT 71.460 103.800 72.980 103.940 ;
        RECT 79.650 103.940 79.970 104.000 ;
        RECT 81.505 103.940 81.795 103.985 ;
        RECT 79.650 103.800 81.795 103.940 ;
        RECT 64.470 103.740 64.790 103.800 ;
        RECT 70.925 103.755 71.215 103.800 ;
        RECT 79.650 103.740 79.970 103.800 ;
        RECT 81.505 103.755 81.795 103.800 ;
        RECT 5.520 103.120 83.260 103.600 ;
        RECT 14.345 102.920 14.635 102.965 ;
        RECT 15.710 102.920 16.030 102.980 ;
        RECT 14.345 102.780 16.030 102.920 ;
        RECT 14.345 102.735 14.635 102.780 ;
        RECT 15.710 102.720 16.030 102.780 ;
        RECT 21.690 102.920 22.010 102.980 ;
        RECT 22.165 102.920 22.455 102.965 ;
        RECT 21.690 102.780 22.455 102.920 ;
        RECT 21.690 102.720 22.010 102.780 ;
        RECT 22.165 102.735 22.455 102.780 ;
        RECT 23.540 102.920 23.830 102.965 ;
        RECT 29.980 102.920 30.270 102.965 ;
        RECT 23.540 102.780 30.270 102.920 ;
        RECT 23.540 102.735 23.830 102.780 ;
        RECT 29.980 102.735 30.270 102.780 ;
        RECT 31.825 102.920 32.115 102.965 ;
        RECT 32.270 102.920 32.590 102.980 ;
        RECT 31.825 102.780 32.590 102.920 ;
        RECT 31.825 102.735 32.115 102.780 ;
        RECT 32.270 102.720 32.590 102.780 ;
        RECT 44.230 102.720 44.550 102.980 ;
        RECT 51.590 102.920 51.910 102.980 ;
        RECT 52.985 102.920 53.275 102.965 ;
        RECT 51.590 102.780 53.275 102.920 ;
        RECT 51.590 102.720 51.910 102.780 ;
        RECT 52.985 102.735 53.275 102.780 ;
        RECT 56.190 102.920 56.510 102.980 ;
        RECT 58.045 102.920 58.335 102.965 ;
        RECT 71.830 102.920 72.150 102.980 ;
        RECT 74.130 102.920 74.450 102.980 ;
        RECT 56.190 102.780 58.335 102.920 ;
        RECT 56.190 102.720 56.510 102.780 ;
        RECT 58.045 102.735 58.335 102.780 ;
        RECT 64.100 102.780 69.300 102.920 ;
        RECT 8.780 102.580 9.070 102.625 ;
        RECT 12.030 102.580 12.350 102.640 ;
        RECT 8.780 102.440 12.350 102.580 ;
        RECT 8.780 102.395 9.070 102.440 ;
        RECT 12.030 102.380 12.350 102.440 ;
        RECT 19.850 102.580 20.170 102.640 ;
        RECT 36.410 102.580 36.730 102.640 ;
        RECT 37.390 102.580 37.680 102.625 ;
        RECT 19.850 102.440 21.460 102.580 ;
        RECT 19.850 102.380 20.170 102.440 ;
        RECT 14.330 102.240 14.650 102.300 ;
        RECT 15.710 102.240 16.030 102.300 ;
        RECT 16.645 102.240 16.935 102.285 ;
        RECT 14.330 102.100 15.480 102.240 ;
        RECT 14.330 102.040 14.650 102.100 ;
        RECT 6.970 101.900 7.290 101.960 ;
        RECT 7.445 101.900 7.735 101.945 ;
        RECT 6.970 101.760 7.735 101.900 ;
        RECT 6.970 101.700 7.290 101.760 ;
        RECT 7.445 101.715 7.735 101.760 ;
        RECT 8.325 101.900 8.615 101.945 ;
        RECT 9.515 101.900 9.805 101.945 ;
        RECT 12.035 101.900 12.325 101.945 ;
        RECT 8.325 101.760 12.325 101.900 ;
        RECT 8.325 101.715 8.615 101.760 ;
        RECT 9.515 101.715 9.805 101.760 ;
        RECT 12.035 101.715 12.325 101.760 ;
        RECT 14.790 101.700 15.110 101.960 ;
        RECT 15.340 101.900 15.480 102.100 ;
        RECT 15.710 102.100 16.935 102.240 ;
        RECT 15.710 102.040 16.030 102.100 ;
        RECT 16.645 102.055 16.935 102.100 ;
        RECT 18.010 102.240 18.330 102.300 ;
        RECT 18.945 102.240 19.235 102.285 ;
        RECT 18.010 102.100 19.235 102.240 ;
        RECT 18.010 102.040 18.330 102.100 ;
        RECT 18.945 102.055 19.235 102.100 ;
        RECT 20.770 102.040 21.090 102.300 ;
        RECT 21.320 102.285 21.460 102.440 ;
        RECT 36.410 102.440 37.680 102.580 ;
        RECT 36.410 102.380 36.730 102.440 ;
        RECT 37.390 102.395 37.680 102.440 ;
        RECT 49.750 102.580 50.070 102.640 ;
        RECT 52.510 102.580 52.830 102.640 ;
        RECT 56.650 102.580 56.970 102.640 ;
        RECT 60.790 102.580 61.110 102.640 ;
        RECT 49.750 102.440 55.960 102.580 ;
        RECT 49.750 102.380 50.070 102.440 ;
        RECT 52.510 102.380 52.830 102.440 ;
        RECT 21.245 102.055 21.535 102.285 ;
        RECT 23.070 102.240 23.390 102.300 ;
        RECT 24.925 102.240 25.215 102.285 ;
        RECT 28.145 102.240 28.435 102.285 ;
        RECT 23.070 102.100 25.215 102.240 ;
        RECT 23.070 102.040 23.390 102.100 ;
        RECT 24.925 102.055 25.215 102.100 ;
        RECT 25.415 102.100 28.435 102.240 ;
        RECT 16.185 101.900 16.475 101.945 ;
        RECT 15.340 101.760 16.475 101.900 ;
        RECT 16.185 101.715 16.475 101.760 ;
        RECT 20.310 101.900 20.630 101.960 ;
        RECT 25.415 101.900 25.555 102.100 ;
        RECT 28.145 102.055 28.435 102.100 ;
        RECT 42.390 102.240 42.710 102.300 ;
        RECT 43.325 102.240 43.615 102.285 ;
        RECT 42.390 102.100 43.615 102.240 ;
        RECT 42.390 102.040 42.710 102.100 ;
        RECT 43.325 102.055 43.615 102.100 ;
        RECT 52.050 102.240 52.370 102.300 ;
        RECT 52.050 102.100 55.040 102.240 ;
        RECT 52.050 102.040 52.370 102.100 ;
        RECT 20.310 101.760 25.555 101.900 ;
        RECT 20.310 101.700 20.630 101.760 ;
        RECT 26.290 101.700 26.610 101.960 ;
        RECT 27.685 101.900 27.975 101.945 ;
        RECT 30.430 101.900 30.750 101.960 ;
        RECT 26.920 101.760 30.750 101.900 ;
        RECT 7.930 101.560 8.220 101.605 ;
        RECT 10.030 101.560 10.320 101.605 ;
        RECT 11.600 101.560 11.890 101.605 ;
        RECT 7.930 101.420 11.890 101.560 ;
        RECT 7.930 101.375 8.220 101.420 ;
        RECT 10.030 101.375 10.320 101.420 ;
        RECT 11.600 101.375 11.890 101.420 ;
        RECT 24.450 101.560 24.770 101.620 ;
        RECT 26.920 101.560 27.060 101.760 ;
        RECT 27.685 101.715 27.975 101.760 ;
        RECT 30.430 101.700 30.750 101.760 ;
        RECT 34.135 101.900 34.425 101.945 ;
        RECT 36.655 101.900 36.945 101.945 ;
        RECT 37.845 101.900 38.135 101.945 ;
        RECT 34.135 101.760 38.135 101.900 ;
        RECT 34.135 101.715 34.425 101.760 ;
        RECT 36.655 101.715 36.945 101.760 ;
        RECT 37.845 101.715 38.135 101.760 ;
        RECT 38.725 101.900 39.015 101.945 ;
        RECT 41.470 101.900 41.790 101.960 ;
        RECT 38.725 101.760 41.790 101.900 ;
        RECT 38.725 101.715 39.015 101.760 ;
        RECT 41.470 101.700 41.790 101.760 ;
        RECT 41.930 101.900 42.250 101.960 ;
        RECT 47.005 101.900 47.295 101.945 ;
        RECT 41.930 101.760 47.295 101.900 ;
        RECT 41.930 101.700 42.250 101.760 ;
        RECT 47.005 101.715 47.295 101.760 ;
        RECT 53.905 101.715 54.195 101.945 ;
        RECT 24.450 101.420 27.060 101.560 ;
        RECT 27.225 101.560 27.515 101.605 ;
        RECT 33.190 101.560 33.510 101.620 ;
        RECT 27.225 101.420 33.510 101.560 ;
        RECT 24.450 101.360 24.770 101.420 ;
        RECT 27.225 101.375 27.515 101.420 ;
        RECT 33.190 101.360 33.510 101.420 ;
        RECT 34.570 101.560 34.860 101.605 ;
        RECT 36.140 101.560 36.430 101.605 ;
        RECT 38.240 101.560 38.530 101.605 ;
        RECT 34.570 101.420 38.530 101.560 ;
        RECT 53.980 101.560 54.120 101.715 ;
        RECT 54.350 101.700 54.670 101.960 ;
        RECT 54.900 101.945 55.040 102.100 ;
        RECT 55.270 102.040 55.590 102.300 ;
        RECT 55.820 102.240 55.960 102.440 ;
        RECT 56.650 102.440 61.110 102.580 ;
        RECT 56.650 102.380 56.970 102.440 ;
        RECT 60.790 102.380 61.110 102.440 ;
        RECT 57.585 102.240 57.875 102.285 ;
        RECT 55.820 102.100 57.875 102.240 ;
        RECT 57.585 102.055 57.875 102.100 ;
        RECT 63.565 102.240 63.855 102.285 ;
        RECT 64.100 102.240 64.240 102.780 ;
        RECT 65.850 102.580 66.170 102.640 ;
        RECT 65.020 102.440 66.170 102.580 ;
        RECT 63.565 102.100 64.240 102.240 ;
        RECT 63.565 102.055 63.855 102.100 ;
        RECT 64.470 102.040 64.790 102.300 ;
        RECT 65.020 102.285 65.160 102.440 ;
        RECT 65.850 102.380 66.170 102.440 ;
        RECT 66.785 102.580 67.075 102.625 ;
        RECT 68.470 102.580 68.760 102.625 ;
        RECT 66.785 102.440 68.760 102.580 ;
        RECT 69.160 102.580 69.300 102.780 ;
        RECT 71.830 102.780 74.450 102.920 ;
        RECT 71.830 102.720 72.150 102.780 ;
        RECT 74.130 102.720 74.450 102.780 ;
        RECT 74.605 102.920 74.895 102.965 ;
        RECT 75.050 102.920 75.370 102.980 ;
        RECT 74.605 102.780 75.370 102.920 ;
        RECT 74.605 102.735 74.895 102.780 ;
        RECT 75.050 102.720 75.370 102.780 ;
        RECT 75.510 102.920 75.830 102.980 ;
        RECT 78.285 102.920 78.575 102.965 ;
        RECT 75.510 102.780 78.575 102.920 ;
        RECT 75.510 102.720 75.830 102.780 ;
        RECT 78.285 102.735 78.575 102.780 ;
        RECT 73.210 102.580 73.530 102.640 ;
        RECT 69.160 102.440 73.530 102.580 ;
        RECT 66.785 102.395 67.075 102.440 ;
        RECT 68.470 102.395 68.760 102.440 ;
        RECT 73.210 102.380 73.530 102.440 ;
        RECT 73.670 102.580 73.990 102.640 ;
        RECT 73.670 102.440 79.420 102.580 ;
        RECT 73.670 102.380 73.990 102.440 ;
        RECT 64.945 102.055 65.235 102.285 ;
        RECT 65.405 102.240 65.695 102.285 ;
        RECT 75.985 102.240 76.275 102.285 ;
        RECT 65.405 102.100 76.275 102.240 ;
        RECT 65.405 102.055 65.695 102.100 ;
        RECT 75.985 102.055 76.275 102.100 ;
        RECT 76.445 102.055 76.735 102.285 ;
        RECT 54.825 101.900 55.115 101.945 ;
        RECT 60.790 101.900 61.110 101.960 ;
        RECT 65.480 101.900 65.620 102.055 ;
        RECT 54.825 101.760 55.500 101.900 ;
        RECT 54.825 101.715 55.115 101.760 ;
        RECT 55.360 101.620 55.500 101.760 ;
        RECT 60.790 101.760 65.620 101.900 ;
        RECT 60.790 101.700 61.110 101.760 ;
        RECT 67.245 101.715 67.535 101.945 ;
        RECT 68.125 101.900 68.415 101.945 ;
        RECT 69.315 101.900 69.605 101.945 ;
        RECT 71.835 101.900 72.125 101.945 ;
        RECT 68.125 101.760 72.125 101.900 ;
        RECT 76.520 101.900 76.660 102.055 ;
        RECT 76.890 102.040 77.210 102.300 ;
        RECT 77.810 102.040 78.130 102.300 ;
        RECT 79.280 102.285 79.420 102.440 ;
        RECT 79.205 102.055 79.495 102.285 ;
        RECT 79.665 102.240 79.955 102.285 ;
        RECT 80.110 102.240 80.430 102.300 ;
        RECT 79.665 102.100 80.430 102.240 ;
        RECT 79.665 102.055 79.955 102.100 ;
        RECT 77.350 101.900 77.670 101.960 ;
        RECT 76.520 101.760 77.670 101.900 ;
        RECT 68.125 101.715 68.415 101.760 ;
        RECT 69.315 101.715 69.605 101.760 ;
        RECT 71.835 101.715 72.125 101.760 ;
        RECT 53.980 101.420 55.040 101.560 ;
        RECT 34.570 101.375 34.860 101.420 ;
        RECT 36.140 101.375 36.430 101.420 ;
        RECT 38.240 101.375 38.530 101.420 ;
        RECT 54.900 101.280 55.040 101.420 ;
        RECT 55.270 101.360 55.590 101.620 ;
        RECT 19.390 101.020 19.710 101.280 ;
        RECT 39.630 101.220 39.950 101.280 ;
        RECT 40.565 101.220 40.855 101.265 ;
        RECT 39.630 101.080 40.855 101.220 ;
        RECT 39.630 101.020 39.950 101.080 ;
        RECT 40.565 101.035 40.855 101.080 ;
        RECT 54.810 101.020 55.130 101.280 ;
        RECT 67.320 101.220 67.460 101.715 ;
        RECT 77.350 101.700 77.670 101.760 ;
        RECT 67.730 101.560 68.020 101.605 ;
        RECT 69.830 101.560 70.120 101.605 ;
        RECT 71.400 101.560 71.690 101.605 ;
        RECT 67.730 101.420 71.690 101.560 ;
        RECT 67.730 101.375 68.020 101.420 ;
        RECT 69.830 101.375 70.120 101.420 ;
        RECT 71.400 101.375 71.690 101.420 ;
        RECT 76.890 101.560 77.210 101.620 ;
        RECT 79.280 101.560 79.420 102.055 ;
        RECT 80.110 102.040 80.430 102.100 ;
        RECT 80.570 102.040 80.890 102.300 ;
        RECT 81.045 102.240 81.335 102.285 ;
        RECT 81.045 102.100 81.720 102.240 ;
        RECT 81.045 102.055 81.335 102.100 ;
        RECT 81.580 101.960 81.720 102.100 ;
        RECT 81.490 101.700 81.810 101.960 ;
        RECT 76.890 101.420 79.420 101.560 ;
        RECT 76.890 101.360 77.210 101.420 ;
        RECT 70.910 101.220 71.230 101.280 ;
        RECT 67.320 101.080 71.230 101.220 ;
        RECT 70.910 101.020 71.230 101.080 ;
        RECT 5.520 100.400 83.260 100.880 ;
        RECT 6.970 100.200 7.290 100.260 ;
        RECT 6.970 100.060 17.780 100.200 ;
        RECT 6.970 100.000 7.290 100.060 ;
        RECT 7.470 99.860 7.760 99.905 ;
        RECT 9.570 99.860 9.860 99.905 ;
        RECT 11.140 99.860 11.430 99.905 ;
        RECT 7.470 99.720 11.430 99.860 ;
        RECT 7.470 99.675 7.760 99.720 ;
        RECT 9.570 99.675 9.860 99.720 ;
        RECT 11.140 99.675 11.430 99.720 ;
        RECT 13.885 99.860 14.175 99.905 ;
        RECT 14.330 99.860 14.650 99.920 ;
        RECT 13.885 99.720 14.650 99.860 ;
        RECT 17.640 99.860 17.780 100.060 ;
        RECT 18.010 100.000 18.330 100.260 ;
        RECT 20.770 100.000 21.090 100.260 ;
        RECT 21.690 100.000 22.010 100.260 ;
        RECT 22.610 100.200 22.930 100.260 ;
        RECT 23.990 100.200 24.310 100.260 ;
        RECT 22.610 100.060 24.310 100.200 ;
        RECT 22.610 100.000 22.930 100.060 ;
        RECT 23.990 100.000 24.310 100.060 ;
        RECT 31.350 100.200 31.670 100.260 ;
        RECT 33.665 100.200 33.955 100.245 ;
        RECT 31.350 100.060 33.955 100.200 ;
        RECT 31.350 100.000 31.670 100.060 ;
        RECT 33.665 100.015 33.955 100.060 ;
        RECT 41.010 100.200 41.330 100.260 ;
        RECT 42.405 100.200 42.695 100.245 ;
        RECT 41.010 100.060 42.695 100.200 ;
        RECT 41.010 100.000 41.330 100.060 ;
        RECT 42.405 100.015 42.695 100.060 ;
        RECT 53.890 100.000 54.210 100.260 ;
        RECT 57.570 100.200 57.890 100.260 ;
        RECT 61.710 100.200 62.030 100.260 ;
        RECT 73.670 100.200 73.990 100.260 ;
        RECT 77.365 100.200 77.655 100.245 ;
        RECT 55.820 100.060 57.890 100.200 ;
        RECT 27.250 99.860 27.540 99.905 ;
        RECT 29.350 99.860 29.640 99.905 ;
        RECT 30.920 99.860 31.210 99.905 ;
        RECT 43.770 99.860 44.090 99.920 ;
        RECT 17.640 99.720 26.520 99.860 ;
        RECT 13.885 99.675 14.175 99.720 ;
        RECT 14.330 99.660 14.650 99.720 ;
        RECT 6.970 99.320 7.290 99.580 ;
        RECT 7.865 99.520 8.155 99.565 ;
        RECT 9.055 99.520 9.345 99.565 ;
        RECT 11.575 99.520 11.865 99.565 ;
        RECT 7.865 99.380 11.865 99.520 ;
        RECT 14.420 99.520 14.560 99.660 ;
        RECT 15.725 99.520 16.015 99.565 ;
        RECT 23.530 99.520 23.850 99.580 ;
        RECT 14.420 99.380 16.015 99.520 ;
        RECT 7.865 99.335 8.155 99.380 ;
        RECT 9.055 99.335 9.345 99.380 ;
        RECT 11.575 99.335 11.865 99.380 ;
        RECT 15.725 99.335 16.015 99.380 ;
        RECT 17.180 99.380 23.850 99.520 ;
        RECT 7.430 99.180 7.750 99.240 ;
        RECT 17.180 99.225 17.320 99.380 ;
        RECT 23.530 99.320 23.850 99.380 ;
        RECT 24.925 99.520 25.215 99.565 ;
        RECT 25.830 99.520 26.150 99.580 ;
        RECT 24.925 99.380 26.150 99.520 ;
        RECT 24.925 99.335 25.215 99.380 ;
        RECT 25.830 99.320 26.150 99.380 ;
        RECT 8.265 99.180 8.555 99.225 ;
        RECT 7.430 99.040 8.555 99.180 ;
        RECT 7.430 98.980 7.750 99.040 ;
        RECT 8.265 98.995 8.555 99.040 ;
        RECT 16.185 98.995 16.475 99.225 ;
        RECT 17.105 98.995 17.395 99.225 ;
        RECT 21.230 99.180 21.550 99.240 ;
        RECT 21.705 99.180 21.995 99.225 ;
        RECT 21.230 99.040 21.995 99.180 ;
        RECT 16.260 98.840 16.400 98.995 ;
        RECT 21.230 98.980 21.550 99.040 ;
        RECT 21.705 98.995 21.995 99.040 ;
        RECT 22.150 98.980 22.470 99.240 ;
        RECT 24.450 98.980 24.770 99.240 ;
        RECT 26.380 99.180 26.520 99.720 ;
        RECT 27.250 99.720 31.210 99.860 ;
        RECT 27.250 99.675 27.540 99.720 ;
        RECT 29.350 99.675 29.640 99.720 ;
        RECT 30.920 99.675 31.210 99.720 ;
        RECT 42.480 99.720 44.090 99.860 ;
        RECT 27.645 99.520 27.935 99.565 ;
        RECT 28.835 99.520 29.125 99.565 ;
        RECT 31.355 99.520 31.645 99.565 ;
        RECT 27.645 99.380 31.645 99.520 ;
        RECT 27.645 99.335 27.935 99.380 ;
        RECT 28.835 99.335 29.125 99.380 ;
        RECT 31.355 99.335 31.645 99.380 ;
        RECT 41.025 99.520 41.315 99.565 ;
        RECT 41.930 99.520 42.250 99.580 ;
        RECT 42.480 99.565 42.620 99.720 ;
        RECT 43.770 99.660 44.090 99.720 ;
        RECT 45.165 99.860 45.455 99.905 ;
        RECT 46.530 99.860 46.850 99.920 ;
        RECT 45.165 99.720 46.850 99.860 ;
        RECT 53.980 99.860 54.120 100.000 ;
        RECT 55.820 99.860 55.960 100.060 ;
        RECT 57.570 100.000 57.890 100.060 ;
        RECT 58.120 100.060 62.030 100.200 ;
        RECT 53.980 99.720 55.960 99.860 ;
        RECT 45.165 99.675 45.455 99.720 ;
        RECT 41.025 99.380 42.250 99.520 ;
        RECT 41.025 99.335 41.315 99.380 ;
        RECT 41.930 99.320 42.250 99.380 ;
        RECT 42.405 99.335 42.695 99.565 ;
        RECT 42.865 99.520 43.155 99.565 ;
        RECT 45.240 99.520 45.380 99.675 ;
        RECT 46.530 99.660 46.850 99.720 ;
        RECT 42.865 99.380 45.380 99.520 ;
        RECT 46.085 99.520 46.375 99.565 ;
        RECT 46.990 99.520 47.310 99.580 ;
        RECT 55.820 99.565 55.960 99.720 ;
        RECT 46.085 99.380 47.310 99.520 ;
        RECT 42.865 99.335 43.155 99.380 ;
        RECT 46.085 99.335 46.375 99.380 ;
        RECT 46.990 99.320 47.310 99.380 ;
        RECT 55.745 99.335 56.035 99.565 ;
        RECT 56.190 99.520 56.510 99.580 ;
        RECT 57.585 99.520 57.875 99.565 ;
        RECT 58.120 99.520 58.260 100.060 ;
        RECT 61.710 100.000 62.030 100.060 ;
        RECT 70.080 100.060 77.655 100.200 ;
        RECT 58.505 99.675 58.795 99.905 ;
        RECT 61.250 99.860 61.570 99.920 ;
        RECT 64.470 99.860 64.790 99.920 ;
        RECT 65.390 99.860 65.710 99.920 ;
        RECT 61.250 99.720 65.710 99.860 ;
        RECT 56.190 99.380 58.260 99.520 ;
        RECT 56.190 99.320 56.510 99.380 ;
        RECT 57.585 99.335 57.875 99.380 ;
        RECT 26.765 99.180 27.055 99.225 ;
        RECT 27.210 99.180 27.530 99.240 ;
        RECT 28.130 99.225 28.450 99.240 ;
        RECT 28.100 99.180 28.450 99.225 ;
        RECT 26.380 99.040 27.530 99.180 ;
        RECT 27.935 99.040 28.450 99.180 ;
        RECT 26.765 98.995 27.055 99.040 ;
        RECT 27.210 98.980 27.530 99.040 ;
        RECT 28.100 98.995 28.450 99.040 ;
        RECT 37.805 98.995 38.095 99.225 ;
        RECT 38.725 98.995 39.015 99.225 ;
        RECT 28.130 98.980 28.450 98.995 ;
        RECT 20.770 98.840 21.090 98.900 ;
        RECT 16.260 98.700 21.090 98.840 ;
        RECT 20.770 98.640 21.090 98.700 ;
        RECT 23.085 98.840 23.375 98.885 ;
        RECT 29.050 98.840 29.370 98.900 ;
        RECT 23.085 98.700 29.370 98.840 ;
        RECT 23.085 98.655 23.375 98.700 ;
        RECT 29.050 98.640 29.370 98.700 ;
        RECT 17.090 98.500 17.410 98.560 ;
        RECT 21.690 98.500 22.010 98.560 ;
        RECT 17.090 98.360 22.010 98.500 ;
        RECT 17.090 98.300 17.410 98.360 ;
        RECT 21.690 98.300 22.010 98.360 ;
        RECT 26.305 98.500 26.595 98.545 ;
        RECT 29.510 98.500 29.830 98.560 ;
        RECT 26.305 98.360 29.830 98.500 ;
        RECT 37.880 98.500 38.020 98.995 ;
        RECT 38.800 98.840 38.940 98.995 ;
        RECT 39.170 98.980 39.490 99.240 ;
        RECT 39.630 98.980 39.950 99.240 ;
        RECT 43.310 98.980 43.630 99.240 ;
        RECT 44.690 98.980 45.010 99.240 ;
        RECT 48.385 99.180 48.675 99.225 ;
        RECT 46.160 99.040 48.675 99.180 ;
        RECT 46.160 98.900 46.300 99.040 ;
        RECT 48.385 98.995 48.675 99.040 ;
        RECT 48.845 99.180 49.135 99.225 ;
        RECT 49.290 99.180 49.610 99.240 ;
        RECT 48.845 99.040 49.610 99.180 ;
        RECT 48.845 98.995 49.135 99.040 ;
        RECT 49.290 98.980 49.610 99.040 ;
        RECT 49.765 98.995 50.055 99.225 ;
        RECT 40.550 98.840 40.870 98.900 ;
        RECT 38.800 98.700 40.870 98.840 ;
        RECT 40.550 98.640 40.870 98.700 ;
        RECT 41.485 98.840 41.775 98.885 ;
        RECT 44.230 98.840 44.550 98.900 ;
        RECT 41.485 98.700 44.550 98.840 ;
        RECT 41.485 98.655 41.775 98.700 ;
        RECT 44.230 98.640 44.550 98.700 ;
        RECT 46.070 98.640 46.390 98.900 ;
        RECT 49.840 98.840 49.980 98.995 ;
        RECT 50.210 98.980 50.530 99.240 ;
        RECT 53.890 99.180 54.210 99.240 ;
        RECT 55.270 99.180 55.590 99.240 ;
        RECT 53.890 99.040 55.590 99.180 ;
        RECT 53.890 98.980 54.210 99.040 ;
        RECT 55.270 98.980 55.590 99.040 ;
        RECT 57.110 98.980 57.430 99.240 ;
        RECT 58.580 99.180 58.720 99.675 ;
        RECT 61.250 99.660 61.570 99.720 ;
        RECT 64.470 99.660 64.790 99.720 ;
        RECT 65.390 99.660 65.710 99.720 ;
        RECT 58.965 99.180 59.255 99.225 ;
        RECT 58.580 99.040 59.255 99.180 ;
        RECT 58.965 98.995 59.255 99.040 ;
        RECT 61.265 98.995 61.555 99.225 ;
        RECT 69.545 99.180 69.835 99.225 ;
        RECT 70.080 99.180 70.220 100.060 ;
        RECT 73.670 100.000 73.990 100.060 ;
        RECT 77.365 100.015 77.655 100.060 ;
        RECT 80.570 100.200 80.890 100.260 ;
        RECT 81.045 100.200 81.335 100.245 ;
        RECT 80.570 100.060 81.335 100.200 ;
        RECT 80.570 100.000 80.890 100.060 ;
        RECT 81.045 100.015 81.335 100.060 ;
        RECT 70.950 99.860 71.240 99.905 ;
        RECT 73.050 99.860 73.340 99.905 ;
        RECT 74.620 99.860 74.910 99.905 ;
        RECT 70.950 99.720 74.910 99.860 ;
        RECT 70.950 99.675 71.240 99.720 ;
        RECT 73.050 99.675 73.340 99.720 ;
        RECT 74.620 99.675 74.910 99.720 ;
        RECT 71.345 99.520 71.635 99.565 ;
        RECT 72.535 99.520 72.825 99.565 ;
        RECT 75.055 99.520 75.345 99.565 ;
        RECT 81.490 99.520 81.810 99.580 ;
        RECT 71.345 99.380 75.345 99.520 ;
        RECT 71.345 99.335 71.635 99.380 ;
        RECT 72.535 99.335 72.825 99.380 ;
        RECT 75.055 99.335 75.345 99.380 ;
        RECT 75.600 99.380 81.810 99.520 ;
        RECT 69.545 99.040 70.220 99.180 ;
        RECT 70.465 99.180 70.755 99.225 ;
        RECT 70.910 99.180 71.230 99.240 ;
        RECT 75.600 99.180 75.740 99.380 ;
        RECT 81.490 99.320 81.810 99.380 ;
        RECT 70.465 99.040 71.230 99.180 ;
        RECT 69.545 98.995 69.835 99.040 ;
        RECT 70.465 98.995 70.755 99.040 ;
        RECT 53.430 98.840 53.750 98.900 ;
        RECT 58.490 98.840 58.810 98.900 ;
        RECT 61.340 98.840 61.480 98.995 ;
        RECT 70.910 98.980 71.230 99.040 ;
        RECT 71.460 99.040 75.740 99.180 ;
        RECT 49.840 98.700 53.750 98.840 ;
        RECT 53.430 98.640 53.750 98.700 ;
        RECT 57.200 98.700 61.480 98.840 ;
        RECT 67.690 98.840 68.010 98.900 ;
        RECT 71.460 98.840 71.600 99.040 ;
        RECT 78.270 98.980 78.590 99.240 ;
        RECT 79.650 98.980 79.970 99.240 ;
        RECT 80.125 99.180 80.415 99.225 ;
        RECT 81.030 99.180 81.350 99.240 ;
        RECT 80.125 99.040 81.350 99.180 ;
        RECT 80.125 98.995 80.415 99.040 ;
        RECT 81.030 98.980 81.350 99.040 ;
        RECT 71.830 98.885 72.150 98.900 ;
        RECT 67.690 98.700 71.600 98.840 ;
        RECT 57.200 98.560 57.340 98.700 ;
        RECT 58.490 98.640 58.810 98.700 ;
        RECT 67.690 98.640 68.010 98.700 ;
        RECT 71.800 98.655 72.150 98.885 ;
        RECT 79.205 98.655 79.495 98.885 ;
        RECT 71.830 98.640 72.150 98.655 ;
        RECT 41.930 98.500 42.250 98.560 ;
        RECT 37.880 98.360 42.250 98.500 ;
        RECT 26.305 98.315 26.595 98.360 ;
        RECT 29.510 98.300 29.830 98.360 ;
        RECT 41.930 98.300 42.250 98.360 ;
        RECT 47.450 98.300 47.770 98.560 ;
        RECT 52.510 98.500 52.830 98.560 ;
        RECT 55.270 98.500 55.590 98.560 ;
        RECT 52.510 98.360 55.590 98.500 ;
        RECT 52.510 98.300 52.830 98.360 ;
        RECT 55.270 98.300 55.590 98.360 ;
        RECT 57.110 98.300 57.430 98.560 ;
        RECT 58.030 98.500 58.350 98.560 ;
        RECT 59.425 98.500 59.715 98.545 ;
        RECT 58.030 98.360 59.715 98.500 ;
        RECT 58.030 98.300 58.350 98.360 ;
        RECT 59.425 98.315 59.715 98.360 ;
        RECT 59.885 98.500 60.175 98.545 ;
        RECT 65.390 98.500 65.710 98.560 ;
        RECT 59.885 98.360 65.710 98.500 ;
        RECT 59.885 98.315 60.175 98.360 ;
        RECT 65.390 98.300 65.710 98.360 ;
        RECT 68.625 98.500 68.915 98.545 ;
        RECT 75.970 98.500 76.290 98.560 ;
        RECT 68.625 98.360 76.290 98.500 ;
        RECT 79.280 98.500 79.420 98.655 ;
        RECT 80.110 98.500 80.430 98.560 ;
        RECT 79.280 98.360 80.430 98.500 ;
        RECT 68.625 98.315 68.915 98.360 ;
        RECT 75.970 98.300 76.290 98.360 ;
        RECT 80.110 98.300 80.430 98.360 ;
        RECT 5.520 97.680 83.260 98.160 ;
        RECT 17.090 97.480 17.410 97.540 ;
        RECT 12.580 97.340 17.410 97.480 ;
        RECT 12.580 97.185 12.720 97.340 ;
        RECT 17.090 97.280 17.410 97.340 ;
        RECT 20.325 97.480 20.615 97.525 ;
        RECT 20.770 97.480 21.090 97.540 ;
        RECT 23.990 97.480 24.310 97.540 ;
        RECT 20.325 97.340 24.310 97.480 ;
        RECT 20.325 97.295 20.615 97.340 ;
        RECT 20.770 97.280 21.090 97.340 ;
        RECT 23.990 97.280 24.310 97.340 ;
        RECT 26.290 97.480 26.610 97.540 ;
        RECT 26.765 97.480 27.055 97.525 ;
        RECT 26.290 97.340 27.055 97.480 ;
        RECT 26.290 97.280 26.610 97.340 ;
        RECT 26.765 97.295 27.055 97.340 ;
        RECT 27.225 97.295 27.515 97.525 ;
        RECT 32.270 97.480 32.590 97.540 ;
        RECT 28.680 97.340 32.590 97.480 ;
        RECT 12.505 96.955 12.795 97.185 ;
        RECT 18.025 97.140 18.315 97.185 ;
        RECT 18.470 97.140 18.790 97.200 ;
        RECT 13.730 97.000 18.790 97.140 ;
        RECT 9.745 96.800 10.035 96.845 ;
        RECT 13.730 96.800 13.870 97.000 ;
        RECT 18.025 96.955 18.315 97.000 ;
        RECT 9.745 96.660 13.870 96.800 ;
        RECT 14.345 96.800 14.635 96.845 ;
        RECT 16.640 96.800 16.930 96.845 ;
        RECT 14.345 96.660 16.930 96.800 ;
        RECT 9.745 96.615 10.035 96.660 ;
        RECT 14.345 96.615 14.635 96.660 ;
        RECT 16.640 96.615 16.930 96.660 ;
        RECT 17.105 96.800 17.395 96.845 ;
        RECT 18.100 96.800 18.240 96.955 ;
        RECT 18.470 96.940 18.790 97.000 ;
        RECT 19.850 97.140 20.170 97.200 ;
        RECT 27.300 97.140 27.440 97.295 ;
        RECT 28.680 97.140 28.820 97.340 ;
        RECT 32.270 97.280 32.590 97.340 ;
        RECT 41.485 97.480 41.775 97.525 ;
        RECT 41.930 97.480 42.250 97.540 ;
        RECT 41.485 97.340 42.250 97.480 ;
        RECT 41.485 97.295 41.775 97.340 ;
        RECT 41.930 97.280 42.250 97.340 ;
        RECT 53.430 97.280 53.750 97.540 ;
        RECT 54.350 97.280 54.670 97.540 ;
        RECT 55.270 97.480 55.590 97.540 ;
        RECT 56.205 97.480 56.495 97.525 ;
        RECT 55.270 97.340 56.495 97.480 ;
        RECT 55.270 97.280 55.590 97.340 ;
        RECT 56.205 97.295 56.495 97.340 ;
        RECT 58.030 97.280 58.350 97.540 ;
        RECT 62.185 97.480 62.475 97.525 ;
        RECT 64.945 97.480 65.235 97.525 ;
        RECT 62.185 97.340 65.235 97.480 ;
        RECT 62.185 97.295 62.475 97.340 ;
        RECT 64.945 97.295 65.235 97.340 ;
        RECT 70.465 97.480 70.755 97.525 ;
        RECT 71.830 97.480 72.150 97.540 ;
        RECT 72.750 97.480 73.070 97.540 ;
        RECT 70.465 97.340 72.150 97.480 ;
        RECT 70.465 97.295 70.755 97.340 ;
        RECT 71.830 97.280 72.150 97.340 ;
        RECT 72.380 97.340 73.070 97.480 ;
        RECT 19.850 97.000 27.440 97.140 ;
        RECT 28.220 97.000 28.820 97.140 ;
        RECT 19.850 96.940 20.170 97.000 ;
        RECT 20.310 96.800 20.630 96.860 ;
        RECT 20.785 96.800 21.075 96.845 ;
        RECT 17.105 96.660 21.075 96.800 ;
        RECT 17.105 96.615 17.395 96.660 ;
        RECT 10.205 96.460 10.495 96.505 ;
        RECT 14.420 96.460 14.560 96.615 ;
        RECT 10.205 96.320 14.560 96.460 ;
        RECT 16.720 96.460 16.860 96.615 ;
        RECT 20.310 96.600 20.630 96.660 ;
        RECT 20.785 96.615 21.075 96.660 ;
        RECT 21.230 96.600 21.550 96.860 ;
        RECT 23.530 96.800 23.850 96.860 ;
        RECT 24.465 96.800 24.755 96.845 ;
        RECT 23.530 96.660 24.755 96.800 ;
        RECT 23.530 96.600 23.850 96.660 ;
        RECT 24.465 96.615 24.755 96.660 ;
        RECT 25.830 96.600 26.150 96.860 ;
        RECT 28.220 96.845 28.360 97.000 ;
        RECT 29.510 96.940 29.830 97.200 ;
        RECT 28.145 96.800 28.435 96.845 ;
        RECT 27.300 96.660 28.435 96.800 ;
        RECT 22.150 96.460 22.470 96.520 ;
        RECT 25.385 96.460 25.675 96.505 ;
        RECT 27.300 96.460 27.440 96.660 ;
        RECT 28.145 96.615 28.435 96.660 ;
        RECT 28.605 96.800 28.895 96.845 ;
        RECT 29.050 96.800 29.370 96.860 ;
        RECT 28.605 96.660 29.370 96.800 ;
        RECT 28.605 96.615 28.895 96.660 ;
        RECT 29.050 96.600 29.370 96.660 ;
        RECT 35.920 96.800 36.210 96.845 ;
        RECT 37.790 96.800 38.110 96.860 ;
        RECT 42.020 96.845 42.160 97.280 ;
        RECT 43.310 97.140 43.630 97.200 ;
        RECT 43.785 97.140 44.075 97.185 ;
        RECT 43.310 97.000 44.075 97.140 ;
        RECT 43.310 96.940 43.630 97.000 ;
        RECT 43.785 96.955 44.075 97.000 ;
        RECT 46.500 97.140 46.790 97.185 ;
        RECT 47.450 97.140 47.770 97.200 ;
        RECT 58.120 97.140 58.260 97.280 ;
        RECT 46.500 97.000 47.770 97.140 ;
        RECT 46.500 96.955 46.790 97.000 ;
        RECT 47.450 96.940 47.770 97.000 ;
        RECT 53.980 97.000 58.260 97.140 ;
        RECT 60.345 97.140 60.635 97.185 ;
        RECT 61.710 97.140 62.030 97.200 ;
        RECT 65.850 97.140 66.170 97.200 ;
        RECT 68.610 97.140 68.930 97.200 ;
        RECT 72.380 97.140 72.520 97.340 ;
        RECT 72.750 97.280 73.070 97.340 ;
        RECT 74.590 97.140 74.910 97.200 ;
        RECT 77.810 97.140 78.130 97.200 ;
        RECT 60.345 97.000 62.170 97.140 ;
        RECT 35.920 96.660 38.110 96.800 ;
        RECT 35.920 96.615 36.210 96.660 ;
        RECT 37.790 96.600 38.110 96.660 ;
        RECT 41.945 96.615 42.235 96.845 ;
        RECT 52.985 96.800 53.275 96.845 ;
        RECT 53.430 96.800 53.750 96.860 ;
        RECT 53.980 96.845 54.120 97.000 ;
        RECT 60.345 96.955 60.635 97.000 ;
        RECT 61.710 96.940 62.170 97.000 ;
        RECT 65.850 97.000 72.520 97.140 ;
        RECT 65.850 96.940 66.170 97.000 ;
        RECT 68.610 96.940 68.930 97.000 ;
        RECT 52.985 96.660 53.750 96.800 ;
        RECT 52.985 96.615 53.275 96.660 ;
        RECT 53.430 96.600 53.750 96.660 ;
        RECT 53.905 96.615 54.195 96.845 ;
        RECT 55.285 96.800 55.575 96.845 ;
        RECT 55.730 96.800 56.050 96.860 ;
        RECT 56.650 96.800 56.970 96.860 ;
        RECT 55.285 96.660 56.050 96.800 ;
        RECT 56.555 96.660 56.970 96.800 ;
        RECT 57.585 96.790 57.875 96.845 ;
        RECT 55.285 96.615 55.575 96.660 ;
        RECT 55.730 96.600 56.050 96.660 ;
        RECT 56.650 96.600 56.970 96.660 ;
        RECT 57.200 96.650 57.875 96.790 ;
        RECT 16.720 96.320 20.080 96.460 ;
        RECT 10.205 96.275 10.495 96.320 ;
        RECT 19.940 96.180 20.080 96.320 ;
        RECT 22.150 96.320 27.440 96.460 ;
        RECT 22.150 96.260 22.470 96.320 ;
        RECT 25.385 96.275 25.675 96.320 ;
        RECT 34.570 96.260 34.890 96.520 ;
        RECT 35.465 96.460 35.755 96.505 ;
        RECT 36.655 96.460 36.945 96.505 ;
        RECT 39.175 96.460 39.465 96.505 ;
        RECT 35.465 96.320 39.465 96.460 ;
        RECT 35.465 96.275 35.755 96.320 ;
        RECT 36.655 96.275 36.945 96.320 ;
        RECT 39.175 96.275 39.465 96.320 ;
        RECT 41.470 96.460 41.790 96.520 ;
        RECT 45.165 96.460 45.455 96.505 ;
        RECT 41.470 96.320 45.455 96.460 ;
        RECT 41.470 96.260 41.790 96.320 ;
        RECT 45.165 96.275 45.455 96.320 ;
        RECT 46.045 96.460 46.335 96.505 ;
        RECT 47.235 96.460 47.525 96.505 ;
        RECT 49.755 96.460 50.045 96.505 ;
        RECT 46.045 96.320 50.045 96.460 ;
        RECT 46.045 96.275 46.335 96.320 ;
        RECT 47.235 96.275 47.525 96.320 ;
        RECT 49.755 96.275 50.045 96.320 ;
        RECT 51.590 96.460 51.910 96.520 ;
        RECT 56.740 96.460 56.880 96.600 ;
        RECT 51.590 96.320 56.880 96.460 ;
        RECT 51.590 96.260 51.910 96.320 ;
        RECT 19.850 95.920 20.170 96.180 ;
        RECT 22.610 96.120 22.930 96.180 ;
        RECT 24.925 96.120 25.215 96.165 ;
        RECT 22.610 95.980 25.215 96.120 ;
        RECT 22.610 95.920 22.930 95.980 ;
        RECT 24.925 95.935 25.215 95.980 ;
        RECT 35.070 96.120 35.360 96.165 ;
        RECT 37.170 96.120 37.460 96.165 ;
        RECT 38.740 96.120 39.030 96.165 ;
        RECT 35.070 95.980 39.030 96.120 ;
        RECT 35.070 95.935 35.360 95.980 ;
        RECT 37.170 95.935 37.460 95.980 ;
        RECT 38.740 95.935 39.030 95.980 ;
        RECT 45.650 96.120 45.940 96.165 ;
        RECT 47.750 96.120 48.040 96.165 ;
        RECT 49.320 96.120 49.610 96.165 ;
        RECT 45.650 95.980 49.610 96.120 ;
        RECT 45.650 95.935 45.940 95.980 ;
        RECT 47.750 95.935 48.040 95.980 ;
        RECT 49.320 95.935 49.610 95.980 ;
        RECT 50.210 96.120 50.530 96.180 ;
        RECT 52.970 96.120 53.290 96.180 ;
        RECT 57.200 96.120 57.340 96.650 ;
        RECT 57.585 96.615 57.875 96.650 ;
        RECT 58.490 96.600 58.810 96.860 ;
        RECT 59.410 96.600 59.730 96.860 ;
        RECT 60.790 96.600 61.110 96.860 ;
        RECT 61.250 96.600 61.570 96.860 ;
        RECT 62.030 96.800 62.170 96.940 ;
        RECT 63.550 96.800 63.870 96.860 ;
        RECT 72.380 96.845 72.520 97.000 ;
        RECT 73.760 97.000 78.130 97.140 ;
        RECT 62.030 96.660 63.870 96.800 ;
        RECT 63.550 96.600 63.870 96.660 ;
        RECT 64.485 96.800 64.775 96.845 ;
        RECT 66.785 96.800 67.075 96.845 ;
        RECT 71.845 96.800 72.135 96.845 ;
        RECT 64.485 96.660 67.075 96.800 ;
        RECT 64.485 96.615 64.775 96.660 ;
        RECT 66.785 96.615 67.075 96.660 ;
        RECT 71.000 96.660 72.135 96.800 ;
        RECT 65.390 96.260 65.710 96.520 ;
        RECT 69.530 96.260 69.850 96.520 ;
        RECT 50.210 95.980 57.340 96.120 ;
        RECT 71.000 96.120 71.140 96.660 ;
        RECT 71.845 96.615 72.135 96.660 ;
        RECT 72.305 96.615 72.595 96.845 ;
        RECT 72.750 96.600 73.070 96.860 ;
        RECT 73.760 96.845 73.900 97.000 ;
        RECT 74.590 96.940 74.910 97.000 ;
        RECT 77.810 96.940 78.130 97.000 ;
        RECT 73.685 96.615 73.975 96.845 ;
        RECT 75.050 96.800 75.370 96.860 ;
        RECT 75.885 96.800 76.175 96.845 ;
        RECT 75.050 96.660 76.175 96.800 ;
        RECT 75.050 96.600 75.370 96.660 ;
        RECT 75.885 96.615 76.175 96.660 ;
        RECT 71.370 96.460 71.690 96.520 ;
        RECT 74.605 96.460 74.895 96.505 ;
        RECT 71.370 96.320 74.895 96.460 ;
        RECT 71.370 96.260 71.690 96.320 ;
        RECT 74.605 96.275 74.895 96.320 ;
        RECT 75.485 96.460 75.775 96.505 ;
        RECT 76.675 96.460 76.965 96.505 ;
        RECT 79.195 96.460 79.485 96.505 ;
        RECT 75.485 96.320 79.485 96.460 ;
        RECT 75.485 96.275 75.775 96.320 ;
        RECT 76.675 96.275 76.965 96.320 ;
        RECT 79.195 96.275 79.485 96.320 ;
        RECT 75.090 96.120 75.380 96.165 ;
        RECT 77.190 96.120 77.480 96.165 ;
        RECT 78.760 96.120 79.050 96.165 ;
        RECT 71.000 95.980 71.600 96.120 ;
        RECT 50.210 95.920 50.530 95.980 ;
        RECT 52.970 95.920 53.290 95.980 ;
        RECT 11.570 95.780 11.890 95.840 ;
        RECT 13.410 95.780 13.730 95.840 ;
        RECT 11.570 95.640 13.730 95.780 ;
        RECT 11.570 95.580 11.890 95.640 ;
        RECT 13.410 95.580 13.730 95.640 ;
        RECT 15.710 95.780 16.030 95.840 ;
        RECT 16.185 95.780 16.475 95.825 ;
        RECT 15.710 95.640 16.475 95.780 ;
        RECT 15.710 95.580 16.030 95.640 ;
        RECT 16.185 95.595 16.475 95.640 ;
        RECT 21.690 95.780 22.010 95.840 ;
        RECT 23.530 95.780 23.850 95.840 ;
        RECT 21.690 95.640 23.850 95.780 ;
        RECT 21.690 95.580 22.010 95.640 ;
        RECT 23.530 95.580 23.850 95.640 ;
        RECT 29.525 95.780 29.815 95.825 ;
        RECT 32.730 95.780 33.050 95.840 ;
        RECT 29.525 95.640 33.050 95.780 ;
        RECT 29.525 95.595 29.815 95.640 ;
        RECT 32.730 95.580 33.050 95.640 ;
        RECT 33.190 95.780 33.510 95.840 ;
        RECT 40.550 95.780 40.870 95.840 ;
        RECT 33.190 95.640 40.870 95.780 ;
        RECT 33.190 95.580 33.510 95.640 ;
        RECT 40.550 95.580 40.870 95.640 ;
        RECT 43.770 95.580 44.090 95.840 ;
        RECT 44.705 95.780 44.995 95.825 ;
        RECT 46.990 95.780 47.310 95.840 ;
        RECT 44.705 95.640 47.310 95.780 ;
        RECT 44.705 95.595 44.995 95.640 ;
        RECT 46.990 95.580 47.310 95.640 ;
        RECT 49.750 95.780 50.070 95.840 ;
        RECT 52.065 95.780 52.355 95.825 ;
        RECT 49.750 95.640 52.355 95.780 ;
        RECT 49.750 95.580 50.070 95.640 ;
        RECT 52.065 95.595 52.355 95.640 ;
        RECT 62.630 95.580 62.950 95.840 ;
        RECT 71.460 95.780 71.600 95.980 ;
        RECT 75.090 95.980 79.050 96.120 ;
        RECT 75.090 95.935 75.380 95.980 ;
        RECT 77.190 95.935 77.480 95.980 ;
        RECT 78.760 95.935 79.050 95.980 ;
        RECT 75.510 95.780 75.830 95.840 ;
        RECT 71.460 95.640 75.830 95.780 ;
        RECT 75.510 95.580 75.830 95.640 ;
        RECT 79.650 95.780 79.970 95.840 ;
        RECT 81.505 95.780 81.795 95.825 ;
        RECT 79.650 95.640 81.795 95.780 ;
        RECT 79.650 95.580 79.970 95.640 ;
        RECT 81.505 95.595 81.795 95.640 ;
        RECT 5.520 94.960 83.260 95.440 ;
        RECT 44.230 94.760 44.550 94.820 ;
        RECT 44.705 94.760 44.995 94.805 ;
        RECT 30.520 94.620 42.620 94.760 ;
        RECT 30.520 93.785 30.660 94.620 ;
        RECT 37.330 94.420 37.620 94.465 ;
        RECT 38.900 94.420 39.190 94.465 ;
        RECT 41.000 94.420 41.290 94.465 ;
        RECT 37.330 94.280 41.290 94.420 ;
        RECT 37.330 94.235 37.620 94.280 ;
        RECT 38.900 94.235 39.190 94.280 ;
        RECT 41.000 94.235 41.290 94.280 ;
        RECT 36.895 94.080 37.185 94.125 ;
        RECT 39.415 94.080 39.705 94.125 ;
        RECT 40.605 94.080 40.895 94.125 ;
        RECT 36.895 93.940 40.895 94.080 ;
        RECT 36.895 93.895 37.185 93.940 ;
        RECT 39.415 93.895 39.705 93.940 ;
        RECT 40.605 93.895 40.895 93.940 ;
        RECT 42.480 94.080 42.620 94.620 ;
        RECT 44.230 94.620 44.995 94.760 ;
        RECT 44.230 94.560 44.550 94.620 ;
        RECT 44.705 94.575 44.995 94.620 ;
        RECT 45.150 94.760 45.470 94.820 ;
        RECT 50.210 94.760 50.530 94.820 ;
        RECT 45.150 94.620 50.530 94.760 ;
        RECT 45.150 94.560 45.470 94.620 ;
        RECT 50.210 94.560 50.530 94.620 ;
        RECT 50.685 94.760 50.975 94.805 ;
        RECT 51.590 94.760 51.910 94.820 ;
        RECT 50.685 94.620 51.910 94.760 ;
        RECT 50.685 94.575 50.975 94.620 ;
        RECT 51.590 94.560 51.910 94.620 ;
        RECT 53.445 94.760 53.735 94.805 ;
        RECT 58.490 94.760 58.810 94.820 ;
        RECT 53.445 94.620 58.810 94.760 ;
        RECT 53.445 94.575 53.735 94.620 ;
        RECT 58.490 94.560 58.810 94.620 ;
        RECT 59.410 94.560 59.730 94.820 ;
        RECT 63.090 94.760 63.410 94.820 ;
        RECT 59.960 94.620 63.410 94.760 ;
        RECT 42.850 94.420 43.170 94.480 ;
        RECT 43.325 94.420 43.615 94.465 ;
        RECT 48.830 94.420 49.150 94.480 ;
        RECT 42.850 94.280 49.150 94.420 ;
        RECT 42.850 94.220 43.170 94.280 ;
        RECT 43.325 94.235 43.615 94.280 ;
        RECT 48.830 94.220 49.150 94.280 ;
        RECT 49.750 94.220 50.070 94.480 ;
        RECT 52.525 94.235 52.815 94.465 ;
        RECT 55.730 94.420 56.050 94.480 ;
        RECT 53.980 94.280 56.050 94.420 ;
        RECT 46.545 94.080 46.835 94.125 ;
        RECT 42.480 93.940 46.835 94.080 ;
        RECT 42.480 93.800 42.620 93.940 ;
        RECT 46.545 93.895 46.835 93.940 ;
        RECT 48.370 94.080 48.690 94.140 ;
        RECT 52.600 94.080 52.740 94.235 ;
        RECT 48.370 93.940 52.740 94.080 ;
        RECT 48.370 93.880 48.690 93.940 ;
        RECT 29.525 93.555 29.815 93.785 ;
        RECT 30.445 93.555 30.735 93.785 ;
        RECT 31.365 93.555 31.655 93.785 ;
        RECT 34.570 93.740 34.890 93.800 ;
        RECT 41.470 93.740 41.790 93.800 ;
        RECT 34.570 93.600 41.790 93.740 ;
        RECT 29.600 93.400 29.740 93.555 ;
        RECT 31.440 93.400 31.580 93.555 ;
        RECT 34.570 93.540 34.890 93.600 ;
        RECT 41.470 93.540 41.790 93.600 ;
        RECT 42.390 93.540 42.710 93.800 ;
        RECT 43.785 93.740 44.075 93.785 ;
        RECT 47.450 93.740 47.770 93.800 ;
        RECT 43.785 93.600 47.770 93.740 ;
        RECT 43.785 93.555 44.075 93.600 ;
        RECT 47.450 93.540 47.770 93.600 ;
        RECT 47.910 93.540 48.230 93.800 ;
        RECT 52.050 93.740 52.370 93.800 ;
        RECT 53.980 93.740 54.120 94.280 ;
        RECT 55.730 94.220 56.050 94.280 ;
        RECT 54.350 94.080 54.670 94.140 ;
        RECT 56.665 94.080 56.955 94.125 ;
        RECT 54.350 93.940 56.955 94.080 ;
        RECT 54.350 93.880 54.670 93.940 ;
        RECT 56.665 93.895 56.955 93.940 ;
        RECT 52.050 93.600 54.120 93.740 ;
        RECT 52.050 93.540 52.370 93.600 ;
        RECT 54.825 93.555 55.115 93.785 ;
        RECT 55.270 93.740 55.590 93.800 ;
        RECT 55.745 93.740 56.035 93.785 ;
        RECT 55.270 93.600 56.035 93.740 ;
        RECT 29.600 93.260 31.580 93.400 ;
        RECT 29.970 92.860 30.290 93.120 ;
        RECT 31.440 93.060 31.580 93.260 ;
        RECT 34.125 93.400 34.415 93.445 ;
        RECT 35.030 93.400 35.350 93.460 ;
        RECT 40.260 93.400 40.550 93.445 ;
        RECT 41.010 93.400 41.330 93.460 ;
        RECT 45.610 93.445 45.930 93.460 ;
        RECT 34.125 93.260 39.400 93.400 ;
        RECT 34.125 93.215 34.415 93.260 ;
        RECT 35.030 93.200 35.350 93.260 ;
        RECT 39.260 93.120 39.400 93.260 ;
        RECT 40.260 93.260 41.330 93.400 ;
        RECT 40.260 93.215 40.550 93.260 ;
        RECT 41.010 93.200 41.330 93.260 ;
        RECT 45.500 93.400 45.930 93.445 ;
        RECT 46.530 93.400 46.850 93.460 ;
        RECT 45.500 93.260 46.850 93.400 ;
        RECT 45.500 93.215 45.930 93.260 ;
        RECT 45.610 93.200 45.930 93.215 ;
        RECT 46.530 93.200 46.850 93.260 ;
        RECT 49.750 93.400 50.070 93.460 ;
        RECT 51.145 93.400 51.435 93.445 ;
        RECT 49.750 93.260 51.435 93.400 ;
        RECT 49.750 93.200 50.070 93.260 ;
        RECT 51.145 93.215 51.435 93.260 ;
        RECT 52.970 93.400 53.290 93.460 ;
        RECT 54.900 93.400 55.040 93.555 ;
        RECT 55.270 93.540 55.590 93.600 ;
        RECT 55.745 93.555 56.035 93.600 ;
        RECT 56.190 93.540 56.510 93.800 ;
        RECT 57.585 93.555 57.875 93.785 ;
        RECT 58.030 93.740 58.350 93.800 ;
        RECT 59.960 93.785 60.100 94.620 ;
        RECT 63.090 94.560 63.410 94.620 ;
        RECT 70.450 94.760 70.770 94.820 ;
        RECT 71.385 94.760 71.675 94.805 ;
        RECT 70.450 94.620 71.675 94.760 ;
        RECT 70.450 94.560 70.770 94.620 ;
        RECT 71.385 94.575 71.675 94.620 ;
        RECT 74.605 94.760 74.895 94.805 ;
        RECT 75.050 94.760 75.370 94.820 ;
        RECT 76.890 94.760 77.210 94.820 ;
        RECT 74.605 94.620 75.370 94.760 ;
        RECT 74.605 94.575 74.895 94.620 ;
        RECT 75.050 94.560 75.370 94.620 ;
        RECT 75.600 94.620 77.210 94.760 ;
        RECT 61.750 94.420 62.040 94.465 ;
        RECT 63.850 94.420 64.140 94.465 ;
        RECT 65.420 94.420 65.710 94.465 ;
        RECT 61.750 94.280 65.710 94.420 ;
        RECT 61.750 94.235 62.040 94.280 ;
        RECT 63.850 94.235 64.140 94.280 ;
        RECT 65.420 94.235 65.710 94.280 ;
        RECT 68.165 94.420 68.455 94.465 ;
        RECT 69.530 94.420 69.850 94.480 ;
        RECT 68.165 94.280 69.850 94.420 ;
        RECT 68.165 94.235 68.455 94.280 ;
        RECT 69.530 94.220 69.850 94.280 ;
        RECT 62.145 94.080 62.435 94.125 ;
        RECT 63.335 94.080 63.625 94.125 ;
        RECT 65.855 94.080 66.145 94.125 ;
        RECT 75.600 94.080 75.740 94.620 ;
        RECT 76.890 94.560 77.210 94.620 ;
        RECT 75.970 94.420 76.290 94.480 ;
        RECT 75.970 94.280 79.420 94.420 ;
        RECT 75.970 94.220 76.290 94.280 ;
        RECT 77.350 94.080 77.670 94.140 ;
        RECT 62.145 93.940 66.145 94.080 ;
        RECT 62.145 93.895 62.435 93.940 ;
        RECT 63.335 93.895 63.625 93.940 ;
        RECT 65.855 93.895 66.145 93.940 ;
        RECT 72.380 93.940 75.740 94.080 ;
        RECT 76.520 93.940 77.670 94.080 ;
        RECT 58.965 93.740 59.255 93.785 ;
        RECT 58.030 93.600 59.255 93.740 ;
        RECT 57.110 93.400 57.430 93.460 ;
        RECT 52.970 93.260 57.430 93.400 ;
        RECT 52.970 93.200 53.290 93.260 ;
        RECT 57.110 93.200 57.430 93.260 ;
        RECT 34.585 93.060 34.875 93.105 ;
        RECT 35.490 93.060 35.810 93.120 ;
        RECT 31.440 92.920 35.810 93.060 ;
        RECT 34.585 92.875 34.875 92.920 ;
        RECT 35.490 92.860 35.810 92.920 ;
        RECT 39.170 92.860 39.490 93.120 ;
        RECT 41.470 93.060 41.790 93.120 ;
        RECT 43.310 93.060 43.630 93.120 ;
        RECT 46.085 93.060 46.375 93.105 ;
        RECT 41.470 92.920 46.375 93.060 ;
        RECT 41.470 92.860 41.790 92.920 ;
        RECT 43.310 92.860 43.630 92.920 ;
        RECT 46.085 92.875 46.375 92.920 ;
        RECT 48.830 93.060 49.150 93.120 ;
        RECT 53.430 93.060 53.750 93.120 ;
        RECT 54.350 93.060 54.670 93.120 ;
        RECT 57.660 93.060 57.800 93.555 ;
        RECT 58.030 93.540 58.350 93.600 ;
        RECT 58.965 93.555 59.255 93.600 ;
        RECT 59.885 93.555 60.175 93.785 ;
        RECT 61.250 93.540 61.570 93.800 ;
        RECT 62.630 93.785 62.950 93.800 ;
        RECT 62.600 93.740 62.950 93.785 ;
        RECT 62.435 93.600 62.950 93.740 ;
        RECT 62.600 93.555 62.950 93.600 ;
        RECT 62.630 93.540 62.950 93.555 ;
        RECT 69.530 93.540 69.850 93.800 ;
        RECT 72.380 93.785 72.520 93.940 ;
        RECT 72.305 93.555 72.595 93.785 ;
        RECT 72.765 93.740 73.055 93.785 ;
        RECT 73.210 93.740 73.530 93.800 ;
        RECT 72.765 93.600 73.530 93.740 ;
        RECT 72.765 93.555 73.055 93.600 ;
        RECT 73.210 93.540 73.530 93.600 ;
        RECT 73.670 93.540 73.990 93.800 ;
        RECT 74.145 93.555 74.435 93.785 ;
        RECT 75.510 93.740 75.830 93.800 ;
        RECT 76.520 93.785 76.660 93.940 ;
        RECT 77.350 93.880 77.670 93.940 ;
        RECT 75.985 93.740 76.275 93.785 ;
        RECT 75.510 93.600 76.275 93.740 ;
        RECT 74.220 93.400 74.360 93.555 ;
        RECT 75.510 93.540 75.830 93.600 ;
        RECT 75.985 93.555 76.275 93.600 ;
        RECT 76.445 93.555 76.735 93.785 ;
        RECT 76.890 93.540 77.210 93.800 ;
        RECT 77.810 93.540 78.130 93.800 ;
        RECT 79.280 93.785 79.420 94.280 ;
        RECT 79.205 93.740 79.495 93.785 ;
        RECT 80.570 93.740 80.890 93.800 ;
        RECT 79.205 93.600 80.890 93.740 ;
        RECT 79.205 93.555 79.495 93.600 ;
        RECT 80.570 93.540 80.890 93.600 ;
        RECT 81.045 93.740 81.335 93.785 ;
        RECT 81.490 93.740 81.810 93.800 ;
        RECT 81.045 93.600 81.810 93.740 ;
        RECT 81.045 93.555 81.335 93.600 ;
        RECT 81.490 93.540 81.810 93.600 ;
        RECT 78.730 93.400 79.050 93.460 ;
        RECT 79.650 93.400 79.970 93.460 ;
        RECT 74.220 93.260 78.500 93.400 ;
        RECT 48.830 92.920 57.800 93.060 ;
        RECT 48.830 92.860 49.150 92.920 ;
        RECT 53.430 92.860 53.750 92.920 ;
        RECT 54.350 92.860 54.670 92.920 ;
        RECT 58.490 92.860 58.810 93.120 ;
        RECT 66.310 93.060 66.630 93.120 ;
        RECT 78.360 93.105 78.500 93.260 ;
        RECT 78.730 93.260 79.970 93.400 ;
        RECT 78.730 93.200 79.050 93.260 ;
        RECT 79.650 93.200 79.970 93.260 ;
        RECT 80.110 93.200 80.430 93.460 ;
        RECT 68.625 93.060 68.915 93.105 ;
        RECT 66.310 92.920 68.915 93.060 ;
        RECT 66.310 92.860 66.630 92.920 ;
        RECT 68.625 92.875 68.915 92.920 ;
        RECT 78.285 92.875 78.575 93.105 ;
        RECT 5.520 92.240 83.260 92.720 ;
        RECT 19.850 92.040 20.170 92.100 ;
        RECT 32.745 92.040 33.035 92.085 ;
        RECT 39.630 92.040 39.950 92.100 ;
        RECT 19.850 91.900 26.060 92.040 ;
        RECT 19.850 91.840 20.170 91.900 ;
        RECT 16.170 91.700 16.490 91.760 ;
        RECT 18.930 91.700 19.250 91.760 ;
        RECT 19.405 91.700 19.695 91.745 ;
        RECT 16.170 91.560 19.695 91.700 ;
        RECT 16.170 91.500 16.490 91.560 ;
        RECT 18.930 91.500 19.250 91.560 ;
        RECT 19.405 91.515 19.695 91.560 ;
        RECT 20.770 91.700 21.090 91.760 ;
        RECT 20.770 91.560 24.220 91.700 ;
        RECT 20.770 91.500 21.090 91.560 ;
        RECT 11.585 91.360 11.875 91.405 ;
        RECT 12.030 91.360 12.350 91.420 ;
        RECT 11.585 91.220 12.350 91.360 ;
        RECT 11.585 91.175 11.875 91.220 ;
        RECT 12.030 91.160 12.350 91.220 ;
        RECT 12.505 91.360 12.795 91.405 ;
        RECT 15.250 91.360 15.570 91.420 ;
        RECT 24.080 91.405 24.220 91.560 ;
        RECT 25.920 91.420 26.060 91.900 ;
        RECT 32.745 91.900 39.950 92.040 ;
        RECT 32.745 91.855 33.035 91.900 ;
        RECT 39.630 91.840 39.950 91.900 ;
        RECT 42.390 92.040 42.710 92.100 ;
        RECT 45.610 92.040 45.930 92.100 ;
        RECT 42.390 91.900 49.060 92.040 ;
        RECT 42.390 91.840 42.710 91.900 ;
        RECT 45.610 91.840 45.930 91.900 ;
        RECT 35.030 91.700 35.350 91.760 ;
        RECT 36.870 91.745 37.190 91.760 ;
        RECT 34.200 91.560 35.350 91.700 ;
        RECT 12.505 91.220 15.570 91.360 ;
        RECT 12.505 91.175 12.795 91.220 ;
        RECT 15.250 91.160 15.570 91.220 ;
        RECT 24.005 91.360 24.295 91.405 ;
        RECT 24.910 91.360 25.230 91.420 ;
        RECT 24.005 91.220 25.230 91.360 ;
        RECT 24.005 91.175 24.295 91.220 ;
        RECT 24.910 91.160 25.230 91.220 ;
        RECT 25.830 91.360 26.150 91.420 ;
        RECT 27.685 91.360 27.975 91.405 ;
        RECT 25.830 91.220 27.975 91.360 ;
        RECT 25.830 91.160 26.150 91.220 ;
        RECT 27.685 91.175 27.975 91.220 ;
        RECT 29.970 91.360 30.290 91.420 ;
        RECT 31.825 91.360 32.115 91.405 ;
        RECT 29.970 91.220 32.115 91.360 ;
        RECT 29.970 91.160 30.290 91.220 ;
        RECT 31.825 91.175 32.115 91.220 ;
        RECT 32.745 91.360 33.035 91.405 ;
        RECT 33.190 91.360 33.510 91.420 ;
        RECT 34.200 91.405 34.340 91.560 ;
        RECT 35.030 91.500 35.350 91.560 ;
        RECT 36.840 91.515 37.190 91.745 ;
        RECT 36.870 91.500 37.190 91.515 ;
        RECT 41.930 91.700 42.250 91.760 ;
        RECT 42.865 91.700 43.155 91.745 ;
        RECT 47.910 91.700 48.230 91.760 ;
        RECT 48.920 91.745 49.060 91.900 ;
        RECT 50.670 91.840 50.990 92.100 ;
        RECT 52.510 92.040 52.830 92.100 ;
        RECT 54.825 92.040 55.115 92.085 ;
        RECT 52.510 91.900 55.115 92.040 ;
        RECT 52.510 91.840 52.830 91.900 ;
        RECT 54.825 91.855 55.115 91.900 ;
        RECT 56.665 92.040 56.955 92.085 ;
        RECT 69.530 92.040 69.850 92.100 ;
        RECT 56.665 91.900 69.850 92.040 ;
        RECT 56.665 91.855 56.955 91.900 ;
        RECT 69.530 91.840 69.850 91.900 ;
        RECT 70.910 91.840 71.230 92.100 ;
        RECT 76.890 92.040 77.210 92.100 ;
        RECT 81.505 92.040 81.795 92.085 ;
        RECT 76.890 91.900 81.795 92.040 ;
        RECT 76.890 91.840 77.210 91.900 ;
        RECT 81.505 91.855 81.795 91.900 ;
        RECT 41.930 91.560 48.230 91.700 ;
        RECT 41.930 91.500 42.250 91.560 ;
        RECT 42.865 91.515 43.155 91.560 ;
        RECT 47.910 91.500 48.230 91.560 ;
        RECT 48.845 91.515 49.135 91.745 ;
        RECT 49.925 91.700 50.215 91.745 ;
        RECT 51.590 91.700 51.910 91.760 ;
        RECT 61.250 91.700 61.570 91.760 ;
        RECT 78.730 91.700 79.050 91.760 ;
        RECT 80.585 91.700 80.875 91.745 ;
        RECT 49.925 91.560 54.580 91.700 ;
        RECT 49.925 91.515 50.215 91.560 ;
        RECT 51.590 91.500 51.910 91.560 ;
        RECT 32.745 91.220 33.510 91.360 ;
        RECT 32.745 91.175 33.035 91.220 ;
        RECT 23.085 91.020 23.375 91.065 ;
        RECT 28.145 91.020 28.435 91.065 ;
        RECT 23.085 90.880 28.435 91.020 ;
        RECT 31.900 91.020 32.040 91.175 ;
        RECT 33.190 91.160 33.510 91.220 ;
        RECT 34.125 91.175 34.415 91.405 ;
        RECT 34.570 91.360 34.890 91.420 ;
        RECT 35.505 91.360 35.795 91.405 ;
        RECT 38.710 91.360 39.030 91.420 ;
        RECT 34.570 91.220 35.795 91.360 ;
        RECT 34.570 91.160 34.890 91.220 ;
        RECT 35.505 91.175 35.795 91.220 ;
        RECT 36.040 91.350 37.100 91.360 ;
        RECT 37.420 91.350 44.460 91.360 ;
        RECT 36.040 91.220 44.460 91.350 ;
        RECT 36.040 91.020 36.180 91.220 ;
        RECT 36.960 91.210 37.560 91.220 ;
        RECT 38.710 91.160 39.030 91.220 ;
        RECT 31.900 90.880 36.180 91.020 ;
        RECT 36.385 91.020 36.675 91.065 ;
        RECT 37.575 91.020 37.865 91.065 ;
        RECT 40.095 91.020 40.385 91.065 ;
        RECT 36.385 90.880 40.385 91.020 ;
        RECT 23.085 90.835 23.375 90.880 ;
        RECT 28.145 90.835 28.435 90.880 ;
        RECT 36.385 90.835 36.675 90.880 ;
        RECT 37.575 90.835 37.865 90.880 ;
        RECT 40.095 90.835 40.385 90.880 ;
        RECT 35.990 90.680 36.280 90.725 ;
        RECT 38.090 90.680 38.380 90.725 ;
        RECT 39.660 90.680 39.950 90.725 ;
        RECT 43.770 90.680 44.090 90.740 ;
        RECT 44.320 90.725 44.460 91.220 ;
        RECT 47.005 91.175 47.295 91.405 ;
        RECT 47.465 91.360 47.755 91.405 ;
        RECT 48.370 91.360 48.690 91.420 ;
        RECT 47.465 91.220 48.690 91.360 ;
        RECT 47.465 91.175 47.755 91.220 ;
        RECT 47.080 91.020 47.220 91.175 ;
        RECT 48.370 91.160 48.690 91.220 ;
        RECT 49.290 91.160 49.610 91.420 ;
        RECT 51.145 91.360 51.435 91.405 ;
        RECT 49.840 91.220 51.435 91.360 ;
        RECT 49.380 91.020 49.520 91.160 ;
        RECT 47.080 90.880 49.520 91.020 ;
        RECT 35.990 90.540 39.950 90.680 ;
        RECT 35.990 90.495 36.280 90.540 ;
        RECT 38.090 90.495 38.380 90.540 ;
        RECT 39.660 90.495 39.950 90.540 ;
        RECT 42.020 90.540 44.090 90.680 ;
        RECT 10.650 90.340 10.970 90.400 ;
        RECT 11.585 90.340 11.875 90.385 ;
        RECT 10.650 90.200 11.875 90.340 ;
        RECT 10.650 90.140 10.970 90.200 ;
        RECT 11.585 90.155 11.875 90.200 ;
        RECT 33.665 90.340 33.955 90.385 ;
        RECT 42.020 90.340 42.160 90.540 ;
        RECT 43.770 90.480 44.090 90.540 ;
        RECT 44.245 90.495 44.535 90.725 ;
        RECT 45.165 90.680 45.455 90.725 ;
        RECT 49.290 90.680 49.610 90.740 ;
        RECT 45.165 90.540 49.610 90.680 ;
        RECT 45.165 90.495 45.455 90.540 ;
        RECT 49.290 90.480 49.610 90.540 ;
        RECT 33.665 90.200 42.160 90.340 ;
        RECT 33.665 90.155 33.955 90.200 ;
        RECT 46.990 90.140 47.310 90.400 ;
        RECT 47.910 90.340 48.230 90.400 ;
        RECT 49.840 90.385 49.980 91.220 ;
        RECT 51.145 91.175 51.435 91.220 ;
        RECT 52.065 91.175 52.355 91.405 ;
        RECT 52.140 91.020 52.280 91.175 ;
        RECT 52.970 91.160 53.290 91.420 ;
        RECT 54.440 91.405 54.580 91.560 ;
        RECT 59.500 91.560 62.170 91.700 ;
        RECT 54.365 91.175 54.655 91.405 ;
        RECT 55.745 91.360 56.035 91.405 ;
        RECT 57.570 91.360 57.890 91.420 ;
        RECT 59.500 91.405 59.640 91.560 ;
        RECT 61.250 91.500 61.570 91.560 ;
        RECT 60.790 91.405 61.110 91.420 ;
        RECT 55.745 91.220 57.890 91.360 ;
        RECT 55.745 91.175 56.035 91.220 ;
        RECT 57.570 91.160 57.890 91.220 ;
        RECT 59.425 91.175 59.715 91.405 ;
        RECT 60.760 91.175 61.110 91.405 ;
        RECT 62.030 91.360 62.170 91.560 ;
        RECT 71.920 91.560 80.875 91.700 ;
        RECT 71.370 91.360 71.690 91.420 ;
        RECT 71.920 91.405 72.060 91.560 ;
        RECT 78.730 91.500 79.050 91.560 ;
        RECT 80.585 91.515 80.875 91.560 ;
        RECT 62.030 91.220 71.690 91.360 ;
        RECT 60.790 91.160 61.110 91.175 ;
        RECT 71.370 91.160 71.690 91.220 ;
        RECT 71.845 91.175 72.135 91.405 ;
        RECT 72.750 91.360 73.070 91.420 ;
        RECT 73.585 91.360 73.875 91.405 ;
        RECT 72.750 91.220 73.875 91.360 ;
        RECT 72.750 91.160 73.070 91.220 ;
        RECT 73.585 91.175 73.875 91.220 ;
        RECT 78.270 91.360 78.590 91.420 ;
        RECT 79.190 91.360 79.510 91.420 ;
        RECT 79.665 91.360 79.955 91.405 ;
        RECT 78.270 91.220 79.955 91.360 ;
        RECT 78.270 91.160 78.590 91.220 ;
        RECT 79.190 91.160 79.510 91.220 ;
        RECT 79.665 91.175 79.955 91.220 ;
        RECT 53.430 91.020 53.750 91.080 ;
        RECT 52.140 90.880 53.750 91.020 ;
        RECT 53.430 90.820 53.750 90.880 ;
        RECT 60.305 91.020 60.595 91.065 ;
        RECT 61.495 91.020 61.785 91.065 ;
        RECT 64.015 91.020 64.305 91.065 ;
        RECT 60.305 90.880 64.305 91.020 ;
        RECT 60.305 90.835 60.595 90.880 ;
        RECT 61.495 90.835 61.785 90.880 ;
        RECT 64.015 90.835 64.305 90.880 ;
        RECT 69.545 90.835 69.835 91.065 ;
        RECT 71.460 91.020 71.600 91.160 ;
        RECT 72.305 91.020 72.595 91.065 ;
        RECT 71.460 90.880 72.595 91.020 ;
        RECT 72.305 90.835 72.595 90.880 ;
        RECT 73.185 91.020 73.475 91.065 ;
        RECT 74.375 91.020 74.665 91.065 ;
        RECT 76.895 91.020 77.185 91.065 ;
        RECT 73.185 90.880 77.185 91.020 ;
        RECT 73.185 90.835 73.475 90.880 ;
        RECT 74.375 90.835 74.665 90.880 ;
        RECT 76.895 90.835 77.185 90.880 ;
        RECT 59.910 90.680 60.200 90.725 ;
        RECT 62.010 90.680 62.300 90.725 ;
        RECT 63.580 90.680 63.870 90.725 ;
        RECT 59.910 90.540 63.870 90.680 ;
        RECT 59.910 90.495 60.200 90.540 ;
        RECT 62.010 90.495 62.300 90.540 ;
        RECT 63.580 90.495 63.870 90.540 ;
        RECT 66.325 90.680 66.615 90.725 ;
        RECT 69.620 90.680 69.760 90.835 ;
        RECT 70.450 90.680 70.770 90.740 ;
        RECT 66.325 90.540 70.770 90.680 ;
        RECT 66.325 90.495 66.615 90.540 ;
        RECT 70.450 90.480 70.770 90.540 ;
        RECT 72.790 90.680 73.080 90.725 ;
        RECT 74.890 90.680 75.180 90.725 ;
        RECT 76.460 90.680 76.750 90.725 ;
        RECT 72.790 90.540 76.750 90.680 ;
        RECT 72.790 90.495 73.080 90.540 ;
        RECT 74.890 90.495 75.180 90.540 ;
        RECT 76.460 90.495 76.750 90.540 ;
        RECT 49.765 90.340 50.055 90.385 ;
        RECT 47.910 90.200 50.055 90.340 ;
        RECT 47.910 90.140 48.230 90.200 ;
        RECT 49.765 90.155 50.055 90.200 ;
        RECT 52.970 90.340 53.290 90.400 ;
        RECT 54.810 90.340 55.130 90.400 ;
        RECT 52.970 90.200 55.130 90.340 ;
        RECT 52.970 90.140 53.290 90.200 ;
        RECT 54.810 90.140 55.130 90.200 ;
        RECT 66.770 90.140 67.090 90.400 ;
        RECT 76.890 90.340 77.210 90.400 ;
        RECT 79.205 90.340 79.495 90.385 ;
        RECT 76.890 90.200 79.495 90.340 ;
        RECT 76.890 90.140 77.210 90.200 ;
        RECT 79.205 90.155 79.495 90.200 ;
        RECT 5.520 89.520 83.260 90.000 ;
        RECT 7.905 89.320 8.195 89.365 ;
        RECT 9.730 89.320 10.050 89.380 ;
        RECT 7.905 89.180 10.050 89.320 ;
        RECT 7.905 89.135 8.195 89.180 ;
        RECT 9.730 89.120 10.050 89.180 ;
        RECT 10.205 89.320 10.495 89.365 ;
        RECT 14.330 89.320 14.650 89.380 ;
        RECT 10.205 89.180 14.650 89.320 ;
        RECT 10.205 89.135 10.495 89.180 ;
        RECT 14.330 89.120 14.650 89.180 ;
        RECT 16.630 89.320 16.950 89.380 ;
        RECT 17.565 89.320 17.855 89.365 ;
        RECT 16.630 89.180 17.855 89.320 ;
        RECT 16.630 89.120 16.950 89.180 ;
        RECT 17.565 89.135 17.855 89.180 ;
        RECT 22.625 89.320 22.915 89.365 ;
        RECT 23.070 89.320 23.390 89.380 ;
        RECT 22.625 89.180 23.390 89.320 ;
        RECT 22.625 89.135 22.915 89.180 ;
        RECT 23.070 89.120 23.390 89.180 ;
        RECT 26.750 89.120 27.070 89.380 ;
        RECT 36.425 89.320 36.715 89.365 ;
        RECT 36.870 89.320 37.190 89.380 ;
        RECT 36.425 89.180 37.190 89.320 ;
        RECT 36.425 89.135 36.715 89.180 ;
        RECT 36.870 89.120 37.190 89.180 ;
        RECT 37.790 89.120 38.110 89.380 ;
        RECT 51.130 89.120 51.450 89.380 ;
        RECT 60.790 89.320 61.110 89.380 ;
        RECT 61.265 89.320 61.555 89.365 ;
        RECT 60.790 89.180 61.555 89.320 ;
        RECT 60.790 89.120 61.110 89.180 ;
        RECT 61.265 89.135 61.555 89.180 ;
        RECT 61.710 89.320 62.030 89.380 ;
        RECT 71.845 89.320 72.135 89.365 ;
        RECT 72.750 89.320 73.070 89.380 ;
        RECT 75.510 89.320 75.830 89.380 ;
        RECT 61.710 89.180 68.380 89.320 ;
        RECT 61.710 89.120 62.030 89.180 ;
        RECT 13.885 88.980 14.175 89.025 ;
        RECT 14.790 88.980 15.110 89.040 ;
        RECT 18.930 88.980 19.250 89.040 ;
        RECT 13.885 88.840 19.250 88.980 ;
        RECT 13.885 88.795 14.175 88.840 ;
        RECT 14.790 88.780 15.110 88.840 ;
        RECT 18.930 88.780 19.250 88.840 ;
        RECT 42.865 88.980 43.155 89.025 ;
        RECT 43.770 88.980 44.090 89.040 ;
        RECT 42.865 88.840 44.090 88.980 ;
        RECT 68.240 88.980 68.380 89.180 ;
        RECT 71.845 89.180 73.070 89.320 ;
        RECT 71.845 89.135 72.135 89.180 ;
        RECT 72.750 89.120 73.070 89.180 ;
        RECT 73.300 89.180 75.830 89.320 ;
        RECT 68.240 88.840 68.840 88.980 ;
        RECT 42.865 88.795 43.155 88.840 ;
        RECT 43.770 88.780 44.090 88.840 ;
        RECT 0.530 88.640 0.850 88.700 ;
        RECT 58.490 88.640 58.810 88.700 ;
        RECT 64.025 88.640 64.315 88.685 ;
        RECT 0.530 88.500 44.920 88.640 ;
        RECT 0.530 88.440 0.850 88.500 ;
        RECT 12.030 88.100 12.350 88.360 ;
        RECT 12.965 88.310 13.255 88.345 ;
        RECT 12.680 88.170 13.255 88.310 ;
        RECT 8.810 87.760 9.130 88.020 ;
        RECT 11.125 87.960 11.415 88.005 ;
        RECT 11.570 87.960 11.890 88.020 ;
        RECT 11.125 87.820 11.890 87.960 ;
        RECT 12.680 87.960 12.820 88.170 ;
        RECT 12.965 88.115 13.255 88.170 ;
        RECT 13.410 88.100 13.730 88.360 ;
        RECT 15.250 88.300 15.570 88.360 ;
        RECT 15.740 88.300 16.030 88.345 ;
        RECT 15.250 88.160 16.030 88.300 ;
        RECT 15.250 88.100 15.570 88.160 ;
        RECT 15.740 88.115 16.030 88.160 ;
        RECT 16.630 88.100 16.950 88.360 ;
        RECT 17.090 88.100 17.410 88.360 ;
        RECT 18.025 88.115 18.315 88.345 ;
        RECT 16.720 87.960 16.860 88.100 ;
        RECT 12.680 87.820 16.860 87.960 ;
        RECT 17.550 87.960 17.870 88.020 ;
        RECT 18.100 87.960 18.240 88.115 ;
        RECT 18.930 88.100 19.250 88.360 ;
        RECT 19.390 88.100 19.710 88.360 ;
        RECT 23.545 88.300 23.835 88.345 ;
        RECT 24.910 88.300 25.230 88.360 ;
        RECT 23.545 88.160 25.230 88.300 ;
        RECT 23.545 88.115 23.835 88.160 ;
        RECT 24.910 88.100 25.230 88.160 ;
        RECT 25.830 88.100 26.150 88.360 ;
        RECT 26.310 88.115 26.600 88.345 ;
        RECT 36.425 88.115 36.715 88.345 ;
        RECT 37.345 88.300 37.635 88.345 ;
        RECT 38.725 88.300 39.015 88.345 ;
        RECT 37.345 88.160 39.015 88.300 ;
        RECT 37.345 88.115 37.635 88.160 ;
        RECT 38.725 88.115 39.015 88.160 ;
        RECT 20.310 87.960 20.630 88.020 ;
        RECT 17.550 87.820 20.630 87.960 ;
        RECT 11.125 87.775 11.415 87.820 ;
        RECT 11.570 87.760 11.890 87.820 ;
        RECT 17.550 87.760 17.870 87.820 ;
        RECT 20.310 87.760 20.630 87.820 ;
        RECT 24.465 87.775 24.755 88.005 ;
        RECT 25.000 87.960 25.140 88.100 ;
        RECT 26.380 87.960 26.520 88.115 ;
        RECT 25.000 87.820 26.520 87.960 ;
        RECT 6.970 87.420 7.290 87.680 ;
        RECT 7.890 87.665 8.210 87.680 ;
        RECT 7.825 87.435 8.210 87.665 ;
        RECT 7.890 87.420 8.210 87.435 ;
        RECT 9.270 87.420 9.590 87.680 ;
        RECT 10.125 87.620 10.415 87.665 ;
        RECT 12.030 87.620 12.350 87.680 ;
        RECT 10.125 87.480 12.350 87.620 ;
        RECT 10.125 87.435 10.415 87.480 ;
        RECT 12.030 87.420 12.350 87.480 ;
        RECT 12.490 87.420 12.810 87.680 ;
        RECT 15.710 87.420 16.030 87.680 ;
        RECT 16.645 87.620 16.935 87.665 ;
        RECT 17.090 87.620 17.410 87.680 ;
        RECT 16.645 87.480 17.410 87.620 ;
        RECT 24.540 87.620 24.680 87.775 ;
        RECT 25.830 87.620 26.150 87.680 ;
        RECT 30.430 87.620 30.750 87.680 ;
        RECT 24.540 87.480 30.750 87.620 ;
        RECT 36.500 87.620 36.640 88.115 ;
        RECT 38.800 87.960 38.940 88.115 ;
        RECT 39.170 88.100 39.490 88.360 ;
        RECT 39.630 88.100 39.950 88.360 ;
        RECT 40.565 88.300 40.855 88.345 ;
        RECT 41.470 88.300 41.790 88.360 ;
        RECT 40.565 88.160 41.790 88.300 ;
        RECT 40.565 88.115 40.855 88.160 ;
        RECT 41.470 88.100 41.790 88.160 ;
        RECT 41.930 88.100 42.250 88.360 ;
        RECT 43.310 88.100 43.630 88.360 ;
        RECT 44.780 88.345 44.920 88.500 ;
        RECT 58.490 88.500 64.315 88.640 ;
        RECT 58.490 88.440 58.810 88.500 ;
        RECT 64.025 88.455 64.315 88.500 ;
        RECT 44.705 88.115 44.995 88.345 ;
        RECT 63.105 88.300 63.395 88.345 ;
        RECT 66.770 88.300 67.090 88.360 ;
        RECT 63.105 88.160 67.090 88.300 ;
        RECT 63.105 88.115 63.395 88.160 ;
        RECT 66.770 88.100 67.090 88.160 ;
        RECT 67.705 88.115 67.995 88.345 ;
        RECT 44.230 87.960 44.550 88.020 ;
        RECT 38.800 87.820 44.550 87.960 ;
        RECT 44.230 87.760 44.550 87.820 ;
        RECT 64.470 87.960 64.790 88.020 ;
        RECT 67.780 87.960 67.920 88.115 ;
        RECT 68.150 88.100 68.470 88.360 ;
        RECT 68.700 88.345 68.840 88.840 ;
        RECT 68.625 88.115 68.915 88.345 ;
        RECT 69.530 88.100 69.850 88.360 ;
        RECT 70.450 88.100 70.770 88.360 ;
        RECT 71.370 88.300 71.690 88.360 ;
        RECT 73.300 88.345 73.440 89.180 ;
        RECT 75.510 89.120 75.830 89.180 ;
        RECT 74.130 88.980 74.450 89.040 ;
        RECT 73.760 88.840 74.450 88.980 ;
        RECT 73.760 88.345 73.900 88.840 ;
        RECT 74.130 88.780 74.450 88.840 ;
        RECT 75.525 88.640 75.815 88.685 ;
        RECT 77.810 88.640 78.130 88.700 ;
        RECT 81.030 88.640 81.350 88.700 ;
        RECT 74.220 88.500 75.815 88.640 ;
        RECT 74.220 88.345 74.360 88.500 ;
        RECT 75.525 88.455 75.815 88.500 ;
        RECT 77.440 88.500 81.350 88.640 ;
        RECT 73.225 88.300 73.515 88.345 ;
        RECT 71.370 88.160 73.515 88.300 ;
        RECT 71.370 88.100 71.690 88.160 ;
        RECT 73.225 88.115 73.515 88.160 ;
        RECT 73.685 88.115 73.975 88.345 ;
        RECT 74.145 88.115 74.435 88.345 ;
        RECT 74.590 88.300 74.910 88.360 ;
        RECT 77.440 88.345 77.580 88.500 ;
        RECT 77.810 88.440 78.130 88.500 ;
        RECT 81.030 88.440 81.350 88.500 ;
        RECT 75.065 88.300 75.355 88.345 ;
        RECT 74.590 88.160 75.355 88.300 ;
        RECT 74.590 88.100 74.910 88.160 ;
        RECT 75.065 88.115 75.355 88.160 ;
        RECT 77.365 88.115 77.655 88.345 ;
        RECT 81.490 88.100 81.810 88.360 ;
        RECT 64.470 87.820 67.920 87.960 ;
        RECT 64.470 87.760 64.790 87.820 ;
        RECT 76.430 87.760 76.750 88.020 ;
        RECT 77.825 87.960 78.115 88.005 ;
        RECT 78.270 87.960 78.590 88.020 ;
        RECT 77.825 87.820 78.590 87.960 ;
        RECT 77.825 87.775 78.115 87.820 ;
        RECT 78.270 87.760 78.590 87.820 ;
        RECT 78.745 87.960 79.035 88.005 ;
        RECT 79.190 87.960 79.510 88.020 ;
        RECT 78.745 87.820 79.510 87.960 ;
        RECT 78.745 87.775 79.035 87.820 ;
        RECT 79.190 87.760 79.510 87.820 ;
        RECT 41.025 87.620 41.315 87.665 ;
        RECT 36.500 87.480 41.315 87.620 ;
        RECT 16.645 87.435 16.935 87.480 ;
        RECT 17.090 87.420 17.410 87.480 ;
        RECT 25.830 87.420 26.150 87.480 ;
        RECT 30.430 87.420 30.750 87.480 ;
        RECT 41.025 87.435 41.315 87.480 ;
        RECT 63.565 87.620 63.855 87.665 ;
        RECT 66.785 87.620 67.075 87.665 ;
        RECT 63.565 87.480 67.075 87.620 ;
        RECT 63.565 87.435 63.855 87.480 ;
        RECT 66.785 87.435 67.075 87.480 ;
        RECT 71.385 87.620 71.675 87.665 ;
        RECT 75.050 87.620 75.370 87.680 ;
        RECT 71.385 87.480 75.370 87.620 ;
        RECT 71.385 87.435 71.675 87.480 ;
        RECT 75.050 87.420 75.370 87.480 ;
        RECT 79.665 87.620 79.955 87.665 ;
        RECT 80.110 87.620 80.430 87.680 ;
        RECT 79.665 87.480 80.430 87.620 ;
        RECT 79.665 87.435 79.955 87.480 ;
        RECT 80.110 87.420 80.430 87.480 ;
        RECT 80.585 87.620 80.875 87.665 ;
        RECT 81.490 87.620 81.810 87.680 ;
        RECT 80.585 87.480 81.810 87.620 ;
        RECT 80.585 87.435 80.875 87.480 ;
        RECT 81.490 87.420 81.810 87.480 ;
        RECT 5.520 86.800 83.260 87.280 ;
        RECT 14.790 86.400 15.110 86.660 ;
        RECT 41.930 86.600 42.250 86.660 ;
        RECT 44.690 86.600 45.010 86.660 ;
        RECT 45.165 86.600 45.455 86.645 ;
        RECT 41.930 86.460 45.455 86.600 ;
        RECT 41.930 86.400 42.250 86.460 ;
        RECT 25.370 86.260 25.690 86.320 ;
        RECT 26.750 86.305 27.070 86.320 ;
        RECT 7.980 86.120 13.870 86.260 ;
        RECT 6.970 85.920 7.290 85.980 ;
        RECT 7.980 85.965 8.120 86.120 ;
        RECT 9.270 85.965 9.590 85.980 ;
        RECT 7.905 85.920 8.195 85.965 ;
        RECT 9.240 85.920 9.590 85.965 ;
        RECT 6.970 85.780 8.195 85.920 ;
        RECT 9.075 85.780 9.590 85.920 ;
        RECT 6.970 85.720 7.290 85.780 ;
        RECT 7.905 85.735 8.195 85.780 ;
        RECT 9.240 85.735 9.590 85.780 ;
        RECT 9.270 85.720 9.590 85.735 ;
        RECT 8.785 85.580 9.075 85.625 ;
        RECT 9.975 85.580 10.265 85.625 ;
        RECT 12.495 85.580 12.785 85.625 ;
        RECT 8.785 85.440 12.785 85.580 ;
        RECT 13.730 85.580 13.870 86.120 ;
        RECT 16.260 86.120 25.690 86.260 ;
        RECT 15.710 85.720 16.030 85.980 ;
        RECT 16.260 85.580 16.400 86.120 ;
        RECT 17.180 85.965 17.320 86.120 ;
        RECT 25.370 86.060 25.690 86.120 ;
        RECT 25.845 86.075 26.135 86.305 ;
        RECT 26.750 86.075 27.135 86.305 ;
        RECT 28.605 86.260 28.895 86.305 ;
        RECT 31.350 86.260 31.670 86.320 ;
        RECT 28.605 86.120 31.670 86.260 ;
        RECT 28.605 86.075 28.895 86.120 ;
        RECT 16.645 85.735 16.935 85.965 ;
        RECT 17.105 85.735 17.395 85.965 ;
        RECT 13.730 85.440 16.400 85.580 ;
        RECT 16.720 85.580 16.860 85.735 ;
        RECT 17.550 85.720 17.870 85.980 ;
        RECT 18.470 85.965 18.790 85.980 ;
        RECT 18.440 85.735 18.790 85.965 ;
        RECT 18.470 85.720 18.790 85.735 ;
        RECT 17.640 85.580 17.780 85.720 ;
        RECT 16.720 85.440 17.780 85.580 ;
        RECT 17.985 85.580 18.275 85.625 ;
        RECT 19.175 85.580 19.465 85.625 ;
        RECT 21.695 85.580 21.985 85.625 ;
        RECT 17.985 85.440 21.985 85.580 ;
        RECT 25.920 85.580 26.060 86.075 ;
        RECT 26.750 86.060 27.070 86.075 ;
        RECT 31.350 86.060 31.670 86.120 ;
        RECT 28.130 85.720 28.450 85.980 ;
        RECT 29.510 85.720 29.830 85.980 ;
        RECT 42.480 85.965 42.620 86.460 ;
        RECT 44.690 86.400 45.010 86.460 ;
        RECT 45.165 86.415 45.455 86.460 ;
        RECT 46.085 86.600 46.375 86.645 ;
        RECT 46.530 86.600 46.850 86.660 ;
        RECT 46.085 86.460 46.850 86.600 ;
        RECT 46.085 86.415 46.375 86.460 ;
        RECT 46.530 86.400 46.850 86.460 ;
        RECT 53.445 86.600 53.735 86.645 ;
        RECT 53.890 86.600 54.210 86.660 ;
        RECT 57.110 86.600 57.430 86.660 ;
        RECT 53.445 86.460 57.430 86.600 ;
        RECT 53.445 86.415 53.735 86.460 ;
        RECT 53.890 86.400 54.210 86.460 ;
        RECT 57.110 86.400 57.430 86.460 ;
        RECT 65.390 86.400 65.710 86.660 ;
        RECT 69.070 86.400 69.390 86.660 ;
        RECT 72.290 86.400 72.610 86.660 ;
        RECT 73.670 86.600 73.990 86.660 ;
        RECT 77.365 86.600 77.655 86.645 ;
        RECT 73.670 86.460 77.655 86.600 ;
        RECT 73.670 86.400 73.990 86.460 ;
        RECT 77.365 86.415 77.655 86.460 ;
        RECT 43.770 86.260 44.090 86.320 ;
        RECT 49.290 86.260 49.610 86.320 ;
        RECT 49.765 86.260 50.055 86.305 ;
        RECT 51.590 86.260 51.910 86.320 ;
        RECT 76.430 86.260 76.750 86.320 ;
        RECT 43.770 86.120 48.600 86.260 ;
        RECT 43.770 86.060 44.090 86.120 ;
        RECT 42.405 85.735 42.695 85.965 ;
        RECT 45.610 85.720 45.930 85.980 ;
        RECT 46.990 85.965 47.310 85.980 ;
        RECT 46.990 85.735 47.445 85.965 ;
        RECT 47.925 85.735 48.215 85.965 ;
        RECT 48.460 85.920 48.600 86.120 ;
        RECT 49.290 86.120 54.580 86.260 ;
        RECT 49.290 86.060 49.610 86.120 ;
        RECT 49.765 86.075 50.055 86.120 ;
        RECT 51.590 86.060 51.910 86.120 ;
        RECT 54.440 85.965 54.580 86.120 ;
        RECT 70.080 86.120 80.340 86.260 ;
        RECT 50.685 85.920 50.975 85.965 ;
        RECT 52.065 85.920 52.355 85.965 ;
        RECT 48.460 85.780 52.355 85.920 ;
        RECT 50.685 85.735 50.975 85.780 ;
        RECT 52.065 85.735 52.355 85.780 ;
        RECT 52.985 85.735 53.275 85.965 ;
        RECT 54.365 85.735 54.655 85.965 ;
        RECT 55.745 85.920 56.035 85.965 ;
        RECT 61.250 85.920 61.570 85.980 ;
        RECT 64.470 85.920 64.790 85.980 ;
        RECT 55.745 85.780 64.790 85.920 ;
        RECT 55.745 85.735 56.035 85.780 ;
        RECT 46.990 85.720 47.310 85.735 ;
        RECT 28.590 85.580 28.910 85.640 ;
        RECT 25.920 85.440 28.910 85.580 ;
        RECT 8.785 85.395 9.075 85.440 ;
        RECT 9.975 85.395 10.265 85.440 ;
        RECT 12.495 85.395 12.785 85.440 ;
        RECT 17.985 85.395 18.275 85.440 ;
        RECT 19.175 85.395 19.465 85.440 ;
        RECT 21.695 85.395 21.985 85.440 ;
        RECT 28.590 85.380 28.910 85.440 ;
        RECT 42.865 85.580 43.155 85.625 ;
        RECT 43.310 85.580 43.630 85.640 ;
        RECT 48.000 85.580 48.140 85.735 ;
        RECT 48.370 85.580 48.690 85.640 ;
        RECT 53.060 85.580 53.200 85.735 ;
        RECT 42.865 85.440 43.630 85.580 ;
        RECT 42.865 85.395 43.155 85.440 ;
        RECT 43.310 85.380 43.630 85.440 ;
        RECT 44.320 85.440 53.200 85.580 ;
        RECT 53.430 85.580 53.750 85.640 ;
        RECT 55.820 85.580 55.960 85.735 ;
        RECT 61.250 85.720 61.570 85.780 ;
        RECT 64.470 85.720 64.790 85.780 ;
        RECT 66.310 85.720 66.630 85.980 ;
        RECT 68.165 85.920 68.455 85.965 ;
        RECT 69.530 85.920 69.850 85.980 ;
        RECT 70.080 85.965 70.220 86.120 ;
        RECT 76.430 86.060 76.750 86.120 ;
        RECT 68.165 85.780 69.850 85.920 ;
        RECT 68.165 85.735 68.455 85.780 ;
        RECT 69.530 85.720 69.850 85.780 ;
        RECT 70.005 85.735 70.295 85.965 ;
        RECT 70.450 85.720 70.770 85.980 ;
        RECT 71.385 85.920 71.675 85.965 ;
        RECT 72.750 85.920 73.070 85.980 ;
        RECT 71.385 85.780 73.070 85.920 ;
        RECT 71.385 85.735 71.675 85.780 ;
        RECT 72.750 85.720 73.070 85.780 ;
        RECT 73.225 85.735 73.515 85.965 ;
        RECT 53.430 85.440 55.960 85.580 ;
        RECT 56.205 85.580 56.495 85.625 ;
        RECT 58.030 85.580 58.350 85.640 ;
        RECT 61.710 85.580 62.030 85.640 ;
        RECT 56.205 85.440 62.030 85.580 ;
        RECT 73.300 85.580 73.440 85.735 ;
        RECT 74.130 85.720 74.450 85.980 ;
        RECT 75.050 85.720 75.370 85.980 ;
        RECT 76.890 85.920 77.210 85.980 ;
        RECT 78.285 85.920 78.575 85.965 ;
        RECT 76.890 85.780 78.575 85.920 ;
        RECT 76.890 85.720 77.210 85.780 ;
        RECT 78.285 85.735 78.575 85.780 ;
        RECT 78.730 85.720 79.050 85.980 ;
        RECT 80.200 85.965 80.340 86.120 ;
        RECT 79.205 85.735 79.495 85.965 ;
        RECT 80.125 85.735 80.415 85.965 ;
        RECT 73.670 85.580 73.990 85.640 ;
        RECT 73.300 85.440 73.990 85.580 ;
        RECT 44.320 85.285 44.460 85.440 ;
        RECT 48.370 85.380 48.690 85.440 ;
        RECT 53.430 85.380 53.750 85.440 ;
        RECT 56.205 85.395 56.495 85.440 ;
        RECT 58.030 85.380 58.350 85.440 ;
        RECT 61.710 85.380 62.030 85.440 ;
        RECT 73.670 85.380 73.990 85.440 ;
        RECT 77.810 85.580 78.130 85.640 ;
        RECT 79.280 85.580 79.420 85.735 ;
        RECT 81.950 85.580 82.270 85.640 ;
        RECT 77.810 85.440 82.270 85.580 ;
        RECT 77.810 85.380 78.130 85.440 ;
        RECT 81.950 85.380 82.270 85.440 ;
        RECT 8.390 85.240 8.680 85.285 ;
        RECT 10.490 85.240 10.780 85.285 ;
        RECT 12.060 85.240 12.350 85.285 ;
        RECT 8.390 85.100 12.350 85.240 ;
        RECT 8.390 85.055 8.680 85.100 ;
        RECT 10.490 85.055 10.780 85.100 ;
        RECT 12.060 85.055 12.350 85.100 ;
        RECT 17.590 85.240 17.880 85.285 ;
        RECT 19.690 85.240 19.980 85.285 ;
        RECT 21.260 85.240 21.550 85.285 ;
        RECT 17.590 85.100 21.550 85.240 ;
        RECT 17.590 85.055 17.880 85.100 ;
        RECT 19.690 85.055 19.980 85.100 ;
        RECT 21.260 85.055 21.550 85.100 ;
        RECT 44.245 85.055 44.535 85.285 ;
        RECT 51.605 85.240 51.895 85.285 ;
        RECT 55.730 85.240 56.050 85.300 ;
        RECT 58.950 85.240 59.270 85.300 ;
        RECT 51.605 85.100 59.270 85.240 ;
        RECT 51.605 85.055 51.895 85.100 ;
        RECT 55.730 85.040 56.050 85.100 ;
        RECT 58.950 85.040 59.270 85.100 ;
        RECT 67.245 85.240 67.535 85.285 ;
        RECT 75.050 85.240 75.370 85.300 ;
        RECT 67.245 85.100 75.370 85.240 ;
        RECT 67.245 85.055 67.535 85.100 ;
        RECT 75.050 85.040 75.370 85.100 ;
        RECT 75.970 85.040 76.290 85.300 ;
        RECT 16.645 84.900 16.935 84.945 ;
        RECT 18.930 84.900 19.250 84.960 ;
        RECT 16.645 84.760 19.250 84.900 ;
        RECT 16.645 84.715 16.935 84.760 ;
        RECT 18.930 84.700 19.250 84.760 ;
        RECT 20.310 84.900 20.630 84.960 ;
        RECT 24.005 84.900 24.295 84.945 ;
        RECT 20.310 84.760 24.295 84.900 ;
        RECT 20.310 84.700 20.630 84.760 ;
        RECT 24.005 84.715 24.295 84.760 ;
        RECT 26.290 84.900 26.610 84.960 ;
        RECT 26.765 84.900 27.055 84.945 ;
        RECT 26.290 84.760 27.055 84.900 ;
        RECT 26.290 84.700 26.610 84.760 ;
        RECT 26.765 84.715 27.055 84.760 ;
        RECT 27.670 84.700 27.990 84.960 ;
        RECT 29.050 84.900 29.370 84.960 ;
        RECT 30.445 84.900 30.735 84.945 ;
        RECT 29.050 84.760 30.735 84.900 ;
        RECT 29.050 84.700 29.370 84.760 ;
        RECT 30.445 84.715 30.735 84.760 ;
        RECT 35.490 84.900 35.810 84.960 ;
        RECT 42.405 84.900 42.695 84.945 ;
        RECT 35.490 84.760 42.695 84.900 ;
        RECT 35.490 84.700 35.810 84.760 ;
        RECT 42.405 84.715 42.695 84.760 ;
        RECT 63.090 84.900 63.410 84.960 ;
        RECT 71.370 84.900 71.690 84.960 ;
        RECT 63.090 84.760 71.690 84.900 ;
        RECT 63.090 84.700 63.410 84.760 ;
        RECT 71.370 84.700 71.690 84.760 ;
        RECT 74.145 84.900 74.435 84.945 ;
        RECT 77.350 84.900 77.670 84.960 ;
        RECT 74.145 84.760 77.670 84.900 ;
        RECT 74.145 84.715 74.435 84.760 ;
        RECT 77.350 84.700 77.670 84.760 ;
        RECT 5.520 84.080 83.260 84.560 ;
        RECT 11.570 83.880 11.890 83.940 ;
        RECT 18.025 83.880 18.315 83.925 ;
        RECT 18.470 83.880 18.790 83.940 ;
        RECT 11.570 83.740 15.480 83.880 ;
        RECT 11.570 83.680 11.890 83.740 ;
        RECT 15.340 83.585 15.480 83.740 ;
        RECT 18.025 83.740 18.790 83.880 ;
        RECT 18.025 83.695 18.315 83.740 ;
        RECT 18.470 83.680 18.790 83.740 ;
        RECT 25.385 83.880 25.675 83.925 ;
        RECT 26.290 83.880 26.610 83.940 ;
        RECT 25.385 83.740 26.610 83.880 ;
        RECT 25.385 83.695 25.675 83.740 ;
        RECT 26.290 83.680 26.610 83.740 ;
        RECT 29.510 83.880 29.830 83.940 ;
        RECT 33.665 83.880 33.955 83.925 ;
        RECT 29.510 83.740 33.955 83.880 ;
        RECT 29.510 83.680 29.830 83.740 ;
        RECT 33.665 83.695 33.955 83.740 ;
        RECT 44.690 83.880 45.010 83.940 ;
        RECT 46.530 83.880 46.850 83.940 ;
        RECT 44.690 83.740 46.850 83.880 ;
        RECT 44.690 83.680 45.010 83.740 ;
        RECT 46.530 83.680 46.850 83.740 ;
        RECT 48.830 83.680 49.150 83.940 ;
        RECT 52.065 83.880 52.355 83.925 ;
        RECT 54.350 83.880 54.670 83.940 ;
        RECT 52.065 83.740 54.670 83.880 ;
        RECT 52.065 83.695 52.355 83.740 ;
        RECT 54.350 83.680 54.670 83.740 ;
        RECT 64.930 83.880 65.250 83.940 ;
        RECT 76.890 83.880 77.210 83.940 ;
        RECT 64.930 83.740 77.210 83.880 ;
        RECT 64.930 83.680 65.250 83.740 ;
        RECT 76.890 83.680 77.210 83.740 ;
        RECT 7.470 83.540 7.760 83.585 ;
        RECT 9.570 83.540 9.860 83.585 ;
        RECT 11.140 83.540 11.430 83.585 ;
        RECT 7.470 83.400 11.430 83.540 ;
        RECT 7.470 83.355 7.760 83.400 ;
        RECT 9.570 83.355 9.860 83.400 ;
        RECT 11.140 83.355 11.430 83.400 ;
        RECT 15.265 83.355 15.555 83.585 ;
        RECT 26.790 83.540 27.080 83.585 ;
        RECT 28.890 83.540 29.180 83.585 ;
        RECT 30.460 83.540 30.750 83.585 ;
        RECT 26.790 83.400 30.750 83.540 ;
        RECT 26.790 83.355 27.080 83.400 ;
        RECT 28.890 83.355 29.180 83.400 ;
        RECT 30.460 83.355 30.750 83.400 ;
        RECT 36.410 83.540 36.700 83.585 ;
        RECT 37.980 83.540 38.270 83.585 ;
        RECT 40.080 83.540 40.370 83.585 ;
        RECT 52.510 83.540 52.830 83.600 ;
        RECT 36.410 83.400 40.370 83.540 ;
        RECT 36.410 83.355 36.700 83.400 ;
        RECT 37.980 83.355 38.270 83.400 ;
        RECT 40.080 83.355 40.370 83.400 ;
        RECT 49.380 83.400 52.830 83.540 ;
        RECT 6.970 83.000 7.290 83.260 ;
        RECT 7.865 83.200 8.155 83.245 ;
        RECT 9.055 83.200 9.345 83.245 ;
        RECT 11.575 83.200 11.865 83.245 ;
        RECT 23.530 83.200 23.850 83.260 ;
        RECT 7.865 83.060 11.865 83.200 ;
        RECT 7.865 83.015 8.155 83.060 ;
        RECT 9.055 83.015 9.345 83.060 ;
        RECT 11.575 83.015 11.865 83.060 ;
        RECT 22.700 83.060 23.850 83.200 ;
        RECT 7.430 82.860 7.750 82.920 ;
        RECT 8.265 82.860 8.555 82.905 ;
        RECT 7.430 82.720 8.555 82.860 ;
        RECT 7.430 82.660 7.750 82.720 ;
        RECT 8.265 82.675 8.555 82.720 ;
        RECT 18.930 82.660 19.250 82.920 ;
        RECT 20.310 82.660 20.630 82.920 ;
        RECT 20.785 82.675 21.075 82.905 ;
        RECT 21.230 82.860 21.550 82.920 ;
        RECT 22.700 82.860 22.840 83.060 ;
        RECT 23.530 83.000 23.850 83.060 ;
        RECT 25.370 83.200 25.690 83.260 ;
        RECT 26.290 83.200 26.610 83.260 ;
        RECT 25.370 83.060 26.610 83.200 ;
        RECT 25.370 83.000 25.690 83.060 ;
        RECT 26.290 83.000 26.610 83.060 ;
        RECT 27.185 83.200 27.475 83.245 ;
        RECT 28.375 83.200 28.665 83.245 ;
        RECT 30.895 83.200 31.185 83.245 ;
        RECT 27.185 83.060 31.185 83.200 ;
        RECT 27.185 83.015 27.475 83.060 ;
        RECT 28.375 83.015 28.665 83.060 ;
        RECT 30.895 83.015 31.185 83.060 ;
        RECT 35.975 83.200 36.265 83.245 ;
        RECT 38.495 83.200 38.785 83.245 ;
        RECT 39.685 83.200 39.975 83.245 ;
        RECT 48.830 83.200 49.150 83.260 ;
        RECT 35.975 83.060 39.975 83.200 ;
        RECT 35.975 83.015 36.265 83.060 ;
        RECT 38.495 83.015 38.785 83.060 ;
        RECT 39.685 83.015 39.975 83.060 ;
        RECT 47.540 83.060 49.150 83.200 ;
        RECT 21.230 82.720 22.840 82.860 ;
        RECT 23.070 82.860 23.390 82.920 ;
        RECT 27.670 82.905 27.990 82.920 ;
        RECT 24.005 82.860 24.295 82.905 ;
        RECT 23.070 82.720 24.295 82.860 ;
        RECT 14.330 82.520 14.650 82.580 ;
        RECT 16.185 82.520 16.475 82.565 ;
        RECT 14.330 82.380 16.475 82.520 ;
        RECT 14.330 82.320 14.650 82.380 ;
        RECT 16.185 82.335 16.475 82.380 ;
        RECT 19.850 82.320 20.170 82.580 ;
        RECT 20.860 82.520 21.000 82.675 ;
        RECT 21.230 82.660 21.550 82.720 ;
        RECT 23.070 82.660 23.390 82.720 ;
        RECT 24.005 82.675 24.295 82.720 ;
        RECT 24.925 82.675 25.215 82.905 ;
        RECT 25.845 82.675 26.135 82.905 ;
        RECT 27.640 82.860 27.990 82.905 ;
        RECT 27.475 82.720 27.990 82.860 ;
        RECT 27.640 82.675 27.990 82.720 ;
        RECT 23.530 82.520 23.850 82.580 ;
        RECT 25.000 82.520 25.140 82.675 ;
        RECT 20.860 82.380 22.840 82.520 ;
        RECT 22.700 82.240 22.840 82.380 ;
        RECT 23.530 82.380 25.140 82.520 ;
        RECT 23.530 82.320 23.850 82.380 ;
        RECT 13.885 82.180 14.175 82.225 ;
        RECT 15.250 82.180 15.570 82.240 ;
        RECT 13.885 82.040 15.570 82.180 ;
        RECT 13.885 81.995 14.175 82.040 ;
        RECT 15.250 81.980 15.570 82.040 ;
        RECT 16.630 81.980 16.950 82.240 ;
        RECT 17.105 82.180 17.395 82.225 ;
        RECT 17.550 82.180 17.870 82.240 ;
        RECT 17.105 82.040 17.870 82.180 ;
        RECT 17.105 81.995 17.395 82.040 ;
        RECT 17.550 81.980 17.870 82.040 ;
        RECT 20.770 82.180 21.090 82.240 ;
        RECT 21.705 82.180 21.995 82.225 ;
        RECT 20.770 82.040 21.995 82.180 ;
        RECT 20.770 81.980 21.090 82.040 ;
        RECT 21.705 81.995 21.995 82.040 ;
        RECT 22.610 81.980 22.930 82.240 ;
        RECT 25.920 82.180 26.060 82.675 ;
        RECT 27.670 82.660 27.990 82.675 ;
        RECT 40.550 82.660 40.870 82.920 ;
        RECT 46.545 82.860 46.835 82.905 ;
        RECT 46.990 82.860 47.310 82.920 ;
        RECT 47.540 82.905 47.680 83.060 ;
        RECT 48.830 83.000 49.150 83.060 ;
        RECT 46.545 82.720 47.310 82.860 ;
        RECT 46.545 82.675 46.835 82.720 ;
        RECT 46.990 82.660 47.310 82.720 ;
        RECT 47.465 82.675 47.755 82.905 ;
        RECT 49.380 82.860 49.520 83.400 ;
        RECT 52.510 83.340 52.830 83.400 ;
        RECT 53.905 83.540 54.195 83.585 ;
        RECT 58.490 83.540 58.810 83.600 ;
        RECT 69.070 83.540 69.390 83.600 ;
        RECT 53.905 83.400 58.810 83.540 ;
        RECT 53.905 83.355 54.195 83.400 ;
        RECT 58.490 83.340 58.810 83.400 ;
        RECT 65.940 83.400 69.390 83.540 ;
        RECT 50.670 83.200 50.990 83.260 ;
        RECT 54.365 83.200 54.655 83.245 ;
        RECT 56.650 83.200 56.970 83.260 ;
        RECT 50.670 83.060 53.200 83.200 ;
        RECT 50.670 83.000 50.990 83.060 ;
        RECT 48.000 82.720 49.520 82.860 ;
        RECT 49.750 82.860 50.070 82.920 ;
        RECT 50.760 82.860 50.900 83.000 ;
        RECT 49.750 82.720 50.900 82.860 ;
        RECT 29.970 82.520 30.290 82.580 ;
        RECT 39.230 82.520 39.520 82.565 ;
        RECT 29.970 82.380 39.520 82.520 ;
        RECT 29.970 82.320 30.290 82.380 ;
        RECT 39.230 82.335 39.520 82.380 ;
        RECT 45.150 82.520 45.470 82.580 ;
        RECT 48.000 82.565 48.140 82.720 ;
        RECT 49.750 82.660 50.070 82.720 ;
        RECT 52.050 82.660 52.370 82.920 ;
        RECT 53.060 82.905 53.200 83.060 ;
        RECT 54.365 83.060 56.970 83.200 ;
        RECT 54.365 83.015 54.655 83.060 ;
        RECT 56.650 83.000 56.970 83.060 ;
        RECT 52.525 82.675 52.815 82.905 ;
        RECT 52.985 82.675 53.275 82.905 ;
        RECT 53.445 82.860 53.735 82.905 ;
        RECT 53.890 82.860 54.210 82.920 ;
        RECT 62.170 82.860 62.490 82.920 ;
        RECT 53.445 82.720 54.210 82.860 ;
        RECT 53.445 82.675 53.735 82.720 ;
        RECT 47.925 82.520 48.215 82.565 ;
        RECT 49.005 82.520 49.295 82.565 ;
        RECT 49.840 82.520 49.980 82.660 ;
        RECT 45.150 82.380 48.215 82.520 ;
        RECT 48.795 82.380 49.980 82.520 ;
        RECT 50.210 82.520 50.530 82.580 ;
        RECT 52.140 82.520 52.280 82.660 ;
        RECT 50.210 82.380 52.280 82.520 ;
        RECT 52.600 82.520 52.740 82.675 ;
        RECT 53.890 82.660 54.210 82.720 ;
        RECT 54.440 82.720 62.490 82.860 ;
        RECT 54.440 82.520 54.580 82.720 ;
        RECT 62.170 82.660 62.490 82.720 ;
        RECT 65.390 82.660 65.710 82.920 ;
        RECT 65.940 82.905 66.080 83.400 ;
        RECT 69.070 83.340 69.390 83.400 ;
        RECT 70.950 83.540 71.240 83.585 ;
        RECT 73.050 83.540 73.340 83.585 ;
        RECT 74.620 83.540 74.910 83.585 ;
        RECT 70.950 83.400 74.910 83.540 ;
        RECT 70.950 83.355 71.240 83.400 ;
        RECT 73.050 83.355 73.340 83.400 ;
        RECT 74.620 83.355 74.910 83.400 ;
        RECT 71.345 83.200 71.635 83.245 ;
        RECT 72.535 83.200 72.825 83.245 ;
        RECT 75.055 83.200 75.345 83.245 ;
        RECT 71.345 83.060 75.345 83.200 ;
        RECT 71.345 83.015 71.635 83.060 ;
        RECT 72.535 83.015 72.825 83.060 ;
        RECT 75.055 83.015 75.345 83.060 ;
        RECT 77.350 83.200 77.670 83.260 ;
        RECT 77.350 83.060 79.880 83.200 ;
        RECT 77.350 83.000 77.670 83.060 ;
        RECT 65.865 82.675 66.155 82.905 ;
        RECT 66.310 82.660 66.630 82.920 ;
        RECT 67.230 82.660 67.550 82.920 ;
        RECT 67.705 82.675 67.995 82.905 ;
        RECT 68.165 82.860 68.455 82.905 ;
        RECT 69.990 82.860 70.310 82.920 ;
        RECT 68.165 82.720 70.310 82.860 ;
        RECT 68.165 82.675 68.455 82.720 ;
        RECT 52.600 82.380 54.580 82.520 ;
        RECT 45.150 82.320 45.470 82.380 ;
        RECT 47.925 82.335 48.215 82.380 ;
        RECT 48.920 82.335 49.295 82.380 ;
        RECT 31.350 82.180 31.670 82.240 ;
        RECT 33.205 82.180 33.495 82.225 ;
        RECT 25.920 82.040 33.495 82.180 ;
        RECT 31.350 81.980 31.670 82.040 ;
        RECT 33.205 81.995 33.495 82.040 ;
        RECT 46.530 82.180 46.850 82.240 ;
        RECT 47.005 82.180 47.295 82.225 ;
        RECT 46.530 82.040 47.295 82.180 ;
        RECT 46.530 81.980 46.850 82.040 ;
        RECT 47.005 81.995 47.295 82.040 ;
        RECT 47.450 82.180 47.770 82.240 ;
        RECT 48.920 82.180 49.060 82.335 ;
        RECT 50.210 82.320 50.530 82.380 ;
        RECT 54.825 82.335 55.115 82.565 ;
        RECT 47.450 82.040 49.060 82.180 ;
        RECT 47.450 81.980 47.770 82.040 ;
        RECT 49.750 81.980 50.070 82.240 ;
        RECT 50.685 82.180 50.975 82.225 ;
        RECT 52.050 82.180 52.370 82.240 ;
        RECT 50.685 82.040 52.370 82.180 ;
        RECT 50.685 81.995 50.975 82.040 ;
        RECT 52.050 81.980 52.370 82.040 ;
        RECT 52.970 82.180 53.290 82.240 ;
        RECT 54.900 82.180 55.040 82.335 ;
        RECT 55.730 82.320 56.050 82.580 ;
        RECT 65.480 82.520 65.620 82.660 ;
        RECT 67.780 82.520 67.920 82.675 ;
        RECT 69.990 82.660 70.310 82.720 ;
        RECT 70.465 82.860 70.755 82.905 ;
        RECT 73.670 82.860 73.990 82.920 ;
        RECT 79.740 82.905 79.880 83.060 ;
        RECT 79.205 82.860 79.495 82.905 ;
        RECT 70.465 82.720 72.980 82.860 ;
        RECT 70.465 82.675 70.755 82.720 ;
        RECT 72.840 82.580 72.980 82.720 ;
        RECT 73.670 82.720 79.495 82.860 ;
        RECT 73.670 82.660 73.990 82.720 ;
        RECT 79.205 82.675 79.495 82.720 ;
        RECT 79.665 82.675 79.955 82.905 ;
        RECT 80.110 82.660 80.430 82.920 ;
        RECT 81.045 82.860 81.335 82.905 ;
        RECT 81.490 82.860 81.810 82.920 ;
        RECT 81.045 82.720 81.810 82.860 ;
        RECT 81.045 82.675 81.335 82.720 ;
        RECT 68.610 82.520 68.930 82.580 ;
        RECT 65.480 82.380 68.930 82.520 ;
        RECT 68.610 82.320 68.930 82.380 ;
        RECT 69.545 82.520 69.835 82.565 ;
        RECT 71.690 82.520 71.980 82.565 ;
        RECT 69.545 82.380 71.980 82.520 ;
        RECT 69.545 82.335 69.835 82.380 ;
        RECT 71.690 82.335 71.980 82.380 ;
        RECT 72.750 82.320 73.070 82.580 ;
        RECT 74.130 82.520 74.450 82.580 ;
        RECT 75.510 82.520 75.830 82.580 ;
        RECT 74.130 82.380 75.830 82.520 ;
        RECT 74.130 82.320 74.450 82.380 ;
        RECT 75.510 82.320 75.830 82.380 ;
        RECT 78.730 82.520 79.050 82.580 ;
        RECT 81.120 82.520 81.260 82.675 ;
        RECT 81.490 82.660 81.810 82.720 ;
        RECT 78.730 82.380 81.260 82.520 ;
        RECT 78.730 82.320 79.050 82.380 ;
        RECT 52.970 82.040 55.040 82.180 ;
        RECT 56.665 82.180 56.955 82.225 ;
        RECT 59.410 82.180 59.730 82.240 ;
        RECT 56.665 82.040 59.730 82.180 ;
        RECT 52.970 81.980 53.290 82.040 ;
        RECT 56.665 81.995 56.955 82.040 ;
        RECT 59.410 81.980 59.730 82.040 ;
        RECT 62.630 82.180 62.950 82.240 ;
        RECT 64.470 82.180 64.790 82.240 ;
        RECT 62.630 82.040 64.790 82.180 ;
        RECT 62.630 81.980 62.950 82.040 ;
        RECT 64.470 81.980 64.790 82.040 ;
        RECT 65.405 82.180 65.695 82.225 ;
        RECT 66.770 82.180 67.090 82.240 ;
        RECT 65.405 82.040 67.090 82.180 ;
        RECT 65.405 81.995 65.695 82.040 ;
        RECT 66.770 81.980 67.090 82.040 ;
        RECT 69.990 82.180 70.310 82.240 ;
        RECT 75.050 82.180 75.370 82.240 ;
        RECT 77.365 82.180 77.655 82.225 ;
        RECT 69.990 82.040 77.655 82.180 ;
        RECT 69.990 81.980 70.310 82.040 ;
        RECT 75.050 81.980 75.370 82.040 ;
        RECT 77.365 81.995 77.655 82.040 ;
        RECT 77.810 81.980 78.130 82.240 ;
        RECT 5.520 81.360 83.260 81.840 ;
        RECT 14.790 81.160 15.110 81.220 ;
        RECT 15.725 81.160 16.015 81.205 ;
        RECT 14.790 81.020 16.015 81.160 ;
        RECT 14.790 80.960 15.110 81.020 ;
        RECT 15.725 80.975 16.015 81.020 ;
        RECT 17.550 80.960 17.870 81.220 ;
        RECT 19.850 80.960 20.170 81.220 ;
        RECT 22.165 81.160 22.455 81.205 ;
        RECT 23.070 81.160 23.390 81.220 ;
        RECT 29.510 81.160 29.830 81.220 ;
        RECT 22.165 81.020 23.390 81.160 ;
        RECT 22.165 80.975 22.455 81.020 ;
        RECT 23.070 80.960 23.390 81.020 ;
        RECT 25.000 81.020 29.830 81.160 ;
        RECT 16.630 80.820 16.950 80.880 ;
        RECT 25.000 80.865 25.140 81.020 ;
        RECT 29.510 80.960 29.830 81.020 ;
        RECT 29.970 80.960 30.290 81.220 ;
        RECT 45.150 81.160 45.470 81.220 ;
        RECT 45.625 81.160 45.915 81.205 ;
        RECT 45.150 81.020 45.915 81.160 ;
        RECT 45.150 80.960 45.470 81.020 ;
        RECT 45.625 80.975 45.915 81.020 ;
        RECT 46.990 80.960 47.310 81.220 ;
        RECT 47.910 80.960 48.230 81.220 ;
        RECT 48.830 81.160 49.150 81.220 ;
        RECT 54.365 81.160 54.655 81.205 ;
        RECT 48.830 81.020 54.655 81.160 ;
        RECT 48.830 80.960 49.150 81.020 ;
        RECT 54.365 80.975 54.655 81.020 ;
        RECT 55.270 81.160 55.590 81.220 ;
        RECT 56.665 81.160 56.955 81.205 ;
        RECT 55.270 81.020 56.955 81.160 ;
        RECT 55.270 80.960 55.590 81.020 ;
        RECT 56.665 80.975 56.955 81.020 ;
        RECT 57.570 80.960 57.890 81.220 ;
        RECT 63.105 81.160 63.395 81.205 ;
        RECT 76.430 81.160 76.750 81.220 ;
        RECT 63.105 81.020 76.750 81.160 ;
        RECT 63.105 80.975 63.395 81.020 ;
        RECT 76.430 80.960 76.750 81.020 ;
        RECT 16.630 80.680 23.300 80.820 ;
        RECT 16.630 80.620 16.950 80.680 ;
        RECT 6.970 80.280 7.290 80.540 ;
        RECT 8.350 80.525 8.670 80.540 ;
        RECT 8.320 80.295 8.670 80.525 ;
        RECT 8.350 80.280 8.670 80.295 ;
        RECT 10.190 80.480 10.510 80.540 ;
        RECT 14.345 80.480 14.635 80.525 ;
        RECT 10.190 80.340 14.635 80.480 ;
        RECT 10.190 80.280 10.510 80.340 ;
        RECT 14.345 80.295 14.635 80.340 ;
        RECT 15.265 80.295 15.555 80.525 ;
        RECT 15.710 80.480 16.030 80.540 ;
        RECT 16.185 80.480 16.475 80.525 ;
        RECT 15.710 80.340 16.475 80.480 ;
        RECT 7.865 80.140 8.155 80.185 ;
        RECT 9.055 80.140 9.345 80.185 ;
        RECT 11.575 80.140 11.865 80.185 ;
        RECT 7.865 80.000 11.865 80.140 ;
        RECT 15.340 80.140 15.480 80.295 ;
        RECT 15.710 80.280 16.030 80.340 ;
        RECT 16.185 80.295 16.475 80.340 ;
        RECT 17.105 80.480 17.395 80.525 ;
        RECT 18.010 80.480 18.330 80.540 ;
        RECT 18.485 80.480 18.775 80.525 ;
        RECT 17.105 80.340 18.775 80.480 ;
        RECT 17.105 80.295 17.395 80.340 ;
        RECT 18.010 80.280 18.330 80.340 ;
        RECT 18.485 80.295 18.775 80.340 ;
        RECT 19.405 80.480 19.695 80.525 ;
        RECT 20.310 80.480 20.630 80.540 ;
        RECT 19.405 80.340 20.630 80.480 ;
        RECT 19.405 80.295 19.695 80.340 ;
        RECT 19.480 80.140 19.620 80.295 ;
        RECT 20.310 80.280 20.630 80.340 ;
        RECT 21.230 80.280 21.550 80.540 ;
        RECT 21.690 80.280 22.010 80.540 ;
        RECT 23.160 80.525 23.300 80.680 ;
        RECT 24.925 80.635 25.215 80.865 ;
        RECT 25.370 80.820 25.690 80.880 ;
        RECT 25.925 80.820 26.215 80.865 ;
        RECT 28.130 80.820 28.450 80.880 ;
        RECT 25.370 80.680 28.450 80.820 ;
        RECT 25.370 80.620 25.690 80.680 ;
        RECT 25.925 80.635 26.215 80.680 ;
        RECT 28.130 80.620 28.450 80.680 ;
        RECT 28.590 80.820 28.910 80.880 ;
        RECT 29.065 80.820 29.355 80.865 ;
        RECT 32.270 80.820 32.590 80.880 ;
        RECT 35.045 80.820 35.335 80.865 ;
        RECT 28.590 80.680 35.335 80.820 ;
        RECT 48.000 80.820 48.140 80.960 ;
        RECT 50.670 80.820 50.990 80.880 ;
        RECT 54.825 80.820 55.115 80.865 ;
        RECT 48.000 80.680 49.520 80.820 ;
        RECT 28.590 80.620 28.910 80.680 ;
        RECT 29.065 80.635 29.355 80.680 ;
        RECT 32.270 80.620 32.590 80.680 ;
        RECT 35.045 80.635 35.335 80.680 ;
        RECT 23.085 80.295 23.375 80.525 ;
        RECT 23.530 80.480 23.850 80.540 ;
        RECT 25.460 80.480 25.600 80.620 ;
        RECT 23.530 80.340 25.600 80.480 ;
        RECT 27.225 80.480 27.515 80.525 ;
        RECT 36.425 80.480 36.715 80.525 ;
        RECT 27.225 80.340 36.715 80.480 ;
        RECT 23.530 80.280 23.850 80.340 ;
        RECT 27.225 80.295 27.515 80.340 ;
        RECT 36.425 80.295 36.715 80.340 ;
        RECT 36.870 80.480 37.190 80.540 ;
        RECT 37.345 80.480 37.635 80.525 ;
        RECT 36.870 80.340 37.635 80.480 ;
        RECT 15.340 80.000 19.620 80.140 ;
        RECT 19.850 80.140 20.170 80.200 ;
        RECT 24.005 80.140 24.295 80.185 ;
        RECT 19.850 80.000 24.295 80.140 ;
        RECT 7.865 79.955 8.155 80.000 ;
        RECT 9.055 79.955 9.345 80.000 ;
        RECT 11.575 79.955 11.865 80.000 ;
        RECT 19.850 79.940 20.170 80.000 ;
        RECT 24.005 79.955 24.295 80.000 ;
        RECT 7.470 79.800 7.760 79.845 ;
        RECT 9.570 79.800 9.860 79.845 ;
        RECT 11.140 79.800 11.430 79.845 ;
        RECT 7.470 79.660 11.430 79.800 ;
        RECT 7.470 79.615 7.760 79.660 ;
        RECT 9.570 79.615 9.860 79.660 ;
        RECT 11.140 79.615 11.430 79.660 ;
        RECT 13.870 79.800 14.190 79.860 ;
        RECT 18.010 79.800 18.330 79.860 ;
        RECT 21.690 79.800 22.010 79.860 ;
        RECT 24.910 79.800 25.230 79.860 ;
        RECT 13.870 79.660 22.010 79.800 ;
        RECT 13.870 79.600 14.190 79.660 ;
        RECT 18.010 79.600 18.330 79.660 ;
        RECT 21.690 79.600 22.010 79.660 ;
        RECT 22.240 79.660 25.230 79.800 ;
        RECT 14.790 79.460 15.110 79.520 ;
        RECT 22.240 79.460 22.380 79.660 ;
        RECT 24.910 79.600 25.230 79.660 ;
        RECT 26.765 79.800 27.055 79.845 ;
        RECT 27.300 79.800 27.440 80.295 ;
        RECT 36.870 80.280 37.190 80.340 ;
        RECT 37.345 80.295 37.635 80.340 ;
        RECT 43.770 80.280 44.090 80.540 ;
        RECT 44.690 80.280 45.010 80.540 ;
        RECT 45.610 80.480 45.930 80.540 ;
        RECT 46.545 80.480 46.835 80.525 ;
        RECT 45.610 80.340 46.835 80.480 ;
        RECT 45.610 80.280 45.930 80.340 ;
        RECT 46.545 80.295 46.835 80.340 ;
        RECT 47.910 80.280 48.230 80.540 ;
        RECT 48.370 80.280 48.690 80.540 ;
        RECT 49.380 80.525 49.520 80.680 ;
        RECT 50.670 80.680 55.115 80.820 ;
        RECT 57.110 80.820 57.430 80.880 ;
        RECT 58.345 80.820 58.635 80.865 ;
        RECT 50.670 80.620 50.990 80.680 ;
        RECT 54.825 80.635 55.115 80.680 ;
        RECT 55.975 80.650 56.265 80.695 ;
        RECT 49.305 80.295 49.595 80.525 ;
        RECT 52.065 80.480 52.355 80.525 ;
        RECT 52.525 80.480 52.815 80.525 ;
        RECT 49.840 80.340 52.815 80.480 ;
        RECT 27.670 79.800 27.990 79.860 ;
        RECT 26.765 79.660 27.990 79.800 ;
        RECT 26.765 79.615 27.055 79.660 ;
        RECT 27.670 79.600 27.990 79.660 ;
        RECT 28.590 79.800 28.910 79.860 ;
        RECT 33.205 79.800 33.495 79.845 ;
        RECT 38.265 79.800 38.555 79.845 ;
        RECT 28.590 79.660 33.495 79.800 ;
        RECT 28.590 79.600 28.910 79.660 ;
        RECT 33.205 79.615 33.495 79.660 ;
        RECT 35.120 79.660 38.555 79.800 ;
        RECT 44.780 79.800 44.920 80.280 ;
        RECT 48.460 79.800 48.600 80.280 ;
        RECT 49.840 80.200 49.980 80.340 ;
        RECT 52.065 80.295 52.355 80.340 ;
        RECT 52.525 80.295 52.815 80.340 ;
        RECT 53.430 80.480 53.750 80.540 ;
        RECT 55.920 80.480 56.265 80.650 ;
        RECT 57.110 80.680 58.635 80.820 ;
        RECT 57.110 80.620 57.430 80.680 ;
        RECT 58.345 80.635 58.635 80.680 ;
        RECT 59.410 80.620 59.730 80.880 ;
        RECT 61.725 80.820 62.015 80.865 ;
        RECT 65.405 80.820 65.695 80.865 ;
        RECT 67.230 80.820 67.550 80.880 ;
        RECT 70.005 80.820 70.295 80.865 ;
        RECT 61.725 80.680 67.000 80.820 ;
        RECT 61.725 80.635 62.015 80.680 ;
        RECT 65.405 80.635 65.695 80.680 ;
        RECT 53.430 80.465 56.265 80.480 ;
        RECT 53.430 80.340 56.060 80.465 ;
        RECT 53.430 80.280 53.750 80.340 ;
        RECT 61.250 80.280 61.570 80.540 ;
        RECT 64.025 80.295 64.315 80.525 ;
        RECT 64.485 80.295 64.775 80.525 ;
        RECT 66.310 80.480 66.630 80.540 ;
        RECT 66.860 80.525 67.000 80.680 ;
        RECT 67.230 80.680 70.295 80.820 ;
        RECT 67.230 80.620 67.550 80.680 ;
        RECT 70.005 80.635 70.295 80.680 ;
        RECT 70.450 80.820 70.770 80.880 ;
        RECT 71.845 80.820 72.135 80.865 ;
        RECT 74.590 80.820 74.910 80.880 ;
        RECT 70.450 80.680 72.135 80.820 ;
        RECT 70.450 80.620 70.770 80.680 ;
        RECT 71.845 80.635 72.135 80.680 ;
        RECT 73.760 80.680 74.910 80.820 ;
        RECT 66.785 80.480 67.075 80.525 ;
        RECT 66.310 80.340 67.075 80.480 ;
        RECT 48.845 80.140 49.135 80.185 ;
        RECT 49.750 80.140 50.070 80.200 ;
        RECT 48.845 80.000 50.070 80.140 ;
        RECT 48.845 79.955 49.135 80.000 ;
        RECT 49.750 79.940 50.070 80.000 ;
        RECT 50.670 80.140 50.990 80.200 ;
        RECT 51.605 80.140 51.895 80.185 ;
        RECT 50.670 80.000 52.740 80.140 ;
        RECT 50.670 79.940 50.990 80.000 ;
        RECT 51.605 79.955 51.895 80.000 ;
        RECT 52.600 79.800 52.740 80.000 ;
        RECT 52.970 79.940 53.290 80.200 ;
        RECT 54.350 80.140 54.670 80.200 ;
        RECT 57.570 80.140 57.890 80.200 ;
        RECT 62.630 80.140 62.950 80.200 ;
        RECT 54.350 80.000 57.890 80.140 ;
        RECT 54.350 79.940 54.670 80.000 ;
        RECT 57.570 79.940 57.890 80.000 ;
        RECT 62.030 80.000 62.950 80.140 ;
        RECT 56.650 79.800 56.970 79.860 ;
        RECT 62.030 79.800 62.170 80.000 ;
        RECT 62.630 79.940 62.950 80.000 ;
        RECT 44.780 79.660 48.140 79.800 ;
        RECT 48.460 79.660 52.280 79.800 ;
        RECT 52.600 79.660 62.170 79.800 ;
        RECT 64.100 79.800 64.240 80.295 ;
        RECT 64.560 80.140 64.700 80.295 ;
        RECT 66.310 80.280 66.630 80.340 ;
        RECT 66.785 80.295 67.075 80.340 ;
        RECT 67.705 80.295 67.995 80.525 ;
        RECT 69.530 80.480 69.850 80.540 ;
        RECT 70.925 80.480 71.215 80.525 ;
        RECT 69.530 80.340 71.215 80.480 ;
        RECT 67.230 80.140 67.550 80.200 ;
        RECT 67.780 80.140 67.920 80.295 ;
        RECT 69.530 80.280 69.850 80.340 ;
        RECT 70.925 80.295 71.215 80.340 ;
        RECT 73.210 80.280 73.530 80.540 ;
        RECT 73.760 80.525 73.900 80.680 ;
        RECT 74.590 80.620 74.910 80.680 ;
        RECT 75.940 80.820 76.230 80.865 ;
        RECT 77.810 80.820 78.130 80.880 ;
        RECT 75.940 80.680 78.130 80.820 ;
        RECT 75.940 80.635 76.230 80.680 ;
        RECT 77.810 80.620 78.130 80.680 ;
        RECT 73.685 80.295 73.975 80.525 ;
        RECT 78.270 80.480 78.590 80.540 ;
        RECT 74.220 80.340 78.590 80.480 ;
        RECT 64.560 80.000 67.920 80.140 ;
        RECT 72.305 80.140 72.595 80.185 ;
        RECT 74.220 80.140 74.360 80.340 ;
        RECT 78.270 80.280 78.590 80.340 ;
        RECT 72.305 80.000 74.360 80.140 ;
        RECT 67.230 79.940 67.550 80.000 ;
        RECT 72.305 79.955 72.595 80.000 ;
        RECT 74.605 79.955 74.895 80.185 ;
        RECT 75.485 80.140 75.775 80.185 ;
        RECT 76.675 80.140 76.965 80.185 ;
        RECT 79.195 80.140 79.485 80.185 ;
        RECT 75.485 80.000 79.485 80.140 ;
        RECT 75.485 79.955 75.775 80.000 ;
        RECT 76.675 79.955 76.965 80.000 ;
        RECT 79.195 79.955 79.485 80.000 ;
        RECT 68.165 79.800 68.455 79.845 ;
        RECT 70.450 79.800 70.770 79.860 ;
        RECT 64.100 79.660 67.920 79.800 ;
        RECT 14.790 79.320 22.380 79.460 ;
        RECT 22.610 79.460 22.930 79.520 ;
        RECT 24.450 79.460 24.770 79.520 ;
        RECT 22.610 79.320 24.770 79.460 ;
        RECT 14.790 79.260 15.110 79.320 ;
        RECT 22.610 79.260 22.930 79.320 ;
        RECT 24.450 79.260 24.770 79.320 ;
        RECT 25.845 79.460 26.135 79.505 ;
        RECT 28.130 79.460 28.450 79.520 ;
        RECT 25.845 79.320 28.450 79.460 ;
        RECT 25.845 79.275 26.135 79.320 ;
        RECT 28.130 79.260 28.450 79.320 ;
        RECT 29.050 79.260 29.370 79.520 ;
        RECT 35.120 79.505 35.260 79.660 ;
        RECT 38.265 79.615 38.555 79.660 ;
        RECT 35.045 79.275 35.335 79.505 ;
        RECT 35.950 79.260 36.270 79.520 ;
        RECT 44.690 79.260 45.010 79.520 ;
        RECT 48.000 79.460 48.140 79.660 ;
        RECT 49.750 79.460 50.070 79.520 ;
        RECT 48.000 79.320 50.070 79.460 ;
        RECT 49.750 79.260 50.070 79.320 ;
        RECT 50.210 79.260 50.530 79.520 ;
        RECT 51.590 79.260 51.910 79.520 ;
        RECT 52.140 79.460 52.280 79.660 ;
        RECT 56.650 79.600 56.970 79.660 ;
        RECT 52.525 79.460 52.815 79.505 ;
        RECT 52.140 79.320 52.815 79.460 ;
        RECT 52.525 79.275 52.815 79.320 ;
        RECT 53.890 79.460 54.210 79.520 ;
        RECT 55.745 79.460 56.035 79.505 ;
        RECT 53.890 79.320 56.035 79.460 ;
        RECT 53.890 79.260 54.210 79.320 ;
        RECT 55.745 79.275 56.035 79.320 ;
        RECT 58.490 79.260 58.810 79.520 ;
        RECT 65.850 79.260 66.170 79.520 ;
        RECT 67.780 79.460 67.920 79.660 ;
        RECT 68.165 79.660 70.770 79.800 ;
        RECT 68.165 79.615 68.455 79.660 ;
        RECT 70.450 79.600 70.770 79.660 ;
        RECT 72.750 79.800 73.070 79.860 ;
        RECT 74.680 79.800 74.820 79.955 ;
        RECT 72.750 79.660 74.820 79.800 ;
        RECT 75.090 79.800 75.380 79.845 ;
        RECT 77.190 79.800 77.480 79.845 ;
        RECT 78.760 79.800 79.050 79.845 ;
        RECT 75.090 79.660 79.050 79.800 ;
        RECT 72.750 79.600 73.070 79.660 ;
        RECT 75.090 79.615 75.380 79.660 ;
        RECT 77.190 79.615 77.480 79.660 ;
        RECT 78.760 79.615 79.050 79.660 ;
        RECT 79.190 79.460 79.510 79.520 ;
        RECT 80.110 79.460 80.430 79.520 ;
        RECT 81.505 79.460 81.795 79.505 ;
        RECT 67.780 79.320 81.795 79.460 ;
        RECT 79.190 79.260 79.510 79.320 ;
        RECT 80.110 79.260 80.430 79.320 ;
        RECT 81.505 79.275 81.795 79.320 ;
        RECT 5.520 78.640 83.260 79.120 ;
        RECT 7.905 78.440 8.195 78.485 ;
        RECT 8.350 78.440 8.670 78.500 ;
        RECT 7.905 78.300 8.670 78.440 ;
        RECT 7.905 78.255 8.195 78.300 ;
        RECT 8.350 78.240 8.670 78.300 ;
        RECT 8.810 78.440 9.130 78.500 ;
        RECT 13.410 78.440 13.730 78.500 ;
        RECT 8.810 78.300 13.730 78.440 ;
        RECT 8.810 78.240 9.130 78.300 ;
        RECT 13.410 78.240 13.730 78.300 ;
        RECT 13.885 78.440 14.175 78.485 ;
        RECT 17.105 78.440 17.395 78.485 ;
        RECT 19.390 78.440 19.710 78.500 ;
        RECT 13.885 78.300 15.400 78.440 ;
        RECT 13.885 78.255 14.175 78.300 ;
        RECT 15.260 78.160 15.400 78.300 ;
        RECT 17.105 78.300 19.710 78.440 ;
        RECT 17.105 78.255 17.395 78.300 ;
        RECT 19.390 78.240 19.710 78.300 ;
        RECT 23.070 78.440 23.390 78.500 ;
        RECT 23.545 78.440 23.835 78.485 ;
        RECT 23.070 78.300 23.835 78.440 ;
        RECT 23.070 78.240 23.390 78.300 ;
        RECT 23.545 78.255 23.835 78.300 ;
        RECT 23.990 78.240 24.310 78.500 ;
        RECT 26.750 78.440 27.070 78.500 ;
        RECT 27.225 78.440 27.515 78.485 ;
        RECT 26.750 78.300 27.515 78.440 ;
        RECT 26.750 78.240 27.070 78.300 ;
        RECT 27.225 78.255 27.515 78.300 ;
        RECT 28.130 78.440 28.450 78.500 ;
        RECT 31.350 78.440 31.670 78.500 ;
        RECT 28.130 78.300 31.670 78.440 ;
        RECT 28.130 78.240 28.450 78.300 ;
        RECT 31.350 78.240 31.670 78.300 ;
        RECT 33.205 78.440 33.495 78.485 ;
        RECT 34.570 78.440 34.890 78.500 ;
        RECT 36.870 78.440 37.190 78.500 ;
        RECT 33.205 78.300 37.190 78.440 ;
        RECT 33.205 78.255 33.495 78.300 ;
        RECT 34.570 78.240 34.890 78.300 ;
        RECT 36.870 78.240 37.190 78.300 ;
        RECT 40.565 78.440 40.855 78.485 ;
        RECT 41.010 78.440 41.330 78.500 ;
        RECT 40.565 78.300 41.330 78.440 ;
        RECT 40.565 78.255 40.855 78.300 ;
        RECT 41.010 78.240 41.330 78.300 ;
        RECT 41.485 78.440 41.775 78.485 ;
        RECT 42.850 78.440 43.170 78.500 ;
        RECT 48.370 78.440 48.690 78.500 ;
        RECT 41.485 78.300 43.170 78.440 ;
        RECT 41.485 78.255 41.775 78.300 ;
        RECT 42.850 78.240 43.170 78.300 ;
        RECT 43.860 78.300 48.690 78.440 ;
        RECT 14.805 77.915 15.095 78.145 ;
        RECT 10.665 77.760 10.955 77.805 ;
        RECT 13.870 77.760 14.190 77.820 ;
        RECT 10.665 77.620 14.190 77.760 ;
        RECT 14.880 77.760 15.020 77.915 ;
        RECT 15.250 77.900 15.570 78.160 ;
        RECT 18.010 78.100 18.330 78.160 ;
        RECT 22.625 78.100 22.915 78.145 ;
        RECT 24.080 78.100 24.220 78.240 ;
        RECT 35.950 78.100 36.240 78.145 ;
        RECT 37.520 78.100 37.810 78.145 ;
        RECT 39.620 78.100 39.910 78.145 ;
        RECT 18.010 77.960 20.540 78.100 ;
        RECT 18.010 77.900 18.330 77.960 ;
        RECT 16.630 77.760 16.950 77.820 ;
        RECT 20.400 77.760 20.540 77.960 ;
        RECT 22.625 77.960 24.220 78.100 ;
        RECT 27.300 77.960 32.040 78.100 ;
        RECT 22.625 77.915 22.915 77.960 ;
        RECT 27.300 77.820 27.440 77.960 ;
        RECT 23.545 77.760 23.835 77.805 ;
        RECT 14.880 77.620 20.080 77.760 ;
        RECT 20.400 77.620 23.835 77.760 ;
        RECT 10.665 77.575 10.955 77.620 ;
        RECT 13.870 77.560 14.190 77.620 ;
        RECT 16.630 77.560 16.950 77.620 ;
        RECT 12.045 77.235 12.335 77.465 ;
        RECT 13.425 77.420 13.715 77.465 ;
        RECT 14.330 77.420 14.650 77.480 ;
        RECT 13.425 77.280 14.650 77.420 ;
        RECT 13.425 77.235 13.715 77.280 ;
        RECT 8.825 77.080 9.115 77.125 ;
        RECT 9.730 77.080 10.050 77.140 ;
        RECT 8.825 76.940 10.050 77.080 ;
        RECT 12.120 77.080 12.260 77.235 ;
        RECT 14.330 77.220 14.650 77.280 ;
        RECT 17.090 77.420 17.410 77.480 ;
        RECT 18.945 77.420 19.235 77.465 ;
        RECT 17.090 77.280 19.235 77.420 ;
        RECT 17.090 77.220 17.410 77.280 ;
        RECT 18.945 77.235 19.235 77.280 ;
        RECT 19.390 77.220 19.710 77.480 ;
        RECT 19.940 77.465 20.080 77.620 ;
        RECT 23.545 77.575 23.835 77.620 ;
        RECT 23.990 77.760 24.310 77.820 ;
        RECT 23.990 77.620 26.520 77.760 ;
        RECT 23.990 77.560 24.310 77.620 ;
        RECT 19.865 77.235 20.155 77.465 ;
        RECT 20.310 77.220 20.630 77.480 ;
        RECT 20.785 77.235 21.075 77.465 ;
        RECT 18.470 77.080 18.790 77.140 ;
        RECT 12.120 76.940 18.790 77.080 ;
        RECT 19.480 77.080 19.620 77.220 ;
        RECT 20.860 77.080 21.000 77.235 ;
        RECT 24.450 77.220 24.770 77.480 ;
        RECT 24.910 77.220 25.230 77.480 ;
        RECT 25.830 77.220 26.150 77.480 ;
        RECT 26.380 77.420 26.520 77.620 ;
        RECT 27.210 77.560 27.530 77.820 ;
        RECT 27.760 77.760 28.820 77.800 ;
        RECT 27.760 77.660 30.205 77.760 ;
        RECT 27.760 77.420 27.900 77.660 ;
        RECT 28.680 77.620 30.205 77.660 ;
        RECT 26.380 77.280 27.900 77.420 ;
        RECT 28.130 77.220 28.450 77.480 ;
        RECT 29.510 77.220 29.830 77.480 ;
        RECT 30.065 77.465 30.205 77.620 ;
        RECT 29.990 77.235 30.280 77.465 ;
        RECT 31.350 77.220 31.670 77.480 ;
        RECT 31.900 77.465 32.040 77.960 ;
        RECT 35.950 77.960 39.910 78.100 ;
        RECT 35.950 77.915 36.240 77.960 ;
        RECT 37.520 77.915 37.810 77.960 ;
        RECT 39.620 77.915 39.910 77.960 ;
        RECT 35.515 77.760 35.805 77.805 ;
        RECT 38.035 77.760 38.325 77.805 ;
        RECT 39.225 77.760 39.515 77.805 ;
        RECT 35.515 77.620 39.515 77.760 ;
        RECT 35.515 77.575 35.805 77.620 ;
        RECT 38.035 77.575 38.325 77.620 ;
        RECT 39.225 77.575 39.515 77.620 ;
        RECT 40.105 77.760 40.395 77.805 ;
        RECT 40.550 77.760 40.870 77.820 ;
        RECT 40.105 77.620 40.870 77.760 ;
        RECT 40.105 77.575 40.395 77.620 ;
        RECT 40.550 77.560 40.870 77.620 ;
        RECT 31.850 77.235 32.140 77.465 ;
        RECT 35.950 77.420 36.270 77.480 ;
        RECT 38.770 77.420 39.060 77.465 ;
        RECT 35.950 77.280 39.060 77.420 ;
        RECT 35.950 77.220 36.270 77.280 ;
        RECT 38.770 77.235 39.060 77.280 ;
        RECT 41.930 77.420 42.250 77.480 ;
        RECT 43.325 77.420 43.615 77.465 ;
        RECT 41.930 77.280 43.615 77.420 ;
        RECT 43.860 77.420 44.000 78.300 ;
        RECT 48.370 78.240 48.690 78.300 ;
        RECT 48.830 78.240 49.150 78.500 ;
        RECT 49.750 78.440 50.070 78.500 ;
        RECT 52.510 78.440 52.830 78.500 ;
        RECT 64.945 78.440 65.235 78.485 ;
        RECT 49.750 78.300 52.830 78.440 ;
        RECT 49.750 78.240 50.070 78.300 ;
        RECT 52.510 78.240 52.830 78.300 ;
        RECT 60.420 78.300 65.235 78.440 ;
        RECT 45.625 78.100 45.915 78.145 ;
        RECT 52.970 78.100 53.290 78.160 ;
        RECT 54.350 78.100 54.670 78.160 ;
        RECT 58.490 78.100 58.810 78.160 ;
        RECT 45.625 77.960 54.670 78.100 ;
        RECT 45.625 77.915 45.915 77.960 ;
        RECT 52.970 77.900 53.290 77.960 ;
        RECT 54.350 77.900 54.670 77.960 ;
        RECT 56.740 77.960 58.810 78.100 ;
        RECT 44.230 77.760 44.550 77.820 ;
        RECT 44.230 77.705 45.840 77.760 ;
        RECT 46.085 77.705 46.375 77.805 ;
        RECT 47.230 77.760 48.140 77.800 ;
        RECT 53.890 77.760 54.210 77.820 ;
        RECT 44.230 77.620 46.375 77.705 ;
        RECT 44.230 77.560 44.550 77.620 ;
        RECT 45.700 77.575 46.375 77.620 ;
        RECT 46.750 77.660 54.210 77.760 ;
        RECT 46.750 77.620 47.370 77.660 ;
        RECT 48.000 77.620 54.210 77.660 ;
        RECT 45.700 77.565 46.300 77.575 ;
        RECT 44.705 77.420 44.995 77.465 ;
        RECT 43.860 77.280 44.995 77.420 ;
        RECT 41.930 77.220 42.250 77.280 ;
        RECT 43.325 77.235 43.615 77.280 ;
        RECT 44.705 77.235 44.995 77.280 ;
        RECT 45.165 77.420 45.455 77.465 ;
        RECT 46.750 77.420 46.890 77.620 ;
        RECT 53.890 77.560 54.210 77.620 ;
        RECT 47.450 77.420 47.770 77.480 ;
        RECT 45.165 77.280 46.890 77.420 ;
        RECT 47.260 77.280 47.770 77.420 ;
        RECT 45.165 77.235 45.455 77.280 ;
        RECT 47.450 77.220 47.770 77.280 ;
        RECT 48.155 77.235 48.445 77.465 ;
        RECT 48.830 77.420 49.150 77.480 ;
        RECT 49.305 77.420 49.595 77.465 ;
        RECT 48.830 77.280 49.595 77.420 ;
        RECT 19.480 76.940 21.000 77.080 ;
        RECT 8.825 76.895 9.115 76.940 ;
        RECT 9.730 76.880 10.050 76.940 ;
        RECT 18.470 76.880 18.790 76.940 ;
        RECT 29.050 76.880 29.370 77.140 ;
        RECT 30.890 76.880 31.210 77.140 ;
        RECT 48.230 77.080 48.370 77.235 ;
        RECT 48.830 77.220 49.150 77.280 ;
        RECT 49.305 77.235 49.595 77.280 ;
        RECT 49.750 77.220 50.070 77.480 ;
        RECT 50.225 77.420 50.515 77.465 ;
        RECT 50.670 77.420 50.990 77.480 ;
        RECT 50.225 77.280 50.990 77.420 ;
        RECT 50.225 77.235 50.515 77.280 ;
        RECT 50.670 77.220 50.990 77.280 ;
        RECT 51.145 77.420 51.435 77.465 ;
        RECT 51.590 77.420 51.910 77.480 ;
        RECT 51.145 77.280 51.910 77.420 ;
        RECT 51.145 77.235 51.435 77.280 ;
        RECT 51.590 77.220 51.910 77.280 ;
        RECT 52.050 77.220 52.370 77.480 ;
        RECT 52.510 77.220 52.830 77.480 ;
        RECT 52.970 77.220 53.290 77.480 ;
        RECT 54.810 77.420 55.130 77.480 ;
        RECT 56.740 77.465 56.880 77.960 ;
        RECT 58.490 77.900 58.810 77.960 ;
        RECT 57.585 77.760 57.875 77.805 ;
        RECT 59.410 77.760 59.730 77.820 ;
        RECT 57.585 77.620 59.730 77.760 ;
        RECT 57.585 77.575 57.875 77.620 ;
        RECT 59.410 77.560 59.730 77.620 ;
        RECT 55.745 77.420 56.035 77.465 ;
        RECT 54.810 77.280 56.035 77.420 ;
        RECT 54.810 77.220 55.130 77.280 ;
        RECT 55.745 77.235 56.035 77.280 ;
        RECT 56.665 77.235 56.955 77.465 ;
        RECT 57.125 77.235 57.415 77.465 ;
        RECT 58.505 77.420 58.795 77.465 ;
        RECT 58.950 77.420 59.270 77.480 ;
        RECT 58.505 77.280 59.270 77.420 ;
        RECT 58.505 77.235 58.795 77.280 ;
        RECT 54.900 77.080 55.040 77.220 ;
        RECT 48.230 76.940 49.060 77.080 ;
        RECT 48.920 76.800 49.060 76.940 ;
        RECT 53.520 76.940 55.040 77.080 ;
        RECT 15.710 76.740 16.030 76.800 ;
        RECT 17.105 76.740 17.395 76.785 ;
        RECT 15.710 76.600 17.395 76.740 ;
        RECT 15.710 76.540 16.030 76.600 ;
        RECT 17.105 76.555 17.395 76.600 ;
        RECT 18.025 76.740 18.315 76.785 ;
        RECT 19.390 76.740 19.710 76.800 ;
        RECT 18.025 76.600 19.710 76.740 ;
        RECT 18.025 76.555 18.315 76.600 ;
        RECT 19.390 76.540 19.710 76.600 ;
        RECT 19.850 76.740 20.170 76.800 ;
        RECT 22.165 76.740 22.455 76.785 ;
        RECT 19.850 76.600 22.455 76.740 ;
        RECT 19.850 76.540 20.170 76.600 ;
        RECT 22.165 76.555 22.455 76.600 ;
        RECT 25.845 76.740 26.135 76.785 ;
        RECT 31.810 76.740 32.130 76.800 ;
        RECT 25.845 76.600 32.130 76.740 ;
        RECT 25.845 76.555 26.135 76.600 ;
        RECT 31.810 76.540 32.130 76.600 ;
        RECT 32.730 76.540 33.050 76.800 ;
        RECT 41.470 76.540 41.790 76.800 ;
        RECT 46.530 76.540 46.850 76.800 ;
        RECT 48.830 76.540 49.150 76.800 ;
        RECT 51.590 76.740 51.910 76.800 ;
        RECT 53.520 76.740 53.660 76.940 ;
        RECT 51.590 76.600 53.660 76.740 ;
        RECT 54.365 76.740 54.655 76.785 ;
        RECT 54.810 76.740 55.130 76.800 ;
        RECT 54.365 76.600 55.130 76.740 ;
        RECT 51.590 76.540 51.910 76.600 ;
        RECT 54.365 76.555 54.655 76.600 ;
        RECT 54.810 76.540 55.130 76.600 ;
        RECT 56.650 76.740 56.970 76.800 ;
        RECT 57.200 76.740 57.340 77.235 ;
        RECT 58.950 77.220 59.270 77.280 ;
        RECT 59.885 77.420 60.175 77.465 ;
        RECT 60.420 77.420 60.560 78.300 ;
        RECT 64.945 78.255 65.235 78.300 ;
        RECT 67.245 78.440 67.535 78.485 ;
        RECT 69.990 78.440 70.310 78.500 ;
        RECT 71.385 78.440 71.675 78.485 ;
        RECT 67.245 78.300 71.675 78.440 ;
        RECT 67.245 78.255 67.535 78.300 ;
        RECT 69.990 78.240 70.310 78.300 ;
        RECT 71.385 78.255 71.675 78.300 ;
        RECT 72.305 78.440 72.595 78.485 ;
        RECT 73.210 78.440 73.530 78.500 ;
        RECT 72.305 78.300 73.530 78.440 ;
        RECT 72.305 78.255 72.595 78.300 ;
        RECT 73.210 78.240 73.530 78.300 ;
        RECT 73.685 78.440 73.975 78.485 ;
        RECT 74.130 78.440 74.450 78.500 ;
        RECT 73.685 78.300 74.450 78.440 ;
        RECT 73.685 78.255 73.975 78.300 ;
        RECT 74.130 78.240 74.450 78.300 ;
        RECT 68.610 78.100 68.930 78.160 ;
        RECT 75.525 78.100 75.815 78.145 ;
        RECT 68.610 77.960 75.815 78.100 ;
        RECT 68.610 77.900 68.930 77.960 ;
        RECT 75.525 77.915 75.815 77.960 ;
        RECT 78.745 77.915 79.035 78.145 ;
        RECT 75.050 77.760 75.370 77.820 ;
        RECT 75.050 77.620 77.120 77.760 ;
        RECT 75.050 77.560 75.370 77.620 ;
        RECT 59.885 77.280 60.560 77.420 ;
        RECT 59.885 77.235 60.175 77.280 ;
        RECT 61.710 77.220 62.030 77.480 ;
        RECT 62.630 77.420 62.950 77.480 ;
        RECT 63.105 77.420 63.395 77.465 ;
        RECT 70.910 77.420 71.230 77.480 ;
        RECT 73.225 77.420 73.515 77.465 ;
        RECT 62.630 77.280 63.395 77.420 ;
        RECT 62.630 77.220 62.950 77.280 ;
        RECT 63.105 77.235 63.395 77.280 ;
        RECT 66.400 77.280 70.680 77.420 ;
        RECT 66.400 77.140 66.540 77.280 ;
        RECT 58.030 77.080 58.350 77.140 ;
        RECT 60.805 77.080 61.095 77.125 ;
        RECT 58.030 76.940 61.095 77.080 ;
        RECT 58.030 76.880 58.350 76.940 ;
        RECT 60.805 76.895 61.095 76.940 ;
        RECT 61.265 77.080 61.555 77.125 ;
        RECT 64.025 77.080 64.315 77.125 ;
        RECT 64.470 77.080 64.790 77.140 ;
        RECT 61.265 76.940 63.320 77.080 ;
        RECT 61.265 76.895 61.555 76.940 ;
        RECT 63.180 76.800 63.320 76.940 ;
        RECT 64.025 76.940 64.790 77.080 ;
        RECT 64.025 76.895 64.315 76.940 ;
        RECT 64.470 76.880 64.790 76.940 ;
        RECT 66.310 76.880 66.630 77.140 ;
        RECT 66.770 77.080 67.090 77.140 ;
        RECT 70.540 77.125 70.680 77.280 ;
        RECT 70.910 77.280 73.515 77.420 ;
        RECT 70.910 77.220 71.230 77.280 ;
        RECT 73.225 77.235 73.515 77.280 ;
        RECT 74.590 77.220 74.910 77.480 ;
        RECT 76.430 77.220 76.750 77.480 ;
        RECT 76.980 77.465 77.120 77.620 ;
        RECT 76.905 77.235 77.195 77.465 ;
        RECT 77.810 77.220 78.130 77.480 ;
        RECT 78.285 77.420 78.575 77.465 ;
        RECT 78.820 77.420 78.960 77.915 ;
        RECT 78.285 77.280 78.960 77.420 ;
        RECT 78.285 77.235 78.575 77.280 ;
        RECT 79.665 77.235 79.955 77.465 ;
        RECT 67.245 77.080 67.535 77.125 ;
        RECT 66.770 76.940 67.535 77.080 ;
        RECT 66.770 76.880 67.090 76.940 ;
        RECT 67.245 76.895 67.535 76.940 ;
        RECT 70.465 76.895 70.755 77.125 ;
        RECT 79.740 77.080 79.880 77.235 ;
        RECT 80.110 77.220 80.430 77.480 ;
        RECT 80.570 77.220 80.890 77.480 ;
        RECT 81.505 77.420 81.795 77.465 ;
        RECT 81.950 77.420 82.270 77.480 ;
        RECT 81.505 77.280 82.270 77.420 ;
        RECT 81.505 77.235 81.795 77.280 ;
        RECT 81.950 77.220 82.270 77.280 ;
        RECT 73.300 76.940 79.880 77.080 ;
        RECT 73.300 76.800 73.440 76.940 ;
        RECT 57.570 76.740 57.890 76.800 ;
        RECT 56.650 76.600 57.890 76.740 ;
        RECT 56.650 76.540 56.970 76.600 ;
        RECT 57.570 76.540 57.890 76.600 ;
        RECT 59.425 76.740 59.715 76.785 ;
        RECT 60.330 76.740 60.650 76.800 ;
        RECT 59.425 76.600 60.650 76.740 ;
        RECT 59.425 76.555 59.715 76.600 ;
        RECT 60.330 76.540 60.650 76.600 ;
        RECT 62.630 76.540 62.950 76.800 ;
        RECT 63.090 76.540 63.410 76.800 ;
        RECT 64.930 76.740 65.250 76.800 ;
        RECT 68.165 76.740 68.455 76.785 ;
        RECT 64.930 76.600 68.455 76.740 ;
        RECT 64.930 76.540 65.250 76.600 ;
        RECT 68.165 76.555 68.455 76.600 ;
        RECT 69.070 76.740 69.390 76.800 ;
        RECT 71.385 76.740 71.675 76.785 ;
        RECT 71.830 76.740 72.150 76.800 ;
        RECT 69.070 76.600 72.150 76.740 ;
        RECT 69.070 76.540 69.390 76.600 ;
        RECT 71.385 76.555 71.675 76.600 ;
        RECT 71.830 76.540 72.150 76.600 ;
        RECT 73.210 76.540 73.530 76.800 ;
        RECT 5.520 75.920 83.260 76.400 ;
        RECT 7.890 75.720 8.210 75.780 ;
        RECT 10.205 75.720 10.495 75.765 ;
        RECT 7.890 75.580 10.495 75.720 ;
        RECT 7.890 75.520 8.210 75.580 ;
        RECT 10.205 75.535 10.495 75.580 ;
        RECT 12.030 75.720 12.350 75.780 ;
        RECT 12.965 75.720 13.255 75.765 ;
        RECT 12.030 75.580 13.255 75.720 ;
        RECT 12.030 75.520 12.350 75.580 ;
        RECT 12.965 75.535 13.255 75.580 ;
        RECT 18.470 75.720 18.790 75.780 ;
        RECT 24.450 75.720 24.770 75.780 ;
        RECT 18.470 75.580 24.770 75.720 ;
        RECT 18.470 75.520 18.790 75.580 ;
        RECT 24.450 75.520 24.770 75.580 ;
        RECT 28.590 75.520 28.910 75.780 ;
        RECT 30.890 75.520 31.210 75.780 ;
        RECT 34.570 75.720 34.890 75.780 ;
        RECT 31.900 75.580 34.890 75.720 ;
        RECT 25.385 75.380 25.675 75.425 ;
        RECT 27.210 75.380 27.530 75.440 ;
        RECT 25.385 75.240 27.530 75.380 ;
        RECT 25.385 75.195 25.675 75.240 ;
        RECT 27.210 75.180 27.530 75.240 ;
        RECT 29.065 75.380 29.355 75.425 ;
        RECT 31.900 75.380 32.040 75.580 ;
        RECT 34.570 75.520 34.890 75.580 ;
        RECT 39.185 75.720 39.475 75.765 ;
        RECT 41.470 75.720 41.790 75.780 ;
        RECT 39.185 75.580 41.790 75.720 ;
        RECT 39.185 75.535 39.475 75.580 ;
        RECT 41.470 75.520 41.790 75.580 ;
        RECT 47.925 75.720 48.215 75.765 ;
        RECT 49.290 75.720 49.610 75.780 ;
        RECT 52.985 75.720 53.275 75.765 ;
        RECT 53.430 75.720 53.750 75.780 ;
        RECT 47.925 75.580 49.610 75.720 ;
        RECT 47.925 75.535 48.215 75.580 ;
        RECT 49.290 75.520 49.610 75.580 ;
        RECT 49.840 75.580 53.750 75.720 ;
        RECT 44.690 75.380 45.010 75.440 ;
        RECT 49.840 75.425 49.980 75.580 ;
        RECT 52.985 75.535 53.275 75.580 ;
        RECT 53.430 75.520 53.750 75.580 ;
        RECT 53.890 75.520 54.210 75.780 ;
        RECT 54.350 75.520 54.670 75.780 ;
        RECT 55.270 75.720 55.590 75.780 ;
        RECT 58.950 75.720 59.270 75.780 ;
        RECT 55.270 75.580 59.270 75.720 ;
        RECT 55.270 75.520 55.590 75.580 ;
        RECT 58.950 75.520 59.270 75.580 ;
        RECT 60.345 75.720 60.635 75.765 ;
        RECT 63.105 75.720 63.395 75.765 ;
        RECT 60.345 75.580 63.395 75.720 ;
        RECT 60.345 75.535 60.635 75.580 ;
        RECT 63.105 75.535 63.395 75.580 ;
        RECT 70.925 75.720 71.215 75.765 ;
        RECT 70.925 75.580 81.260 75.720 ;
        RECT 70.925 75.535 71.215 75.580 ;
        RECT 29.065 75.240 32.040 75.380 ;
        RECT 32.360 75.240 40.780 75.380 ;
        RECT 29.065 75.195 29.355 75.240 ;
        RECT 9.745 75.040 10.035 75.085 ;
        RECT 10.190 75.040 10.510 75.100 ;
        RECT 9.745 74.900 10.510 75.040 ;
        RECT 9.745 74.855 10.035 74.900 ;
        RECT 10.190 74.840 10.510 74.900 ;
        RECT 10.650 74.840 10.970 75.100 ;
        RECT 12.490 74.840 12.810 75.100 ;
        RECT 13.425 75.040 13.715 75.085 ;
        RECT 23.530 75.040 23.850 75.100 ;
        RECT 13.425 74.900 23.850 75.040 ;
        RECT 13.425 74.855 13.715 74.900 ;
        RECT 23.530 74.840 23.850 74.900 ;
        RECT 25.830 75.040 26.150 75.100 ;
        RECT 26.305 75.040 26.595 75.085 ;
        RECT 25.830 74.900 26.595 75.040 ;
        RECT 25.830 74.840 26.150 74.900 ;
        RECT 26.305 74.855 26.595 74.900 ;
        RECT 27.670 74.840 27.990 75.100 ;
        RECT 26.765 74.700 27.055 74.745 ;
        RECT 29.140 74.700 29.280 75.195 ;
        RECT 29.970 74.840 30.290 75.100 ;
        RECT 32.360 75.085 32.500 75.240 ;
        RECT 40.640 75.100 40.780 75.240 ;
        RECT 44.690 75.240 49.520 75.380 ;
        RECT 44.690 75.180 45.010 75.240 ;
        RECT 32.285 74.855 32.575 75.085 ;
        RECT 33.565 75.040 33.855 75.085 ;
        RECT 32.820 74.900 33.855 75.040 ;
        RECT 26.765 74.560 29.280 74.700 ;
        RECT 31.810 74.700 32.130 74.760 ;
        RECT 32.820 74.700 32.960 74.900 ;
        RECT 33.565 74.855 33.855 74.900 ;
        RECT 40.550 75.040 40.870 75.100 ;
        RECT 49.380 75.085 49.520 75.240 ;
        RECT 49.765 75.195 50.055 75.425 ;
        RECT 50.225 75.380 50.515 75.425 ;
        RECT 52.510 75.380 52.830 75.440 ;
        RECT 53.980 75.380 54.120 75.520 ;
        RECT 50.225 75.240 54.120 75.380 ;
        RECT 54.440 75.380 54.580 75.520 ;
        RECT 81.120 75.440 81.260 75.580 ;
        RECT 57.110 75.380 57.430 75.440 ;
        RECT 54.440 75.240 55.960 75.380 ;
        RECT 50.225 75.195 50.515 75.240 ;
        RECT 52.510 75.180 52.830 75.240 ;
        RECT 41.025 75.040 41.315 75.085 ;
        RECT 40.550 74.900 41.315 75.040 ;
        RECT 40.550 74.840 40.870 74.900 ;
        RECT 41.025 74.855 41.315 74.900 ;
        RECT 42.360 75.040 42.650 75.085 ;
        RECT 48.385 75.040 48.675 75.085 ;
        RECT 42.360 74.900 48.675 75.040 ;
        RECT 42.360 74.855 42.650 74.900 ;
        RECT 48.385 74.855 48.675 74.900 ;
        RECT 49.305 74.855 49.595 75.085 ;
        RECT 50.815 75.040 51.105 75.085 ;
        RECT 50.760 74.855 51.105 75.040 ;
        RECT 52.065 74.855 52.355 75.085 ;
        RECT 31.810 74.560 32.960 74.700 ;
        RECT 33.165 74.700 33.455 74.745 ;
        RECT 34.355 74.700 34.645 74.745 ;
        RECT 36.875 74.700 37.165 74.745 ;
        RECT 33.165 74.560 37.165 74.700 ;
        RECT 26.765 74.515 27.055 74.560 ;
        RECT 31.810 74.500 32.130 74.560 ;
        RECT 33.165 74.515 33.455 74.560 ;
        RECT 34.355 74.515 34.645 74.560 ;
        RECT 36.875 74.515 37.165 74.560 ;
        RECT 41.905 74.700 42.195 74.745 ;
        RECT 43.095 74.700 43.385 74.745 ;
        RECT 45.615 74.700 45.905 74.745 ;
        RECT 41.905 74.560 45.905 74.700 ;
        RECT 41.905 74.515 42.195 74.560 ;
        RECT 43.095 74.515 43.385 74.560 ;
        RECT 45.615 74.515 45.905 74.560 ;
        RECT 46.070 74.700 46.390 74.760 ;
        RECT 50.760 74.700 50.900 74.855 ;
        RECT 46.070 74.560 50.900 74.700 ;
        RECT 51.605 74.700 51.895 74.745 ;
        RECT 52.140 74.700 52.280 74.855 ;
        RECT 52.970 74.840 53.290 75.100 ;
        RECT 53.445 75.040 53.735 75.085 ;
        RECT 53.890 75.040 54.210 75.100 ;
        RECT 53.445 74.900 54.210 75.040 ;
        RECT 53.445 74.855 53.735 74.900 ;
        RECT 53.890 74.840 54.210 74.900 ;
        RECT 54.365 74.855 54.655 75.085 ;
        RECT 54.825 74.855 55.115 75.085 ;
        RECT 54.440 74.700 54.580 74.855 ;
        RECT 51.605 74.560 52.280 74.700 ;
        RECT 52.600 74.560 54.580 74.700 ;
        RECT 46.070 74.500 46.390 74.560 ;
        RECT 51.605 74.515 51.895 74.560 ;
        RECT 32.770 74.360 33.060 74.405 ;
        RECT 34.870 74.360 35.160 74.405 ;
        RECT 36.440 74.360 36.730 74.405 ;
        RECT 32.770 74.220 36.730 74.360 ;
        RECT 32.770 74.175 33.060 74.220 ;
        RECT 34.870 74.175 35.160 74.220 ;
        RECT 36.440 74.175 36.730 74.220 ;
        RECT 41.510 74.360 41.800 74.405 ;
        RECT 43.610 74.360 43.900 74.405 ;
        RECT 45.180 74.360 45.470 74.405 ;
        RECT 41.510 74.220 45.470 74.360 ;
        RECT 41.510 74.175 41.800 74.220 ;
        RECT 43.610 74.175 43.900 74.220 ;
        RECT 45.180 74.175 45.470 74.220 ;
        RECT 49.290 74.360 49.610 74.420 ;
        RECT 50.670 74.360 50.990 74.420 ;
        RECT 51.680 74.360 51.820 74.515 ;
        RECT 49.290 74.220 51.820 74.360 ;
        RECT 52.050 74.360 52.370 74.420 ;
        RECT 52.600 74.360 52.740 74.560 ;
        RECT 52.050 74.220 52.740 74.360 ;
        RECT 54.350 74.360 54.670 74.420 ;
        RECT 54.900 74.360 55.040 74.855 ;
        RECT 55.270 74.840 55.590 75.100 ;
        RECT 55.820 75.040 55.960 75.240 ;
        RECT 57.110 75.240 72.520 75.380 ;
        RECT 57.110 75.180 57.430 75.240 ;
        RECT 72.380 75.100 72.520 75.240 ;
        RECT 73.760 75.240 77.580 75.380 ;
        RECT 73.760 75.100 73.900 75.240 ;
        RECT 57.585 75.040 57.875 75.085 ;
        RECT 55.820 74.900 57.875 75.040 ;
        RECT 57.585 74.855 57.875 74.900 ;
        RECT 58.490 74.840 58.810 75.100 ;
        RECT 58.950 74.840 59.270 75.100 ;
        RECT 59.425 75.040 59.715 75.085 ;
        RECT 61.710 75.040 62.030 75.100 ;
        RECT 59.425 74.900 62.030 75.040 ;
        RECT 59.425 74.855 59.715 74.900 ;
        RECT 58.030 74.700 58.350 74.760 ;
        RECT 59.500 74.700 59.640 74.855 ;
        RECT 61.710 74.840 62.030 74.900 ;
        RECT 62.645 75.040 62.935 75.085 ;
        RECT 64.945 75.040 65.235 75.085 ;
        RECT 62.645 74.900 65.235 75.040 ;
        RECT 62.645 74.855 62.935 74.900 ;
        RECT 64.945 74.855 65.235 74.900 ;
        RECT 70.005 75.040 70.295 75.085 ;
        RECT 70.450 75.040 70.770 75.100 ;
        RECT 70.005 74.900 70.770 75.040 ;
        RECT 70.005 74.855 70.295 74.900 ;
        RECT 70.450 74.840 70.770 74.900 ;
        RECT 72.290 75.040 72.610 75.100 ;
        RECT 73.225 75.040 73.515 75.085 ;
        RECT 72.290 74.900 73.515 75.040 ;
        RECT 72.290 74.840 72.610 74.900 ;
        RECT 73.225 74.855 73.515 74.900 ;
        RECT 58.030 74.560 59.640 74.700 ;
        RECT 60.330 74.700 60.650 74.760 ;
        RECT 60.330 74.560 62.860 74.700 ;
        RECT 58.030 74.500 58.350 74.560 ;
        RECT 60.330 74.500 60.650 74.560 ;
        RECT 54.350 74.220 55.040 74.360 ;
        RECT 56.665 74.360 56.955 74.405 ;
        RECT 62.170 74.360 62.490 74.420 ;
        RECT 56.665 74.220 62.490 74.360 ;
        RECT 62.720 74.360 62.860 74.560 ;
        RECT 63.565 74.515 63.855 74.745 ;
        RECT 66.310 74.700 66.630 74.760 ;
        RECT 67.705 74.700 67.995 74.745 ;
        RECT 66.310 74.560 67.995 74.700 ;
        RECT 63.640 74.360 63.780 74.515 ;
        RECT 66.310 74.500 66.630 74.560 ;
        RECT 67.705 74.515 67.995 74.560 ;
        RECT 69.070 74.500 69.390 74.760 ;
        RECT 62.720 74.220 63.780 74.360 ;
        RECT 73.300 74.360 73.440 74.855 ;
        RECT 73.670 74.840 73.990 75.100 ;
        RECT 74.145 74.855 74.435 75.085 ;
        RECT 74.220 74.700 74.360 74.855 ;
        RECT 75.050 74.840 75.370 75.100 ;
        RECT 76.890 74.840 77.210 75.100 ;
        RECT 77.440 75.085 77.580 75.240 ;
        RECT 81.030 75.180 81.350 75.440 ;
        RECT 77.365 74.855 77.655 75.085 ;
        RECT 77.825 75.040 78.115 75.085 ;
        RECT 78.270 75.040 78.590 75.100 ;
        RECT 77.825 74.900 78.590 75.040 ;
        RECT 77.825 74.855 78.115 74.900 ;
        RECT 78.270 74.840 78.590 74.900 ;
        RECT 78.745 75.040 79.035 75.085 ;
        RECT 79.650 75.040 79.970 75.100 ;
        RECT 78.745 74.900 79.970 75.040 ;
        RECT 78.745 74.855 79.035 74.900 ;
        RECT 79.650 74.840 79.970 74.900 ;
        RECT 80.110 74.840 80.430 75.100 ;
        RECT 79.205 74.700 79.495 74.745 ;
        RECT 74.220 74.560 79.495 74.700 ;
        RECT 79.205 74.515 79.495 74.560 ;
        RECT 74.130 74.360 74.450 74.420 ;
        RECT 73.300 74.220 74.450 74.360 ;
        RECT 49.290 74.160 49.610 74.220 ;
        RECT 50.670 74.160 50.990 74.220 ;
        RECT 52.050 74.160 52.370 74.220 ;
        RECT 54.350 74.160 54.670 74.220 ;
        RECT 56.665 74.175 56.955 74.220 ;
        RECT 62.170 74.160 62.490 74.220 ;
        RECT 74.130 74.160 74.450 74.220 ;
        RECT 75.050 74.360 75.370 74.420 ;
        RECT 79.650 74.360 79.970 74.420 ;
        RECT 75.050 74.220 79.970 74.360 ;
        RECT 75.050 74.160 75.370 74.220 ;
        RECT 79.650 74.160 79.970 74.220 ;
        RECT 23.530 74.020 23.850 74.080 ;
        RECT 24.465 74.020 24.755 74.065 ;
        RECT 23.530 73.880 24.755 74.020 ;
        RECT 23.530 73.820 23.850 73.880 ;
        RECT 24.465 73.835 24.755 73.880 ;
        RECT 47.450 74.020 47.770 74.080 ;
        RECT 52.970 74.020 53.290 74.080 ;
        RECT 47.450 73.880 53.290 74.020 ;
        RECT 47.450 73.820 47.770 73.880 ;
        RECT 52.970 73.820 53.290 73.880 ;
        RECT 60.790 73.820 61.110 74.080 ;
        RECT 61.710 74.020 62.030 74.080 ;
        RECT 68.610 74.020 68.930 74.080 ;
        RECT 61.710 73.880 68.930 74.020 ;
        RECT 61.710 73.820 62.030 73.880 ;
        RECT 68.610 73.820 68.930 73.880 ;
        RECT 71.845 74.020 72.135 74.065 ;
        RECT 73.670 74.020 73.990 74.080 ;
        RECT 71.845 73.880 73.990 74.020 ;
        RECT 71.845 73.835 72.135 73.880 ;
        RECT 73.670 73.820 73.990 73.880 ;
        RECT 75.510 73.820 75.830 74.080 ;
        RECT 5.520 73.200 83.260 73.680 ;
        RECT 28.130 72.800 28.450 73.060 ;
        RECT 52.065 73.000 52.355 73.045 ;
        RECT 52.510 73.000 52.830 73.060 ;
        RECT 52.065 72.860 52.830 73.000 ;
        RECT 52.065 72.815 52.355 72.860 ;
        RECT 52.510 72.800 52.830 72.860 ;
        RECT 53.445 72.815 53.735 73.045 ;
        RECT 53.890 73.000 54.210 73.060 ;
        RECT 55.285 73.000 55.575 73.045 ;
        RECT 68.165 73.000 68.455 73.045 ;
        RECT 53.890 72.860 55.575 73.000 ;
        RECT 31.350 72.460 31.670 72.720 ;
        RECT 43.770 72.460 44.090 72.720 ;
        RECT 45.150 72.660 45.470 72.720 ;
        RECT 47.450 72.660 47.770 72.720 ;
        RECT 48.370 72.660 48.690 72.720 ;
        RECT 50.225 72.660 50.515 72.705 ;
        RECT 45.150 72.520 48.140 72.660 ;
        RECT 45.150 72.460 45.470 72.520 ;
        RECT 47.450 72.460 47.770 72.520 ;
        RECT 20.310 72.320 20.630 72.380 ;
        RECT 21.245 72.320 21.535 72.365 ;
        RECT 20.310 72.180 21.535 72.320 ;
        RECT 20.310 72.120 20.630 72.180 ;
        RECT 21.245 72.135 21.535 72.180 ;
        RECT 24.450 72.320 24.770 72.380 ;
        RECT 28.605 72.320 28.895 72.365 ;
        RECT 31.440 72.320 31.580 72.460 ;
        RECT 34.570 72.320 34.890 72.380 ;
        RECT 35.950 72.320 36.270 72.380 ;
        RECT 24.450 72.180 31.580 72.320 ;
        RECT 32.360 72.180 36.270 72.320 ;
        RECT 24.450 72.120 24.770 72.180 ;
        RECT 28.605 72.135 28.895 72.180 ;
        RECT 16.630 71.780 16.950 72.040 ;
        RECT 21.690 71.980 22.010 72.040 ;
        RECT 22.165 71.980 22.455 72.025 ;
        RECT 21.690 71.840 22.455 71.980 ;
        RECT 21.690 71.780 22.010 71.840 ;
        RECT 22.165 71.795 22.455 71.840 ;
        RECT 22.625 71.980 22.915 72.025 ;
        RECT 23.070 71.980 23.390 72.040 ;
        RECT 22.625 71.840 23.390 71.980 ;
        RECT 22.625 71.795 22.915 71.840 ;
        RECT 23.070 71.780 23.390 71.840 ;
        RECT 25.385 71.980 25.675 72.025 ;
        RECT 26.290 71.980 26.610 72.040 ;
        RECT 25.385 71.840 26.610 71.980 ;
        RECT 25.385 71.795 25.675 71.840 ;
        RECT 26.290 71.780 26.610 71.840 ;
        RECT 27.210 71.780 27.530 72.040 ;
        RECT 29.985 71.980 30.275 72.025 ;
        RECT 30.430 71.980 30.750 72.040 ;
        RECT 29.985 71.840 30.750 71.980 ;
        RECT 29.985 71.795 30.275 71.840 ;
        RECT 30.430 71.780 30.750 71.840 ;
        RECT 30.890 71.780 31.210 72.040 ;
        RECT 31.365 71.980 31.655 72.025 ;
        RECT 31.810 71.980 32.130 72.040 ;
        RECT 32.360 72.025 32.500 72.180 ;
        RECT 34.570 72.120 34.890 72.180 ;
        RECT 35.950 72.120 36.270 72.180 ;
        RECT 46.070 72.320 46.390 72.380 ;
        RECT 48.000 72.365 48.140 72.520 ;
        RECT 48.370 72.520 50.515 72.660 ;
        RECT 48.370 72.460 48.690 72.520 ;
        RECT 50.225 72.475 50.515 72.520 ;
        RECT 52.970 72.460 53.290 72.720 ;
        RECT 53.520 72.660 53.660 72.815 ;
        RECT 53.890 72.800 54.210 72.860 ;
        RECT 55.285 72.815 55.575 72.860 ;
        RECT 55.820 72.860 68.455 73.000 ;
        RECT 53.520 72.520 55.500 72.660 ;
        RECT 55.360 72.380 55.500 72.520 ;
        RECT 47.005 72.320 47.295 72.365 ;
        RECT 46.070 72.180 47.295 72.320 ;
        RECT 46.070 72.120 46.390 72.180 ;
        RECT 47.005 72.135 47.295 72.180 ;
        RECT 47.925 72.135 48.215 72.365 ;
        RECT 49.750 72.320 50.070 72.380 ;
        RECT 53.905 72.320 54.195 72.365 ;
        RECT 49.750 72.180 54.195 72.320 ;
        RECT 49.750 72.120 50.070 72.180 ;
        RECT 53.905 72.135 54.195 72.180 ;
        RECT 55.270 72.120 55.590 72.380 ;
        RECT 31.365 71.840 32.130 71.980 ;
        RECT 31.365 71.795 31.655 71.840 ;
        RECT 31.810 71.780 32.130 71.840 ;
        RECT 32.285 71.795 32.575 72.025 ;
        RECT 33.665 71.795 33.955 72.025 ;
        RECT 39.185 71.980 39.475 72.025 ;
        RECT 40.090 71.980 40.410 72.040 ;
        RECT 39.185 71.840 40.410 71.980 ;
        RECT 39.185 71.795 39.475 71.840 ;
        RECT 23.990 71.640 24.310 71.700 ;
        RECT 33.740 71.640 33.880 71.795 ;
        RECT 40.090 71.780 40.410 71.840 ;
        RECT 40.565 71.795 40.855 72.025 ;
        RECT 36.410 71.640 36.730 71.700 ;
        RECT 23.990 71.500 36.730 71.640 ;
        RECT 40.640 71.640 40.780 71.795 ;
        RECT 41.470 71.780 41.790 72.040 ;
        RECT 42.850 71.780 43.170 72.040 ;
        RECT 44.690 71.980 45.010 72.040 ;
        RECT 55.820 72.025 55.960 72.860 ;
        RECT 68.165 72.815 68.455 72.860 ;
        RECT 71.385 73.000 71.675 73.045 ;
        RECT 75.970 73.000 76.290 73.060 ;
        RECT 78.270 73.000 78.590 73.060 ;
        RECT 81.505 73.000 81.795 73.045 ;
        RECT 71.385 72.860 77.120 73.000 ;
        RECT 71.385 72.815 71.675 72.860 ;
        RECT 75.970 72.800 76.290 72.860 ;
        RECT 56.650 72.660 56.970 72.720 ;
        RECT 56.280 72.520 56.970 72.660 ;
        RECT 46.545 71.980 46.835 72.025 ;
        RECT 44.690 71.840 46.835 71.980 ;
        RECT 44.690 71.780 45.010 71.840 ;
        RECT 46.545 71.795 46.835 71.840 ;
        RECT 53.445 71.795 53.735 72.025 ;
        RECT 55.745 71.795 56.035 72.025 ;
        RECT 41.930 71.640 42.250 71.700 ;
        RECT 40.640 71.500 42.250 71.640 ;
        RECT 53.520 71.640 53.660 71.795 ;
        RECT 56.280 71.640 56.420 72.520 ;
        RECT 56.650 72.460 56.970 72.520 ;
        RECT 59.450 72.660 59.740 72.705 ;
        RECT 61.550 72.660 61.840 72.705 ;
        RECT 63.120 72.660 63.410 72.705 ;
        RECT 59.450 72.520 63.410 72.660 ;
        RECT 59.450 72.475 59.740 72.520 ;
        RECT 61.550 72.475 61.840 72.520 ;
        RECT 63.120 72.475 63.410 72.520 ;
        RECT 69.990 72.660 70.310 72.720 ;
        RECT 70.925 72.660 71.215 72.705 ;
        RECT 69.990 72.520 71.215 72.660 ;
        RECT 69.990 72.460 70.310 72.520 ;
        RECT 70.925 72.475 71.215 72.520 ;
        RECT 72.790 72.660 73.080 72.705 ;
        RECT 74.890 72.660 75.180 72.705 ;
        RECT 76.460 72.660 76.750 72.705 ;
        RECT 72.790 72.520 76.750 72.660 ;
        RECT 76.980 72.660 77.120 72.860 ;
        RECT 78.270 72.860 81.795 73.000 ;
        RECT 78.270 72.800 78.590 72.860 ;
        RECT 81.505 72.815 81.795 72.860 ;
        RECT 80.570 72.660 80.890 72.720 ;
        RECT 76.980 72.520 80.890 72.660 ;
        RECT 72.790 72.475 73.080 72.520 ;
        RECT 74.890 72.475 75.180 72.520 ;
        RECT 76.460 72.475 76.750 72.520 ;
        RECT 80.570 72.460 80.890 72.520 ;
        RECT 58.490 72.320 58.810 72.380 ;
        RECT 56.740 72.180 58.810 72.320 ;
        RECT 56.740 72.025 56.880 72.180 ;
        RECT 58.490 72.120 58.810 72.180 ;
        RECT 59.845 72.320 60.135 72.365 ;
        RECT 61.035 72.320 61.325 72.365 ;
        RECT 63.555 72.320 63.845 72.365 ;
        RECT 59.845 72.180 63.845 72.320 ;
        RECT 59.845 72.135 60.135 72.180 ;
        RECT 61.035 72.135 61.325 72.180 ;
        RECT 63.555 72.135 63.845 72.180 ;
        RECT 66.770 72.320 67.090 72.380 ;
        RECT 69.530 72.320 69.850 72.380 ;
        RECT 73.185 72.320 73.475 72.365 ;
        RECT 74.375 72.320 74.665 72.365 ;
        RECT 76.895 72.320 77.185 72.365 ;
        RECT 66.770 72.180 69.300 72.320 ;
        RECT 66.770 72.120 67.090 72.180 ;
        RECT 56.665 71.795 56.955 72.025 ;
        RECT 57.110 71.780 57.430 72.040 ;
        RECT 57.585 71.980 57.875 72.025 ;
        RECT 58.030 71.980 58.350 72.040 ;
        RECT 57.585 71.840 58.350 71.980 ;
        RECT 57.585 71.795 57.875 71.840 ;
        RECT 58.030 71.780 58.350 71.840 ;
        RECT 58.965 71.980 59.255 72.025 ;
        RECT 59.410 71.980 59.730 72.040 ;
        RECT 66.325 71.980 66.615 72.025 ;
        RECT 68.625 71.980 68.915 72.025 ;
        RECT 58.965 71.840 59.730 71.980 ;
        RECT 58.965 71.795 59.255 71.840 ;
        RECT 59.410 71.780 59.730 71.840 ;
        RECT 59.960 71.840 66.615 71.980 ;
        RECT 59.960 71.640 60.100 71.840 ;
        RECT 66.325 71.795 66.615 71.840 ;
        RECT 67.780 71.840 68.915 71.980 ;
        RECT 69.160 71.980 69.300 72.180 ;
        RECT 69.530 72.180 72.060 72.320 ;
        RECT 69.530 72.120 69.850 72.180 ;
        RECT 69.160 71.950 70.220 71.980 ;
        RECT 70.410 71.950 70.700 71.995 ;
        RECT 69.160 71.840 70.700 71.950 ;
        RECT 53.520 71.500 56.420 71.640 ;
        RECT 58.120 71.500 60.100 71.640 ;
        RECT 60.300 71.640 60.590 71.685 ;
        RECT 60.790 71.640 61.110 71.700 ;
        RECT 60.300 71.500 61.110 71.640 ;
        RECT 23.990 71.440 24.310 71.500 ;
        RECT 36.410 71.440 36.730 71.500 ;
        RECT 41.930 71.440 42.250 71.500 ;
        RECT 17.090 71.100 17.410 71.360 ;
        RECT 21.230 71.300 21.550 71.360 ;
        RECT 22.625 71.300 22.915 71.345 ;
        RECT 21.230 71.160 22.915 71.300 ;
        RECT 21.230 71.100 21.550 71.160 ;
        RECT 22.625 71.115 22.915 71.160 ;
        RECT 23.070 71.300 23.390 71.360 ;
        RECT 25.830 71.300 26.150 71.360 ;
        RECT 23.070 71.160 26.150 71.300 ;
        RECT 23.070 71.100 23.390 71.160 ;
        RECT 25.830 71.100 26.150 71.160 ;
        RECT 26.305 71.300 26.595 71.345 ;
        RECT 27.670 71.300 27.990 71.360 ;
        RECT 26.305 71.160 27.990 71.300 ;
        RECT 26.305 71.115 26.595 71.160 ;
        RECT 27.670 71.100 27.990 71.160 ;
        RECT 28.130 71.300 28.450 71.360 ;
        RECT 29.065 71.300 29.355 71.345 ;
        RECT 28.130 71.160 29.355 71.300 ;
        RECT 28.130 71.100 28.450 71.160 ;
        RECT 29.065 71.115 29.355 71.160 ;
        RECT 29.970 71.300 30.290 71.360 ;
        RECT 32.745 71.300 33.035 71.345 ;
        RECT 29.970 71.160 33.035 71.300 ;
        RECT 29.970 71.100 30.290 71.160 ;
        RECT 32.745 71.115 33.035 71.160 ;
        RECT 34.570 71.100 34.890 71.360 ;
        RECT 41.470 71.300 41.790 71.360 ;
        RECT 44.705 71.300 44.995 71.345 ;
        RECT 41.470 71.160 44.995 71.300 ;
        RECT 41.470 71.100 41.790 71.160 ;
        RECT 44.705 71.115 44.995 71.160 ;
        RECT 52.065 71.300 52.355 71.345 ;
        RECT 53.430 71.300 53.750 71.360 ;
        RECT 52.065 71.160 53.750 71.300 ;
        RECT 52.065 71.115 52.355 71.160 ;
        RECT 53.430 71.100 53.750 71.160 ;
        RECT 55.270 71.300 55.590 71.360 ;
        RECT 58.120 71.300 58.260 71.500 ;
        RECT 60.300 71.455 60.590 71.500 ;
        RECT 60.790 71.440 61.110 71.500 ;
        RECT 64.470 71.640 64.790 71.700 ;
        RECT 67.245 71.640 67.535 71.685 ;
        RECT 64.470 71.500 67.535 71.640 ;
        RECT 64.470 71.440 64.790 71.500 ;
        RECT 67.245 71.455 67.535 71.500 ;
        RECT 55.270 71.160 58.260 71.300 ;
        RECT 58.505 71.300 58.795 71.345 ;
        RECT 64.010 71.300 64.330 71.360 ;
        RECT 58.505 71.160 64.330 71.300 ;
        RECT 55.270 71.100 55.590 71.160 ;
        RECT 58.505 71.115 58.795 71.160 ;
        RECT 64.010 71.100 64.330 71.160 ;
        RECT 65.865 71.300 66.155 71.345 ;
        RECT 66.310 71.300 66.630 71.360 ;
        RECT 65.865 71.160 66.630 71.300 ;
        RECT 65.865 71.115 66.155 71.160 ;
        RECT 66.310 71.100 66.630 71.160 ;
        RECT 66.770 71.300 67.090 71.360 ;
        RECT 67.780 71.300 67.920 71.840 ;
        RECT 68.625 71.795 68.915 71.840 ;
        RECT 70.080 71.810 70.700 71.840 ;
        RECT 70.410 71.765 70.700 71.810 ;
        RECT 71.920 71.685 72.060 72.180 ;
        RECT 73.185 72.180 77.185 72.320 ;
        RECT 73.185 72.135 73.475 72.180 ;
        RECT 74.375 72.135 74.665 72.180 ;
        RECT 76.895 72.135 77.185 72.180 ;
        RECT 72.305 71.980 72.595 72.025 ;
        RECT 72.750 71.980 73.070 72.040 ;
        RECT 73.670 72.025 73.990 72.040 ;
        RECT 73.640 71.980 73.990 72.025 ;
        RECT 72.305 71.840 73.070 71.980 ;
        RECT 73.475 71.840 73.990 71.980 ;
        RECT 72.305 71.795 72.595 71.840 ;
        RECT 72.750 71.780 73.070 71.840 ;
        RECT 73.640 71.795 73.990 71.840 ;
        RECT 73.670 71.780 73.990 71.795 ;
        RECT 78.270 71.980 78.590 72.040 ;
        RECT 80.585 71.980 80.875 72.025 ;
        RECT 78.270 71.840 80.875 71.980 ;
        RECT 78.270 71.780 78.590 71.840 ;
        RECT 80.585 71.795 80.875 71.840 ;
        RECT 71.845 71.640 72.135 71.685 ;
        RECT 76.430 71.640 76.750 71.700 ;
        RECT 71.845 71.500 76.750 71.640 ;
        RECT 71.845 71.455 72.135 71.500 ;
        RECT 76.430 71.440 76.750 71.500 ;
        RECT 79.665 71.640 79.955 71.685 ;
        RECT 81.030 71.640 81.350 71.700 ;
        RECT 79.665 71.500 81.350 71.640 ;
        RECT 79.665 71.455 79.955 71.500 ;
        RECT 81.030 71.440 81.350 71.500 ;
        RECT 66.770 71.160 67.920 71.300 ;
        RECT 69.070 71.300 69.390 71.360 ;
        RECT 74.590 71.300 74.910 71.360 ;
        RECT 69.070 71.160 74.910 71.300 ;
        RECT 66.770 71.100 67.090 71.160 ;
        RECT 69.070 71.100 69.390 71.160 ;
        RECT 74.590 71.100 74.910 71.160 ;
        RECT 79.205 71.300 79.495 71.345 ;
        RECT 80.110 71.300 80.430 71.360 ;
        RECT 79.205 71.160 80.430 71.300 ;
        RECT 79.205 71.115 79.495 71.160 ;
        RECT 80.110 71.100 80.430 71.160 ;
        RECT 5.520 70.480 83.260 70.960 ;
        RECT 14.330 70.280 14.650 70.340 ;
        RECT 15.710 70.280 16.030 70.340 ;
        RECT 23.085 70.280 23.375 70.325 ;
        RECT 25.830 70.280 26.150 70.340 ;
        RECT 27.210 70.280 27.530 70.340 ;
        RECT 14.330 70.140 21.920 70.280 ;
        RECT 14.330 70.080 14.650 70.140 ;
        RECT 15.710 70.080 16.030 70.140 ;
        RECT 18.485 69.940 18.775 69.985 ;
        RECT 18.930 69.940 19.250 70.000 ;
        RECT 18.485 69.800 19.250 69.940 ;
        RECT 18.485 69.755 18.775 69.800 ;
        RECT 18.930 69.740 19.250 69.800 ;
        RECT 19.635 69.770 19.925 69.815 ;
        RECT 9.285 69.415 9.575 69.645 ;
        RECT 9.360 69.260 9.500 69.415 ;
        RECT 10.190 69.400 10.510 69.660 ;
        RECT 17.105 69.415 17.395 69.645 ;
        RECT 12.030 69.260 12.350 69.320 ;
        RECT 9.360 69.120 12.350 69.260 ;
        RECT 17.180 69.260 17.320 69.415 ;
        RECT 18.010 69.400 18.330 69.660 ;
        RECT 19.610 69.600 19.925 69.770 ;
        RECT 21.230 69.600 21.550 69.660 ;
        RECT 21.780 69.645 21.920 70.140 ;
        RECT 23.085 70.140 27.530 70.280 ;
        RECT 23.085 70.095 23.375 70.140 ;
        RECT 25.830 70.080 26.150 70.140 ;
        RECT 27.210 70.080 27.530 70.140 ;
        RECT 34.585 70.280 34.875 70.325 ;
        RECT 35.490 70.280 35.810 70.340 ;
        RECT 34.585 70.140 35.810 70.280 ;
        RECT 34.585 70.095 34.875 70.140 ;
        RECT 35.490 70.080 35.810 70.140 ;
        RECT 45.610 70.280 45.930 70.340 ;
        RECT 47.005 70.280 47.295 70.325 ;
        RECT 45.610 70.140 47.295 70.280 ;
        RECT 45.610 70.080 45.930 70.140 ;
        RECT 47.005 70.095 47.295 70.140 ;
        RECT 48.845 70.280 49.135 70.325 ;
        RECT 52.510 70.280 52.830 70.340 ;
        RECT 48.845 70.140 52.830 70.280 ;
        RECT 48.845 70.095 49.135 70.140 ;
        RECT 52.510 70.080 52.830 70.140 ;
        RECT 53.905 70.280 54.195 70.325 ;
        RECT 55.270 70.280 55.590 70.340 ;
        RECT 53.905 70.140 55.590 70.280 ;
        RECT 53.905 70.095 54.195 70.140 ;
        RECT 55.270 70.080 55.590 70.140 ;
        RECT 64.010 70.080 64.330 70.340 ;
        RECT 70.910 70.080 71.230 70.340 ;
        RECT 72.305 70.280 72.595 70.325 ;
        RECT 75.970 70.280 76.290 70.340 ;
        RECT 72.305 70.140 76.290 70.280 ;
        RECT 72.305 70.095 72.595 70.140 ;
        RECT 75.970 70.080 76.290 70.140 ;
        RECT 81.030 70.080 81.350 70.340 ;
        RECT 40.550 69.940 40.870 70.000 ;
        RECT 51.130 69.940 51.450 70.000 ;
        RECT 22.700 69.800 29.280 69.940 ;
        RECT 19.610 69.460 21.550 69.600 ;
        RECT 21.230 69.400 21.550 69.460 ;
        RECT 21.705 69.600 21.995 69.645 ;
        RECT 22.150 69.600 22.470 69.660 ;
        RECT 22.700 69.645 22.840 69.800 ;
        RECT 21.705 69.460 22.470 69.600 ;
        RECT 21.705 69.415 21.995 69.460 ;
        RECT 22.150 69.400 22.470 69.460 ;
        RECT 22.625 69.415 22.915 69.645 ;
        RECT 25.830 69.600 26.150 69.660 ;
        RECT 23.620 69.460 26.150 69.600 ;
        RECT 20.310 69.260 20.630 69.320 ;
        RECT 17.180 69.120 20.630 69.260 ;
        RECT 12.030 69.060 12.350 69.120 ;
        RECT 20.310 69.060 20.630 69.120 ;
        RECT 20.785 69.260 21.075 69.305 ;
        RECT 23.620 69.260 23.760 69.460 ;
        RECT 25.830 69.400 26.150 69.460 ;
        RECT 28.590 69.645 28.910 69.660 ;
        RECT 28.590 69.415 28.940 69.645 ;
        RECT 29.140 69.600 29.280 69.800 ;
        RECT 30.060 69.800 39.400 69.940 ;
        RECT 30.060 69.645 30.200 69.800 ;
        RECT 29.140 69.460 29.740 69.600 ;
        RECT 28.590 69.400 28.910 69.415 ;
        RECT 20.785 69.120 23.760 69.260 ;
        RECT 25.395 69.260 25.685 69.305 ;
        RECT 27.915 69.260 28.205 69.305 ;
        RECT 29.105 69.260 29.395 69.305 ;
        RECT 25.395 69.120 29.395 69.260 ;
        RECT 29.600 69.260 29.740 69.460 ;
        RECT 29.985 69.415 30.275 69.645 ;
        RECT 31.825 69.600 32.115 69.645 ;
        RECT 34.110 69.600 34.430 69.660 ;
        RECT 31.825 69.460 34.430 69.600 ;
        RECT 31.825 69.415 32.115 69.460 ;
        RECT 34.110 69.400 34.430 69.460 ;
        RECT 34.570 69.400 34.890 69.660 ;
        RECT 35.030 69.400 35.350 69.660 ;
        RECT 39.260 69.645 39.400 69.800 ;
        RECT 40.550 69.800 51.450 69.940 ;
        RECT 40.550 69.740 40.870 69.800 ;
        RECT 51.130 69.740 51.450 69.800 ;
        RECT 66.310 69.940 66.630 70.000 ;
        RECT 74.100 69.940 74.390 69.985 ;
        RECT 75.510 69.940 75.830 70.000 ;
        RECT 66.310 69.800 71.600 69.940 ;
        RECT 66.310 69.740 66.630 69.800 ;
        RECT 39.185 69.600 39.475 69.645 ;
        RECT 40.090 69.600 40.410 69.660 ;
        RECT 41.470 69.645 41.790 69.660 ;
        RECT 41.440 69.600 41.790 69.645 ;
        RECT 39.185 69.460 40.410 69.600 ;
        RECT 41.275 69.460 41.790 69.600 ;
        RECT 39.185 69.415 39.475 69.460 ;
        RECT 40.090 69.400 40.410 69.460 ;
        RECT 41.440 69.415 41.790 69.460 ;
        RECT 41.470 69.400 41.790 69.415 ;
        RECT 47.450 69.600 47.770 69.660 ;
        RECT 49.765 69.600 50.055 69.645 ;
        RECT 47.450 69.460 50.055 69.600 ;
        RECT 47.450 69.400 47.770 69.460 ;
        RECT 49.765 69.415 50.055 69.460 ;
        RECT 40.985 69.260 41.275 69.305 ;
        RECT 42.175 69.260 42.465 69.305 ;
        RECT 44.695 69.260 44.985 69.305 ;
        RECT 29.600 69.120 33.880 69.260 ;
        RECT 20.785 69.075 21.075 69.120 ;
        RECT 25.395 69.075 25.685 69.120 ;
        RECT 27.915 69.075 28.205 69.120 ;
        RECT 29.105 69.075 29.395 69.120 ;
        RECT 18.010 68.920 18.330 68.980 ;
        RECT 21.690 68.920 22.010 68.980 ;
        RECT 24.450 68.920 24.770 68.980 ;
        RECT 18.010 68.780 24.770 68.920 ;
        RECT 18.010 68.720 18.330 68.780 ;
        RECT 21.690 68.720 22.010 68.780 ;
        RECT 24.450 68.720 24.770 68.780 ;
        RECT 25.830 68.920 26.120 68.965 ;
        RECT 27.400 68.920 27.690 68.965 ;
        RECT 29.500 68.920 29.790 68.965 ;
        RECT 25.830 68.780 29.790 68.920 ;
        RECT 25.830 68.735 26.120 68.780 ;
        RECT 27.400 68.735 27.690 68.780 ;
        RECT 29.500 68.735 29.790 68.780 ;
        RECT 33.190 68.720 33.510 68.980 ;
        RECT 33.740 68.965 33.880 69.120 ;
        RECT 40.985 69.120 44.985 69.260 ;
        RECT 49.840 69.260 49.980 69.415 ;
        RECT 50.670 69.400 50.990 69.660 ;
        RECT 52.970 69.400 53.290 69.660 ;
        RECT 54.825 69.600 55.115 69.645 ;
        RECT 56.190 69.600 56.510 69.660 ;
        RECT 53.520 69.460 56.510 69.600 ;
        RECT 52.065 69.260 52.355 69.305 ;
        RECT 49.840 69.120 52.355 69.260 ;
        RECT 40.985 69.075 41.275 69.120 ;
        RECT 42.175 69.075 42.465 69.120 ;
        RECT 44.695 69.075 44.985 69.120 ;
        RECT 52.065 69.075 52.355 69.120 ;
        RECT 52.510 69.260 52.830 69.320 ;
        RECT 53.520 69.260 53.660 69.460 ;
        RECT 54.825 69.415 55.115 69.460 ;
        RECT 56.190 69.400 56.510 69.460 ;
        RECT 56.665 69.600 56.955 69.645 ;
        RECT 60.330 69.600 60.650 69.660 ;
        RECT 56.665 69.460 60.650 69.600 ;
        RECT 56.665 69.415 56.955 69.460 ;
        RECT 60.330 69.400 60.650 69.460 ;
        RECT 63.565 69.600 63.855 69.645 ;
        RECT 65.865 69.600 66.155 69.645 ;
        RECT 63.565 69.460 66.155 69.600 ;
        RECT 63.565 69.415 63.855 69.460 ;
        RECT 65.865 69.415 66.155 69.460 ;
        RECT 69.530 69.400 69.850 69.660 ;
        RECT 71.460 69.645 71.600 69.800 ;
        RECT 74.100 69.800 75.830 69.940 ;
        RECT 74.100 69.755 74.390 69.800 ;
        RECT 75.510 69.740 75.830 69.800 ;
        RECT 70.925 69.415 71.215 69.645 ;
        RECT 71.385 69.415 71.675 69.645 ;
        RECT 52.510 69.120 53.660 69.260 ;
        RECT 53.890 69.260 54.210 69.320 ;
        RECT 57.585 69.260 57.875 69.305 ;
        RECT 53.890 69.120 57.875 69.260 ;
        RECT 52.510 69.060 52.830 69.120 ;
        RECT 53.890 69.060 54.210 69.120 ;
        RECT 57.585 69.075 57.875 69.120 ;
        RECT 62.170 69.260 62.490 69.320 ;
        RECT 64.485 69.260 64.775 69.305 ;
        RECT 62.170 69.120 64.775 69.260 ;
        RECT 62.170 69.060 62.490 69.120 ;
        RECT 64.485 69.075 64.775 69.120 ;
        RECT 69.070 69.060 69.390 69.320 ;
        RECT 71.000 69.260 71.140 69.415 ;
        RECT 80.110 69.400 80.430 69.660 ;
        RECT 71.830 69.260 72.150 69.320 ;
        RECT 71.000 69.120 72.150 69.260 ;
        RECT 71.830 69.060 72.150 69.120 ;
        RECT 72.750 69.060 73.070 69.320 ;
        RECT 73.645 69.260 73.935 69.305 ;
        RECT 74.835 69.260 75.125 69.305 ;
        RECT 77.355 69.260 77.645 69.305 ;
        RECT 73.645 69.120 77.645 69.260 ;
        RECT 73.645 69.075 73.935 69.120 ;
        RECT 74.835 69.075 75.125 69.120 ;
        RECT 77.355 69.075 77.645 69.120 ;
        RECT 33.665 68.735 33.955 68.965 ;
        RECT 40.590 68.920 40.880 68.965 ;
        RECT 42.690 68.920 42.980 68.965 ;
        RECT 44.260 68.920 44.550 68.965 ;
        RECT 40.590 68.780 44.550 68.920 ;
        RECT 40.590 68.735 40.880 68.780 ;
        RECT 42.690 68.735 42.980 68.780 ;
        RECT 44.260 68.735 44.550 68.780 ;
        RECT 69.990 68.920 70.310 68.980 ;
        RECT 70.465 68.920 70.755 68.965 ;
        RECT 69.990 68.780 70.755 68.920 ;
        RECT 69.990 68.720 70.310 68.780 ;
        RECT 70.465 68.735 70.755 68.780 ;
        RECT 73.250 68.920 73.540 68.965 ;
        RECT 75.350 68.920 75.640 68.965 ;
        RECT 76.920 68.920 77.210 68.965 ;
        RECT 73.250 68.780 77.210 68.920 ;
        RECT 73.250 68.735 73.540 68.780 ;
        RECT 75.350 68.735 75.640 68.780 ;
        RECT 76.920 68.735 77.210 68.780 ;
        RECT 9.730 68.380 10.050 68.640 ;
        RECT 17.565 68.580 17.855 68.625 ;
        RECT 18.470 68.580 18.790 68.640 ;
        RECT 17.565 68.440 18.790 68.580 ;
        RECT 17.565 68.395 17.855 68.440 ;
        RECT 18.470 68.380 18.790 68.440 ;
        RECT 19.405 68.580 19.695 68.625 ;
        RECT 19.850 68.580 20.170 68.640 ;
        RECT 19.405 68.440 20.170 68.580 ;
        RECT 19.405 68.395 19.695 68.440 ;
        RECT 19.850 68.380 20.170 68.440 ;
        RECT 20.310 68.380 20.630 68.640 ;
        RECT 22.150 68.580 22.470 68.640 ;
        RECT 26.750 68.580 27.070 68.640 ;
        RECT 22.150 68.440 27.070 68.580 ;
        RECT 22.150 68.380 22.470 68.440 ;
        RECT 26.750 68.380 27.070 68.440 ;
        RECT 29.050 68.580 29.370 68.640 ;
        RECT 32.515 68.580 32.805 68.625 ;
        RECT 29.050 68.440 32.805 68.580 ;
        RECT 29.050 68.380 29.370 68.440 ;
        RECT 32.515 68.395 32.805 68.440 ;
        RECT 60.790 68.380 61.110 68.640 ;
        RECT 61.250 68.580 61.570 68.640 ;
        RECT 61.725 68.580 62.015 68.625 ;
        RECT 61.250 68.440 62.015 68.580 ;
        RECT 61.250 68.380 61.570 68.440 ;
        RECT 61.725 68.395 62.015 68.440 ;
        RECT 78.270 68.580 78.590 68.640 ;
        RECT 79.665 68.580 79.955 68.625 ;
        RECT 78.270 68.440 79.955 68.580 ;
        RECT 78.270 68.380 78.590 68.440 ;
        RECT 79.665 68.395 79.955 68.440 ;
        RECT 5.520 67.760 83.260 68.240 ;
        RECT 23.990 67.560 24.310 67.620 ;
        RECT 26.290 67.560 26.610 67.620 ;
        RECT 7.060 67.420 26.610 67.560 ;
        RECT 7.060 66.925 7.200 67.420 ;
        RECT 23.990 67.360 24.310 67.420 ;
        RECT 26.290 67.360 26.610 67.420 ;
        RECT 35.950 67.360 36.270 67.620 ;
        RECT 64.930 67.560 65.250 67.620 ;
        RECT 69.530 67.560 69.850 67.620 ;
        RECT 75.510 67.560 75.830 67.620 ;
        RECT 64.930 67.420 76.660 67.560 ;
        RECT 64.930 67.360 65.250 67.420 ;
        RECT 69.530 67.360 69.850 67.420 ;
        RECT 75.510 67.360 75.830 67.420 ;
        RECT 7.470 67.220 7.760 67.265 ;
        RECT 9.570 67.220 9.860 67.265 ;
        RECT 11.140 67.220 11.430 67.265 ;
        RECT 7.470 67.080 11.430 67.220 ;
        RECT 7.470 67.035 7.760 67.080 ;
        RECT 9.570 67.035 9.860 67.080 ;
        RECT 11.140 67.035 11.430 67.080 ;
        RECT 12.030 67.220 12.350 67.280 ;
        RECT 13.885 67.220 14.175 67.265 ;
        RECT 12.030 67.080 14.175 67.220 ;
        RECT 12.030 67.020 12.350 67.080 ;
        RECT 13.885 67.035 14.175 67.080 ;
        RECT 15.710 67.220 16.030 67.280 ;
        RECT 16.185 67.220 16.475 67.265 ;
        RECT 20.785 67.220 21.075 67.265 ;
        RECT 21.230 67.220 21.550 67.280 ;
        RECT 36.410 67.220 36.730 67.280 ;
        RECT 57.570 67.220 57.890 67.280 ;
        RECT 60.370 67.220 60.660 67.265 ;
        RECT 62.470 67.220 62.760 67.265 ;
        RECT 64.040 67.220 64.330 67.265 ;
        RECT 15.710 67.080 20.080 67.220 ;
        RECT 6.985 66.695 7.275 66.925 ;
        RECT 7.865 66.880 8.155 66.925 ;
        RECT 9.055 66.880 9.345 66.925 ;
        RECT 11.575 66.880 11.865 66.925 ;
        RECT 7.865 66.740 11.865 66.880 ;
        RECT 13.960 66.880 14.100 67.035 ;
        RECT 15.710 67.020 16.030 67.080 ;
        RECT 16.185 67.035 16.475 67.080 ;
        RECT 16.645 66.880 16.935 66.925 ;
        RECT 13.960 66.740 16.935 66.880 ;
        RECT 7.865 66.695 8.155 66.740 ;
        RECT 9.055 66.695 9.345 66.740 ;
        RECT 11.575 66.695 11.865 66.740 ;
        RECT 16.645 66.695 16.935 66.740 ;
        RECT 14.330 66.540 14.650 66.600 ;
        RECT 14.805 66.540 15.095 66.585 ;
        RECT 14.330 66.400 15.095 66.540 ;
        RECT 14.330 66.340 14.650 66.400 ;
        RECT 14.805 66.355 15.095 66.400 ;
        RECT 15.250 66.540 15.570 66.600 ;
        RECT 17.565 66.540 17.855 66.585 ;
        RECT 15.250 66.400 17.855 66.540 ;
        RECT 15.250 66.340 15.570 66.400 ;
        RECT 17.565 66.355 17.855 66.400 ;
        RECT 18.010 66.340 18.330 66.600 ;
        RECT 19.940 66.585 20.080 67.080 ;
        RECT 20.785 67.080 21.550 67.220 ;
        RECT 20.785 67.035 21.075 67.080 ;
        RECT 21.230 67.020 21.550 67.080 ;
        RECT 36.040 67.080 36.730 67.220 ;
        RECT 20.325 66.880 20.615 66.925 ;
        RECT 24.450 66.880 24.770 66.940 ;
        RECT 20.325 66.740 24.770 66.880 ;
        RECT 20.325 66.695 20.615 66.740 ;
        RECT 24.450 66.680 24.770 66.740 ;
        RECT 26.290 66.880 26.610 66.940 ;
        RECT 26.765 66.880 27.055 66.925 ;
        RECT 26.290 66.740 27.055 66.880 ;
        RECT 26.290 66.680 26.610 66.740 ;
        RECT 26.765 66.695 27.055 66.740 ;
        RECT 29.970 66.880 30.290 66.940 ;
        RECT 36.040 66.925 36.180 67.080 ;
        RECT 36.410 67.020 36.730 67.080 ;
        RECT 54.900 67.080 58.720 67.220 ;
        RECT 30.445 66.880 30.735 66.925 ;
        RECT 29.970 66.740 30.735 66.880 ;
        RECT 29.970 66.680 30.290 66.740 ;
        RECT 30.445 66.695 30.735 66.740 ;
        RECT 35.965 66.695 36.255 66.925 ;
        RECT 18.945 66.540 19.235 66.585 ;
        RECT 18.515 66.400 19.235 66.540 ;
        RECT 8.350 66.245 8.670 66.260 ;
        RECT 8.320 66.015 8.670 66.245 ;
        RECT 8.350 66.000 8.670 66.015 ;
        RECT 16.170 66.000 16.490 66.260 ;
        RECT 16.645 66.200 16.935 66.245 ;
        RECT 17.090 66.200 17.410 66.260 ;
        RECT 16.645 66.060 17.410 66.200 ;
        RECT 16.645 66.015 16.935 66.060 ;
        RECT 17.090 66.000 17.410 66.060 ;
        RECT 14.330 65.860 14.650 65.920 ;
        RECT 15.265 65.860 15.555 65.905 ;
        RECT 14.330 65.720 15.555 65.860 ;
        RECT 14.330 65.660 14.650 65.720 ;
        RECT 15.265 65.675 15.555 65.720 ;
        RECT 17.550 65.860 17.870 65.920 ;
        RECT 18.515 65.860 18.655 66.400 ;
        RECT 18.945 66.355 19.235 66.400 ;
        RECT 19.865 66.355 20.155 66.585 ;
        RECT 21.230 66.340 21.550 66.600 ;
        RECT 23.085 66.540 23.375 66.585 ;
        RECT 35.030 66.540 35.350 66.600 ;
        RECT 23.085 66.400 35.350 66.540 ;
        RECT 23.085 66.355 23.375 66.400 ;
        RECT 35.030 66.340 35.350 66.400 ;
        RECT 36.410 66.340 36.730 66.600 ;
        RECT 37.330 66.540 37.650 66.600 ;
        RECT 41.010 66.540 41.330 66.600 ;
        RECT 37.330 66.400 41.330 66.540 ;
        RECT 37.330 66.340 37.650 66.400 ;
        RECT 41.010 66.340 41.330 66.400 ;
        RECT 41.470 66.540 41.790 66.600 ;
        RECT 41.945 66.540 42.235 66.585 ;
        RECT 41.470 66.400 42.235 66.540 ;
        RECT 41.470 66.340 41.790 66.400 ;
        RECT 41.945 66.355 42.235 66.400 ;
        RECT 48.370 66.540 48.690 66.600 ;
        RECT 49.290 66.540 49.610 66.600 ;
        RECT 48.370 66.400 49.610 66.540 ;
        RECT 48.370 66.340 48.690 66.400 ;
        RECT 49.290 66.340 49.610 66.400 ;
        RECT 49.750 66.540 50.070 66.600 ;
        RECT 51.145 66.540 51.435 66.585 ;
        RECT 49.750 66.400 51.435 66.540 ;
        RECT 49.750 66.340 50.070 66.400 ;
        RECT 51.145 66.355 51.435 66.400 ;
        RECT 51.605 66.540 51.895 66.585 ;
        RECT 52.970 66.540 53.290 66.600 ;
        RECT 51.605 66.400 53.290 66.540 ;
        RECT 51.605 66.355 51.895 66.400 ;
        RECT 52.970 66.340 53.290 66.400 ;
        RECT 53.430 66.340 53.750 66.600 ;
        RECT 34.110 66.000 34.430 66.260 ;
        RECT 52.525 66.200 52.815 66.245 ;
        RECT 54.900 66.200 55.040 67.080 ;
        RECT 57.570 67.020 57.890 67.080 ;
        RECT 55.270 66.880 55.590 66.940 ;
        RECT 55.270 66.740 58.260 66.880 ;
        RECT 55.270 66.680 55.590 66.740 ;
        RECT 58.120 66.585 58.260 66.740 ;
        RECT 58.580 66.585 58.720 67.080 ;
        RECT 60.370 67.080 64.330 67.220 ;
        RECT 60.370 67.035 60.660 67.080 ;
        RECT 62.470 67.035 62.760 67.080 ;
        RECT 64.040 67.035 64.330 67.080 ;
        RECT 66.785 67.220 67.075 67.265 ;
        RECT 69.070 67.220 69.390 67.280 ;
        RECT 70.910 67.220 71.230 67.280 ;
        RECT 66.785 67.080 71.230 67.220 ;
        RECT 76.520 67.220 76.660 67.420 ;
        RECT 76.890 67.360 77.210 67.620 ;
        RECT 77.810 67.360 78.130 67.620 ;
        RECT 76.520 67.080 77.120 67.220 ;
        RECT 66.785 67.035 67.075 67.080 ;
        RECT 69.070 67.020 69.390 67.080 ;
        RECT 70.910 67.020 71.230 67.080 ;
        RECT 60.765 66.880 61.055 66.925 ;
        RECT 61.955 66.880 62.245 66.925 ;
        RECT 64.475 66.880 64.765 66.925 ;
        RECT 60.765 66.740 64.765 66.880 ;
        RECT 60.765 66.695 61.055 66.740 ;
        RECT 61.955 66.695 62.245 66.740 ;
        RECT 64.475 66.695 64.765 66.740 ;
        RECT 71.830 66.880 72.150 66.940 ;
        RECT 73.225 66.880 73.515 66.925 ;
        RECT 76.430 66.880 76.750 66.940 ;
        RECT 71.830 66.740 73.515 66.880 ;
        RECT 71.830 66.680 72.150 66.740 ;
        RECT 73.225 66.695 73.515 66.740 ;
        RECT 75.140 66.740 76.750 66.880 ;
        RECT 56.205 66.540 56.495 66.585 ;
        RECT 56.665 66.540 56.955 66.585 ;
        RECT 56.205 66.400 56.955 66.540 ;
        RECT 56.205 66.355 56.495 66.400 ;
        RECT 56.665 66.355 56.955 66.400 ;
        RECT 58.045 66.355 58.335 66.585 ;
        RECT 58.505 66.355 58.795 66.585 ;
        RECT 59.870 66.340 60.190 66.600 ;
        RECT 61.250 66.585 61.570 66.600 ;
        RECT 61.220 66.540 61.570 66.585 ;
        RECT 61.055 66.400 61.570 66.540 ;
        RECT 61.220 66.355 61.570 66.400 ;
        RECT 69.545 66.540 69.835 66.585 ;
        RECT 70.450 66.540 70.770 66.600 ;
        RECT 75.140 66.585 75.280 66.740 ;
        RECT 76.430 66.680 76.750 66.740 ;
        RECT 69.545 66.400 70.770 66.540 ;
        RECT 69.545 66.355 69.835 66.400 ;
        RECT 61.250 66.340 61.570 66.355 ;
        RECT 70.450 66.340 70.770 66.400 ;
        RECT 75.065 66.355 75.355 66.585 ;
        RECT 75.970 66.340 76.290 66.600 ;
        RECT 76.980 66.540 77.120 67.080 ;
        RECT 78.745 66.540 79.035 66.585 ;
        RECT 76.980 66.400 79.035 66.540 ;
        RECT 78.745 66.355 79.035 66.400 ;
        RECT 80.570 66.340 80.890 66.600 ;
        RECT 52.525 66.060 55.040 66.200 ;
        RECT 52.525 66.015 52.815 66.060 ;
        RECT 57.585 66.015 57.875 66.245 ;
        RECT 73.670 66.200 73.990 66.260 ;
        RECT 74.145 66.200 74.435 66.245 ;
        RECT 68.700 66.060 73.440 66.200 ;
        RECT 17.550 65.720 18.655 65.860 ;
        RECT 20.770 65.860 21.090 65.920 ;
        RECT 22.165 65.860 22.455 65.905 ;
        RECT 20.770 65.720 22.455 65.860 ;
        RECT 17.550 65.660 17.870 65.720 ;
        RECT 20.770 65.660 21.090 65.720 ;
        RECT 22.165 65.675 22.455 65.720 ;
        RECT 32.730 65.860 33.050 65.920 ;
        RECT 33.665 65.860 33.955 65.905 ;
        RECT 32.730 65.720 33.955 65.860 ;
        RECT 32.730 65.660 33.050 65.720 ;
        RECT 33.665 65.675 33.955 65.720 ;
        RECT 36.870 65.860 37.190 65.920 ;
        RECT 37.345 65.860 37.635 65.905 ;
        RECT 36.870 65.720 37.635 65.860 ;
        RECT 36.870 65.660 37.190 65.720 ;
        RECT 37.345 65.675 37.635 65.720 ;
        RECT 38.710 65.860 39.030 65.920 ;
        RECT 39.185 65.860 39.475 65.905 ;
        RECT 38.710 65.720 39.475 65.860 ;
        RECT 38.710 65.660 39.030 65.720 ;
        RECT 39.185 65.675 39.475 65.720 ;
        RECT 48.830 65.860 49.150 65.920 ;
        RECT 50.225 65.860 50.515 65.905 ;
        RECT 48.830 65.720 50.515 65.860 ;
        RECT 48.830 65.660 49.150 65.720 ;
        RECT 50.225 65.675 50.515 65.720 ;
        RECT 52.065 65.860 52.355 65.905 ;
        RECT 57.660 65.860 57.800 66.015 ;
        RECT 52.065 65.720 57.800 65.860 ;
        RECT 58.950 65.860 59.270 65.920 ;
        RECT 68.700 65.905 68.840 66.060 ;
        RECT 73.300 65.920 73.440 66.060 ;
        RECT 73.670 66.060 74.435 66.200 ;
        RECT 73.670 66.000 73.990 66.060 ;
        RECT 74.145 66.015 74.435 66.060 ;
        RECT 76.430 66.200 76.750 66.260 ;
        RECT 79.205 66.200 79.495 66.245 ;
        RECT 76.430 66.060 79.495 66.200 ;
        RECT 76.430 66.000 76.750 66.060 ;
        RECT 79.205 66.015 79.495 66.060 ;
        RECT 79.665 66.015 79.955 66.245 ;
        RECT 59.425 65.860 59.715 65.905 ;
        RECT 58.950 65.720 59.715 65.860 ;
        RECT 52.065 65.675 52.355 65.720 ;
        RECT 58.950 65.660 59.270 65.720 ;
        RECT 59.425 65.675 59.715 65.720 ;
        RECT 68.625 65.675 68.915 65.905 ;
        RECT 70.450 65.660 70.770 65.920 ;
        RECT 73.210 65.860 73.530 65.920 ;
        RECT 78.730 65.860 79.050 65.920 ;
        RECT 79.740 65.860 79.880 66.015 ;
        RECT 73.210 65.720 79.880 65.860 ;
        RECT 73.210 65.660 73.530 65.720 ;
        RECT 78.730 65.660 79.050 65.720 ;
        RECT 5.520 65.040 83.260 65.520 ;
        RECT 7.905 64.840 8.195 64.885 ;
        RECT 8.350 64.840 8.670 64.900 ;
        RECT 7.905 64.700 8.670 64.840 ;
        RECT 7.905 64.655 8.195 64.700 ;
        RECT 8.350 64.640 8.670 64.700 ;
        RECT 9.285 64.840 9.575 64.885 ;
        RECT 9.730 64.840 10.050 64.900 ;
        RECT 9.285 64.700 10.050 64.840 ;
        RECT 9.285 64.655 9.575 64.700 ;
        RECT 9.730 64.640 10.050 64.700 ;
        RECT 17.105 64.840 17.395 64.885 ;
        RECT 18.930 64.840 19.250 64.900 ;
        RECT 24.925 64.840 25.215 64.885 ;
        RECT 28.590 64.840 28.910 64.900 ;
        RECT 17.105 64.700 19.620 64.840 ;
        RECT 17.105 64.655 17.395 64.700 ;
        RECT 18.930 64.640 19.250 64.700 ;
        RECT 8.825 64.500 9.115 64.545 ;
        RECT 11.125 64.500 11.415 64.545 ;
        RECT 8.825 64.360 11.415 64.500 ;
        RECT 8.825 64.315 9.115 64.360 ;
        RECT 11.125 64.315 11.415 64.360 ;
        RECT 12.030 64.300 12.350 64.560 ;
        RECT 13.885 64.500 14.175 64.545 ;
        RECT 14.330 64.500 14.650 64.560 ;
        RECT 19.480 64.545 19.620 64.700 ;
        RECT 24.925 64.700 28.910 64.840 ;
        RECT 24.925 64.655 25.215 64.700 ;
        RECT 28.590 64.640 28.910 64.700 ;
        RECT 29.050 64.640 29.370 64.900 ;
        RECT 32.285 64.840 32.575 64.885 ;
        RECT 36.410 64.840 36.730 64.900 ;
        RECT 41.025 64.840 41.315 64.885 ;
        RECT 32.285 64.700 41.315 64.840 ;
        RECT 32.285 64.655 32.575 64.700 ;
        RECT 36.410 64.640 36.730 64.700 ;
        RECT 41.025 64.655 41.315 64.700 ;
        RECT 41.470 64.640 41.790 64.900 ;
        RECT 52.065 64.655 52.355 64.885 ;
        RECT 53.430 64.840 53.750 64.900 ;
        RECT 54.365 64.840 54.655 64.885 ;
        RECT 53.430 64.700 54.655 64.840 ;
        RECT 13.885 64.360 16.860 64.500 ;
        RECT 13.885 64.315 14.175 64.360 ;
        RECT 14.330 64.300 14.650 64.360 ;
        RECT 9.270 64.160 9.590 64.220 ;
        RECT 9.745 64.160 10.035 64.205 ;
        RECT 9.270 64.020 10.035 64.160 ;
        RECT 9.270 63.960 9.590 64.020 ;
        RECT 9.745 63.975 10.035 64.020 ;
        RECT 10.190 64.160 10.510 64.220 ;
        RECT 12.965 64.160 13.255 64.205 ;
        RECT 10.190 64.020 13.255 64.160 ;
        RECT 10.190 63.960 10.510 64.020 ;
        RECT 12.580 63.880 12.720 64.020 ;
        RECT 12.965 63.975 13.255 64.020 ;
        RECT 13.425 64.160 13.715 64.205 ;
        RECT 14.805 64.160 15.095 64.205 ;
        RECT 15.710 64.160 16.030 64.220 ;
        RECT 16.185 64.160 16.475 64.205 ;
        RECT 13.425 64.020 14.100 64.160 ;
        RECT 13.425 63.975 13.715 64.020 ;
        RECT 13.960 63.880 14.100 64.020 ;
        RECT 14.805 64.020 15.205 64.160 ;
        RECT 15.710 64.020 16.475 64.160 ;
        RECT 14.805 63.975 15.095 64.020 ;
        RECT 10.665 63.820 10.955 63.865 ;
        RECT 11.570 63.820 11.890 63.880 ;
        RECT 10.665 63.680 11.890 63.820 ;
        RECT 10.665 63.635 10.955 63.680 ;
        RECT 11.570 63.620 11.890 63.680 ;
        RECT 12.490 63.620 12.810 63.880 ;
        RECT 13.870 63.620 14.190 63.880 ;
        RECT 14.880 63.820 15.020 63.975 ;
        RECT 15.710 63.960 16.030 64.020 ;
        RECT 16.185 63.975 16.475 64.020 ;
        RECT 15.265 63.820 15.555 63.865 ;
        RECT 14.420 63.680 15.555 63.820 ;
        RECT 16.720 63.820 16.860 64.360 ;
        RECT 19.405 64.315 19.695 64.545 ;
        RECT 24.005 64.500 24.295 64.545 ;
        RECT 34.110 64.500 34.430 64.560 ;
        RECT 52.140 64.500 52.280 64.655 ;
        RECT 53.430 64.640 53.750 64.700 ;
        RECT 54.365 64.655 54.655 64.700 ;
        RECT 59.425 64.840 59.715 64.885 ;
        RECT 60.790 64.840 61.110 64.900 ;
        RECT 59.425 64.700 61.110 64.840 ;
        RECT 59.425 64.655 59.715 64.700 ;
        RECT 60.790 64.640 61.110 64.700 ;
        RECT 64.025 64.840 64.315 64.885 ;
        RECT 68.165 64.840 68.455 64.885 ;
        RECT 70.450 64.840 70.770 64.900 ;
        RECT 64.025 64.700 67.460 64.840 ;
        RECT 64.025 64.655 64.315 64.700 ;
        RECT 24.005 64.360 25.140 64.500 ;
        RECT 24.005 64.315 24.295 64.360 ;
        RECT 25.000 64.220 25.140 64.360 ;
        RECT 25.460 64.360 28.820 64.500 ;
        RECT 18.470 63.960 18.790 64.220 ;
        RECT 18.945 64.160 19.235 64.205 ;
        RECT 19.850 64.160 20.170 64.220 ;
        RECT 18.945 64.020 20.170 64.160 ;
        RECT 18.945 63.975 19.235 64.020 ;
        RECT 19.850 63.960 20.170 64.020 ;
        RECT 20.325 63.975 20.615 64.205 ;
        RECT 19.390 63.820 19.710 63.880 ;
        RECT 16.720 63.680 19.710 63.820 ;
        RECT 11.660 63.480 11.800 63.620 ;
        RECT 12.950 63.480 13.270 63.540 ;
        RECT 11.660 63.340 13.270 63.480 ;
        RECT 12.950 63.280 13.270 63.340 ;
        RECT 14.420 63.140 14.560 63.680 ;
        RECT 15.265 63.635 15.555 63.680 ;
        RECT 19.390 63.620 19.710 63.680 ;
        RECT 14.805 63.480 15.095 63.525 ;
        RECT 20.400 63.480 20.540 63.975 ;
        RECT 20.770 63.960 21.090 64.220 ;
        RECT 24.910 63.960 25.230 64.220 ;
        RECT 25.460 64.205 25.600 64.360 ;
        RECT 28.680 64.220 28.820 64.360 ;
        RECT 30.980 64.360 34.430 64.500 ;
        RECT 25.385 63.975 25.675 64.205 ;
        RECT 26.305 64.160 26.595 64.205 ;
        RECT 27.670 64.160 27.990 64.220 ;
        RECT 26.305 64.020 27.990 64.160 ;
        RECT 26.305 63.975 26.595 64.020 ;
        RECT 27.670 63.960 27.990 64.020 ;
        RECT 28.130 63.960 28.450 64.220 ;
        RECT 28.590 63.960 28.910 64.220 ;
        RECT 29.510 64.160 29.830 64.220 ;
        RECT 30.980 64.205 31.120 64.360 ;
        RECT 34.110 64.300 34.430 64.360 ;
        RECT 35.120 64.360 40.780 64.500 ;
        RECT 29.985 64.160 30.275 64.205 ;
        RECT 29.510 64.020 30.275 64.160 ;
        RECT 29.510 63.960 29.830 64.020 ;
        RECT 29.985 63.975 30.275 64.020 ;
        RECT 30.905 63.975 31.195 64.205 ;
        RECT 32.730 63.960 33.050 64.220 ;
        RECT 26.750 63.620 27.070 63.880 ;
        RECT 27.225 63.635 27.515 63.865 ;
        RECT 30.445 63.820 30.735 63.865 ;
        RECT 34.570 63.820 34.890 63.880 ;
        RECT 35.120 63.820 35.260 64.360 ;
        RECT 38.710 64.205 39.030 64.220 ;
        RECT 38.710 64.160 39.060 64.205 ;
        RECT 38.710 64.020 39.225 64.160 ;
        RECT 38.710 63.975 39.060 64.020 ;
        RECT 38.710 63.960 39.030 63.975 ;
        RECT 40.090 63.960 40.410 64.220 ;
        RECT 40.640 64.205 40.780 64.360 ;
        RECT 41.100 64.360 52.280 64.500 ;
        RECT 41.100 64.220 41.240 64.360 ;
        RECT 53.890 64.300 54.210 64.560 ;
        RECT 60.330 64.500 60.650 64.560 ;
        RECT 67.320 64.500 67.460 64.700 ;
        RECT 68.165 64.700 70.770 64.840 ;
        RECT 68.165 64.655 68.455 64.700 ;
        RECT 70.450 64.640 70.770 64.700 ;
        RECT 75.510 64.840 75.830 64.900 ;
        RECT 77.365 64.840 77.655 64.885 ;
        RECT 80.110 64.840 80.430 64.900 ;
        RECT 75.510 64.700 77.120 64.840 ;
        RECT 75.510 64.640 75.830 64.700 ;
        RECT 70.910 64.500 71.230 64.560 ;
        RECT 76.980 64.500 77.120 64.700 ;
        RECT 77.365 64.700 80.430 64.840 ;
        RECT 77.365 64.655 77.655 64.700 ;
        RECT 80.110 64.640 80.430 64.700 ;
        RECT 60.330 64.360 65.620 64.500 ;
        RECT 67.320 64.360 70.680 64.500 ;
        RECT 60.330 64.300 60.650 64.360 ;
        RECT 40.565 63.975 40.855 64.205 ;
        RECT 41.010 63.960 41.330 64.220 ;
        RECT 45.165 64.160 45.455 64.205 ;
        RECT 47.465 64.160 47.755 64.205 ;
        RECT 45.165 64.020 47.755 64.160 ;
        RECT 45.165 63.975 45.455 64.020 ;
        RECT 47.465 63.975 47.755 64.020 ;
        RECT 59.885 64.160 60.175 64.205 ;
        RECT 61.710 64.160 62.030 64.220 ;
        RECT 59.885 64.020 62.030 64.160 ;
        RECT 59.885 63.975 60.175 64.020 ;
        RECT 61.710 63.960 62.030 64.020 ;
        RECT 65.480 64.160 65.620 64.360 ;
        RECT 70.540 64.205 70.680 64.360 ;
        RECT 70.910 64.360 76.660 64.500 ;
        RECT 76.980 64.360 79.880 64.500 ;
        RECT 70.910 64.300 71.230 64.360 ;
        RECT 65.480 64.020 69.300 64.160 ;
        RECT 30.445 63.680 35.260 63.820 ;
        RECT 35.515 63.820 35.805 63.865 ;
        RECT 38.035 63.820 38.325 63.865 ;
        RECT 39.225 63.820 39.515 63.865 ;
        RECT 42.865 63.820 43.155 63.865 ;
        RECT 35.515 63.680 39.515 63.820 ;
        RECT 30.445 63.635 30.735 63.680 ;
        RECT 14.805 63.340 20.540 63.480 ;
        RECT 22.165 63.480 22.455 63.525 ;
        RECT 24.450 63.480 24.770 63.540 ;
        RECT 22.165 63.340 24.770 63.480 ;
        RECT 14.805 63.295 15.095 63.340 ;
        RECT 22.165 63.295 22.455 63.340 ;
        RECT 24.450 63.280 24.770 63.340 ;
        RECT 15.710 63.140 16.030 63.200 ;
        RECT 17.090 63.140 17.410 63.200 ;
        RECT 14.420 63.000 17.410 63.140 ;
        RECT 15.710 62.940 16.030 63.000 ;
        RECT 17.090 62.940 17.410 63.000 ;
        RECT 17.565 63.140 17.855 63.185 ;
        RECT 18.010 63.140 18.330 63.200 ;
        RECT 17.565 63.000 18.330 63.140 ;
        RECT 17.565 62.955 17.855 63.000 ;
        RECT 18.010 62.940 18.330 63.000 ;
        RECT 23.530 63.140 23.850 63.200 ;
        RECT 24.005 63.140 24.295 63.185 ;
        RECT 23.530 63.000 24.295 63.140 ;
        RECT 23.530 62.940 23.850 63.000 ;
        RECT 24.005 62.955 24.295 63.000 ;
        RECT 26.750 63.140 27.070 63.200 ;
        RECT 27.300 63.140 27.440 63.635 ;
        RECT 34.570 63.620 34.890 63.680 ;
        RECT 35.515 63.635 35.805 63.680 ;
        RECT 38.035 63.635 38.325 63.680 ;
        RECT 39.225 63.635 39.515 63.680 ;
        RECT 41.100 63.680 43.155 63.820 ;
        RECT 41.100 63.540 41.240 63.680 ;
        RECT 42.865 63.635 43.155 63.680 ;
        RECT 45.610 63.620 45.930 63.880 ;
        RECT 46.530 63.620 46.850 63.880 ;
        RECT 49.750 63.820 50.070 63.880 ;
        RECT 50.225 63.820 50.515 63.865 ;
        RECT 49.750 63.680 50.515 63.820 ;
        RECT 49.750 63.620 50.070 63.680 ;
        RECT 50.225 63.635 50.515 63.680 ;
        RECT 54.825 63.635 55.115 63.865 ;
        RECT 29.970 63.480 30.290 63.540 ;
        RECT 33.205 63.480 33.495 63.525 ;
        RECT 29.970 63.340 33.495 63.480 ;
        RECT 29.970 63.280 30.290 63.340 ;
        RECT 33.205 63.295 33.495 63.340 ;
        RECT 35.950 63.480 36.240 63.525 ;
        RECT 37.520 63.480 37.810 63.525 ;
        RECT 39.620 63.480 39.910 63.525 ;
        RECT 35.950 63.340 39.910 63.480 ;
        RECT 35.950 63.295 36.240 63.340 ;
        RECT 37.520 63.295 37.810 63.340 ;
        RECT 39.620 63.295 39.910 63.340 ;
        RECT 41.010 63.280 41.330 63.540 ;
        RECT 49.290 63.480 49.610 63.540 ;
        RECT 54.900 63.480 55.040 63.635 ;
        RECT 60.330 63.620 60.650 63.880 ;
        RECT 63.090 63.820 63.410 63.880 ;
        RECT 65.480 63.865 65.620 64.020 ;
        RECT 64.485 63.820 64.775 63.865 ;
        RECT 63.090 63.680 64.775 63.820 ;
        RECT 63.090 63.620 63.410 63.680 ;
        RECT 64.485 63.635 64.775 63.680 ;
        RECT 65.405 63.635 65.695 63.865 ;
        RECT 68.150 63.820 68.470 63.880 ;
        RECT 69.160 63.865 69.300 64.020 ;
        RECT 70.465 63.975 70.755 64.205 ;
        RECT 71.830 64.160 72.150 64.220 ;
        RECT 74.145 64.160 74.435 64.205 ;
        RECT 71.830 64.020 74.435 64.160 ;
        RECT 71.830 63.960 72.150 64.020 ;
        RECT 74.145 63.975 74.435 64.020 ;
        RECT 74.590 63.960 74.910 64.220 ;
        RECT 76.520 64.205 76.660 64.360 ;
        RECT 75.525 63.975 75.815 64.205 ;
        RECT 76.445 63.975 76.735 64.205 ;
        RECT 77.825 64.160 78.115 64.205 ;
        RECT 78.270 64.160 78.590 64.220 ;
        RECT 77.825 64.020 78.590 64.160 ;
        RECT 77.825 63.975 78.115 64.020 ;
        RECT 68.625 63.820 68.915 63.865 ;
        RECT 68.150 63.680 68.915 63.820 ;
        RECT 68.150 63.620 68.470 63.680 ;
        RECT 68.625 63.635 68.915 63.680 ;
        RECT 69.085 63.635 69.375 63.865 ;
        RECT 73.210 63.620 73.530 63.880 ;
        RECT 73.670 63.820 73.990 63.880 ;
        RECT 75.600 63.820 75.740 63.975 ;
        RECT 73.670 63.680 75.740 63.820 ;
        RECT 75.970 63.820 76.290 63.880 ;
        RECT 77.900 63.820 78.040 63.975 ;
        RECT 78.270 63.960 78.590 64.020 ;
        RECT 78.730 63.960 79.050 64.220 ;
        RECT 79.190 63.960 79.510 64.220 ;
        RECT 79.740 64.205 79.880 64.360 ;
        RECT 79.665 63.975 79.955 64.205 ;
        RECT 75.970 63.680 78.040 63.820 ;
        RECT 73.670 63.620 73.990 63.680 ;
        RECT 75.970 63.620 76.290 63.680 ;
        RECT 49.290 63.340 55.040 63.480 ;
        RECT 61.710 63.480 62.030 63.540 ;
        RECT 66.325 63.480 66.615 63.525 ;
        RECT 61.710 63.340 66.615 63.480 ;
        RECT 49.290 63.280 49.610 63.340 ;
        RECT 61.710 63.280 62.030 63.340 ;
        RECT 66.325 63.295 66.615 63.340 ;
        RECT 67.690 63.480 68.010 63.540 ;
        RECT 80.585 63.480 80.875 63.525 ;
        RECT 67.690 63.340 80.875 63.480 ;
        RECT 67.690 63.280 68.010 63.340 ;
        RECT 80.585 63.295 80.875 63.340 ;
        RECT 26.750 63.000 27.440 63.140 ;
        RECT 27.670 63.140 27.990 63.200 ;
        RECT 35.030 63.140 35.350 63.200 ;
        RECT 40.550 63.140 40.870 63.200 ;
        RECT 27.670 63.000 40.870 63.140 ;
        RECT 26.750 62.940 27.070 63.000 ;
        RECT 27.670 62.940 27.990 63.000 ;
        RECT 35.030 62.940 35.350 63.000 ;
        RECT 40.550 62.940 40.870 63.000 ;
        RECT 41.470 63.140 41.790 63.200 ;
        RECT 43.325 63.140 43.615 63.185 ;
        RECT 41.470 63.000 43.615 63.140 ;
        RECT 41.470 62.940 41.790 63.000 ;
        RECT 43.325 62.955 43.615 63.000 ;
        RECT 57.570 62.940 57.890 63.200 ;
        RECT 61.250 63.140 61.570 63.200 ;
        RECT 62.185 63.140 62.475 63.185 ;
        RECT 61.250 63.000 62.475 63.140 ;
        RECT 61.250 62.940 61.570 63.000 ;
        RECT 62.185 62.955 62.475 63.000 ;
        RECT 70.910 63.140 71.230 63.200 ;
        RECT 74.130 63.140 74.450 63.200 ;
        RECT 70.910 63.000 74.450 63.140 ;
        RECT 70.910 62.940 71.230 63.000 ;
        RECT 74.130 62.940 74.450 63.000 ;
        RECT 5.520 62.320 83.260 62.800 ;
        RECT 10.205 62.120 10.495 62.165 ;
        RECT 15.725 62.120 16.015 62.165 ;
        RECT 16.170 62.120 16.490 62.180 ;
        RECT 25.830 62.120 26.150 62.180 ;
        RECT 10.205 61.980 13.180 62.120 ;
        RECT 10.205 61.935 10.495 61.980 ;
        RECT 10.280 61.440 10.420 61.935 ;
        RECT 8.440 61.300 10.420 61.440 ;
        RECT 13.040 61.440 13.180 61.980 ;
        RECT 15.725 61.980 16.490 62.120 ;
        RECT 15.725 61.935 16.015 61.980 ;
        RECT 16.170 61.920 16.490 61.980 ;
        RECT 24.080 61.980 26.150 62.120 ;
        RECT 15.250 61.780 15.570 61.840 ;
        RECT 17.565 61.780 17.855 61.825 ;
        RECT 15.250 61.640 17.855 61.780 ;
        RECT 15.250 61.580 15.570 61.640 ;
        RECT 17.565 61.595 17.855 61.640 ;
        RECT 20.785 61.780 21.075 61.825 ;
        RECT 24.080 61.780 24.220 61.980 ;
        RECT 25.830 61.920 26.150 61.980 ;
        RECT 28.590 62.120 28.910 62.180 ;
        RECT 31.365 62.120 31.655 62.165 ;
        RECT 28.590 61.980 31.655 62.120 ;
        RECT 28.590 61.920 28.910 61.980 ;
        RECT 31.365 61.935 31.655 61.980 ;
        RECT 34.110 62.120 34.430 62.180 ;
        RECT 41.025 62.120 41.315 62.165 ;
        RECT 34.110 61.980 41.315 62.120 ;
        RECT 34.110 61.920 34.430 61.980 ;
        RECT 41.025 61.935 41.315 61.980 ;
        RECT 45.610 62.120 45.930 62.180 ;
        RECT 46.085 62.120 46.375 62.165 ;
        RECT 45.610 61.980 46.375 62.120 ;
        RECT 20.785 61.640 24.220 61.780 ;
        RECT 24.490 61.780 24.780 61.825 ;
        RECT 26.590 61.780 26.880 61.825 ;
        RECT 28.160 61.780 28.450 61.825 ;
        RECT 24.490 61.640 28.450 61.780 ;
        RECT 20.785 61.595 21.075 61.640 ;
        RECT 24.490 61.595 24.780 61.640 ;
        RECT 26.590 61.595 26.880 61.640 ;
        RECT 28.160 61.595 28.450 61.640 ;
        RECT 34.610 61.780 34.900 61.825 ;
        RECT 36.710 61.780 37.000 61.825 ;
        RECT 38.280 61.780 38.570 61.825 ;
        RECT 34.610 61.640 38.570 61.780 ;
        RECT 34.610 61.595 34.900 61.640 ;
        RECT 36.710 61.595 37.000 61.640 ;
        RECT 38.280 61.595 38.570 61.640 ;
        RECT 13.410 61.440 13.730 61.500 ;
        RECT 13.040 61.300 13.730 61.440 ;
        RECT 8.440 61.145 8.580 61.300 ;
        RECT 8.365 60.915 8.655 61.145 ;
        RECT 8.825 61.100 9.115 61.145 ;
        RECT 12.490 61.100 12.810 61.160 ;
        RECT 13.040 61.145 13.180 61.300 ;
        RECT 13.410 61.240 13.730 61.300 ;
        RECT 8.825 60.960 12.810 61.100 ;
        RECT 8.825 60.915 9.115 60.960 ;
        RECT 7.430 60.760 7.750 60.820 ;
        RECT 10.280 60.805 10.420 60.960 ;
        RECT 12.490 60.900 12.810 60.960 ;
        RECT 12.965 60.915 13.255 61.145 ;
        RECT 15.340 61.100 15.480 61.580 ;
        RECT 17.090 61.440 17.410 61.500 ;
        RECT 18.025 61.440 18.315 61.485 ;
        RECT 17.090 61.300 18.315 61.440 ;
        RECT 17.090 61.240 17.410 61.300 ;
        RECT 18.025 61.255 18.315 61.300 ;
        RECT 24.885 61.440 25.175 61.485 ;
        RECT 26.075 61.440 26.365 61.485 ;
        RECT 28.595 61.440 28.885 61.485 ;
        RECT 24.885 61.300 28.885 61.440 ;
        RECT 24.885 61.255 25.175 61.300 ;
        RECT 26.075 61.255 26.365 61.300 ;
        RECT 28.595 61.255 28.885 61.300 ;
        RECT 30.890 61.440 31.210 61.500 ;
        RECT 35.005 61.440 35.295 61.485 ;
        RECT 36.195 61.440 36.485 61.485 ;
        RECT 38.715 61.440 39.005 61.485 ;
        RECT 30.890 61.300 33.880 61.440 ;
        RECT 30.890 61.240 31.210 61.300 ;
        RECT 13.500 60.960 15.480 61.100 ;
        RECT 13.500 60.805 13.640 60.960 ;
        RECT 16.645 60.915 16.935 61.145 ;
        RECT 22.625 61.100 22.915 61.145 ;
        RECT 23.070 61.100 23.390 61.160 ;
        RECT 22.625 60.960 23.390 61.100 ;
        RECT 22.625 60.915 22.915 60.960 ;
        RECT 9.285 60.760 9.575 60.805 ;
        RECT 7.430 60.620 9.575 60.760 ;
        RECT 10.280 60.620 10.575 60.805 ;
        RECT 13.425 60.760 13.715 60.805 ;
        RECT 7.430 60.560 7.750 60.620 ;
        RECT 9.285 60.575 9.575 60.620 ;
        RECT 10.285 60.575 10.575 60.620 ;
        RECT 10.740 60.620 13.715 60.760 ;
        RECT 7.935 60.420 8.225 60.465 ;
        RECT 8.810 60.420 9.130 60.480 ;
        RECT 7.935 60.280 9.130 60.420 ;
        RECT 9.360 60.420 9.500 60.575 ;
        RECT 10.740 60.420 10.880 60.620 ;
        RECT 13.425 60.575 13.715 60.620 ;
        RECT 13.870 60.760 14.190 60.820 ;
        RECT 14.345 60.760 14.635 60.805 ;
        RECT 16.720 60.760 16.860 60.915 ;
        RECT 23.070 60.900 23.390 60.960 ;
        RECT 23.990 60.900 24.310 61.160 ;
        RECT 30.430 61.100 30.750 61.160 ;
        RECT 33.740 61.145 33.880 61.300 ;
        RECT 35.005 61.300 39.005 61.440 ;
        RECT 35.005 61.255 35.295 61.300 ;
        RECT 36.195 61.255 36.485 61.300 ;
        RECT 38.715 61.255 39.005 61.300 ;
        RECT 32.285 61.100 32.575 61.145 ;
        RECT 29.600 60.960 32.575 61.100 ;
        RECT 19.390 60.760 19.710 60.820 ;
        RECT 13.870 60.620 19.710 60.760 ;
        RECT 13.870 60.560 14.190 60.620 ;
        RECT 14.345 60.575 14.635 60.620 ;
        RECT 19.390 60.560 19.710 60.620 ;
        RECT 21.705 60.760 21.995 60.805 ;
        RECT 23.545 60.760 23.835 60.805 ;
        RECT 24.450 60.760 24.770 60.820 ;
        RECT 21.705 60.620 23.300 60.760 ;
        RECT 21.705 60.575 21.995 60.620 ;
        RECT 9.360 60.280 10.880 60.420 ;
        RECT 7.935 60.235 8.225 60.280 ;
        RECT 8.810 60.220 9.130 60.280 ;
        RECT 11.110 60.220 11.430 60.480 ;
        RECT 11.570 60.220 11.890 60.480 ;
        RECT 15.710 60.420 16.030 60.480 ;
        RECT 19.850 60.420 20.170 60.480 ;
        RECT 15.710 60.280 20.170 60.420 ;
        RECT 15.710 60.220 16.030 60.280 ;
        RECT 19.850 60.220 20.170 60.280 ;
        RECT 22.150 60.220 22.470 60.480 ;
        RECT 23.160 60.420 23.300 60.620 ;
        RECT 23.545 60.620 24.770 60.760 ;
        RECT 23.545 60.575 23.835 60.620 ;
        RECT 24.450 60.560 24.770 60.620 ;
        RECT 25.340 60.760 25.630 60.805 ;
        RECT 26.290 60.760 26.610 60.820 ;
        RECT 25.340 60.620 26.610 60.760 ;
        RECT 25.340 60.575 25.630 60.620 ;
        RECT 26.290 60.560 26.610 60.620 ;
        RECT 29.050 60.420 29.370 60.480 ;
        RECT 29.600 60.420 29.740 60.960 ;
        RECT 30.430 60.900 30.750 60.960 ;
        RECT 32.285 60.915 32.575 60.960 ;
        RECT 33.665 60.915 33.955 61.145 ;
        RECT 34.125 61.100 34.415 61.145 ;
        RECT 40.090 61.100 40.410 61.160 ;
        RECT 34.125 60.960 40.410 61.100 ;
        RECT 41.100 61.100 41.240 61.935 ;
        RECT 45.610 61.920 45.930 61.980 ;
        RECT 46.085 61.935 46.375 61.980 ;
        RECT 50.225 62.120 50.515 62.165 ;
        RECT 53.430 62.120 53.750 62.180 ;
        RECT 50.225 61.980 53.750 62.120 ;
        RECT 50.225 61.935 50.515 61.980 ;
        RECT 53.430 61.920 53.750 61.980 ;
        RECT 58.505 62.120 58.795 62.165 ;
        RECT 75.050 62.120 75.370 62.180 ;
        RECT 58.505 61.980 75.370 62.120 ;
        RECT 58.505 61.935 58.795 61.980 ;
        RECT 75.050 61.920 75.370 61.980 ;
        RECT 52.970 61.780 53.260 61.825 ;
        RECT 54.540 61.780 54.830 61.825 ;
        RECT 56.640 61.780 56.930 61.825 ;
        RECT 52.970 61.640 56.930 61.780 ;
        RECT 52.970 61.595 53.260 61.640 ;
        RECT 54.540 61.595 54.830 61.640 ;
        RECT 56.640 61.595 56.930 61.640 ;
        RECT 60.370 61.780 60.660 61.825 ;
        RECT 62.470 61.780 62.760 61.825 ;
        RECT 64.040 61.780 64.330 61.825 ;
        RECT 60.370 61.640 64.330 61.780 ;
        RECT 60.370 61.595 60.660 61.640 ;
        RECT 62.470 61.595 62.760 61.640 ;
        RECT 64.040 61.595 64.330 61.640 ;
        RECT 66.785 61.780 67.075 61.825 ;
        RECT 69.990 61.780 70.310 61.840 ;
        RECT 73.210 61.780 73.530 61.840 ;
        RECT 66.785 61.640 73.530 61.780 ;
        RECT 66.785 61.595 67.075 61.640 ;
        RECT 69.990 61.580 70.310 61.640 ;
        RECT 73.210 61.580 73.530 61.640 ;
        RECT 48.830 61.240 49.150 61.500 ;
        RECT 52.535 61.440 52.825 61.485 ;
        RECT 55.055 61.440 55.345 61.485 ;
        RECT 56.245 61.440 56.535 61.485 ;
        RECT 58.950 61.440 59.270 61.500 ;
        RECT 52.535 61.300 56.535 61.440 ;
        RECT 52.535 61.255 52.825 61.300 ;
        RECT 55.055 61.255 55.345 61.300 ;
        RECT 56.245 61.255 56.535 61.300 ;
        RECT 56.740 61.300 59.270 61.440 ;
        RECT 42.405 61.100 42.695 61.145 ;
        RECT 41.100 60.960 42.695 61.100 ;
        RECT 34.125 60.915 34.415 60.960 ;
        RECT 40.090 60.900 40.410 60.960 ;
        RECT 42.405 60.915 42.695 60.960 ;
        RECT 45.610 60.900 45.930 61.160 ;
        RECT 47.925 61.100 48.215 61.145 ;
        RECT 50.210 61.100 50.530 61.160 ;
        RECT 47.925 60.960 50.530 61.100 ;
        RECT 47.925 60.915 48.215 60.960 ;
        RECT 50.210 60.900 50.530 60.960 ;
        RECT 55.845 61.100 56.135 61.145 ;
        RECT 56.740 61.100 56.880 61.300 ;
        RECT 58.950 61.240 59.270 61.300 ;
        RECT 59.870 61.240 60.190 61.500 ;
        RECT 60.765 61.440 61.055 61.485 ;
        RECT 61.955 61.440 62.245 61.485 ;
        RECT 64.475 61.440 64.765 61.485 ;
        RECT 60.765 61.300 64.765 61.440 ;
        RECT 60.765 61.255 61.055 61.300 ;
        RECT 61.955 61.255 62.245 61.300 ;
        RECT 64.475 61.255 64.765 61.300 ;
        RECT 67.690 61.440 68.010 61.500 ;
        RECT 76.430 61.440 76.750 61.500 ;
        RECT 79.650 61.440 79.970 61.500 ;
        RECT 67.690 61.300 79.970 61.440 ;
        RECT 67.690 61.240 68.010 61.300 ;
        RECT 76.430 61.240 76.750 61.300 ;
        RECT 79.650 61.240 79.970 61.300 ;
        RECT 55.845 60.960 56.880 61.100 ;
        RECT 55.845 60.915 56.135 60.960 ;
        RECT 57.110 60.900 57.430 61.160 ;
        RECT 59.410 60.900 59.730 61.160 ;
        RECT 59.960 61.100 60.100 61.240 ;
        RECT 67.245 61.100 67.535 61.145 ;
        RECT 69.530 61.100 69.850 61.160 ;
        RECT 70.465 61.100 70.755 61.145 ;
        RECT 59.960 60.960 68.840 61.100 ;
        RECT 67.245 60.915 67.535 60.960 ;
        RECT 29.970 60.760 30.290 60.820 ;
        RECT 35.460 60.760 35.750 60.805 ;
        RECT 36.410 60.760 36.730 60.820 ;
        RECT 61.250 60.805 61.570 60.820 ;
        RECT 29.970 60.620 33.880 60.760 ;
        RECT 29.970 60.560 30.290 60.620 ;
        RECT 30.905 60.420 31.195 60.465 ;
        RECT 23.160 60.280 31.195 60.420 ;
        RECT 29.050 60.220 29.370 60.280 ;
        RECT 30.905 60.235 31.195 60.280 ;
        RECT 33.190 60.220 33.510 60.480 ;
        RECT 33.740 60.420 33.880 60.620 ;
        RECT 35.460 60.620 36.730 60.760 ;
        RECT 35.460 60.575 35.750 60.620 ;
        RECT 36.410 60.560 36.730 60.620 ;
        RECT 41.485 60.575 41.775 60.805 ;
        RECT 61.220 60.575 61.570 60.805 ;
        RECT 68.700 60.760 68.840 60.960 ;
        RECT 69.530 60.960 70.755 61.100 ;
        RECT 69.530 60.900 69.850 60.960 ;
        RECT 70.465 60.915 70.755 60.960 ;
        RECT 70.910 61.100 71.230 61.160 ;
        RECT 76.905 61.100 77.195 61.145 ;
        RECT 70.910 60.960 77.195 61.100 ;
        RECT 70.910 60.900 71.230 60.960 ;
        RECT 76.905 60.915 77.195 60.960 ;
        RECT 77.350 60.900 77.670 61.160 ;
        RECT 77.825 61.100 78.115 61.145 ;
        RECT 78.270 61.100 78.590 61.160 ;
        RECT 77.825 60.960 78.590 61.100 ;
        RECT 77.825 60.915 78.115 60.960 ;
        RECT 78.270 60.900 78.590 60.960 ;
        RECT 78.730 60.900 79.050 61.160 ;
        RECT 72.750 60.760 73.070 60.820 ;
        RECT 74.145 60.760 74.435 60.805 ;
        RECT 74.590 60.760 74.910 60.820 ;
        RECT 68.700 60.620 74.910 60.760 ;
        RECT 41.560 60.420 41.700 60.575 ;
        RECT 61.250 60.560 61.570 60.575 ;
        RECT 72.750 60.560 73.070 60.620 ;
        RECT 74.145 60.575 74.435 60.620 ;
        RECT 74.590 60.560 74.910 60.620 ;
        RECT 79.205 60.575 79.495 60.805 ;
        RECT 80.110 60.760 80.430 60.820 ;
        RECT 81.950 60.760 82.270 60.820 ;
        RECT 80.110 60.620 82.270 60.760 ;
        RECT 33.740 60.280 41.700 60.420 ;
        RECT 43.310 60.220 43.630 60.480 ;
        RECT 45.150 60.220 45.470 60.480 ;
        RECT 48.385 60.420 48.675 60.465 ;
        RECT 53.430 60.420 53.750 60.480 ;
        RECT 48.385 60.280 53.750 60.420 ;
        RECT 48.385 60.235 48.675 60.280 ;
        RECT 53.430 60.220 53.750 60.280 ;
        RECT 58.490 60.420 58.810 60.480 ;
        RECT 69.530 60.420 69.850 60.480 ;
        RECT 58.490 60.280 69.850 60.420 ;
        RECT 58.490 60.220 58.810 60.280 ;
        RECT 69.530 60.220 69.850 60.280 ;
        RECT 70.450 60.420 70.770 60.480 ;
        RECT 73.670 60.420 73.990 60.480 ;
        RECT 70.450 60.280 73.990 60.420 ;
        RECT 70.450 60.220 70.770 60.280 ;
        RECT 73.670 60.220 73.990 60.280 ;
        RECT 75.525 60.420 75.815 60.465 ;
        RECT 75.970 60.420 76.290 60.480 ;
        RECT 75.525 60.280 76.290 60.420 ;
        RECT 75.525 60.235 75.815 60.280 ;
        RECT 75.970 60.220 76.290 60.280 ;
        RECT 77.810 60.420 78.130 60.480 ;
        RECT 79.280 60.420 79.420 60.575 ;
        RECT 80.110 60.560 80.430 60.620 ;
        RECT 81.950 60.560 82.270 60.620 ;
        RECT 77.810 60.280 79.420 60.420 ;
        RECT 77.810 60.220 78.130 60.280 ;
        RECT 81.030 60.220 81.350 60.480 ;
        RECT 5.520 59.600 83.260 60.080 ;
        RECT 6.985 59.400 7.275 59.445 ;
        RECT 7.430 59.400 7.750 59.460 ;
        RECT 6.985 59.260 7.750 59.400 ;
        RECT 6.985 59.215 7.275 59.260 ;
        RECT 7.430 59.200 7.750 59.260 ;
        RECT 11.110 59.400 11.430 59.460 ;
        RECT 14.330 59.400 14.650 59.460 ;
        RECT 17.565 59.400 17.855 59.445 ;
        RECT 11.110 59.260 14.650 59.400 ;
        RECT 11.110 59.200 11.430 59.260 ;
        RECT 14.330 59.200 14.650 59.260 ;
        RECT 14.880 59.260 17.855 59.400 ;
        RECT 9.270 59.060 9.590 59.120 ;
        RECT 14.880 59.060 15.020 59.260 ;
        RECT 17.565 59.215 17.855 59.260 ;
        RECT 19.850 59.400 20.170 59.460 ;
        RECT 21.705 59.400 21.995 59.445 ;
        RECT 19.850 59.260 21.995 59.400 ;
        RECT 19.850 59.200 20.170 59.260 ;
        RECT 21.705 59.215 21.995 59.260 ;
        RECT 22.150 59.400 22.470 59.460 ;
        RECT 24.450 59.400 24.770 59.460 ;
        RECT 22.150 59.260 24.770 59.400 ;
        RECT 22.150 59.200 22.470 59.260 ;
        RECT 24.450 59.200 24.770 59.260 ;
        RECT 24.925 59.400 25.215 59.445 ;
        RECT 26.290 59.400 26.610 59.460 ;
        RECT 24.925 59.260 26.610 59.400 ;
        RECT 24.925 59.215 25.215 59.260 ;
        RECT 26.290 59.200 26.610 59.260 ;
        RECT 29.985 59.400 30.275 59.445 ;
        RECT 30.890 59.400 31.210 59.460 ;
        RECT 29.985 59.260 31.210 59.400 ;
        RECT 29.985 59.215 30.275 59.260 ;
        RECT 30.890 59.200 31.210 59.260 ;
        RECT 35.635 59.400 35.925 59.445 ;
        RECT 43.310 59.400 43.630 59.460 ;
        RECT 35.635 59.260 43.630 59.400 ;
        RECT 35.635 59.215 35.925 59.260 ;
        RECT 43.310 59.200 43.630 59.260 ;
        RECT 49.765 59.400 50.055 59.445 ;
        RECT 53.890 59.400 54.210 59.460 ;
        RECT 49.765 59.260 54.210 59.400 ;
        RECT 49.765 59.215 50.055 59.260 ;
        RECT 53.890 59.200 54.210 59.260 ;
        RECT 59.410 59.400 59.730 59.460 ;
        RECT 67.690 59.400 68.010 59.460 ;
        RECT 59.410 59.260 68.010 59.400 ;
        RECT 59.410 59.200 59.730 59.260 ;
        RECT 67.690 59.200 68.010 59.260 ;
        RECT 68.165 59.400 68.455 59.445 ;
        RECT 68.610 59.400 68.930 59.460 ;
        RECT 75.510 59.400 75.830 59.460 ;
        RECT 68.165 59.260 68.930 59.400 ;
        RECT 68.165 59.215 68.455 59.260 ;
        RECT 68.610 59.200 68.930 59.260 ;
        RECT 69.160 59.260 75.830 59.400 ;
        RECT 9.270 58.920 15.020 59.060 ;
        RECT 15.185 59.060 15.475 59.105 ;
        RECT 15.710 59.060 16.030 59.120 ;
        RECT 15.185 58.920 16.030 59.060 ;
        RECT 9.270 58.860 9.590 58.920 ;
        RECT 15.185 58.875 15.475 58.920 ;
        RECT 15.710 58.860 16.030 58.920 ;
        RECT 16.170 58.860 16.490 59.120 ;
        RECT 23.990 59.060 24.310 59.120 ;
        RECT 16.720 58.920 24.310 59.060 ;
        RECT 12.605 58.720 12.895 58.765 ;
        RECT 13.885 58.740 14.175 58.765 ;
        RECT 13.885 58.720 15.020 58.740 ;
        RECT 16.720 58.720 16.860 58.920 ;
        RECT 23.990 58.860 24.310 58.920 ;
        RECT 25.370 59.060 25.690 59.120 ;
        RECT 25.845 59.060 26.135 59.105 ;
        RECT 25.370 58.920 26.135 59.060 ;
        RECT 25.370 58.860 25.690 58.920 ;
        RECT 25.845 58.875 26.135 58.920 ;
        RECT 32.270 59.060 32.590 59.120 ;
        RECT 34.585 59.060 34.875 59.105 ;
        RECT 32.270 58.920 34.875 59.060 ;
        RECT 32.270 58.860 32.590 58.920 ;
        RECT 34.585 58.875 34.875 58.920 ;
        RECT 40.520 59.060 40.810 59.105 ;
        RECT 41.470 59.060 41.790 59.120 ;
        RECT 40.520 58.920 41.790 59.060 ;
        RECT 40.520 58.875 40.810 58.920 ;
        RECT 41.470 58.860 41.790 58.920 ;
        RECT 49.290 58.860 49.610 59.120 ;
        RECT 55.440 59.060 55.730 59.105 ;
        RECT 57.570 59.060 57.890 59.120 ;
        RECT 61.710 59.105 62.030 59.120 ;
        RECT 61.680 59.060 62.030 59.105 ;
        RECT 55.440 58.920 57.890 59.060 ;
        RECT 61.515 58.920 62.030 59.060 ;
        RECT 55.440 58.875 55.730 58.920 ;
        RECT 57.570 58.860 57.890 58.920 ;
        RECT 61.680 58.875 62.030 58.920 ;
        RECT 61.710 58.860 62.030 58.875 ;
        RECT 12.605 58.580 13.640 58.720 ;
        RECT 12.605 58.535 12.895 58.580 ;
        RECT 9.295 58.380 9.585 58.425 ;
        RECT 11.815 58.380 12.105 58.425 ;
        RECT 13.005 58.380 13.295 58.425 ;
        RECT 9.295 58.240 13.295 58.380 ;
        RECT 13.500 58.380 13.640 58.580 ;
        RECT 13.885 58.600 16.860 58.720 ;
        RECT 13.885 58.535 14.175 58.600 ;
        RECT 14.880 58.580 16.860 58.600 ;
        RECT 17.090 58.520 17.410 58.780 ;
        RECT 17.550 58.720 17.870 58.780 ;
        RECT 18.945 58.720 19.235 58.765 ;
        RECT 17.550 58.580 19.235 58.720 ;
        RECT 17.550 58.520 17.870 58.580 ;
        RECT 18.945 58.535 19.235 58.580 ;
        RECT 19.850 58.720 20.170 58.780 ;
        RECT 20.325 58.720 20.615 58.765 ;
        RECT 19.850 58.580 20.615 58.720 ;
        RECT 19.850 58.520 20.170 58.580 ;
        RECT 20.325 58.535 20.615 58.580 ;
        RECT 20.770 58.520 21.090 58.780 ;
        RECT 22.165 58.535 22.455 58.765 ;
        RECT 23.085 58.720 23.375 58.765 ;
        RECT 22.700 58.580 23.375 58.720 ;
        RECT 22.240 58.380 22.380 58.535 ;
        RECT 13.500 58.240 14.560 58.380 ;
        RECT 9.295 58.195 9.585 58.240 ;
        RECT 11.815 58.195 12.105 58.240 ;
        RECT 13.005 58.195 13.295 58.240 ;
        RECT 14.420 58.085 14.560 58.240 ;
        RECT 14.880 58.240 22.380 58.380 ;
        RECT 9.730 58.040 10.020 58.085 ;
        RECT 11.300 58.040 11.590 58.085 ;
        RECT 13.400 58.040 13.690 58.085 ;
        RECT 9.730 57.900 13.690 58.040 ;
        RECT 9.730 57.855 10.020 57.900 ;
        RECT 11.300 57.855 11.590 57.900 ;
        RECT 13.400 57.855 13.690 57.900 ;
        RECT 14.345 57.855 14.635 58.085 ;
        RECT 14.880 57.760 15.020 58.240 ;
        RECT 19.390 58.040 19.710 58.100 ;
        RECT 22.700 58.040 22.840 58.580 ;
        RECT 23.085 58.535 23.375 58.580 ;
        RECT 23.530 58.520 23.850 58.780 ;
        RECT 27.685 58.720 27.975 58.765 ;
        RECT 26.380 58.580 27.975 58.720 ;
        RECT 19.390 57.900 22.840 58.040 ;
        RECT 23.620 58.040 23.760 58.520 ;
        RECT 26.380 58.100 26.520 58.580 ;
        RECT 27.685 58.535 27.975 58.580 ;
        RECT 29.050 58.520 29.370 58.780 ;
        RECT 30.445 58.535 30.735 58.765 ;
        RECT 33.205 58.720 33.495 58.765 ;
        RECT 35.490 58.720 35.810 58.780 ;
        RECT 33.205 58.580 35.810 58.720 ;
        RECT 33.205 58.535 33.495 58.580 ;
        RECT 28.130 58.380 28.450 58.440 ;
        RECT 30.520 58.380 30.660 58.535 ;
        RECT 35.490 58.520 35.810 58.580 ;
        RECT 39.185 58.720 39.475 58.765 ;
        RECT 39.630 58.720 39.950 58.780 ;
        RECT 39.185 58.580 39.950 58.720 ;
        RECT 39.185 58.535 39.475 58.580 ;
        RECT 39.630 58.520 39.950 58.580 ;
        RECT 41.930 58.720 42.250 58.780 ;
        RECT 41.930 58.580 44.460 58.720 ;
        RECT 41.930 58.520 42.250 58.580 ;
        RECT 44.320 58.440 44.460 58.580 ;
        RECT 46.530 58.520 46.850 58.780 ;
        RECT 47.450 58.520 47.770 58.780 ;
        RECT 56.665 58.720 56.955 58.765 ;
        RECT 57.110 58.720 57.430 58.780 ;
        RECT 60.330 58.720 60.650 58.780 ;
        RECT 69.160 58.765 69.300 59.260 ;
        RECT 75.510 59.200 75.830 59.260 ;
        RECT 74.130 59.060 74.450 59.120 ;
        RECT 70.080 58.920 74.450 59.060 ;
        RECT 56.665 58.580 60.650 58.720 ;
        RECT 56.665 58.535 56.955 58.580 ;
        RECT 57.110 58.520 57.430 58.580 ;
        RECT 60.330 58.520 60.650 58.580 ;
        RECT 69.085 58.535 69.375 58.765 ;
        RECT 69.530 58.720 69.850 58.780 ;
        RECT 70.080 58.765 70.220 58.920 ;
        RECT 74.130 58.860 74.450 58.920 ;
        RECT 70.005 58.720 70.295 58.765 ;
        RECT 69.530 58.580 70.295 58.720 ;
        RECT 69.530 58.520 69.850 58.580 ;
        RECT 70.005 58.535 70.295 58.580 ;
        RECT 70.450 58.520 70.770 58.780 ;
        RECT 71.830 58.720 72.150 58.780 ;
        RECT 71.000 58.580 72.150 58.720 ;
        RECT 28.130 58.240 30.660 58.380 ;
        RECT 40.065 58.380 40.355 58.425 ;
        RECT 41.255 58.380 41.545 58.425 ;
        RECT 43.775 58.380 44.065 58.425 ;
        RECT 40.065 58.240 44.065 58.380 ;
        RECT 28.130 58.180 28.450 58.240 ;
        RECT 40.065 58.195 40.355 58.240 ;
        RECT 41.255 58.195 41.545 58.240 ;
        RECT 43.775 58.195 44.065 58.240 ;
        RECT 44.230 58.380 44.550 58.440 ;
        RECT 47.540 58.380 47.680 58.520 ;
        RECT 44.230 58.240 47.680 58.380 ;
        RECT 52.075 58.380 52.365 58.425 ;
        RECT 54.595 58.380 54.885 58.425 ;
        RECT 55.785 58.380 56.075 58.425 ;
        RECT 52.075 58.240 56.075 58.380 ;
        RECT 44.230 58.180 44.550 58.240 ;
        RECT 52.075 58.195 52.365 58.240 ;
        RECT 54.595 58.195 54.885 58.240 ;
        RECT 55.785 58.195 56.075 58.240 ;
        RECT 61.225 58.380 61.515 58.425 ;
        RECT 62.415 58.380 62.705 58.425 ;
        RECT 64.935 58.380 65.225 58.425 ;
        RECT 61.225 58.240 65.225 58.380 ;
        RECT 61.225 58.195 61.515 58.240 ;
        RECT 62.415 58.195 62.705 58.240 ;
        RECT 64.935 58.195 65.225 58.240 ;
        RECT 26.290 58.040 26.610 58.100 ;
        RECT 23.620 57.900 26.610 58.040 ;
        RECT 19.390 57.840 19.710 57.900 ;
        RECT 26.290 57.840 26.610 57.900 ;
        RECT 34.125 58.040 34.415 58.085 ;
        RECT 35.950 58.040 36.270 58.100 ;
        RECT 34.125 57.900 36.270 58.040 ;
        RECT 34.125 57.855 34.415 57.900 ;
        RECT 35.950 57.840 36.270 57.900 ;
        RECT 36.410 57.840 36.730 58.100 ;
        RECT 39.670 58.040 39.960 58.085 ;
        RECT 41.770 58.040 42.060 58.085 ;
        RECT 43.340 58.040 43.630 58.085 ;
        RECT 39.670 57.900 43.630 58.040 ;
        RECT 39.670 57.855 39.960 57.900 ;
        RECT 41.770 57.855 42.060 57.900 ;
        RECT 43.340 57.855 43.630 57.900 ;
        RECT 52.510 58.040 52.800 58.085 ;
        RECT 54.080 58.040 54.370 58.085 ;
        RECT 56.180 58.040 56.470 58.085 ;
        RECT 52.510 57.900 56.470 58.040 ;
        RECT 52.510 57.855 52.800 57.900 ;
        RECT 54.080 57.855 54.370 57.900 ;
        RECT 56.180 57.855 56.470 57.900 ;
        RECT 60.830 58.040 61.120 58.085 ;
        RECT 62.930 58.040 63.220 58.085 ;
        RECT 64.500 58.040 64.790 58.085 ;
        RECT 60.830 57.900 64.790 58.040 ;
        RECT 60.830 57.855 61.120 57.900 ;
        RECT 62.930 57.855 63.220 57.900 ;
        RECT 64.500 57.855 64.790 57.900 ;
        RECT 67.245 58.040 67.535 58.085 ;
        RECT 69.990 58.040 70.310 58.100 ;
        RECT 67.245 57.900 70.310 58.040 ;
        RECT 67.245 57.855 67.535 57.900 ;
        RECT 69.990 57.840 70.310 57.900 ;
        RECT 14.790 57.500 15.110 57.760 ;
        RECT 15.250 57.700 15.570 57.760 ;
        RECT 17.090 57.700 17.410 57.760 ;
        RECT 15.250 57.560 17.410 57.700 ;
        RECT 15.250 57.500 15.570 57.560 ;
        RECT 17.090 57.500 17.410 57.560 ;
        RECT 17.550 57.700 17.870 57.760 ;
        RECT 22.165 57.700 22.455 57.745 ;
        RECT 17.550 57.560 22.455 57.700 ;
        RECT 17.550 57.500 17.870 57.560 ;
        RECT 22.165 57.515 22.455 57.560 ;
        RECT 25.845 57.700 26.135 57.745 ;
        RECT 28.145 57.700 28.435 57.745 ;
        RECT 25.845 57.560 28.435 57.700 ;
        RECT 25.845 57.515 26.135 57.560 ;
        RECT 28.145 57.515 28.435 57.560 ;
        RECT 34.570 57.700 34.890 57.760 ;
        RECT 35.505 57.700 35.795 57.745 ;
        RECT 34.570 57.560 35.795 57.700 ;
        RECT 34.570 57.500 34.890 57.560 ;
        RECT 35.505 57.515 35.795 57.560 ;
        RECT 46.070 57.700 46.390 57.760 ;
        RECT 49.750 57.700 50.070 57.760 ;
        RECT 46.070 57.560 50.070 57.700 ;
        RECT 71.000 57.700 71.140 58.580 ;
        RECT 71.830 58.520 72.150 58.580 ;
        RECT 72.765 58.535 73.055 58.765 ;
        RECT 71.370 58.380 71.690 58.440 ;
        RECT 72.840 58.380 72.980 58.535 ;
        RECT 74.590 58.520 74.910 58.780 ;
        RECT 75.885 58.720 76.175 58.765 ;
        RECT 75.140 58.580 76.175 58.720 ;
        RECT 71.370 58.240 72.980 58.380 ;
        RECT 74.130 58.380 74.450 58.440 ;
        RECT 75.140 58.380 75.280 58.580 ;
        RECT 75.885 58.535 76.175 58.580 ;
        RECT 74.130 58.240 75.280 58.380 ;
        RECT 75.485 58.380 75.775 58.425 ;
        RECT 76.675 58.380 76.965 58.425 ;
        RECT 79.195 58.380 79.485 58.425 ;
        RECT 75.485 58.240 79.485 58.380 ;
        RECT 71.370 58.180 71.690 58.240 ;
        RECT 74.130 58.180 74.450 58.240 ;
        RECT 75.485 58.195 75.775 58.240 ;
        RECT 76.675 58.195 76.965 58.240 ;
        RECT 79.195 58.195 79.485 58.240 ;
        RECT 75.090 58.040 75.380 58.085 ;
        RECT 77.190 58.040 77.480 58.085 ;
        RECT 78.760 58.040 79.050 58.085 ;
        RECT 75.090 57.900 79.050 58.040 ;
        RECT 75.090 57.855 75.380 57.900 ;
        RECT 77.190 57.855 77.480 57.900 ;
        RECT 78.760 57.855 79.050 57.900 ;
        RECT 71.385 57.700 71.675 57.745 ;
        RECT 71.000 57.560 71.675 57.700 ;
        RECT 46.070 57.500 46.390 57.560 ;
        RECT 49.750 57.500 50.070 57.560 ;
        RECT 71.385 57.515 71.675 57.560 ;
        RECT 71.830 57.700 72.150 57.760 ;
        RECT 73.685 57.700 73.975 57.745 ;
        RECT 71.830 57.560 73.975 57.700 ;
        RECT 71.830 57.500 72.150 57.560 ;
        RECT 73.685 57.515 73.975 57.560 ;
        RECT 75.510 57.700 75.830 57.760 ;
        RECT 80.110 57.700 80.430 57.760 ;
        RECT 81.505 57.700 81.795 57.745 ;
        RECT 75.510 57.560 81.795 57.700 ;
        RECT 75.510 57.500 75.830 57.560 ;
        RECT 80.110 57.500 80.430 57.560 ;
        RECT 81.505 57.515 81.795 57.560 ;
        RECT 5.520 56.880 83.260 57.360 ;
        RECT 8.810 56.680 9.130 56.740 ;
        RECT 8.810 56.540 12.260 56.680 ;
        RECT 8.810 56.480 9.130 56.540 ;
        RECT 7.470 56.340 7.760 56.385 ;
        RECT 9.570 56.340 9.860 56.385 ;
        RECT 11.140 56.340 11.430 56.385 ;
        RECT 7.470 56.200 11.430 56.340 ;
        RECT 7.470 56.155 7.760 56.200 ;
        RECT 9.570 56.155 9.860 56.200 ;
        RECT 11.140 56.155 11.430 56.200 ;
        RECT 7.865 56.000 8.155 56.045 ;
        RECT 9.055 56.000 9.345 56.045 ;
        RECT 11.575 56.000 11.865 56.045 ;
        RECT 7.865 55.860 11.865 56.000 ;
        RECT 12.120 56.000 12.260 56.540 ;
        RECT 13.870 56.480 14.190 56.740 ;
        RECT 14.345 56.680 14.635 56.725 ;
        RECT 15.710 56.680 16.030 56.740 ;
        RECT 14.345 56.540 16.030 56.680 ;
        RECT 14.345 56.495 14.635 56.540 ;
        RECT 15.710 56.480 16.030 56.540 ;
        RECT 26.290 56.480 26.610 56.740 ;
        RECT 27.225 56.680 27.515 56.725 ;
        RECT 28.590 56.680 28.910 56.740 ;
        RECT 30.890 56.680 31.210 56.740 ;
        RECT 27.225 56.540 31.210 56.680 ;
        RECT 27.225 56.495 27.515 56.540 ;
        RECT 28.590 56.480 28.910 56.540 ;
        RECT 30.890 56.480 31.210 56.540 ;
        RECT 42.850 56.680 43.170 56.740 ;
        RECT 42.850 56.540 43.540 56.680 ;
        RECT 42.850 56.480 43.170 56.540 ;
        RECT 22.165 56.340 22.455 56.385 ;
        RECT 23.070 56.340 23.390 56.400 ;
        RECT 22.165 56.200 23.390 56.340 ;
        RECT 22.165 56.155 22.455 56.200 ;
        RECT 23.070 56.140 23.390 56.200 ;
        RECT 23.545 56.000 23.835 56.045 ;
        RECT 32.730 56.000 33.050 56.060 ;
        RECT 12.120 55.860 14.560 56.000 ;
        RECT 7.865 55.815 8.155 55.860 ;
        RECT 9.055 55.815 9.345 55.860 ;
        RECT 11.575 55.815 11.865 55.860 ;
        RECT 6.985 55.660 7.275 55.705 ;
        RECT 13.870 55.660 14.190 55.720 ;
        RECT 14.420 55.705 14.560 55.860 ;
        RECT 23.545 55.860 33.050 56.000 ;
        RECT 43.400 56.000 43.540 56.540 ;
        RECT 44.690 56.480 45.010 56.740 ;
        RECT 45.610 56.680 45.930 56.740 ;
        RECT 48.845 56.680 49.135 56.725 ;
        RECT 45.610 56.540 49.135 56.680 ;
        RECT 45.610 56.480 45.930 56.540 ;
        RECT 48.845 56.495 49.135 56.540 ;
        RECT 49.765 56.680 50.055 56.725 ;
        RECT 52.510 56.680 52.830 56.740 ;
        RECT 66.310 56.680 66.630 56.740 ;
        RECT 49.765 56.540 52.830 56.680 ;
        RECT 49.765 56.495 50.055 56.540 ;
        RECT 52.510 56.480 52.830 56.540 ;
        RECT 54.440 56.540 66.630 56.680 ;
        RECT 43.785 56.340 44.075 56.385 ;
        RECT 48.370 56.340 48.690 56.400 ;
        RECT 43.785 56.200 48.690 56.340 ;
        RECT 43.785 56.155 44.075 56.200 ;
        RECT 48.370 56.140 48.690 56.200 ;
        RECT 46.675 56.000 46.965 56.045 ;
        RECT 54.440 56.000 54.580 56.540 ;
        RECT 66.310 56.480 66.630 56.540 ;
        RECT 66.785 56.680 67.075 56.725 ;
        RECT 67.230 56.680 67.550 56.740 ;
        RECT 66.785 56.540 67.550 56.680 ;
        RECT 66.785 56.495 67.075 56.540 ;
        RECT 67.230 56.480 67.550 56.540 ;
        RECT 70.910 56.680 71.230 56.740 ;
        RECT 72.750 56.680 73.070 56.740 ;
        RECT 70.910 56.540 73.070 56.680 ;
        RECT 70.910 56.480 71.230 56.540 ;
        RECT 72.750 56.480 73.070 56.540 ;
        RECT 74.130 56.480 74.450 56.740 ;
        RECT 81.030 56.680 81.350 56.740 ;
        RECT 74.680 56.540 81.350 56.680 ;
        RECT 74.680 56.340 74.820 56.540 ;
        RECT 81.030 56.480 81.350 56.540 ;
        RECT 71.920 56.200 74.820 56.340 ;
        RECT 75.090 56.340 75.380 56.385 ;
        RECT 77.190 56.340 77.480 56.385 ;
        RECT 78.760 56.340 79.050 56.385 ;
        RECT 75.090 56.200 79.050 56.340 ;
        RECT 69.530 56.000 69.850 56.060 ;
        RECT 43.400 55.860 45.840 56.000 ;
        RECT 23.545 55.815 23.835 55.860 ;
        RECT 32.730 55.800 33.050 55.860 ;
        RECT 6.985 55.520 14.190 55.660 ;
        RECT 6.985 55.475 7.275 55.520 ;
        RECT 13.870 55.460 14.190 55.520 ;
        RECT 14.345 55.475 14.635 55.705 ;
        RECT 15.265 55.475 15.555 55.705 ;
        RECT 20.770 55.660 21.090 55.720 ;
        RECT 21.705 55.660 21.995 55.705 ;
        RECT 20.770 55.520 21.995 55.660 ;
        RECT 8.350 55.365 8.670 55.380 ;
        RECT 8.320 55.135 8.670 55.365 ;
        RECT 8.350 55.120 8.670 55.135 ;
        RECT 11.110 55.320 11.430 55.380 ;
        RECT 15.340 55.320 15.480 55.475 ;
        RECT 20.770 55.460 21.090 55.520 ;
        RECT 21.705 55.475 21.995 55.520 ;
        RECT 22.610 55.460 22.930 55.720 ;
        RECT 23.085 55.475 23.375 55.705 ;
        RECT 24.005 55.660 24.295 55.705 ;
        RECT 24.450 55.660 24.770 55.720 ;
        RECT 28.590 55.660 28.910 55.720 ;
        RECT 45.700 55.705 45.840 55.860 ;
        RECT 46.675 55.860 54.580 56.000 ;
        RECT 66.400 55.860 69.850 56.000 ;
        RECT 46.675 55.815 46.965 55.860 ;
        RECT 24.005 55.520 28.910 55.660 ;
        RECT 24.005 55.475 24.295 55.520 ;
        RECT 11.110 55.180 15.480 55.320 ;
        RECT 15.710 55.320 16.030 55.380 ;
        RECT 18.930 55.320 19.250 55.380 ;
        RECT 15.710 55.180 19.250 55.320 ;
        RECT 23.160 55.320 23.300 55.475 ;
        RECT 24.450 55.460 24.770 55.520 ;
        RECT 28.590 55.460 28.910 55.520 ;
        RECT 45.625 55.660 45.915 55.705 ;
        RECT 46.070 55.660 46.390 55.720 ;
        RECT 45.625 55.520 46.390 55.660 ;
        RECT 45.625 55.475 45.915 55.520 ;
        RECT 46.070 55.460 46.390 55.520 ;
        RECT 47.450 55.460 47.770 55.720 ;
        RECT 51.130 55.660 51.450 55.720 ;
        RECT 58.490 55.660 58.810 55.720 ;
        RECT 66.400 55.705 66.540 55.860 ;
        RECT 69.530 55.800 69.850 55.860 ;
        RECT 51.130 55.520 58.810 55.660 ;
        RECT 51.130 55.460 51.450 55.520 ;
        RECT 58.490 55.460 58.810 55.520 ;
        RECT 66.325 55.475 66.615 55.705 ;
        RECT 67.245 55.660 67.535 55.705 ;
        RECT 68.625 55.660 68.915 55.705 ;
        RECT 69.070 55.660 69.390 55.720 ;
        RECT 71.920 55.705 72.060 56.200 ;
        RECT 75.090 56.155 75.380 56.200 ;
        RECT 77.190 56.155 77.480 56.200 ;
        RECT 78.760 56.155 79.050 56.200 ;
        RECT 79.650 56.340 79.970 56.400 ;
        RECT 81.505 56.340 81.795 56.385 ;
        RECT 79.650 56.200 81.795 56.340 ;
        RECT 79.650 56.140 79.970 56.200 ;
        RECT 81.505 56.155 81.795 56.200 ;
        RECT 74.590 55.800 74.910 56.060 ;
        RECT 75.485 56.000 75.775 56.045 ;
        RECT 76.675 56.000 76.965 56.045 ;
        RECT 79.195 56.000 79.485 56.045 ;
        RECT 75.485 55.860 79.485 56.000 ;
        RECT 75.485 55.815 75.775 55.860 ;
        RECT 76.675 55.815 76.965 55.860 ;
        RECT 79.195 55.815 79.485 55.860 ;
        RECT 67.245 55.520 69.390 55.660 ;
        RECT 67.245 55.475 67.535 55.520 ;
        RECT 68.625 55.475 68.915 55.520 ;
        RECT 69.070 55.460 69.390 55.520 ;
        RECT 70.925 55.475 71.215 55.705 ;
        RECT 71.845 55.475 72.135 55.705 ;
        RECT 23.530 55.320 23.850 55.380 ;
        RECT 27.145 55.320 27.435 55.365 ;
        RECT 27.670 55.320 27.990 55.380 ;
        RECT 23.160 55.180 27.990 55.320 ;
        RECT 11.110 55.120 11.430 55.180 ;
        RECT 15.710 55.120 16.030 55.180 ;
        RECT 18.930 55.120 19.250 55.180 ;
        RECT 23.530 55.120 23.850 55.180 ;
        RECT 27.145 55.135 27.435 55.180 ;
        RECT 27.670 55.120 27.990 55.180 ;
        RECT 28.145 55.320 28.435 55.365 ;
        RECT 29.050 55.320 29.370 55.380 ;
        RECT 28.145 55.180 29.370 55.320 ;
        RECT 28.145 55.135 28.435 55.180 ;
        RECT 29.050 55.120 29.370 55.180 ;
        RECT 41.945 55.320 42.235 55.365 ;
        RECT 44.230 55.320 44.550 55.380 ;
        RECT 41.945 55.180 44.550 55.320 ;
        RECT 41.945 55.135 42.235 55.180 ;
        RECT 44.230 55.120 44.550 55.180 ;
        RECT 45.150 55.320 45.470 55.380 ;
        RECT 47.925 55.320 48.215 55.365 ;
        RECT 60.330 55.320 60.650 55.380 ;
        RECT 62.185 55.320 62.475 55.365 ;
        RECT 45.150 55.180 47.680 55.320 ;
        RECT 45.150 55.120 45.470 55.180 ;
        RECT 10.190 54.980 10.510 55.040 ;
        RECT 12.950 54.980 13.270 55.040 ;
        RECT 10.190 54.840 13.270 54.980 ;
        RECT 10.190 54.780 10.510 54.840 ;
        RECT 12.950 54.780 13.270 54.840 ;
        RECT 23.990 54.980 24.310 55.040 ;
        RECT 25.370 54.980 25.690 55.040 ;
        RECT 40.550 54.980 40.870 55.040 ;
        RECT 23.990 54.840 40.870 54.980 ;
        RECT 23.990 54.780 24.310 54.840 ;
        RECT 25.370 54.780 25.690 54.840 ;
        RECT 40.550 54.780 40.870 54.840 ;
        RECT 42.995 54.980 43.285 55.025 ;
        RECT 43.770 54.980 44.090 55.040 ;
        RECT 45.610 54.980 45.930 55.040 ;
        RECT 42.995 54.840 45.930 54.980 ;
        RECT 47.540 54.980 47.680 55.180 ;
        RECT 47.925 55.180 58.260 55.320 ;
        RECT 47.925 55.135 48.215 55.180 ;
        RECT 48.925 54.980 49.215 55.025 ;
        RECT 47.540 54.840 49.215 54.980 ;
        RECT 58.120 54.980 58.260 55.180 ;
        RECT 60.330 55.180 62.475 55.320 ;
        RECT 60.330 55.120 60.650 55.180 ;
        RECT 62.185 55.135 62.475 55.180 ;
        RECT 67.705 55.320 67.995 55.365 ;
        RECT 69.530 55.320 69.850 55.380 ;
        RECT 67.705 55.180 69.850 55.320 ;
        RECT 67.705 55.135 67.995 55.180 ;
        RECT 69.530 55.120 69.850 55.180 ;
        RECT 63.550 54.980 63.870 55.040 ;
        RECT 70.450 54.980 70.770 55.040 ;
        RECT 71.000 54.980 71.140 55.475 ;
        RECT 72.290 55.460 72.610 55.720 ;
        RECT 72.750 55.460 73.070 55.720 ;
        RECT 75.970 55.705 76.290 55.720 ;
        RECT 75.940 55.660 76.290 55.705 ;
        RECT 75.775 55.520 76.290 55.660 ;
        RECT 75.940 55.475 76.290 55.520 ;
        RECT 75.970 55.460 76.290 55.475 ;
        RECT 71.370 55.320 71.690 55.380 ;
        RECT 76.430 55.320 76.750 55.380 ;
        RECT 71.370 55.180 76.750 55.320 ;
        RECT 71.370 55.120 71.690 55.180 ;
        RECT 76.430 55.120 76.750 55.180 ;
        RECT 78.730 54.980 79.050 55.040 ;
        RECT 58.120 54.840 79.050 54.980 ;
        RECT 42.995 54.795 43.285 54.840 ;
        RECT 43.770 54.780 44.090 54.840 ;
        RECT 45.610 54.780 45.930 54.840 ;
        RECT 48.925 54.795 49.215 54.840 ;
        RECT 63.550 54.780 63.870 54.840 ;
        RECT 70.450 54.780 70.770 54.840 ;
        RECT 78.730 54.780 79.050 54.840 ;
        RECT 5.520 54.160 83.260 54.640 ;
        RECT 8.350 53.760 8.670 54.020 ;
        RECT 16.170 53.960 16.490 54.020 ;
        RECT 11.200 53.820 16.490 53.960 ;
        RECT 9.205 53.620 9.495 53.665 ;
        RECT 9.205 53.480 9.960 53.620 ;
        RECT 9.205 53.435 9.495 53.480 ;
        RECT 9.820 52.940 9.960 53.480 ;
        RECT 10.190 53.420 10.510 53.680 ;
        RECT 11.200 53.325 11.340 53.820 ;
        RECT 16.170 53.760 16.490 53.820 ;
        RECT 35.950 53.960 36.270 54.020 ;
        RECT 37.345 53.960 37.635 54.005 ;
        RECT 35.950 53.820 37.635 53.960 ;
        RECT 35.950 53.760 36.270 53.820 ;
        RECT 37.345 53.775 37.635 53.820 ;
        RECT 68.150 53.760 68.470 54.020 ;
        RECT 75.050 53.960 75.370 54.020 ;
        RECT 69.160 53.820 75.370 53.960 ;
        RECT 12.045 53.620 12.335 53.665 ;
        RECT 12.950 53.620 13.270 53.680 ;
        RECT 12.045 53.480 13.270 53.620 ;
        RECT 12.045 53.435 12.335 53.480 ;
        RECT 12.950 53.420 13.270 53.480 ;
        RECT 28.590 53.420 28.910 53.680 ;
        RECT 38.265 53.620 38.555 53.665 ;
        RECT 43.310 53.620 43.630 53.680 ;
        RECT 38.265 53.480 43.630 53.620 ;
        RECT 38.265 53.435 38.555 53.480 ;
        RECT 43.310 53.420 43.630 53.480 ;
        RECT 45.625 53.620 45.915 53.665 ;
        RECT 45.625 53.480 48.600 53.620 ;
        RECT 45.625 53.435 45.915 53.480 ;
        RECT 11.125 53.095 11.415 53.325 ;
        RECT 11.570 53.280 11.890 53.340 ;
        RECT 12.505 53.280 12.795 53.325 ;
        RECT 11.570 53.140 12.795 53.280 ;
        RECT 11.570 53.080 11.890 53.140 ;
        RECT 12.505 53.095 12.795 53.140 ;
        RECT 13.425 53.280 13.715 53.325 ;
        RECT 17.550 53.280 17.870 53.340 ;
        RECT 13.425 53.140 17.870 53.280 ;
        RECT 13.425 53.095 13.715 53.140 ;
        RECT 17.550 53.080 17.870 53.140 ;
        RECT 20.310 53.080 20.630 53.340 ;
        RECT 23.530 53.080 23.850 53.340 ;
        RECT 24.910 53.080 25.230 53.340 ;
        RECT 26.765 53.095 27.055 53.325 ;
        RECT 27.685 53.280 27.975 53.325 ;
        RECT 28.130 53.280 28.450 53.340 ;
        RECT 27.685 53.140 28.450 53.280 ;
        RECT 27.685 53.095 27.975 53.140 ;
        RECT 12.965 52.940 13.255 52.985 ;
        RECT 9.820 52.800 13.255 52.940 ;
        RECT 25.000 52.940 25.140 53.080 ;
        RECT 26.290 52.940 26.610 53.000 ;
        RECT 25.000 52.800 26.610 52.940 ;
        RECT 12.965 52.755 13.255 52.800 ;
        RECT 26.290 52.740 26.610 52.800 ;
        RECT 17.090 52.600 17.410 52.660 ;
        RECT 20.325 52.600 20.615 52.645 ;
        RECT 17.090 52.460 20.615 52.600 ;
        RECT 17.090 52.400 17.410 52.460 ;
        RECT 20.325 52.415 20.615 52.460 ;
        RECT 22.610 52.600 22.930 52.660 ;
        RECT 23.990 52.600 24.310 52.660 ;
        RECT 26.840 52.600 26.980 53.095 ;
        RECT 28.130 53.080 28.450 53.140 ;
        RECT 36.870 53.080 37.190 53.340 ;
        RECT 41.485 53.095 41.775 53.325 ;
        RECT 42.405 53.280 42.695 53.325 ;
        RECT 45.150 53.280 45.470 53.340 ;
        RECT 48.460 53.325 48.600 53.480 ;
        RECT 42.405 53.140 45.470 53.280 ;
        RECT 42.405 53.095 42.695 53.140 ;
        RECT 41.560 52.940 41.700 53.095 ;
        RECT 45.150 53.080 45.470 53.140 ;
        RECT 46.545 53.280 46.835 53.325 ;
        RECT 48.385 53.280 48.675 53.325 ;
        RECT 48.830 53.280 49.150 53.340 ;
        RECT 46.545 53.140 48.140 53.280 ;
        RECT 46.545 53.095 46.835 53.140 ;
        RECT 42.850 52.940 43.170 53.000 ;
        RECT 41.560 52.800 43.170 52.940 ;
        RECT 42.850 52.740 43.170 52.800 ;
        RECT 44.230 52.940 44.550 53.000 ;
        RECT 47.005 52.940 47.295 52.985 ;
        RECT 44.230 52.800 47.295 52.940 ;
        RECT 48.000 52.940 48.140 53.140 ;
        RECT 48.385 53.140 49.150 53.280 ;
        RECT 48.385 53.095 48.675 53.140 ;
        RECT 48.830 53.080 49.150 53.140 ;
        RECT 60.330 53.080 60.650 53.340 ;
        RECT 69.160 53.325 69.300 53.820 ;
        RECT 75.050 53.760 75.370 53.820 ;
        RECT 76.430 53.960 76.750 54.020 ;
        RECT 79.190 53.960 79.510 54.020 ;
        RECT 81.505 53.960 81.795 54.005 ;
        RECT 76.430 53.820 81.795 53.960 ;
        RECT 76.430 53.760 76.750 53.820 ;
        RECT 79.190 53.760 79.510 53.820 ;
        RECT 81.505 53.775 81.795 53.820 ;
        RECT 74.145 53.620 74.435 53.665 ;
        RECT 75.830 53.620 76.120 53.665 ;
        RECT 74.145 53.480 76.120 53.620 ;
        RECT 74.145 53.435 74.435 53.480 ;
        RECT 75.830 53.435 76.120 53.480 ;
        RECT 67.245 53.095 67.535 53.325 ;
        RECT 69.085 53.095 69.375 53.325 ;
        RECT 70.450 53.280 70.770 53.340 ;
        RECT 70.925 53.280 71.215 53.325 ;
        RECT 70.450 53.140 71.215 53.280 ;
        RECT 52.510 52.940 52.830 53.000 ;
        RECT 48.000 52.800 52.830 52.940 ;
        RECT 67.320 52.940 67.460 53.095 ;
        RECT 70.450 53.080 70.770 53.140 ;
        RECT 70.925 53.095 71.215 53.140 ;
        RECT 71.830 53.080 72.150 53.340 ;
        RECT 72.290 53.080 72.610 53.340 ;
        RECT 72.765 53.280 73.055 53.325 ;
        RECT 77.350 53.280 77.670 53.340 ;
        RECT 72.765 53.140 77.670 53.280 ;
        RECT 72.765 53.095 73.055 53.140 ;
        RECT 77.350 53.080 77.670 53.140 ;
        RECT 74.130 52.940 74.450 53.000 ;
        RECT 67.320 52.800 74.450 52.940 ;
        RECT 44.230 52.740 44.550 52.800 ;
        RECT 47.005 52.755 47.295 52.800 ;
        RECT 52.510 52.740 52.830 52.800 ;
        RECT 74.130 52.740 74.450 52.800 ;
        RECT 74.590 52.740 74.910 53.000 ;
        RECT 75.485 52.940 75.775 52.985 ;
        RECT 76.675 52.940 76.965 52.985 ;
        RECT 79.195 52.940 79.485 52.985 ;
        RECT 75.485 52.800 79.485 52.940 ;
        RECT 75.485 52.755 75.775 52.800 ;
        RECT 76.675 52.755 76.965 52.800 ;
        RECT 79.195 52.755 79.485 52.800 ;
        RECT 22.610 52.460 26.980 52.600 ;
        RECT 41.010 52.600 41.330 52.660 ;
        RECT 47.465 52.600 47.755 52.645 ;
        RECT 41.010 52.460 47.755 52.600 ;
        RECT 22.610 52.400 22.930 52.460 ;
        RECT 23.990 52.400 24.310 52.460 ;
        RECT 41.010 52.400 41.330 52.460 ;
        RECT 47.465 52.415 47.755 52.460 ;
        RECT 66.325 52.600 66.615 52.645 ;
        RECT 75.090 52.600 75.380 52.645 ;
        RECT 77.190 52.600 77.480 52.645 ;
        RECT 78.760 52.600 79.050 52.645 ;
        RECT 66.325 52.460 74.820 52.600 ;
        RECT 66.325 52.415 66.615 52.460 ;
        RECT 9.270 52.060 9.590 52.320 ;
        RECT 29.510 52.060 29.830 52.320 ;
        RECT 38.250 52.060 38.570 52.320 ;
        RECT 42.390 52.060 42.710 52.320 ;
        RECT 44.705 52.260 44.995 52.305 ;
        RECT 45.610 52.260 45.930 52.320 ;
        RECT 44.705 52.120 45.930 52.260 ;
        RECT 44.705 52.075 44.995 52.120 ;
        RECT 45.610 52.060 45.930 52.120 ;
        RECT 47.925 52.260 48.215 52.305 ;
        RECT 54.810 52.260 55.130 52.320 ;
        RECT 47.925 52.120 55.130 52.260 ;
        RECT 47.925 52.075 48.215 52.120 ;
        RECT 54.810 52.060 55.130 52.120 ;
        RECT 69.545 52.260 69.835 52.305 ;
        RECT 69.990 52.260 70.310 52.320 ;
        RECT 69.545 52.120 70.310 52.260 ;
        RECT 74.680 52.260 74.820 52.460 ;
        RECT 75.090 52.460 79.050 52.600 ;
        RECT 75.090 52.415 75.380 52.460 ;
        RECT 77.190 52.415 77.480 52.460 ;
        RECT 78.760 52.415 79.050 52.460 ;
        RECT 75.970 52.260 76.290 52.320 ;
        RECT 74.680 52.120 76.290 52.260 ;
        RECT 69.545 52.075 69.835 52.120 ;
        RECT 69.990 52.060 70.310 52.120 ;
        RECT 75.970 52.060 76.290 52.120 ;
        RECT 5.520 51.440 83.260 51.920 ;
        RECT 15.725 51.240 16.015 51.285 ;
        RECT 16.170 51.240 16.490 51.300 ;
        RECT 15.725 51.100 16.490 51.240 ;
        RECT 15.725 51.055 16.015 51.100 ;
        RECT 16.170 51.040 16.490 51.100 ;
        RECT 26.305 51.240 26.595 51.285 ;
        RECT 28.590 51.240 28.910 51.300 ;
        RECT 26.305 51.100 28.910 51.240 ;
        RECT 26.305 51.055 26.595 51.100 ;
        RECT 28.590 51.040 28.910 51.100 ;
        RECT 35.505 51.240 35.795 51.285 ;
        RECT 35.950 51.240 36.270 51.300 ;
        RECT 35.505 51.100 36.270 51.240 ;
        RECT 35.505 51.055 35.795 51.100 ;
        RECT 35.950 51.040 36.270 51.100 ;
        RECT 36.425 51.240 36.715 51.285 ;
        RECT 39.630 51.240 39.950 51.300 ;
        RECT 36.425 51.100 39.950 51.240 ;
        RECT 36.425 51.055 36.715 51.100 ;
        RECT 39.630 51.040 39.950 51.100 ;
        RECT 40.105 51.240 40.395 51.285 ;
        RECT 43.310 51.240 43.630 51.300 ;
        RECT 40.105 51.100 43.630 51.240 ;
        RECT 40.105 51.055 40.395 51.100 ;
        RECT 43.310 51.040 43.630 51.100 ;
        RECT 43.770 51.040 44.090 51.300 ;
        RECT 64.945 51.240 65.235 51.285 ;
        RECT 76.430 51.240 76.750 51.300 ;
        RECT 64.945 51.100 76.750 51.240 ;
        RECT 64.945 51.055 65.235 51.100 ;
        RECT 76.430 51.040 76.750 51.100 ;
        RECT 81.045 51.240 81.335 51.285 ;
        RECT 81.490 51.240 81.810 51.300 ;
        RECT 81.045 51.100 81.810 51.240 ;
        RECT 81.045 51.055 81.335 51.100 ;
        RECT 81.490 51.040 81.810 51.100 ;
        RECT 29.050 50.900 29.340 50.945 ;
        RECT 30.620 50.900 30.910 50.945 ;
        RECT 32.720 50.900 33.010 50.945 ;
        RECT 29.050 50.760 33.010 50.900 ;
        RECT 29.050 50.715 29.340 50.760 ;
        RECT 30.620 50.715 30.910 50.760 ;
        RECT 32.720 50.715 33.010 50.760 ;
        RECT 40.550 50.700 40.870 50.960 ;
        RECT 44.705 50.900 44.995 50.945 ;
        RECT 42.020 50.760 44.995 50.900 ;
        RECT 13.870 50.560 14.190 50.620 ;
        RECT 19.850 50.560 20.170 50.620 ;
        RECT 21.705 50.560 21.995 50.605 ;
        RECT 13.870 50.420 21.995 50.560 ;
        RECT 13.870 50.360 14.190 50.420 ;
        RECT 19.850 50.360 20.170 50.420 ;
        RECT 21.705 50.375 21.995 50.420 ;
        RECT 28.615 50.560 28.905 50.605 ;
        RECT 31.135 50.560 31.425 50.605 ;
        RECT 32.325 50.560 32.615 50.605 ;
        RECT 28.615 50.420 32.615 50.560 ;
        RECT 28.615 50.375 28.905 50.420 ;
        RECT 31.135 50.375 31.425 50.420 ;
        RECT 32.325 50.375 32.615 50.420 ;
        RECT 16.630 50.020 16.950 50.280 ;
        RECT 18.010 50.020 18.330 50.280 ;
        RECT 23.530 50.220 23.850 50.280 ;
        RECT 19.480 50.080 23.850 50.220 ;
        RECT 17.565 49.880 17.855 49.925 ;
        RECT 19.480 49.880 19.620 50.080 ;
        RECT 23.530 50.020 23.850 50.080 ;
        RECT 25.845 50.220 26.135 50.265 ;
        RECT 27.210 50.220 27.530 50.280 ;
        RECT 25.845 50.080 27.530 50.220 ;
        RECT 25.845 50.035 26.135 50.080 ;
        RECT 27.210 50.020 27.530 50.080 ;
        RECT 33.190 50.020 33.510 50.280 ;
        RECT 33.665 50.220 33.955 50.265 ;
        RECT 34.570 50.220 34.890 50.280 ;
        RECT 36.885 50.220 37.175 50.265 ;
        RECT 33.665 50.080 37.175 50.220 ;
        RECT 33.665 50.035 33.955 50.080 ;
        RECT 34.570 50.020 34.890 50.080 ;
        RECT 36.885 50.035 37.175 50.080 ;
        RECT 40.565 50.220 40.855 50.265 ;
        RECT 41.470 50.220 41.790 50.280 ;
        RECT 42.020 50.265 42.160 50.760 ;
        RECT 44.705 50.715 44.995 50.760 ;
        RECT 56.230 50.900 56.520 50.945 ;
        RECT 58.330 50.900 58.620 50.945 ;
        RECT 59.900 50.900 60.190 50.945 ;
        RECT 70.450 50.900 70.770 50.960 ;
        RECT 56.230 50.760 60.190 50.900 ;
        RECT 56.230 50.715 56.520 50.760 ;
        RECT 58.330 50.715 58.620 50.760 ;
        RECT 59.900 50.715 60.190 50.760 ;
        RECT 68.240 50.760 70.770 50.900 ;
        RECT 42.390 50.560 42.710 50.620 ;
        RECT 47.465 50.560 47.755 50.605 ;
        RECT 42.390 50.420 47.755 50.560 ;
        RECT 42.390 50.360 42.710 50.420 ;
        RECT 47.465 50.375 47.755 50.420 ;
        RECT 56.625 50.560 56.915 50.605 ;
        RECT 57.815 50.560 58.105 50.605 ;
        RECT 60.335 50.560 60.625 50.605 ;
        RECT 56.625 50.420 60.625 50.560 ;
        RECT 56.625 50.375 56.915 50.420 ;
        RECT 57.815 50.375 58.105 50.420 ;
        RECT 60.335 50.375 60.625 50.420 ;
        RECT 64.470 50.560 64.790 50.620 ;
        RECT 64.470 50.420 67.920 50.560 ;
        RECT 64.470 50.360 64.790 50.420 ;
        RECT 40.565 50.080 41.790 50.220 ;
        RECT 40.565 50.035 40.855 50.080 ;
        RECT 41.470 50.020 41.790 50.080 ;
        RECT 41.945 50.035 42.235 50.265 ;
        RECT 42.850 50.020 43.170 50.280 ;
        RECT 43.785 50.220 44.075 50.265 ;
        RECT 45.610 50.220 45.930 50.280 ;
        RECT 43.400 50.080 45.930 50.220 ;
        RECT 17.565 49.740 19.620 49.880 ;
        RECT 19.865 49.880 20.155 49.925 ;
        RECT 24.450 49.880 24.770 49.940 ;
        RECT 19.865 49.740 24.770 49.880 ;
        RECT 17.565 49.695 17.855 49.740 ;
        RECT 19.865 49.695 20.155 49.740 ;
        RECT 24.450 49.680 24.770 49.740 ;
        RECT 31.810 49.925 32.130 49.940 ;
        RECT 31.810 49.695 32.160 49.925 ;
        RECT 35.505 49.880 35.795 49.925 ;
        RECT 35.505 49.740 37.100 49.880 ;
        RECT 35.505 49.695 35.795 49.740 ;
        RECT 31.810 49.680 32.130 49.695 ;
        RECT 36.960 49.600 37.100 49.740 ;
        RECT 20.325 49.540 20.615 49.585 ;
        RECT 22.610 49.540 22.930 49.600 ;
        RECT 32.270 49.540 32.590 49.600 ;
        RECT 20.325 49.400 32.590 49.540 ;
        RECT 20.325 49.355 20.615 49.400 ;
        RECT 22.610 49.340 22.930 49.400 ;
        RECT 32.270 49.340 32.590 49.400 ;
        RECT 36.870 49.340 37.190 49.600 ;
        RECT 41.485 49.540 41.775 49.585 ;
        RECT 43.400 49.540 43.540 50.080 ;
        RECT 43.785 50.035 44.075 50.080 ;
        RECT 45.610 50.020 45.930 50.080 ;
        RECT 52.510 50.020 52.830 50.280 ;
        RECT 55.745 50.220 56.035 50.265 ;
        RECT 55.745 50.080 60.560 50.220 ;
        RECT 55.745 50.035 56.035 50.080 ;
        RECT 57.660 49.940 57.800 50.080 ;
        RECT 60.420 49.940 60.560 50.080 ;
        RECT 65.850 50.020 66.170 50.280 ;
        RECT 67.780 50.265 67.920 50.420 ;
        RECT 68.240 50.265 68.380 50.760 ;
        RECT 70.450 50.700 70.770 50.760 ;
        RECT 70.950 50.900 71.240 50.945 ;
        RECT 73.050 50.900 73.340 50.945 ;
        RECT 74.620 50.900 74.910 50.945 ;
        RECT 70.950 50.760 74.910 50.900 ;
        RECT 70.950 50.715 71.240 50.760 ;
        RECT 73.050 50.715 73.340 50.760 ;
        RECT 74.620 50.715 74.910 50.760 ;
        RECT 71.345 50.560 71.635 50.605 ;
        RECT 72.535 50.560 72.825 50.605 ;
        RECT 75.055 50.560 75.345 50.605 ;
        RECT 68.700 50.420 71.140 50.560 ;
        RECT 68.700 50.265 68.840 50.420 ;
        RECT 67.705 50.035 67.995 50.265 ;
        RECT 68.165 50.035 68.455 50.265 ;
        RECT 68.625 50.035 68.915 50.265 ;
        RECT 69.545 50.220 69.835 50.265 ;
        RECT 69.990 50.220 70.310 50.280 ;
        RECT 69.545 50.080 70.310 50.220 ;
        RECT 69.545 50.035 69.835 50.080 ;
        RECT 69.990 50.020 70.310 50.080 ;
        RECT 70.465 50.035 70.755 50.265 ;
        RECT 71.000 50.220 71.140 50.420 ;
        RECT 71.345 50.420 75.345 50.560 ;
        RECT 71.345 50.375 71.635 50.420 ;
        RECT 72.535 50.375 72.825 50.420 ;
        RECT 75.055 50.375 75.345 50.420 ;
        RECT 77.825 50.220 78.115 50.265 ;
        RECT 71.000 50.080 78.115 50.220 ;
        RECT 77.825 50.035 78.115 50.080 ;
        RECT 80.125 50.220 80.415 50.265 ;
        RECT 80.570 50.220 80.890 50.280 ;
        RECT 80.125 50.080 80.890 50.220 ;
        RECT 80.125 50.035 80.415 50.080 ;
        RECT 57.110 49.925 57.430 49.940 ;
        RECT 57.080 49.695 57.430 49.925 ;
        RECT 57.110 49.680 57.430 49.695 ;
        RECT 57.570 49.680 57.890 49.940 ;
        RECT 60.330 49.880 60.650 49.940 ;
        RECT 65.390 49.880 65.710 49.940 ;
        RECT 70.540 49.880 70.680 50.035 ;
        RECT 80.570 50.020 80.890 50.080 ;
        RECT 71.690 49.880 71.980 49.925 ;
        RECT 78.745 49.880 79.035 49.925 ;
        RECT 60.330 49.740 70.680 49.880 ;
        RECT 71.000 49.740 71.980 49.880 ;
        RECT 60.330 49.680 60.650 49.740 ;
        RECT 65.390 49.680 65.710 49.740 ;
        RECT 41.485 49.400 43.540 49.540 ;
        RECT 43.770 49.540 44.090 49.600 ;
        RECT 49.305 49.540 49.595 49.585 ;
        RECT 43.770 49.400 49.595 49.540 ;
        RECT 41.485 49.355 41.775 49.400 ;
        RECT 43.770 49.340 44.090 49.400 ;
        RECT 49.305 49.355 49.595 49.400 ;
        RECT 62.170 49.540 62.490 49.600 ;
        RECT 62.645 49.540 62.935 49.585 ;
        RECT 62.170 49.400 62.935 49.540 ;
        RECT 62.170 49.340 62.490 49.400 ;
        RECT 62.645 49.355 62.935 49.400 ;
        RECT 66.325 49.540 66.615 49.585 ;
        RECT 71.000 49.540 71.140 49.740 ;
        RECT 71.690 49.695 71.980 49.740 ;
        RECT 77.440 49.740 79.035 49.880 ;
        RECT 66.325 49.400 71.140 49.540 ;
        RECT 74.130 49.540 74.450 49.600 ;
        RECT 77.440 49.585 77.580 49.740 ;
        RECT 78.745 49.695 79.035 49.740 ;
        RECT 79.665 49.695 79.955 49.925 ;
        RECT 77.365 49.540 77.655 49.585 ;
        RECT 74.130 49.400 77.655 49.540 ;
        RECT 66.325 49.355 66.615 49.400 ;
        RECT 74.130 49.340 74.450 49.400 ;
        RECT 77.365 49.355 77.655 49.400 ;
        RECT 77.810 49.540 78.130 49.600 ;
        RECT 79.740 49.540 79.880 49.695 ;
        RECT 80.570 49.540 80.890 49.600 ;
        RECT 77.810 49.400 80.890 49.540 ;
        RECT 77.810 49.340 78.130 49.400 ;
        RECT 80.570 49.340 80.890 49.400 ;
        RECT 5.520 48.720 83.260 49.200 ;
        RECT 15.265 48.520 15.555 48.565 ;
        RECT 16.630 48.520 16.950 48.580 ;
        RECT 15.265 48.380 16.950 48.520 ;
        RECT 15.265 48.335 15.555 48.380 ;
        RECT 16.630 48.320 16.950 48.380 ;
        RECT 18.485 48.520 18.775 48.565 ;
        RECT 20.785 48.520 21.075 48.565 ;
        RECT 18.485 48.380 21.075 48.520 ;
        RECT 18.485 48.335 18.775 48.380 ;
        RECT 20.785 48.335 21.075 48.380 ;
        RECT 22.165 48.520 22.455 48.565 ;
        RECT 23.530 48.520 23.850 48.580 ;
        RECT 22.165 48.380 23.850 48.520 ;
        RECT 22.165 48.335 22.455 48.380 ;
        RECT 23.530 48.320 23.850 48.380 ;
        RECT 31.810 48.320 32.130 48.580 ;
        RECT 34.570 48.320 34.890 48.580 ;
        RECT 42.850 48.520 43.170 48.580 ;
        RECT 45.150 48.520 45.470 48.580 ;
        RECT 42.850 48.380 45.470 48.520 ;
        RECT 42.850 48.320 43.170 48.380 ;
        RECT 45.150 48.320 45.470 48.380 ;
        RECT 64.470 48.320 64.790 48.580 ;
        RECT 72.750 48.520 73.070 48.580 ;
        RECT 68.700 48.380 73.070 48.520 ;
        RECT 19.390 48.180 19.710 48.240 ;
        RECT 20.325 48.180 20.615 48.225 ;
        RECT 14.420 48.040 20.615 48.180 ;
        RECT 14.420 47.885 14.560 48.040 ;
        RECT 19.390 47.980 19.710 48.040 ;
        RECT 20.325 47.995 20.615 48.040 ;
        RECT 21.370 48.180 21.660 48.225 ;
        RECT 23.070 48.180 23.390 48.240 ;
        RECT 21.370 48.040 23.390 48.180 ;
        RECT 21.370 47.995 21.660 48.040 ;
        RECT 23.070 47.980 23.390 48.040 ;
        RECT 29.510 48.180 29.830 48.240 ;
        RECT 32.585 48.180 32.875 48.225 ;
        RECT 29.510 48.040 32.875 48.180 ;
        RECT 29.510 47.980 29.830 48.040 ;
        RECT 32.585 47.995 32.875 48.040 ;
        RECT 33.665 47.995 33.955 48.225 ;
        RECT 62.170 48.180 62.490 48.240 ;
        RECT 68.700 48.180 68.840 48.380 ;
        RECT 72.750 48.320 73.070 48.380 ;
        RECT 73.760 48.380 74.820 48.520 ;
        RECT 41.560 48.040 49.060 48.180 ;
        RECT 13.885 47.655 14.175 47.885 ;
        RECT 14.345 47.655 14.635 47.885 ;
        RECT 13.960 47.500 14.100 47.655 ;
        RECT 16.630 47.640 16.950 47.900 ;
        RECT 19.850 47.840 20.170 47.900 ;
        RECT 24.005 47.840 24.295 47.885 ;
        RECT 17.180 47.700 19.620 47.840 ;
        RECT 14.790 47.500 15.110 47.560 ;
        RECT 17.180 47.545 17.320 47.700 ;
        RECT 13.960 47.360 15.110 47.500 ;
        RECT 14.790 47.300 15.110 47.360 ;
        RECT 15.265 47.315 15.555 47.545 ;
        RECT 17.105 47.315 17.395 47.545 ;
        RECT 18.010 47.500 18.330 47.560 ;
        RECT 18.945 47.500 19.235 47.545 ;
        RECT 18.010 47.360 19.235 47.500 ;
        RECT 19.480 47.500 19.620 47.700 ;
        RECT 19.850 47.700 24.295 47.840 ;
        RECT 19.850 47.640 20.170 47.700 ;
        RECT 24.005 47.655 24.295 47.700 ;
        RECT 29.985 47.840 30.275 47.885 ;
        RECT 31.350 47.840 31.670 47.900 ;
        RECT 33.740 47.840 33.880 47.995 ;
        RECT 41.560 47.885 41.700 48.040 ;
        RECT 29.985 47.700 31.670 47.840 ;
        RECT 29.985 47.655 30.275 47.700 ;
        RECT 31.350 47.640 31.670 47.700 ;
        RECT 32.360 47.700 33.880 47.840 ;
        RECT 40.205 47.840 40.495 47.885 ;
        RECT 40.205 47.700 41.240 47.840 ;
        RECT 32.360 47.560 32.500 47.700 ;
        RECT 40.205 47.655 40.495 47.700 ;
        RECT 27.210 47.500 27.530 47.560 ;
        RECT 27.685 47.500 27.975 47.545 ;
        RECT 19.480 47.360 27.975 47.500 ;
        RECT 15.340 46.820 15.480 47.315 ;
        RECT 18.010 47.300 18.330 47.360 ;
        RECT 18.945 47.315 19.235 47.360 ;
        RECT 27.210 47.300 27.530 47.360 ;
        RECT 27.685 47.315 27.975 47.360 ;
        RECT 32.270 47.300 32.590 47.560 ;
        RECT 36.895 47.500 37.185 47.545 ;
        RECT 39.415 47.500 39.705 47.545 ;
        RECT 40.605 47.500 40.895 47.545 ;
        RECT 36.895 47.360 40.895 47.500 ;
        RECT 41.100 47.500 41.240 47.700 ;
        RECT 41.485 47.655 41.775 47.885 ;
        RECT 43.310 47.840 43.630 47.900 ;
        RECT 48.920 47.885 49.060 48.040 ;
        RECT 62.170 48.040 68.840 48.180 ;
        RECT 69.070 48.180 69.390 48.240 ;
        RECT 70.910 48.180 71.230 48.240 ;
        RECT 73.760 48.180 73.900 48.380 ;
        RECT 69.070 48.040 73.900 48.180 ;
        RECT 62.170 47.980 62.490 48.040 ;
        RECT 69.070 47.980 69.390 48.040 ;
        RECT 70.910 47.980 71.230 48.040 ;
        RECT 74.130 47.980 74.450 48.240 ;
        RECT 74.680 48.180 74.820 48.380 ;
        RECT 76.905 48.180 77.195 48.225 ;
        RECT 74.680 48.040 74.850 48.180 ;
        RECT 46.545 47.840 46.835 47.885 ;
        RECT 43.310 47.700 46.835 47.840 ;
        RECT 43.310 47.640 43.630 47.700 ;
        RECT 46.545 47.655 46.835 47.700 ;
        RECT 48.845 47.840 49.135 47.885 ;
        RECT 49.290 47.840 49.610 47.900 ;
        RECT 48.845 47.700 49.610 47.840 ;
        RECT 48.845 47.655 49.135 47.700 ;
        RECT 49.290 47.640 49.610 47.700 ;
        RECT 50.180 47.840 50.470 47.885 ;
        RECT 52.050 47.840 52.370 47.900 ;
        RECT 50.180 47.700 52.370 47.840 ;
        RECT 50.180 47.655 50.470 47.700 ;
        RECT 52.050 47.640 52.370 47.700 ;
        RECT 57.570 47.640 57.890 47.900 ;
        RECT 58.920 47.840 59.210 47.885 ;
        RECT 63.090 47.840 63.410 47.900 ;
        RECT 58.920 47.700 63.410 47.840 ;
        RECT 58.920 47.655 59.210 47.700 ;
        RECT 63.090 47.640 63.410 47.700 ;
        RECT 65.390 47.640 65.710 47.900 ;
        RECT 66.770 47.885 67.090 47.900 ;
        RECT 66.740 47.655 67.090 47.885 ;
        RECT 66.770 47.640 67.090 47.655 ;
        RECT 73.670 47.640 73.990 47.900 ;
        RECT 74.710 47.885 74.850 48.040 ;
        RECT 75.140 48.040 77.195 48.180 ;
        RECT 75.140 47.900 75.280 48.040 ;
        RECT 76.905 47.995 77.195 48.040 ;
        RECT 78.270 48.180 78.590 48.240 ;
        RECT 78.745 48.180 79.035 48.225 ;
        RECT 78.270 48.040 79.035 48.180 ;
        RECT 78.270 47.980 78.590 48.040 ;
        RECT 78.745 47.995 79.035 48.040 ;
        RECT 79.205 48.180 79.495 48.225 ;
        RECT 80.570 48.180 80.890 48.240 ;
        RECT 79.205 48.040 80.890 48.180 ;
        RECT 79.205 47.995 79.495 48.040 ;
        RECT 80.570 47.980 80.890 48.040 ;
        RECT 74.605 47.655 74.895 47.885 ;
        RECT 75.050 47.640 75.370 47.900 ;
        RECT 75.525 47.655 75.815 47.885 ;
        RECT 77.825 47.655 78.115 47.885 ;
        RECT 41.100 47.360 41.700 47.500 ;
        RECT 36.895 47.315 37.185 47.360 ;
        RECT 39.415 47.315 39.705 47.360 ;
        RECT 40.605 47.315 40.895 47.360 ;
        RECT 28.605 47.160 28.895 47.205 ;
        RECT 33.650 47.160 33.970 47.220 ;
        RECT 28.605 47.020 33.970 47.160 ;
        RECT 28.605 46.975 28.895 47.020 ;
        RECT 33.650 46.960 33.970 47.020 ;
        RECT 37.330 47.160 37.620 47.205 ;
        RECT 38.900 47.160 39.190 47.205 ;
        RECT 41.000 47.160 41.290 47.205 ;
        RECT 37.330 47.020 41.290 47.160 ;
        RECT 41.560 47.160 41.700 47.360 ;
        RECT 41.930 47.300 42.250 47.560 ;
        RECT 47.910 47.300 48.230 47.560 ;
        RECT 49.725 47.500 50.015 47.545 ;
        RECT 50.915 47.500 51.205 47.545 ;
        RECT 53.435 47.500 53.725 47.545 ;
        RECT 49.725 47.360 53.725 47.500 ;
        RECT 49.725 47.315 50.015 47.360 ;
        RECT 50.915 47.315 51.205 47.360 ;
        RECT 53.435 47.315 53.725 47.360 ;
        RECT 58.465 47.500 58.755 47.545 ;
        RECT 59.655 47.500 59.945 47.545 ;
        RECT 62.175 47.500 62.465 47.545 ;
        RECT 58.465 47.360 62.465 47.500 ;
        RECT 58.465 47.315 58.755 47.360 ;
        RECT 59.655 47.315 59.945 47.360 ;
        RECT 62.175 47.315 62.465 47.360 ;
        RECT 66.285 47.500 66.575 47.545 ;
        RECT 67.475 47.500 67.765 47.545 ;
        RECT 69.995 47.500 70.285 47.545 ;
        RECT 75.600 47.500 75.740 47.655 ;
        RECT 66.285 47.360 70.285 47.500 ;
        RECT 66.285 47.315 66.575 47.360 ;
        RECT 67.475 47.315 67.765 47.360 ;
        RECT 69.995 47.315 70.285 47.360 ;
        RECT 72.380 47.360 75.740 47.500 ;
        RECT 77.900 47.500 78.040 47.655 ;
        RECT 80.110 47.640 80.430 47.900 ;
        RECT 79.650 47.500 79.970 47.560 ;
        RECT 77.900 47.360 79.970 47.500 ;
        RECT 45.625 47.160 45.915 47.205 ;
        RECT 41.560 47.020 45.915 47.160 ;
        RECT 37.330 46.975 37.620 47.020 ;
        RECT 38.900 46.975 39.190 47.020 ;
        RECT 41.000 46.975 41.290 47.020 ;
        RECT 45.625 46.975 45.915 47.020 ;
        RECT 49.330 47.160 49.620 47.205 ;
        RECT 51.430 47.160 51.720 47.205 ;
        RECT 53.000 47.160 53.290 47.205 ;
        RECT 49.330 47.020 53.290 47.160 ;
        RECT 49.330 46.975 49.620 47.020 ;
        RECT 51.430 46.975 51.720 47.020 ;
        RECT 53.000 46.975 53.290 47.020 ;
        RECT 58.070 47.160 58.360 47.205 ;
        RECT 60.170 47.160 60.460 47.205 ;
        RECT 61.740 47.160 62.030 47.205 ;
        RECT 58.070 47.020 62.030 47.160 ;
        RECT 58.070 46.975 58.360 47.020 ;
        RECT 60.170 46.975 60.460 47.020 ;
        RECT 61.740 46.975 62.030 47.020 ;
        RECT 65.890 47.160 66.180 47.205 ;
        RECT 67.990 47.160 68.280 47.205 ;
        RECT 69.560 47.160 69.850 47.205 ;
        RECT 65.890 47.020 69.850 47.160 ;
        RECT 65.890 46.975 66.180 47.020 ;
        RECT 67.990 46.975 68.280 47.020 ;
        RECT 69.560 46.975 69.850 47.020 ;
        RECT 72.380 46.880 72.520 47.360 ;
        RECT 79.650 47.300 79.970 47.360 ;
        RECT 72.750 46.960 73.070 47.220 ;
        RECT 20.310 46.820 20.630 46.880 ;
        RECT 15.340 46.680 20.630 46.820 ;
        RECT 20.310 46.620 20.630 46.680 ;
        RECT 32.730 46.620 33.050 46.880 ;
        RECT 46.070 46.820 46.390 46.880 ;
        RECT 47.465 46.820 47.755 46.865 ;
        RECT 46.070 46.680 47.755 46.820 ;
        RECT 46.070 46.620 46.390 46.680 ;
        RECT 47.465 46.635 47.755 46.680 ;
        RECT 53.890 46.820 54.210 46.880 ;
        RECT 55.745 46.820 56.035 46.865 ;
        RECT 61.250 46.820 61.570 46.880 ;
        RECT 66.310 46.820 66.630 46.880 ;
        RECT 53.890 46.680 66.630 46.820 ;
        RECT 53.890 46.620 54.210 46.680 ;
        RECT 55.745 46.635 56.035 46.680 ;
        RECT 61.250 46.620 61.570 46.680 ;
        RECT 66.310 46.620 66.630 46.680 ;
        RECT 72.290 46.620 72.610 46.880 ;
        RECT 73.210 46.820 73.530 46.880 ;
        RECT 81.045 46.820 81.335 46.865 ;
        RECT 73.210 46.680 81.335 46.820 ;
        RECT 73.210 46.620 73.530 46.680 ;
        RECT 81.045 46.635 81.335 46.680 ;
        RECT 5.520 46.000 83.260 46.480 ;
        RECT 9.270 45.800 9.590 45.860 ;
        RECT 9.745 45.800 10.035 45.845 ;
        RECT 9.270 45.660 10.035 45.800 ;
        RECT 9.270 45.600 9.590 45.660 ;
        RECT 9.745 45.615 10.035 45.660 ;
        RECT 18.010 45.600 18.330 45.860 ;
        RECT 19.865 45.615 20.155 45.845 ;
        RECT 20.310 45.800 20.630 45.860 ;
        RECT 22.625 45.800 22.915 45.845 ;
        RECT 20.310 45.660 22.915 45.800 ;
        RECT 7.890 45.460 8.210 45.520 ;
        RECT 12.505 45.460 12.795 45.505 ;
        RECT 7.890 45.320 12.795 45.460 ;
        RECT 7.890 45.260 8.210 45.320 ;
        RECT 12.505 45.275 12.795 45.320 ;
        RECT 11.570 45.120 11.890 45.180 ;
        RECT 11.200 44.980 11.890 45.120 ;
        RECT 11.200 44.825 11.340 44.980 ;
        RECT 11.570 44.920 11.890 44.980 ;
        RECT 11.125 44.595 11.415 44.825 ;
        RECT 15.710 44.780 16.030 44.840 ;
        RECT 11.660 44.640 16.030 44.780 ;
        RECT 7.430 44.440 7.750 44.500 ;
        RECT 9.585 44.440 9.875 44.485 ;
        RECT 7.430 44.300 9.875 44.440 ;
        RECT 7.430 44.240 7.750 44.300 ;
        RECT 9.585 44.255 9.875 44.300 ;
        RECT 10.190 44.440 10.510 44.500 ;
        RECT 10.665 44.440 10.955 44.485 ;
        RECT 10.190 44.300 10.955 44.440 ;
        RECT 10.190 44.240 10.510 44.300 ;
        RECT 10.665 44.255 10.955 44.300 ;
        RECT 11.660 44.160 11.800 44.640 ;
        RECT 15.710 44.580 16.030 44.640 ;
        RECT 16.185 44.780 16.475 44.825 ;
        RECT 17.550 44.780 17.870 44.840 ;
        RECT 16.185 44.640 17.870 44.780 ;
        RECT 18.100 44.780 18.240 45.600 ;
        RECT 19.940 45.460 20.080 45.615 ;
        RECT 20.310 45.600 20.630 45.660 ;
        RECT 22.625 45.615 22.915 45.660 ;
        RECT 23.990 45.800 24.310 45.860 ;
        RECT 24.925 45.800 25.215 45.845 ;
        RECT 23.990 45.660 25.215 45.800 ;
        RECT 23.990 45.600 24.310 45.660 ;
        RECT 24.925 45.615 25.215 45.660 ;
        RECT 41.485 45.800 41.775 45.845 ;
        RECT 41.930 45.800 42.250 45.860 ;
        RECT 41.485 45.660 42.250 45.800 ;
        RECT 41.485 45.615 41.775 45.660 ;
        RECT 41.930 45.600 42.250 45.660 ;
        RECT 42.850 45.600 43.170 45.860 ;
        RECT 57.110 45.600 57.430 45.860 ;
        RECT 67.230 45.600 67.550 45.860 ;
        RECT 81.030 45.600 81.350 45.860 ;
        RECT 31.350 45.460 31.670 45.520 ;
        RECT 19.940 45.320 31.670 45.460 ;
        RECT 31.350 45.260 31.670 45.320 ;
        RECT 35.070 45.460 35.360 45.505 ;
        RECT 37.170 45.460 37.460 45.505 ;
        RECT 38.740 45.460 39.030 45.505 ;
        RECT 35.070 45.320 39.030 45.460 ;
        RECT 35.070 45.275 35.360 45.320 ;
        RECT 37.170 45.275 37.460 45.320 ;
        RECT 38.740 45.275 39.030 45.320 ;
        RECT 43.785 45.275 44.075 45.505 ;
        RECT 45.190 45.460 45.480 45.505 ;
        RECT 47.290 45.460 47.580 45.505 ;
        RECT 48.860 45.460 49.150 45.505 ;
        RECT 45.190 45.320 49.150 45.460 ;
        RECT 45.190 45.275 45.480 45.320 ;
        RECT 47.290 45.275 47.580 45.320 ;
        RECT 48.860 45.275 49.150 45.320 ;
        RECT 61.250 45.460 61.570 45.520 ;
        RECT 72.290 45.460 72.610 45.520 ;
        RECT 61.250 45.320 72.610 45.460 ;
        RECT 18.470 45.120 18.790 45.180 ;
        RECT 18.470 44.980 19.620 45.120 ;
        RECT 18.470 44.920 18.790 44.980 ;
        RECT 18.945 44.780 19.235 44.825 ;
        RECT 18.100 44.640 19.235 44.780 ;
        RECT 19.480 44.780 19.620 44.980 ;
        RECT 19.850 44.920 20.170 45.180 ;
        RECT 35.465 45.120 35.755 45.165 ;
        RECT 36.655 45.120 36.945 45.165 ;
        RECT 39.175 45.120 39.465 45.165 ;
        RECT 20.860 44.980 24.220 45.120 ;
        RECT 20.325 44.780 20.615 44.825 ;
        RECT 19.480 44.640 20.615 44.780 ;
        RECT 16.185 44.595 16.475 44.640 ;
        RECT 17.550 44.580 17.870 44.640 ;
        RECT 18.945 44.595 19.235 44.640 ;
        RECT 20.325 44.595 20.615 44.640 ;
        RECT 12.505 44.440 12.795 44.485 ;
        RECT 14.790 44.440 15.110 44.500 ;
        RECT 17.090 44.440 17.410 44.500 ;
        RECT 12.505 44.300 13.870 44.440 ;
        RECT 12.505 44.255 12.795 44.300 ;
        RECT 8.810 43.900 9.130 44.160 ;
        RECT 11.570 43.900 11.890 44.160 ;
        RECT 13.730 44.100 13.870 44.300 ;
        RECT 14.790 44.300 17.410 44.440 ;
        RECT 14.790 44.240 15.110 44.300 ;
        RECT 17.090 44.240 17.410 44.300 ;
        RECT 14.330 44.100 14.650 44.160 ;
        RECT 16.630 44.100 16.950 44.160 ;
        RECT 20.860 44.100 21.000 44.980 ;
        RECT 24.080 44.825 24.220 44.980 ;
        RECT 35.465 44.980 39.465 45.120 ;
        RECT 35.465 44.935 35.755 44.980 ;
        RECT 36.655 44.935 36.945 44.980 ;
        RECT 39.175 44.935 39.465 44.980 ;
        RECT 41.470 45.120 41.790 45.180 ;
        RECT 43.860 45.120 44.000 45.275 ;
        RECT 61.250 45.260 61.570 45.320 ;
        RECT 41.470 44.980 44.000 45.120 ;
        RECT 41.470 44.920 41.790 44.980 ;
        RECT 23.545 44.780 23.835 44.825 ;
        RECT 21.320 44.640 23.835 44.780 ;
        RECT 21.320 44.145 21.460 44.640 ;
        RECT 23.545 44.595 23.835 44.640 ;
        RECT 24.005 44.595 24.295 44.825 ;
        RECT 25.385 44.780 25.675 44.825 ;
        RECT 26.290 44.780 26.610 44.840 ;
        RECT 25.385 44.640 26.610 44.780 ;
        RECT 25.385 44.595 25.675 44.640 ;
        RECT 26.290 44.580 26.610 44.640 ;
        RECT 27.225 44.595 27.515 44.825 ;
        RECT 27.670 44.780 27.990 44.840 ;
        RECT 34.125 44.780 34.415 44.825 ;
        RECT 27.670 44.640 34.415 44.780 ;
        RECT 27.300 44.440 27.440 44.595 ;
        RECT 27.670 44.580 27.990 44.640 ;
        RECT 34.125 44.595 34.415 44.640 ;
        RECT 34.585 44.595 34.875 44.825 ;
        RECT 35.920 44.780 36.210 44.825 ;
        RECT 38.250 44.780 38.570 44.840 ;
        RECT 35.920 44.640 38.570 44.780 ;
        RECT 35.920 44.595 36.210 44.640 ;
        RECT 30.445 44.440 30.735 44.485 ;
        RECT 31.810 44.440 32.130 44.500 ;
        RECT 33.190 44.440 33.510 44.500 ;
        RECT 34.660 44.440 34.800 44.595 ;
        RECT 38.250 44.580 38.570 44.640 ;
        RECT 27.300 44.300 34.800 44.440 ;
        RECT 30.445 44.255 30.735 44.300 ;
        RECT 31.810 44.240 32.130 44.300 ;
        RECT 33.190 44.240 33.510 44.300 ;
        RECT 41.930 44.240 42.250 44.500 ;
        RECT 43.860 44.440 44.000 44.980 ;
        RECT 45.585 45.120 45.875 45.165 ;
        RECT 46.775 45.120 47.065 45.165 ;
        RECT 49.295 45.120 49.585 45.165 ;
        RECT 45.585 44.980 49.585 45.120 ;
        RECT 45.585 44.935 45.875 44.980 ;
        RECT 46.775 44.935 47.065 44.980 ;
        RECT 49.295 44.935 49.585 44.980 ;
        RECT 59.870 44.920 60.190 45.180 ;
        RECT 60.790 45.120 61.110 45.180 ;
        RECT 60.790 44.980 67.460 45.120 ;
        RECT 60.790 44.920 61.110 44.980 ;
        RECT 44.705 44.780 44.995 44.825 ;
        RECT 56.665 44.780 56.955 44.825 ;
        RECT 58.490 44.780 58.810 44.840 ;
        RECT 67.320 44.825 67.460 44.980 ;
        RECT 66.785 44.780 67.075 44.825 ;
        RECT 44.705 44.640 49.520 44.780 ;
        RECT 44.705 44.595 44.995 44.640 ;
        RECT 49.380 44.500 49.520 44.640 ;
        RECT 56.665 44.640 67.075 44.780 ;
        RECT 56.665 44.595 56.955 44.640 ;
        RECT 58.490 44.580 58.810 44.640 ;
        RECT 66.785 44.595 67.075 44.640 ;
        RECT 67.245 44.595 67.535 44.825 ;
        RECT 67.690 44.580 68.010 44.840 ;
        RECT 69.070 44.580 69.390 44.840 ;
        RECT 71.460 44.825 71.600 45.320 ;
        RECT 72.290 45.260 72.610 45.320 ;
        RECT 71.385 44.595 71.675 44.825 ;
        RECT 74.590 44.780 74.910 44.840 ;
        RECT 75.525 44.780 75.815 44.825 ;
        RECT 74.590 44.640 75.815 44.780 ;
        RECT 74.590 44.580 74.910 44.640 ;
        RECT 75.525 44.595 75.815 44.640 ;
        RECT 75.970 44.580 76.290 44.840 ;
        RECT 76.445 44.595 76.735 44.825 ;
        RECT 76.890 44.780 77.210 44.840 ;
        RECT 77.365 44.780 77.655 44.825 ;
        RECT 76.890 44.640 77.655 44.780 ;
        RECT 45.930 44.440 46.220 44.485 ;
        RECT 43.860 44.300 46.220 44.440 ;
        RECT 45.930 44.255 46.220 44.300 ;
        RECT 49.290 44.440 49.610 44.500 ;
        RECT 52.525 44.440 52.815 44.485 ;
        RECT 49.290 44.300 52.815 44.440 ;
        RECT 49.290 44.240 49.610 44.300 ;
        RECT 52.525 44.255 52.815 44.300 ;
        RECT 58.965 44.440 59.255 44.485 ;
        RECT 62.170 44.440 62.490 44.500 ;
        RECT 58.965 44.300 62.490 44.440 ;
        RECT 58.965 44.255 59.255 44.300 ;
        RECT 62.170 44.240 62.490 44.300 ;
        RECT 62.630 44.240 62.950 44.500 ;
        RECT 69.160 44.440 69.300 44.580 ;
        RECT 72.305 44.440 72.595 44.485 ;
        RECT 75.050 44.440 75.370 44.500 ;
        RECT 69.160 44.300 75.370 44.440 ;
        RECT 76.520 44.440 76.660 44.595 ;
        RECT 76.890 44.580 77.210 44.640 ;
        RECT 77.365 44.595 77.655 44.640 ;
        RECT 78.730 44.580 79.050 44.840 ;
        RECT 79.190 44.780 79.510 44.840 ;
        RECT 80.125 44.780 80.415 44.825 ;
        RECT 79.190 44.640 80.415 44.780 ;
        RECT 79.190 44.580 79.510 44.640 ;
        RECT 80.125 44.595 80.415 44.640 ;
        RECT 77.825 44.440 78.115 44.485 ;
        RECT 76.520 44.300 78.115 44.440 ;
        RECT 72.305 44.255 72.595 44.300 ;
        RECT 75.050 44.240 75.370 44.300 ;
        RECT 77.825 44.255 78.115 44.300 ;
        RECT 79.650 44.440 79.970 44.500 ;
        RECT 80.570 44.440 80.890 44.500 ;
        RECT 79.650 44.300 80.890 44.440 ;
        RECT 79.650 44.240 79.970 44.300 ;
        RECT 80.570 44.240 80.890 44.300 ;
        RECT 13.730 43.960 21.000 44.100 ;
        RECT 14.330 43.900 14.650 43.960 ;
        RECT 16.630 43.900 16.950 43.960 ;
        RECT 21.245 43.915 21.535 44.145 ;
        RECT 41.470 44.100 41.790 44.160 ;
        RECT 42.945 44.100 43.235 44.145 ;
        RECT 45.150 44.100 45.470 44.160 ;
        RECT 41.470 43.960 45.470 44.100 ;
        RECT 41.470 43.900 41.790 43.960 ;
        RECT 42.945 43.915 43.235 43.960 ;
        RECT 45.150 43.900 45.470 43.960 ;
        RECT 51.605 44.100 51.895 44.145 ;
        RECT 55.730 44.100 56.050 44.160 ;
        RECT 51.605 43.960 56.050 44.100 ;
        RECT 51.605 43.915 51.895 43.960 ;
        RECT 55.730 43.900 56.050 43.960 ;
        RECT 59.410 43.900 59.730 44.160 ;
        RECT 61.710 44.100 62.030 44.160 ;
        RECT 69.085 44.100 69.375 44.145 ;
        RECT 61.710 43.960 69.375 44.100 ;
        RECT 61.710 43.900 62.030 43.960 ;
        RECT 69.085 43.915 69.375 43.960 ;
        RECT 69.530 44.100 69.850 44.160 ;
        RECT 70.465 44.100 70.755 44.145 ;
        RECT 69.530 43.960 70.755 44.100 ;
        RECT 69.530 43.900 69.850 43.960 ;
        RECT 70.465 43.915 70.755 43.960 ;
        RECT 74.130 43.900 74.450 44.160 ;
        RECT 5.520 43.280 83.260 43.760 ;
        RECT 6.985 43.080 7.275 43.125 ;
        RECT 11.570 43.080 11.890 43.140 ;
        RECT 6.985 42.940 11.890 43.080 ;
        RECT 6.985 42.895 7.275 42.940 ;
        RECT 11.570 42.880 11.890 42.940 ;
        RECT 19.390 43.080 19.710 43.140 ;
        RECT 21.705 43.080 21.995 43.125 ;
        RECT 19.390 42.940 21.995 43.080 ;
        RECT 19.390 42.880 19.710 42.940 ;
        RECT 21.705 42.895 21.995 42.940 ;
        RECT 23.530 43.080 23.850 43.140 ;
        RECT 25.005 43.080 25.295 43.125 ;
        RECT 23.530 42.940 25.295 43.080 ;
        RECT 23.530 42.880 23.850 42.940 ;
        RECT 25.005 42.895 25.295 42.940 ;
        RECT 26.305 43.080 26.595 43.125 ;
        RECT 26.750 43.080 27.070 43.140 ;
        RECT 26.305 42.940 27.070 43.080 ;
        RECT 26.305 42.895 26.595 42.940 ;
        RECT 26.750 42.880 27.070 42.940 ;
        RECT 41.485 43.080 41.775 43.125 ;
        RECT 42.390 43.080 42.710 43.140 ;
        RECT 41.485 42.940 42.710 43.080 ;
        RECT 41.485 42.895 41.775 42.940 ;
        RECT 42.390 42.880 42.710 42.940 ;
        RECT 48.830 42.880 49.150 43.140 ;
        RECT 52.050 42.880 52.370 43.140 ;
        RECT 53.890 42.880 54.210 43.140 ;
        RECT 62.645 43.080 62.935 43.125 ;
        RECT 63.090 43.080 63.410 43.140 ;
        RECT 62.645 42.940 63.410 43.080 ;
        RECT 62.645 42.895 62.935 42.940 ;
        RECT 63.090 42.880 63.410 42.940 ;
        RECT 64.470 43.080 64.790 43.140 ;
        RECT 64.945 43.080 65.235 43.125 ;
        RECT 64.470 42.940 65.235 43.080 ;
        RECT 64.470 42.880 64.790 42.940 ;
        RECT 64.945 42.895 65.235 42.940 ;
        RECT 12.030 42.740 12.350 42.800 ;
        RECT 12.030 42.600 13.640 42.740 ;
        RECT 12.030 42.540 12.350 42.600 ;
        RECT 12.490 42.445 12.810 42.460 ;
        RECT 12.490 42.215 12.840 42.445 ;
        RECT 12.490 42.200 12.810 42.215 ;
        RECT 9.295 42.060 9.585 42.105 ;
        RECT 11.815 42.060 12.105 42.105 ;
        RECT 13.005 42.060 13.295 42.105 ;
        RECT 9.295 41.920 13.295 42.060 ;
        RECT 13.500 42.060 13.640 42.600 ;
        RECT 14.330 42.540 14.650 42.800 ;
        RECT 15.345 42.740 15.635 42.785 ;
        RECT 14.880 42.600 15.635 42.740 ;
        RECT 13.870 42.200 14.190 42.460 ;
        RECT 14.880 42.060 15.020 42.600 ;
        RECT 15.345 42.555 15.635 42.600 ;
        RECT 19.850 42.740 20.170 42.800 ;
        RECT 22.625 42.740 22.915 42.785 ;
        RECT 19.850 42.600 22.915 42.740 ;
        RECT 19.850 42.540 20.170 42.600 ;
        RECT 22.625 42.555 22.915 42.600 ;
        RECT 24.005 42.740 24.295 42.785 ;
        RECT 27.670 42.740 27.990 42.800 ;
        RECT 31.825 42.740 32.115 42.785 ;
        RECT 24.005 42.600 27.990 42.740 ;
        RECT 24.005 42.555 24.295 42.600 ;
        RECT 27.670 42.540 27.990 42.600 ;
        RECT 28.220 42.600 32.115 42.740 ;
        RECT 16.645 42.400 16.935 42.445 ;
        RECT 13.500 41.920 15.020 42.060 ;
        RECT 16.260 42.260 16.935 42.400 ;
        RECT 9.295 41.875 9.585 41.920 ;
        RECT 11.815 41.875 12.105 41.920 ;
        RECT 13.005 41.875 13.295 41.920 ;
        RECT 9.730 41.720 10.020 41.765 ;
        RECT 11.300 41.720 11.590 41.765 ;
        RECT 13.400 41.720 13.690 41.765 ;
        RECT 9.730 41.580 13.690 41.720 ;
        RECT 9.730 41.535 10.020 41.580 ;
        RECT 11.300 41.535 11.590 41.580 ;
        RECT 13.400 41.535 13.690 41.580 ;
        RECT 14.790 41.720 15.110 41.780 ;
        RECT 16.260 41.765 16.400 42.260 ;
        RECT 16.645 42.215 16.935 42.260 ;
        RECT 17.550 42.200 17.870 42.460 ;
        RECT 23.545 42.215 23.835 42.445 ;
        RECT 23.620 42.060 23.760 42.215 ;
        RECT 27.210 42.200 27.530 42.460 ;
        RECT 28.220 42.445 28.360 42.600 ;
        RECT 31.825 42.555 32.115 42.600 ;
        RECT 35.920 42.740 36.210 42.785 ;
        RECT 40.550 42.740 40.870 42.800 ;
        RECT 60.805 42.740 61.095 42.785 ;
        RECT 64.010 42.740 64.330 42.800 ;
        RECT 35.920 42.600 40.870 42.740 ;
        RECT 35.920 42.555 36.210 42.600 ;
        RECT 40.550 42.540 40.870 42.600 ;
        RECT 42.020 42.600 49.520 42.740 ;
        RECT 28.145 42.215 28.435 42.445 ;
        RECT 28.590 42.200 28.910 42.460 ;
        RECT 31.350 42.400 31.670 42.460 ;
        RECT 42.020 42.445 42.160 42.600 ;
        RECT 49.380 42.460 49.520 42.600 ;
        RECT 60.805 42.600 64.330 42.740 ;
        RECT 60.805 42.555 61.095 42.600 ;
        RECT 64.010 42.540 64.330 42.600 ;
        RECT 32.745 42.400 33.035 42.445 ;
        RECT 31.350 42.260 33.035 42.400 ;
        RECT 31.350 42.200 31.670 42.260 ;
        RECT 32.745 42.215 33.035 42.260 ;
        RECT 41.945 42.215 42.235 42.445 ;
        RECT 42.390 42.400 42.710 42.460 ;
        RECT 43.225 42.400 43.515 42.445 ;
        RECT 42.390 42.260 43.515 42.400 ;
        RECT 42.390 42.200 42.710 42.260 ;
        RECT 43.225 42.215 43.515 42.260 ;
        RECT 49.290 42.200 49.610 42.460 ;
        RECT 54.365 42.400 54.655 42.445 ;
        RECT 59.410 42.400 59.730 42.460 ;
        RECT 60.345 42.400 60.635 42.445 ;
        RECT 64.485 42.400 64.775 42.445 ;
        RECT 54.365 42.260 64.775 42.400 ;
        RECT 65.020 42.400 65.160 42.895 ;
        RECT 66.770 42.880 67.090 43.140 ;
        RECT 68.610 43.080 68.930 43.140 ;
        RECT 78.730 43.080 79.050 43.140 ;
        RECT 81.505 43.080 81.795 43.125 ;
        RECT 68.610 42.940 73.900 43.080 ;
        RECT 68.610 42.880 68.930 42.940 ;
        RECT 73.210 42.740 73.530 42.800 ;
        RECT 71.920 42.600 73.530 42.740 ;
        RECT 68.165 42.400 68.455 42.445 ;
        RECT 65.020 42.260 68.455 42.400 ;
        RECT 54.365 42.215 54.655 42.260 ;
        RECT 23.990 42.060 24.310 42.120 ;
        RECT 29.510 42.060 29.830 42.120 ;
        RECT 23.620 41.920 24.310 42.060 ;
        RECT 23.990 41.860 24.310 41.920 ;
        RECT 25.920 41.920 29.830 42.060 ;
        RECT 16.185 41.720 16.475 41.765 ;
        RECT 14.790 41.580 16.475 41.720 ;
        RECT 14.790 41.520 15.110 41.580 ;
        RECT 16.185 41.535 16.475 41.580 ;
        RECT 16.645 41.720 16.935 41.765 ;
        RECT 20.310 41.720 20.630 41.780 ;
        RECT 25.920 41.765 26.060 41.920 ;
        RECT 29.510 41.860 29.830 41.920 ;
        RECT 33.650 41.860 33.970 42.120 ;
        RECT 34.585 41.875 34.875 42.105 ;
        RECT 35.465 42.060 35.755 42.105 ;
        RECT 36.655 42.060 36.945 42.105 ;
        RECT 39.175 42.060 39.465 42.105 ;
        RECT 35.465 41.920 39.465 42.060 ;
        RECT 35.465 41.875 35.755 41.920 ;
        RECT 36.655 41.875 36.945 41.920 ;
        RECT 39.175 41.875 39.465 41.920 ;
        RECT 42.825 42.060 43.115 42.105 ;
        RECT 44.015 42.060 44.305 42.105 ;
        RECT 46.535 42.060 46.825 42.105 ;
        RECT 42.825 41.920 46.825 42.060 ;
        RECT 42.825 41.875 43.115 41.920 ;
        RECT 44.015 41.875 44.305 41.920 ;
        RECT 46.535 41.875 46.825 41.920 ;
        RECT 47.910 42.060 48.230 42.120 ;
        RECT 54.440 42.060 54.580 42.215 ;
        RECT 59.410 42.200 59.730 42.260 ;
        RECT 60.345 42.215 60.635 42.260 ;
        RECT 64.485 42.215 64.775 42.260 ;
        RECT 68.165 42.215 68.455 42.260 ;
        RECT 68.610 42.200 68.930 42.460 ;
        RECT 69.085 42.400 69.375 42.445 ;
        RECT 69.530 42.400 69.850 42.460 ;
        RECT 69.085 42.260 69.850 42.400 ;
        RECT 69.085 42.215 69.375 42.260 ;
        RECT 69.530 42.200 69.850 42.260 ;
        RECT 69.990 42.400 70.310 42.460 ;
        RECT 71.920 42.445 72.060 42.600 ;
        RECT 73.210 42.540 73.530 42.600 ;
        RECT 70.925 42.400 71.215 42.445 ;
        RECT 69.990 42.260 71.215 42.400 ;
        RECT 69.990 42.200 70.310 42.260 ;
        RECT 70.925 42.215 71.215 42.260 ;
        RECT 71.845 42.215 72.135 42.445 ;
        RECT 72.305 42.215 72.595 42.445 ;
        RECT 72.765 42.400 73.055 42.445 ;
        RECT 73.760 42.400 73.900 42.940 ;
        RECT 78.730 42.940 81.795 43.080 ;
        RECT 78.730 42.880 79.050 42.940 ;
        RECT 81.505 42.895 81.795 42.940 ;
        RECT 74.130 42.740 74.450 42.800 ;
        RECT 75.830 42.740 76.120 42.785 ;
        RECT 74.130 42.600 76.120 42.740 ;
        RECT 74.130 42.540 74.450 42.600 ;
        RECT 75.830 42.555 76.120 42.600 ;
        RECT 78.730 42.400 79.050 42.460 ;
        RECT 72.765 42.260 79.050 42.400 ;
        RECT 72.765 42.215 73.055 42.260 ;
        RECT 47.910 41.920 54.580 42.060 ;
        RECT 16.645 41.580 20.630 41.720 ;
        RECT 16.645 41.535 16.935 41.580 ;
        RECT 20.310 41.520 20.630 41.580 ;
        RECT 25.845 41.535 26.135 41.765 ;
        RECT 27.670 41.520 27.990 41.780 ;
        RECT 31.810 41.720 32.130 41.780 ;
        RECT 34.660 41.720 34.800 41.875 ;
        RECT 47.910 41.860 48.230 41.920 ;
        RECT 54.810 41.860 55.130 42.120 ;
        RECT 61.710 41.860 62.030 42.120 ;
        RECT 65.390 41.860 65.710 42.120 ;
        RECT 66.770 42.060 67.090 42.120 ;
        RECT 68.700 42.060 68.840 42.200 ;
        RECT 72.380 42.060 72.520 42.215 ;
        RECT 66.770 41.920 68.840 42.060 ;
        RECT 71.920 41.920 72.520 42.060 ;
        RECT 66.770 41.860 67.090 41.920 ;
        RECT 71.920 41.780 72.060 41.920 ;
        RECT 31.810 41.580 34.800 41.720 ;
        RECT 35.070 41.720 35.360 41.765 ;
        RECT 37.170 41.720 37.460 41.765 ;
        RECT 38.740 41.720 39.030 41.765 ;
        RECT 35.070 41.580 39.030 41.720 ;
        RECT 31.810 41.520 32.130 41.580 ;
        RECT 35.070 41.535 35.360 41.580 ;
        RECT 37.170 41.535 37.460 41.580 ;
        RECT 38.740 41.535 39.030 41.580 ;
        RECT 42.430 41.720 42.720 41.765 ;
        RECT 44.530 41.720 44.820 41.765 ;
        RECT 46.100 41.720 46.390 41.765 ;
        RECT 42.430 41.580 46.390 41.720 ;
        RECT 42.430 41.535 42.720 41.580 ;
        RECT 44.530 41.535 44.820 41.580 ;
        RECT 46.100 41.535 46.390 41.580 ;
        RECT 71.830 41.520 72.150 41.780 ;
        RECT 15.265 41.380 15.555 41.425 ;
        RECT 15.710 41.380 16.030 41.440 ;
        RECT 15.265 41.240 16.030 41.380 ;
        RECT 15.265 41.195 15.555 41.240 ;
        RECT 15.710 41.180 16.030 41.240 ;
        RECT 23.070 41.380 23.390 41.440 ;
        RECT 24.925 41.380 25.215 41.425 ;
        RECT 26.750 41.380 27.070 41.440 ;
        RECT 23.070 41.240 27.070 41.380 ;
        RECT 23.070 41.180 23.390 41.240 ;
        RECT 24.925 41.195 25.215 41.240 ;
        RECT 26.750 41.180 27.070 41.240 ;
        RECT 48.830 41.380 49.150 41.440 ;
        RECT 53.430 41.380 53.750 41.440 ;
        RECT 56.190 41.380 56.510 41.440 ;
        RECT 48.830 41.240 56.510 41.380 ;
        RECT 48.830 41.180 49.150 41.240 ;
        RECT 53.430 41.180 53.750 41.240 ;
        RECT 56.190 41.180 56.510 41.240 ;
        RECT 58.505 41.380 58.795 41.425 ;
        RECT 58.950 41.380 59.270 41.440 ;
        RECT 58.505 41.240 59.270 41.380 ;
        RECT 58.505 41.195 58.795 41.240 ;
        RECT 58.950 41.180 59.270 41.240 ;
        RECT 64.930 41.380 65.250 41.440 ;
        RECT 72.840 41.380 72.980 42.215 ;
        RECT 78.730 42.200 79.050 42.260 ;
        RECT 74.590 41.860 74.910 42.120 ;
        RECT 75.485 42.060 75.775 42.105 ;
        RECT 76.675 42.060 76.965 42.105 ;
        RECT 79.195 42.060 79.485 42.105 ;
        RECT 75.485 41.920 79.485 42.060 ;
        RECT 75.485 41.875 75.775 41.920 ;
        RECT 76.675 41.875 76.965 41.920 ;
        RECT 79.195 41.875 79.485 41.920 ;
        RECT 74.145 41.720 74.435 41.765 ;
        RECT 75.090 41.720 75.380 41.765 ;
        RECT 77.190 41.720 77.480 41.765 ;
        RECT 78.760 41.720 79.050 41.765 ;
        RECT 74.145 41.580 74.820 41.720 ;
        RECT 74.145 41.535 74.435 41.580 ;
        RECT 64.930 41.240 72.980 41.380 ;
        RECT 74.680 41.380 74.820 41.580 ;
        RECT 75.090 41.580 79.050 41.720 ;
        RECT 75.090 41.535 75.380 41.580 ;
        RECT 77.190 41.535 77.480 41.580 ;
        RECT 78.760 41.535 79.050 41.580 ;
        RECT 75.970 41.380 76.290 41.440 ;
        RECT 74.680 41.240 76.290 41.380 ;
        RECT 64.930 41.180 65.250 41.240 ;
        RECT 75.970 41.180 76.290 41.240 ;
        RECT 5.520 40.560 83.260 41.040 ;
        RECT 13.870 40.360 14.190 40.420 ;
        RECT 7.980 40.220 14.190 40.360 ;
        RECT 7.980 39.725 8.120 40.220 ;
        RECT 13.870 40.160 14.190 40.220 ;
        RECT 14.330 40.360 14.650 40.420 ;
        RECT 14.805 40.360 15.095 40.405 ;
        RECT 26.765 40.360 27.055 40.405 ;
        RECT 32.285 40.360 32.575 40.405 ;
        RECT 14.330 40.220 18.240 40.360 ;
        RECT 14.330 40.160 14.650 40.220 ;
        RECT 14.805 40.175 15.095 40.220 ;
        RECT 8.390 40.020 8.680 40.065 ;
        RECT 10.490 40.020 10.780 40.065 ;
        RECT 12.060 40.020 12.350 40.065 ;
        RECT 8.390 39.880 12.350 40.020 ;
        RECT 8.390 39.835 8.680 39.880 ;
        RECT 10.490 39.835 10.780 39.880 ;
        RECT 12.060 39.835 12.350 39.880 ;
        RECT 12.950 40.020 13.270 40.080 ;
        RECT 18.100 40.065 18.240 40.220 ;
        RECT 26.765 40.220 32.575 40.360 ;
        RECT 26.765 40.175 27.055 40.220 ;
        RECT 32.285 40.175 32.575 40.220 ;
        RECT 40.565 40.360 40.855 40.405 ;
        RECT 41.930 40.360 42.250 40.420 ;
        RECT 40.565 40.220 42.250 40.360 ;
        RECT 40.565 40.175 40.855 40.220 ;
        RECT 41.930 40.160 42.250 40.220 ;
        RECT 44.690 40.160 45.010 40.420 ;
        RECT 46.545 40.175 46.835 40.405 ;
        RECT 47.465 40.360 47.755 40.405 ;
        RECT 55.270 40.360 55.590 40.420 ;
        RECT 47.465 40.220 55.590 40.360 ;
        RECT 47.465 40.175 47.755 40.220 ;
        RECT 15.265 40.020 15.555 40.065 ;
        RECT 12.950 39.880 15.555 40.020 ;
        RECT 12.950 39.820 13.270 39.880 ;
        RECT 15.265 39.835 15.555 39.880 ;
        RECT 18.025 39.835 18.315 40.065 ;
        RECT 20.325 40.020 20.615 40.065 ;
        RECT 27.210 40.020 27.530 40.080 ;
        RECT 20.325 39.880 27.530 40.020 ;
        RECT 20.325 39.835 20.615 39.880 ;
        RECT 7.905 39.495 8.195 39.725 ;
        RECT 8.785 39.680 9.075 39.725 ;
        RECT 9.975 39.680 10.265 39.725 ;
        RECT 12.495 39.680 12.785 39.725 ;
        RECT 8.785 39.540 12.785 39.680 ;
        RECT 15.340 39.680 15.480 39.835 ;
        RECT 27.210 39.820 27.530 39.880 ;
        RECT 28.130 40.020 28.450 40.080 ;
        RECT 28.605 40.020 28.895 40.065 ;
        RECT 29.065 40.020 29.355 40.065 ;
        RECT 28.130 39.880 29.355 40.020 ;
        RECT 28.130 39.820 28.450 39.880 ;
        RECT 28.605 39.835 28.895 39.880 ;
        RECT 29.065 39.835 29.355 39.880 ;
        RECT 31.350 40.020 31.670 40.080 ;
        RECT 46.620 40.020 46.760 40.175 ;
        RECT 55.270 40.160 55.590 40.220 ;
        RECT 56.665 40.360 56.955 40.405 ;
        RECT 58.490 40.360 58.810 40.420 ;
        RECT 60.790 40.360 61.110 40.420 ;
        RECT 56.665 40.220 61.110 40.360 ;
        RECT 56.665 40.175 56.955 40.220 ;
        RECT 58.490 40.160 58.810 40.220 ;
        RECT 60.790 40.160 61.110 40.220 ;
        RECT 63.550 40.360 63.870 40.420 ;
        RECT 66.325 40.360 66.615 40.405 ;
        RECT 67.230 40.360 67.550 40.420 ;
        RECT 63.550 40.220 67.550 40.360 ;
        RECT 63.550 40.160 63.870 40.220 ;
        RECT 66.325 40.175 66.615 40.220 ;
        RECT 67.230 40.160 67.550 40.220 ;
        RECT 80.110 40.360 80.430 40.420 ;
        RECT 81.505 40.360 81.795 40.405 ;
        RECT 80.110 40.220 81.795 40.360 ;
        RECT 80.110 40.160 80.430 40.220 ;
        RECT 81.505 40.175 81.795 40.220 ;
        RECT 48.830 40.020 49.150 40.080 ;
        RECT 31.350 39.880 37.560 40.020 ;
        RECT 46.620 39.880 49.150 40.020 ;
        RECT 31.350 39.820 31.670 39.880 ;
        RECT 34.585 39.680 34.875 39.725 ;
        RECT 15.340 39.540 21.920 39.680 ;
        RECT 8.785 39.495 9.075 39.540 ;
        RECT 9.975 39.495 10.265 39.540 ;
        RECT 12.495 39.495 12.785 39.540 ;
        RECT 7.980 39.340 8.120 39.495 ;
        RECT 8.350 39.340 8.670 39.400 ;
        RECT 9.270 39.385 9.590 39.400 ;
        RECT 9.240 39.340 9.590 39.385 ;
        RECT 7.980 39.200 8.670 39.340 ;
        RECT 9.075 39.200 9.590 39.340 ;
        RECT 8.350 39.140 8.670 39.200 ;
        RECT 9.240 39.155 9.590 39.200 ;
        RECT 9.270 39.140 9.590 39.155 ;
        RECT 15.250 39.340 15.570 39.400 ;
        RECT 17.105 39.340 17.395 39.385 ;
        RECT 17.550 39.340 17.870 39.400 ;
        RECT 19.020 39.385 19.160 39.540 ;
        RECT 15.250 39.200 17.870 39.340 ;
        RECT 15.250 39.140 15.570 39.200 ;
        RECT 17.105 39.155 17.395 39.200 ;
        RECT 17.550 39.140 17.870 39.200 ;
        RECT 18.945 39.155 19.235 39.385 ;
        RECT 19.405 39.340 19.695 39.385 ;
        RECT 19.850 39.340 20.170 39.400 ;
        RECT 19.405 39.200 20.170 39.340 ;
        RECT 19.405 39.155 19.695 39.200 ;
        RECT 19.850 39.140 20.170 39.200 ;
        RECT 20.770 39.140 21.090 39.400 ;
        RECT 21.780 39.385 21.920 39.540 ;
        RECT 30.980 39.540 34.875 39.680 ;
        RECT 21.705 39.155 21.995 39.385 ;
        RECT 28.590 39.340 28.910 39.400 ;
        RECT 30.430 39.340 30.750 39.400 ;
        RECT 30.980 39.385 31.120 39.540 ;
        RECT 34.585 39.495 34.875 39.540 ;
        RECT 30.905 39.340 31.195 39.385 ;
        RECT 28.590 39.200 31.195 39.340 ;
        RECT 28.590 39.140 28.910 39.200 ;
        RECT 30.430 39.140 30.750 39.200 ;
        RECT 30.905 39.155 31.195 39.200 ;
        RECT 31.350 39.340 31.670 39.400 ;
        RECT 33.205 39.340 33.495 39.385 ;
        RECT 31.350 39.200 33.495 39.340 ;
        RECT 31.350 39.140 31.670 39.200 ;
        RECT 33.205 39.155 33.495 39.200 ;
        RECT 33.650 39.140 33.970 39.400 ;
        RECT 37.420 39.385 37.560 39.880 ;
        RECT 48.830 39.820 49.150 39.880 ;
        RECT 50.210 40.020 50.500 40.065 ;
        RECT 51.780 40.020 52.070 40.065 ;
        RECT 53.880 40.020 54.170 40.065 ;
        RECT 50.210 39.880 54.170 40.020 ;
        RECT 50.210 39.835 50.500 39.880 ;
        RECT 51.780 39.835 52.070 39.880 ;
        RECT 53.880 39.835 54.170 39.880 ;
        RECT 58.070 40.020 58.360 40.065 ;
        RECT 60.170 40.020 60.460 40.065 ;
        RECT 61.740 40.020 62.030 40.065 ;
        RECT 58.070 39.880 62.030 40.020 ;
        RECT 58.070 39.835 58.360 39.880 ;
        RECT 60.170 39.835 60.460 39.880 ;
        RECT 61.740 39.835 62.030 39.880 ;
        RECT 64.010 40.020 64.330 40.080 ;
        RECT 64.485 40.020 64.775 40.065 ;
        RECT 74.130 40.020 74.450 40.080 ;
        RECT 64.010 39.880 74.450 40.020 ;
        RECT 64.010 39.820 64.330 39.880 ;
        RECT 64.485 39.835 64.775 39.880 ;
        RECT 74.130 39.820 74.450 39.880 ;
        RECT 75.090 40.020 75.380 40.065 ;
        RECT 77.190 40.020 77.480 40.065 ;
        RECT 78.760 40.020 79.050 40.065 ;
        RECT 75.090 39.880 79.050 40.020 ;
        RECT 75.090 39.835 75.380 39.880 ;
        RECT 77.190 39.835 77.480 39.880 ;
        RECT 78.760 39.835 79.050 39.880 ;
        RECT 42.850 39.680 43.170 39.740 ;
        RECT 43.325 39.680 43.615 39.725 ;
        RECT 46.085 39.680 46.375 39.725 ;
        RECT 42.850 39.540 46.375 39.680 ;
        RECT 42.850 39.480 43.170 39.540 ;
        RECT 43.325 39.495 43.615 39.540 ;
        RECT 46.085 39.495 46.375 39.540 ;
        RECT 49.775 39.680 50.065 39.725 ;
        RECT 52.295 39.680 52.585 39.725 ;
        RECT 53.485 39.680 53.775 39.725 ;
        RECT 57.585 39.680 57.875 39.725 ;
        RECT 49.775 39.540 53.775 39.680 ;
        RECT 49.775 39.495 50.065 39.540 ;
        RECT 52.295 39.495 52.585 39.540 ;
        RECT 53.485 39.495 53.775 39.540 ;
        RECT 54.440 39.540 57.875 39.680 ;
        RECT 34.125 39.155 34.415 39.385 ;
        RECT 37.345 39.155 37.635 39.385 ;
        RECT 39.185 39.155 39.475 39.385 ;
        RECT 40.105 39.340 40.395 39.385 ;
        RECT 46.545 39.340 46.835 39.385 ;
        RECT 40.105 39.200 46.835 39.340 ;
        RECT 40.105 39.155 40.395 39.200 ;
        RECT 46.545 39.155 46.835 39.200 ;
        RECT 49.290 39.340 49.610 39.400 ;
        RECT 54.440 39.385 54.580 39.540 ;
        RECT 57.585 39.495 57.875 39.540 ;
        RECT 58.465 39.680 58.755 39.725 ;
        RECT 59.655 39.680 59.945 39.725 ;
        RECT 62.175 39.680 62.465 39.725 ;
        RECT 58.465 39.540 62.465 39.680 ;
        RECT 58.465 39.495 58.755 39.540 ;
        RECT 59.655 39.495 59.945 39.540 ;
        RECT 62.175 39.495 62.465 39.540 ;
        RECT 62.630 39.680 62.950 39.740 ;
        RECT 74.590 39.680 74.910 39.740 ;
        RECT 62.630 39.540 74.910 39.680 ;
        RECT 62.630 39.480 62.950 39.540 ;
        RECT 74.590 39.480 74.910 39.540 ;
        RECT 75.485 39.680 75.775 39.725 ;
        RECT 76.675 39.680 76.965 39.725 ;
        RECT 79.195 39.680 79.485 39.725 ;
        RECT 75.485 39.540 79.485 39.680 ;
        RECT 75.485 39.495 75.775 39.540 ;
        RECT 76.675 39.495 76.965 39.540 ;
        RECT 79.195 39.495 79.485 39.540 ;
        RECT 54.365 39.340 54.655 39.385 ;
        RECT 49.290 39.200 54.655 39.340 ;
        RECT 12.030 39.000 12.350 39.060 ;
        RECT 16.185 39.000 16.475 39.045 ;
        RECT 20.325 39.000 20.615 39.045 ;
        RECT 12.030 38.860 16.475 39.000 ;
        RECT 12.030 38.800 12.350 38.860 ;
        RECT 16.185 38.815 16.475 38.860 ;
        RECT 17.180 38.860 20.615 39.000 ;
        RECT 17.180 38.720 17.320 38.860 ;
        RECT 20.325 38.815 20.615 38.860 ;
        RECT 23.990 39.000 24.310 39.060 ;
        RECT 31.825 39.000 32.115 39.045 ;
        RECT 34.200 39.000 34.340 39.155 ;
        RECT 34.570 39.000 34.890 39.060 ;
        RECT 36.425 39.000 36.715 39.045 ;
        RECT 23.990 38.860 36.715 39.000 ;
        RECT 39.260 39.000 39.400 39.155 ;
        RECT 45.610 39.000 45.930 39.060 ;
        RECT 39.260 38.860 45.930 39.000 ;
        RECT 46.620 39.000 46.760 39.155 ;
        RECT 49.290 39.140 49.610 39.200 ;
        RECT 54.365 39.155 54.655 39.200 ;
        RECT 54.825 39.155 55.115 39.385 ;
        RECT 55.745 39.340 56.035 39.385 ;
        RECT 56.190 39.340 56.510 39.400 ;
        RECT 58.950 39.385 59.270 39.400 ;
        RECT 58.920 39.340 59.270 39.385 ;
        RECT 55.745 39.200 56.510 39.340 ;
        RECT 58.755 39.200 59.270 39.340 ;
        RECT 55.745 39.155 56.035 39.200 ;
        RECT 52.050 39.000 52.370 39.060 ;
        RECT 46.620 38.860 52.370 39.000 ;
        RECT 23.990 38.800 24.310 38.860 ;
        RECT 31.825 38.815 32.115 38.860 ;
        RECT 34.570 38.800 34.890 38.860 ;
        RECT 36.425 38.815 36.715 38.860 ;
        RECT 45.610 38.800 45.930 38.860 ;
        RECT 52.050 38.800 52.370 38.860 ;
        RECT 52.970 39.045 53.290 39.060 ;
        RECT 52.970 39.000 53.320 39.045 ;
        RECT 52.970 38.860 53.485 39.000 ;
        RECT 52.970 38.815 53.320 38.860 ;
        RECT 52.970 38.800 53.290 38.815 ;
        RECT 14.330 38.660 14.650 38.720 ;
        RECT 15.710 38.660 16.030 38.720 ;
        RECT 16.645 38.660 16.935 38.705 ;
        RECT 14.330 38.520 16.935 38.660 ;
        RECT 14.330 38.460 14.650 38.520 ;
        RECT 15.710 38.460 16.030 38.520 ;
        RECT 16.645 38.475 16.935 38.520 ;
        RECT 17.090 38.460 17.410 38.720 ;
        RECT 21.230 38.460 21.550 38.720 ;
        RECT 25.845 38.660 26.135 38.705 ;
        RECT 26.290 38.660 26.610 38.720 ;
        RECT 25.845 38.520 26.610 38.660 ;
        RECT 25.845 38.475 26.135 38.520 ;
        RECT 26.290 38.460 26.610 38.520 ;
        RECT 26.750 38.660 27.070 38.720 ;
        RECT 28.590 38.660 28.910 38.720 ;
        RECT 26.750 38.520 28.910 38.660 ;
        RECT 26.750 38.460 27.070 38.520 ;
        RECT 28.590 38.460 28.910 38.520 ;
        RECT 29.970 38.460 30.290 38.720 ;
        RECT 30.430 38.660 30.750 38.720 ;
        RECT 33.650 38.660 33.970 38.720 ;
        RECT 30.430 38.520 33.970 38.660 ;
        RECT 30.430 38.460 30.750 38.520 ;
        RECT 33.650 38.460 33.970 38.520 ;
        RECT 35.490 38.460 35.810 38.720 ;
        RECT 40.105 38.660 40.395 38.705 ;
        RECT 49.750 38.660 50.070 38.720 ;
        RECT 54.900 38.660 55.040 39.155 ;
        RECT 56.190 39.140 56.510 39.200 ;
        RECT 58.920 39.155 59.270 39.200 ;
        RECT 58.950 39.140 59.270 39.155 ;
        RECT 64.470 39.340 64.790 39.400 ;
        RECT 66.325 39.340 66.615 39.385 ;
        RECT 67.690 39.340 68.010 39.400 ;
        RECT 64.470 39.200 68.010 39.340 ;
        RECT 64.470 39.140 64.790 39.200 ;
        RECT 66.325 39.155 66.615 39.200 ;
        RECT 67.690 39.140 68.010 39.200 ;
        RECT 68.150 39.140 68.470 39.400 ;
        RECT 68.610 39.340 68.930 39.400 ;
        RECT 69.990 39.340 70.310 39.400 ;
        RECT 70.465 39.340 70.755 39.385 ;
        RECT 68.610 39.200 70.755 39.340 ;
        RECT 68.610 39.140 68.930 39.200 ;
        RECT 69.990 39.140 70.310 39.200 ;
        RECT 70.465 39.155 70.755 39.200 ;
        RECT 71.370 39.140 71.690 39.400 ;
        RECT 71.830 39.140 72.150 39.400 ;
        RECT 72.290 39.140 72.610 39.400 ;
        RECT 75.970 39.385 76.290 39.400 ;
        RECT 75.940 39.340 76.290 39.385 ;
        RECT 75.775 39.200 76.290 39.340 ;
        RECT 75.940 39.155 76.290 39.200 ;
        RECT 75.970 39.140 76.290 39.155 ;
        RECT 60.790 39.000 61.110 39.060 ;
        RECT 71.920 39.000 72.060 39.140 ;
        RECT 75.510 39.000 75.830 39.060 ;
        RECT 60.790 38.860 65.620 39.000 ;
        RECT 71.920 38.860 75.830 39.000 ;
        RECT 60.790 38.800 61.110 38.860 ;
        RECT 65.480 38.705 65.620 38.860 ;
        RECT 75.510 38.800 75.830 38.860 ;
        RECT 40.105 38.520 55.040 38.660 ;
        RECT 40.105 38.475 40.395 38.520 ;
        RECT 49.750 38.460 50.070 38.520 ;
        RECT 65.405 38.475 65.695 38.705 ;
        RECT 73.670 38.460 73.990 38.720 ;
        RECT 74.130 38.660 74.450 38.720 ;
        RECT 75.050 38.660 75.370 38.720 ;
        RECT 81.490 38.660 81.810 38.720 ;
        RECT 74.130 38.520 81.810 38.660 ;
        RECT 74.130 38.460 74.450 38.520 ;
        RECT 75.050 38.460 75.370 38.520 ;
        RECT 81.490 38.460 81.810 38.520 ;
        RECT 5.520 37.840 83.260 38.320 ;
        RECT 14.790 37.640 15.110 37.700 ;
        RECT 7.060 37.500 15.110 37.640 ;
        RECT 7.060 37.005 7.200 37.500 ;
        RECT 14.790 37.440 15.110 37.500 ;
        RECT 15.250 37.440 15.570 37.700 ;
        RECT 15.725 37.455 16.015 37.685 ;
        RECT 16.565 37.640 16.855 37.685 ;
        RECT 21.230 37.640 21.550 37.700 ;
        RECT 16.565 37.500 21.550 37.640 ;
        RECT 16.565 37.455 16.855 37.500 ;
        RECT 7.430 37.100 7.750 37.360 ;
        RECT 9.700 37.300 9.990 37.345 ;
        RECT 15.800 37.300 15.940 37.455 ;
        RECT 21.230 37.440 21.550 37.500 ;
        RECT 23.530 37.440 23.850 37.700 ;
        RECT 30.430 37.640 30.750 37.700 ;
        RECT 24.540 37.500 30.750 37.640 ;
        RECT 9.700 37.160 15.940 37.300 ;
        RECT 9.700 37.115 9.990 37.160 ;
        RECT 17.565 37.115 17.855 37.345 ;
        RECT 23.085 37.300 23.375 37.345 ;
        RECT 24.540 37.300 24.680 37.500 ;
        RECT 30.430 37.440 30.750 37.500 ;
        RECT 30.890 37.440 31.210 37.700 ;
        RECT 40.565 37.640 40.855 37.685 ;
        RECT 42.390 37.640 42.710 37.700 ;
        RECT 47.910 37.640 48.230 37.700 ;
        RECT 40.565 37.500 42.710 37.640 ;
        RECT 40.565 37.455 40.855 37.500 ;
        RECT 42.390 37.440 42.710 37.500 ;
        RECT 42.940 37.500 48.230 37.640 ;
        RECT 42.940 37.300 43.080 37.500 ;
        RECT 47.910 37.440 48.230 37.500 ;
        RECT 56.650 37.640 56.970 37.700 ;
        RECT 68.150 37.640 68.470 37.700 ;
        RECT 56.650 37.500 68.470 37.640 ;
        RECT 56.650 37.440 56.970 37.500 ;
        RECT 68.150 37.440 68.470 37.500 ;
        RECT 81.030 37.440 81.350 37.700 ;
        RECT 49.290 37.300 49.610 37.360 ;
        RECT 62.630 37.300 62.950 37.360 ;
        RECT 74.590 37.300 74.910 37.360 ;
        RECT 23.085 37.160 24.680 37.300 ;
        RECT 25.000 37.160 28.360 37.300 ;
        RECT 23.085 37.115 23.375 37.160 ;
        RECT 6.985 36.775 7.275 37.005 ;
        RECT 7.890 36.760 8.210 37.020 ;
        RECT 8.350 36.760 8.670 37.020 ;
        RECT 11.110 36.960 11.430 37.020 ;
        RECT 17.640 36.960 17.780 37.115 ;
        RECT 18.485 36.960 18.775 37.005 ;
        RECT 11.110 36.820 18.775 36.960 ;
        RECT 11.110 36.760 11.430 36.820 ;
        RECT 18.485 36.775 18.775 36.820 ;
        RECT 19.405 36.775 19.695 37.005 ;
        RECT 9.245 36.620 9.535 36.665 ;
        RECT 10.435 36.620 10.725 36.665 ;
        RECT 12.955 36.620 13.245 36.665 ;
        RECT 19.480 36.620 19.620 36.775 ;
        RECT 19.850 36.760 20.170 37.020 ;
        RECT 20.310 36.760 20.630 37.020 ;
        RECT 22.165 36.775 22.455 37.005 ;
        RECT 9.245 36.480 13.245 36.620 ;
        RECT 9.245 36.435 9.535 36.480 ;
        RECT 10.435 36.435 10.725 36.480 ;
        RECT 12.955 36.435 13.245 36.480 ;
        RECT 16.720 36.480 19.620 36.620 ;
        RECT 22.240 36.620 22.380 36.775 ;
        RECT 23.530 36.760 23.850 37.020 ;
        RECT 24.005 36.960 24.295 37.005 ;
        RECT 25.000 36.960 25.140 37.160 ;
        RECT 28.220 37.020 28.360 37.160 ;
        RECT 39.260 37.160 43.080 37.300 ;
        RECT 45.240 37.160 49.610 37.300 ;
        RECT 24.005 36.820 25.140 36.960 ;
        RECT 25.340 36.960 25.630 37.005 ;
        RECT 26.750 36.960 27.070 37.020 ;
        RECT 25.340 36.820 27.070 36.960 ;
        RECT 24.005 36.775 24.295 36.820 ;
        RECT 25.340 36.775 25.630 36.820 ;
        RECT 26.750 36.760 27.070 36.820 ;
        RECT 28.130 36.960 28.450 37.020 ;
        RECT 31.810 36.960 32.130 37.020 ;
        RECT 28.130 36.820 32.130 36.960 ;
        RECT 28.130 36.760 28.450 36.820 ;
        RECT 31.810 36.760 32.130 36.820 ;
        RECT 33.160 36.960 33.450 37.005 ;
        RECT 35.030 36.960 35.350 37.020 ;
        RECT 39.260 37.005 39.400 37.160 ;
        RECT 33.160 36.820 35.350 36.960 ;
        RECT 33.160 36.775 33.450 36.820 ;
        RECT 35.030 36.760 35.350 36.820 ;
        RECT 39.185 36.775 39.475 37.005 ;
        RECT 39.645 36.960 39.935 37.005 ;
        RECT 41.470 36.960 41.790 37.020 ;
        RECT 39.645 36.820 41.790 36.960 ;
        RECT 39.645 36.775 39.935 36.820 ;
        RECT 41.470 36.760 41.790 36.820 ;
        RECT 41.945 36.960 42.235 37.005 ;
        RECT 43.770 36.960 44.090 37.020 ;
        RECT 45.240 37.005 45.380 37.160 ;
        RECT 49.290 37.100 49.610 37.160 ;
        RECT 57.660 37.160 65.620 37.300 ;
        RECT 41.945 36.820 44.090 36.960 ;
        RECT 41.945 36.775 42.235 36.820 ;
        RECT 43.770 36.760 44.090 36.820 ;
        RECT 45.165 36.775 45.455 37.005 ;
        RECT 46.445 36.960 46.735 37.005 ;
        RECT 45.700 36.820 46.735 36.960 ;
        RECT 24.885 36.620 25.175 36.665 ;
        RECT 26.075 36.620 26.365 36.665 ;
        RECT 28.595 36.620 28.885 36.665 ;
        RECT 22.240 36.480 24.220 36.620 ;
        RECT 8.850 36.280 9.140 36.325 ;
        RECT 10.950 36.280 11.240 36.325 ;
        RECT 12.520 36.280 12.810 36.325 ;
        RECT 8.850 36.140 12.810 36.280 ;
        RECT 8.850 36.095 9.140 36.140 ;
        RECT 10.950 36.095 11.240 36.140 ;
        RECT 12.520 36.095 12.810 36.140 ;
        RECT 9.730 35.940 10.050 36.000 ;
        RECT 11.570 35.940 11.890 36.000 ;
        RECT 16.720 35.985 16.860 36.480 ;
        RECT 21.705 36.280 21.995 36.325 ;
        RECT 23.070 36.280 23.390 36.340 ;
        RECT 21.705 36.140 23.390 36.280 ;
        RECT 21.705 36.095 21.995 36.140 ;
        RECT 23.070 36.080 23.390 36.140 ;
        RECT 16.645 35.940 16.935 35.985 ;
        RECT 9.730 35.800 16.935 35.940 ;
        RECT 24.080 35.940 24.220 36.480 ;
        RECT 24.885 36.480 28.885 36.620 ;
        RECT 24.885 36.435 25.175 36.480 ;
        RECT 26.075 36.435 26.365 36.480 ;
        RECT 28.595 36.435 28.885 36.480 ;
        RECT 32.705 36.620 32.995 36.665 ;
        RECT 33.895 36.620 34.185 36.665 ;
        RECT 36.415 36.620 36.705 36.665 ;
        RECT 32.705 36.480 36.705 36.620 ;
        RECT 32.705 36.435 32.995 36.480 ;
        RECT 33.895 36.435 34.185 36.480 ;
        RECT 36.415 36.435 36.705 36.480 ;
        RECT 40.565 36.620 40.855 36.665 ;
        RECT 41.010 36.620 41.330 36.680 ;
        RECT 40.565 36.480 41.330 36.620 ;
        RECT 40.565 36.435 40.855 36.480 ;
        RECT 41.010 36.420 41.330 36.480 ;
        RECT 42.405 36.620 42.695 36.665 ;
        RECT 43.310 36.620 43.630 36.680 ;
        RECT 45.700 36.620 45.840 36.820 ;
        RECT 46.445 36.775 46.735 36.820 ;
        RECT 48.370 36.960 48.690 37.020 ;
        RECT 52.525 36.960 52.815 37.005 ;
        RECT 48.370 36.820 52.815 36.960 ;
        RECT 48.370 36.760 48.690 36.820 ;
        RECT 52.525 36.775 52.815 36.820 ;
        RECT 55.730 36.760 56.050 37.020 ;
        RECT 57.660 37.005 57.800 37.160 ;
        RECT 62.630 37.100 62.950 37.160 ;
        RECT 57.585 36.775 57.875 37.005 ;
        RECT 58.030 36.960 58.350 37.020 ;
        RECT 65.480 37.005 65.620 37.160 ;
        RECT 74.590 37.160 79.880 37.300 ;
        RECT 74.590 37.100 74.910 37.160 ;
        RECT 58.865 36.960 59.155 37.005 ;
        RECT 58.030 36.820 59.155 36.960 ;
        RECT 58.030 36.760 58.350 36.820 ;
        RECT 58.865 36.775 59.155 36.820 ;
        RECT 65.405 36.775 65.695 37.005 ;
        RECT 65.850 36.960 66.170 37.020 ;
        RECT 66.685 36.960 66.975 37.005 ;
        RECT 65.850 36.820 66.975 36.960 ;
        RECT 65.850 36.760 66.170 36.820 ;
        RECT 66.685 36.775 66.975 36.820 ;
        RECT 73.670 36.960 73.990 37.020 ;
        RECT 79.740 37.005 79.880 37.160 ;
        RECT 78.330 36.960 78.620 37.005 ;
        RECT 73.670 36.820 78.620 36.960 ;
        RECT 73.670 36.760 73.990 36.820 ;
        RECT 78.330 36.775 78.620 36.820 ;
        RECT 79.665 36.775 79.955 37.005 ;
        RECT 80.110 36.760 80.430 37.020 ;
        RECT 42.405 36.480 43.630 36.620 ;
        RECT 42.405 36.435 42.695 36.480 ;
        RECT 43.310 36.420 43.630 36.480 ;
        RECT 43.860 36.480 45.840 36.620 ;
        RECT 46.045 36.620 46.335 36.665 ;
        RECT 47.235 36.620 47.525 36.665 ;
        RECT 49.755 36.620 50.045 36.665 ;
        RECT 46.045 36.480 50.045 36.620 ;
        RECT 43.860 36.325 44.000 36.480 ;
        RECT 46.045 36.435 46.335 36.480 ;
        RECT 47.235 36.435 47.525 36.480 ;
        RECT 49.755 36.435 50.045 36.480 ;
        RECT 58.465 36.620 58.755 36.665 ;
        RECT 59.655 36.620 59.945 36.665 ;
        RECT 62.175 36.620 62.465 36.665 ;
        RECT 58.465 36.480 62.465 36.620 ;
        RECT 58.465 36.435 58.755 36.480 ;
        RECT 59.655 36.435 59.945 36.480 ;
        RECT 62.175 36.435 62.465 36.480 ;
        RECT 66.285 36.620 66.575 36.665 ;
        RECT 67.475 36.620 67.765 36.665 ;
        RECT 69.995 36.620 70.285 36.665 ;
        RECT 66.285 36.480 70.285 36.620 ;
        RECT 66.285 36.435 66.575 36.480 ;
        RECT 67.475 36.435 67.765 36.480 ;
        RECT 69.995 36.435 70.285 36.480 ;
        RECT 75.075 36.620 75.365 36.665 ;
        RECT 77.595 36.620 77.885 36.665 ;
        RECT 78.785 36.620 79.075 36.665 ;
        RECT 75.075 36.480 79.075 36.620 ;
        RECT 75.075 36.435 75.365 36.480 ;
        RECT 77.595 36.435 77.885 36.480 ;
        RECT 78.785 36.435 79.075 36.480 ;
        RECT 24.490 36.280 24.780 36.325 ;
        RECT 26.590 36.280 26.880 36.325 ;
        RECT 28.160 36.280 28.450 36.325 ;
        RECT 24.490 36.140 28.450 36.280 ;
        RECT 24.490 36.095 24.780 36.140 ;
        RECT 26.590 36.095 26.880 36.140 ;
        RECT 28.160 36.095 28.450 36.140 ;
        RECT 32.310 36.280 32.600 36.325 ;
        RECT 34.410 36.280 34.700 36.325 ;
        RECT 35.980 36.280 36.270 36.325 ;
        RECT 32.310 36.140 36.270 36.280 ;
        RECT 32.310 36.095 32.600 36.140 ;
        RECT 34.410 36.095 34.700 36.140 ;
        RECT 35.980 36.095 36.270 36.140 ;
        RECT 43.785 36.095 44.075 36.325 ;
        RECT 45.650 36.280 45.940 36.325 ;
        RECT 47.750 36.280 48.040 36.325 ;
        RECT 49.320 36.280 49.610 36.325 ;
        RECT 45.650 36.140 49.610 36.280 ;
        RECT 45.650 36.095 45.940 36.140 ;
        RECT 47.750 36.095 48.040 36.140 ;
        RECT 49.320 36.095 49.610 36.140 ;
        RECT 58.070 36.280 58.360 36.325 ;
        RECT 60.170 36.280 60.460 36.325 ;
        RECT 61.740 36.280 62.030 36.325 ;
        RECT 58.070 36.140 62.030 36.280 ;
        RECT 58.070 36.095 58.360 36.140 ;
        RECT 60.170 36.095 60.460 36.140 ;
        RECT 61.740 36.095 62.030 36.140 ;
        RECT 64.485 36.280 64.775 36.325 ;
        RECT 64.930 36.280 65.250 36.340 ;
        RECT 64.485 36.140 65.250 36.280 ;
        RECT 64.485 36.095 64.775 36.140 ;
        RECT 64.930 36.080 65.250 36.140 ;
        RECT 65.890 36.280 66.180 36.325 ;
        RECT 67.990 36.280 68.280 36.325 ;
        RECT 69.560 36.280 69.850 36.325 ;
        RECT 65.890 36.140 69.850 36.280 ;
        RECT 65.890 36.095 66.180 36.140 ;
        RECT 67.990 36.095 68.280 36.140 ;
        RECT 69.560 36.095 69.850 36.140 ;
        RECT 75.510 36.280 75.800 36.325 ;
        RECT 77.080 36.280 77.370 36.325 ;
        RECT 79.180 36.280 79.470 36.325 ;
        RECT 75.510 36.140 79.470 36.280 ;
        RECT 75.510 36.095 75.800 36.140 ;
        RECT 77.080 36.095 77.370 36.140 ;
        RECT 79.180 36.095 79.470 36.140 ;
        RECT 29.970 35.940 30.290 36.000 ;
        RECT 33.190 35.940 33.510 36.000 ;
        RECT 38.725 35.940 39.015 35.985 ;
        RECT 40.090 35.940 40.410 36.000 ;
        RECT 24.080 35.800 40.410 35.940 ;
        RECT 9.730 35.740 10.050 35.800 ;
        RECT 11.570 35.740 11.890 35.800 ;
        RECT 16.645 35.755 16.935 35.800 ;
        RECT 29.970 35.740 30.290 35.800 ;
        RECT 33.190 35.740 33.510 35.800 ;
        RECT 38.725 35.755 39.015 35.800 ;
        RECT 40.090 35.740 40.410 35.800 ;
        RECT 52.050 35.940 52.370 36.000 ;
        RECT 53.890 35.940 54.210 36.000 ;
        RECT 52.050 35.800 54.210 35.940 ;
        RECT 52.050 35.740 52.370 35.800 ;
        RECT 53.890 35.740 54.210 35.800 ;
        RECT 69.990 35.940 70.310 36.000 ;
        RECT 72.305 35.940 72.595 35.985 ;
        RECT 69.990 35.800 72.595 35.940 ;
        RECT 69.990 35.740 70.310 35.800 ;
        RECT 72.305 35.755 72.595 35.800 ;
        RECT 72.750 35.740 73.070 36.000 ;
        RECT 5.520 35.120 83.260 35.600 ;
        RECT 11.570 34.920 11.890 34.980 ;
        RECT 14.805 34.920 15.095 34.965 ;
        RECT 11.570 34.780 15.095 34.920 ;
        RECT 11.570 34.720 11.890 34.780 ;
        RECT 14.805 34.735 15.095 34.780 ;
        RECT 12.030 34.580 12.350 34.640 ;
        RECT 8.900 34.440 12.350 34.580 ;
        RECT 14.880 34.580 15.020 34.735 ;
        RECT 15.710 34.720 16.030 34.980 ;
        RECT 17.090 34.720 17.410 34.980 ;
        RECT 23.990 34.920 24.310 34.980 ;
        RECT 17.640 34.780 24.310 34.920 ;
        RECT 17.640 34.580 17.780 34.780 ;
        RECT 23.990 34.720 24.310 34.780 ;
        RECT 25.830 34.720 26.150 34.980 ;
        RECT 28.590 34.920 28.910 34.980 ;
        RECT 30.890 34.920 31.210 34.980 ;
        RECT 33.650 34.920 33.970 34.980 ;
        RECT 34.585 34.920 34.875 34.965 ;
        RECT 28.590 34.780 33.420 34.920 ;
        RECT 28.590 34.720 28.910 34.780 ;
        RECT 30.890 34.720 31.210 34.780 ;
        RECT 14.880 34.440 17.780 34.580 ;
        RECT 19.430 34.580 19.720 34.625 ;
        RECT 21.530 34.580 21.820 34.625 ;
        RECT 23.100 34.580 23.390 34.625 ;
        RECT 19.430 34.440 23.390 34.580 ;
        RECT 8.900 34.285 9.040 34.440 ;
        RECT 12.030 34.380 12.350 34.440 ;
        RECT 19.430 34.395 19.720 34.440 ;
        RECT 21.530 34.395 21.820 34.440 ;
        RECT 23.100 34.395 23.390 34.440 ;
        RECT 28.170 34.580 28.460 34.625 ;
        RECT 30.270 34.580 30.560 34.625 ;
        RECT 31.840 34.580 32.130 34.625 ;
        RECT 28.170 34.440 32.130 34.580 ;
        RECT 33.280 34.580 33.420 34.780 ;
        RECT 33.650 34.780 34.875 34.920 ;
        RECT 33.650 34.720 33.970 34.780 ;
        RECT 34.585 34.735 34.875 34.780 ;
        RECT 35.030 34.720 35.350 34.980 ;
        RECT 35.965 34.735 36.255 34.965 ;
        RECT 36.040 34.580 36.180 34.735 ;
        RECT 56.650 34.720 56.970 34.980 ;
        RECT 57.585 34.920 57.875 34.965 ;
        RECT 58.030 34.920 58.350 34.980 ;
        RECT 57.585 34.780 58.350 34.920 ;
        RECT 57.585 34.735 57.875 34.780 ;
        RECT 58.030 34.720 58.350 34.780 ;
        RECT 64.945 34.920 65.235 34.965 ;
        RECT 65.850 34.920 66.170 34.980 ;
        RECT 64.945 34.780 66.170 34.920 ;
        RECT 64.945 34.735 65.235 34.780 ;
        RECT 65.850 34.720 66.170 34.780 ;
        RECT 72.290 34.920 72.610 34.980 ;
        RECT 73.225 34.920 73.515 34.965 ;
        RECT 72.290 34.780 73.515 34.920 ;
        RECT 72.290 34.720 72.610 34.780 ;
        RECT 73.225 34.735 73.515 34.780 ;
        RECT 33.280 34.440 36.180 34.580 ;
        RECT 75.090 34.580 75.380 34.625 ;
        RECT 77.190 34.580 77.480 34.625 ;
        RECT 78.760 34.580 79.050 34.625 ;
        RECT 75.090 34.440 79.050 34.580 ;
        RECT 28.170 34.395 28.460 34.440 ;
        RECT 30.270 34.395 30.560 34.440 ;
        RECT 31.840 34.395 32.130 34.440 ;
        RECT 75.090 34.395 75.380 34.440 ;
        RECT 77.190 34.395 77.480 34.440 ;
        RECT 78.760 34.395 79.050 34.440 ;
        RECT 8.825 34.055 9.115 34.285 ;
        RECT 10.205 34.240 10.495 34.285 ;
        RECT 11.570 34.240 11.890 34.300 ;
        RECT 10.205 34.100 11.890 34.240 ;
        RECT 10.205 34.055 10.495 34.100 ;
        RECT 11.570 34.040 11.890 34.100 ;
        RECT 13.870 34.240 14.190 34.300 ;
        RECT 16.170 34.240 16.490 34.300 ;
        RECT 18.945 34.240 19.235 34.285 ;
        RECT 13.870 34.100 19.235 34.240 ;
        RECT 13.870 34.040 14.190 34.100 ;
        RECT 16.170 34.040 16.490 34.100 ;
        RECT 18.945 34.055 19.235 34.100 ;
        RECT 19.825 34.240 20.115 34.285 ;
        RECT 21.015 34.240 21.305 34.285 ;
        RECT 23.535 34.240 23.825 34.285 ;
        RECT 19.825 34.100 23.825 34.240 ;
        RECT 19.825 34.055 20.115 34.100 ;
        RECT 21.015 34.055 21.305 34.100 ;
        RECT 23.535 34.055 23.825 34.100 ;
        RECT 28.565 34.240 28.855 34.285 ;
        RECT 29.755 34.240 30.045 34.285 ;
        RECT 32.275 34.240 32.565 34.285 ;
        RECT 28.565 34.100 32.565 34.240 ;
        RECT 28.565 34.055 28.855 34.100 ;
        RECT 29.755 34.055 30.045 34.100 ;
        RECT 32.275 34.055 32.565 34.100 ;
        RECT 45.610 34.240 45.930 34.300 ;
        RECT 46.085 34.240 46.375 34.285 ;
        RECT 45.610 34.100 46.375 34.240 ;
        RECT 45.610 34.040 45.930 34.100 ;
        RECT 46.085 34.055 46.375 34.100 ;
        RECT 52.985 34.240 53.275 34.285 ;
        RECT 55.270 34.240 55.590 34.300 ;
        RECT 55.870 34.240 56.160 34.285 ;
        RECT 52.985 34.100 56.160 34.240 ;
        RECT 52.985 34.055 53.275 34.100 ;
        RECT 55.270 34.040 55.590 34.100 ;
        RECT 55.870 34.055 56.160 34.100 ;
        RECT 60.790 34.040 61.110 34.300 ;
        RECT 74.590 34.040 74.910 34.300 ;
        RECT 75.485 34.240 75.775 34.285 ;
        RECT 76.675 34.240 76.965 34.285 ;
        RECT 79.195 34.240 79.485 34.285 ;
        RECT 75.485 34.100 79.485 34.240 ;
        RECT 75.485 34.055 75.775 34.100 ;
        RECT 76.675 34.055 76.965 34.100 ;
        RECT 79.195 34.055 79.485 34.100 ;
        RECT 8.365 33.900 8.655 33.945 ;
        RECT 14.330 33.900 14.650 33.960 ;
        RECT 19.390 33.900 19.710 33.960 ;
        RECT 8.365 33.760 14.650 33.900 ;
        RECT 8.365 33.715 8.655 33.760 ;
        RECT 14.330 33.700 14.650 33.760 ;
        RECT 16.390 33.760 19.710 33.900 ;
        RECT 16.390 33.730 16.530 33.760 ;
        RECT 10.665 33.560 10.955 33.605 ;
        RECT 11.110 33.560 11.430 33.620 ;
        RECT 10.665 33.420 11.430 33.560 ;
        RECT 10.665 33.375 10.955 33.420 ;
        RECT 11.110 33.360 11.430 33.420 ;
        RECT 11.570 33.605 11.890 33.620 ;
        RECT 11.570 33.375 11.955 33.605 ;
        RECT 13.410 33.560 13.730 33.620 ;
        RECT 14.790 33.605 15.110 33.620 ;
        RECT 16.260 33.605 16.530 33.730 ;
        RECT 19.390 33.700 19.710 33.760 ;
        RECT 20.280 33.900 20.570 33.945 ;
        RECT 23.070 33.900 23.390 33.960 ;
        RECT 26.305 33.900 26.595 33.945 ;
        RECT 20.280 33.760 23.390 33.900 ;
        RECT 20.280 33.715 20.570 33.760 ;
        RECT 23.070 33.700 23.390 33.760 ;
        RECT 24.540 33.760 26.595 33.900 ;
        RECT 13.885 33.560 14.175 33.605 ;
        RECT 12.120 33.420 14.175 33.560 ;
        RECT 11.570 33.360 11.890 33.375 ;
        RECT 11.200 33.220 11.340 33.360 ;
        RECT 12.120 33.220 12.260 33.420 ;
        RECT 13.410 33.360 13.730 33.420 ;
        RECT 13.885 33.375 14.175 33.420 ;
        RECT 14.790 33.375 15.175 33.605 ;
        RECT 16.185 33.590 16.530 33.605 ;
        RECT 16.185 33.375 16.475 33.590 ;
        RECT 14.790 33.360 15.110 33.375 ;
        RECT 11.200 33.080 12.260 33.220 ;
        RECT 12.490 33.020 12.810 33.280 ;
        RECT 12.950 33.220 13.270 33.280 ;
        RECT 14.330 33.220 14.650 33.280 ;
        RECT 17.185 33.220 17.475 33.265 ;
        RECT 12.950 33.080 17.475 33.220 ;
        RECT 12.950 33.020 13.270 33.080 ;
        RECT 14.330 33.020 14.650 33.080 ;
        RECT 17.185 33.035 17.475 33.080 ;
        RECT 18.025 33.220 18.315 33.265 ;
        RECT 19.850 33.220 20.170 33.280 ;
        RECT 24.540 33.220 24.680 33.760 ;
        RECT 26.305 33.715 26.595 33.760 ;
        RECT 27.210 33.700 27.530 33.960 ;
        RECT 27.685 33.900 27.975 33.945 ;
        RECT 28.130 33.900 28.450 33.960 ;
        RECT 27.685 33.760 28.450 33.900 ;
        RECT 27.685 33.715 27.975 33.760 ;
        RECT 28.130 33.700 28.450 33.760 ;
        RECT 34.570 33.900 34.890 33.960 ;
        RECT 39.185 33.900 39.475 33.945 ;
        RECT 34.570 33.760 39.475 33.900 ;
        RECT 34.570 33.700 34.890 33.760 ;
        RECT 39.185 33.715 39.475 33.760 ;
        RECT 40.090 33.700 40.410 33.960 ;
        RECT 49.305 33.715 49.595 33.945 ;
        RECT 26.750 33.360 27.070 33.620 ;
        RECT 29.020 33.560 29.310 33.605 ;
        RECT 29.510 33.560 29.830 33.620 ;
        RECT 29.020 33.420 29.830 33.560 ;
        RECT 29.020 33.375 29.310 33.420 ;
        RECT 29.510 33.360 29.830 33.420 ;
        RECT 35.490 33.605 35.810 33.620 ;
        RECT 35.490 33.375 36.095 33.605 ;
        RECT 36.885 33.560 37.175 33.605 ;
        RECT 39.645 33.560 39.935 33.605 ;
        RECT 36.885 33.420 39.935 33.560 ;
        RECT 49.380 33.560 49.520 33.715 ;
        RECT 53.430 33.700 53.750 33.960 ;
        RECT 53.890 33.900 54.210 33.960 ;
        RECT 54.825 33.900 55.115 33.945 ;
        RECT 53.890 33.760 55.115 33.900 ;
        RECT 53.890 33.700 54.210 33.760 ;
        RECT 54.825 33.715 55.115 33.760 ;
        RECT 63.090 33.900 63.410 33.960 ;
        RECT 64.485 33.900 64.775 33.945 ;
        RECT 63.090 33.760 64.775 33.900 ;
        RECT 63.090 33.700 63.410 33.760 ;
        RECT 64.485 33.715 64.775 33.760 ;
        RECT 66.310 33.700 66.630 33.960 ;
        RECT 66.770 33.700 67.090 33.960 ;
        RECT 67.245 33.900 67.535 33.945 ;
        RECT 67.690 33.900 68.010 33.960 ;
        RECT 67.245 33.760 68.010 33.900 ;
        RECT 67.245 33.715 67.535 33.760 ;
        RECT 67.690 33.700 68.010 33.760 ;
        RECT 68.165 33.900 68.455 33.945 ;
        RECT 68.610 33.900 68.930 33.960 ;
        RECT 68.165 33.760 68.930 33.900 ;
        RECT 68.165 33.715 68.455 33.760 ;
        RECT 68.610 33.700 68.930 33.760 ;
        RECT 69.990 33.900 70.310 33.960 ;
        RECT 70.465 33.900 70.755 33.945 ;
        RECT 69.990 33.760 70.755 33.900 ;
        RECT 69.990 33.700 70.310 33.760 ;
        RECT 70.465 33.715 70.755 33.760 ;
        RECT 70.910 33.900 71.230 33.960 ;
        RECT 71.385 33.900 71.675 33.945 ;
        RECT 70.910 33.760 71.675 33.900 ;
        RECT 70.910 33.700 71.230 33.760 ;
        RECT 71.385 33.715 71.675 33.760 ;
        RECT 72.305 33.900 72.595 33.945 ;
        RECT 73.210 33.900 73.530 33.960 ;
        RECT 72.305 33.760 73.530 33.900 ;
        RECT 72.305 33.715 72.595 33.760 ;
        RECT 73.210 33.700 73.530 33.760 ;
        RECT 55.285 33.560 55.575 33.605 ;
        RECT 55.730 33.560 56.050 33.620 ;
        RECT 49.380 33.420 56.050 33.560 ;
        RECT 36.885 33.375 37.175 33.420 ;
        RECT 39.645 33.375 39.935 33.420 ;
        RECT 55.285 33.375 55.575 33.420 ;
        RECT 35.490 33.360 35.810 33.375 ;
        RECT 55.730 33.360 56.050 33.420 ;
        RECT 59.885 33.560 60.175 33.605 ;
        RECT 64.930 33.560 65.250 33.620 ;
        RECT 59.885 33.420 65.250 33.560 ;
        RECT 59.885 33.375 60.175 33.420 ;
        RECT 64.930 33.360 65.250 33.420 ;
        RECT 71.830 33.560 72.150 33.620 ;
        RECT 72.750 33.560 73.070 33.620 ;
        RECT 71.830 33.420 73.070 33.560 ;
        RECT 71.830 33.360 72.150 33.420 ;
        RECT 72.750 33.360 73.070 33.420 ;
        RECT 75.940 33.560 76.230 33.605 ;
        RECT 77.810 33.560 78.130 33.620 ;
        RECT 75.940 33.420 78.130 33.560 ;
        RECT 75.940 33.375 76.230 33.420 ;
        RECT 77.810 33.360 78.130 33.420 ;
        RECT 18.025 33.080 24.680 33.220 ;
        RECT 49.765 33.220 50.055 33.265 ;
        RECT 50.210 33.220 50.530 33.280 ;
        RECT 49.765 33.080 50.530 33.220 ;
        RECT 18.025 33.035 18.315 33.080 ;
        RECT 19.850 33.020 20.170 33.080 ;
        RECT 49.765 33.035 50.055 33.080 ;
        RECT 50.210 33.020 50.530 33.080 ;
        RECT 59.410 33.020 59.730 33.280 ;
        RECT 63.565 33.220 63.855 33.265 ;
        RECT 65.850 33.220 66.170 33.280 ;
        RECT 63.565 33.080 66.170 33.220 ;
        RECT 63.565 33.035 63.855 33.080 ;
        RECT 65.850 33.020 66.170 33.080 ;
        RECT 68.150 33.220 68.470 33.280 ;
        RECT 72.290 33.220 72.610 33.280 ;
        RECT 79.650 33.220 79.970 33.280 ;
        RECT 68.150 33.080 79.970 33.220 ;
        RECT 68.150 33.020 68.470 33.080 ;
        RECT 72.290 33.020 72.610 33.080 ;
        RECT 79.650 33.020 79.970 33.080 ;
        RECT 81.030 33.220 81.350 33.280 ;
        RECT 81.505 33.220 81.795 33.265 ;
        RECT 81.030 33.080 81.795 33.220 ;
        RECT 81.030 33.020 81.350 33.080 ;
        RECT 81.505 33.035 81.795 33.080 ;
        RECT 5.520 32.400 83.260 32.880 ;
        RECT 19.390 32.200 19.710 32.260 ;
        RECT 15.420 32.060 19.710 32.200 ;
        RECT 13.885 31.520 14.175 31.565 ;
        RECT 15.420 31.520 15.560 32.060 ;
        RECT 19.390 32.000 19.710 32.060 ;
        RECT 27.670 32.200 27.990 32.260 ;
        RECT 31.825 32.200 32.115 32.245 ;
        RECT 27.670 32.060 32.115 32.200 ;
        RECT 27.670 32.000 27.990 32.060 ;
        RECT 31.825 32.015 32.115 32.060 ;
        RECT 33.665 32.200 33.955 32.245 ;
        RECT 34.570 32.200 34.890 32.260 ;
        RECT 33.665 32.060 34.890 32.200 ;
        RECT 33.665 32.015 33.955 32.060 ;
        RECT 15.710 31.860 16.030 31.920 ;
        RECT 17.410 31.860 17.700 31.905 ;
        RECT 24.305 31.860 24.595 31.905 ;
        RECT 15.710 31.720 17.700 31.860 ;
        RECT 15.710 31.660 16.030 31.720 ;
        RECT 17.410 31.675 17.700 31.720 ;
        RECT 18.100 31.720 24.595 31.860 ;
        RECT 13.885 31.380 15.560 31.520 ;
        RECT 13.885 31.335 14.175 31.380 ;
        RECT 16.170 31.320 16.490 31.580 ;
        RECT 18.100 31.520 18.240 31.720 ;
        RECT 24.305 31.675 24.595 31.720 ;
        RECT 25.385 31.675 25.675 31.905 ;
        RECT 29.525 31.860 29.815 31.905 ;
        RECT 33.740 31.860 33.880 32.015 ;
        RECT 34.570 32.000 34.890 32.060 ;
        RECT 44.230 32.200 44.550 32.260 ;
        RECT 47.465 32.200 47.755 32.245 ;
        RECT 44.230 32.060 47.755 32.200 ;
        RECT 44.230 32.000 44.550 32.060 ;
        RECT 47.465 32.015 47.755 32.060 ;
        RECT 51.605 32.200 51.895 32.245 ;
        RECT 54.810 32.200 55.130 32.260 ;
        RECT 51.605 32.060 55.130 32.200 ;
        RECT 51.605 32.015 51.895 32.060 ;
        RECT 54.810 32.000 55.130 32.060 ;
        RECT 55.745 32.200 56.035 32.245 ;
        RECT 56.190 32.200 56.510 32.260 ;
        RECT 55.745 32.060 56.510 32.200 ;
        RECT 55.745 32.015 56.035 32.060 ;
        RECT 56.190 32.000 56.510 32.060 ;
        RECT 56.665 32.200 56.955 32.245 ;
        RECT 59.870 32.200 60.190 32.260 ;
        RECT 56.665 32.060 60.190 32.200 ;
        RECT 56.665 32.015 56.955 32.060 ;
        RECT 59.870 32.000 60.190 32.060 ;
        RECT 60.345 32.200 60.635 32.245 ;
        RECT 65.390 32.200 65.710 32.260 ;
        RECT 60.345 32.060 65.710 32.200 ;
        RECT 60.345 32.015 60.635 32.060 ;
        RECT 65.390 32.000 65.710 32.060 ;
        RECT 67.690 32.000 68.010 32.260 ;
        RECT 70.465 32.200 70.755 32.245 ;
        RECT 71.370 32.200 71.690 32.260 ;
        RECT 70.465 32.060 71.690 32.200 ;
        RECT 70.465 32.015 70.755 32.060 ;
        RECT 71.370 32.000 71.690 32.060 ;
        RECT 73.685 32.200 73.975 32.245 ;
        RECT 75.970 32.200 76.290 32.260 ;
        RECT 73.685 32.060 76.290 32.200 ;
        RECT 73.685 32.015 73.975 32.060 ;
        RECT 75.970 32.000 76.290 32.060 ;
        RECT 77.810 32.000 78.130 32.260 ;
        RECT 78.270 32.000 78.590 32.260 ;
        RECT 80.110 32.200 80.430 32.260 ;
        RECT 79.740 32.060 80.430 32.200 ;
        RECT 29.525 31.720 33.880 31.860 ;
        RECT 52.445 31.860 52.735 31.905 ;
        RECT 52.445 31.720 53.200 31.860 ;
        RECT 29.525 31.675 29.815 31.720 ;
        RECT 52.445 31.675 52.735 31.720 ;
        RECT 16.720 31.380 18.240 31.520 ;
        RECT 20.310 31.520 20.630 31.580 ;
        RECT 25.460 31.520 25.600 31.675 ;
        RECT 20.310 31.380 25.600 31.520 ;
        RECT 32.745 31.520 33.035 31.565 ;
        RECT 33.650 31.520 33.970 31.580 ;
        RECT 32.745 31.380 33.970 31.520 ;
        RECT 14.330 30.980 14.650 31.240 ;
        RECT 15.725 31.180 16.015 31.225 ;
        RECT 16.720 31.180 16.860 31.380 ;
        RECT 20.310 31.320 20.630 31.380 ;
        RECT 32.745 31.335 33.035 31.380 ;
        RECT 33.650 31.320 33.970 31.380 ;
        RECT 34.125 31.335 34.415 31.565 ;
        RECT 47.465 31.335 47.755 31.565 ;
        RECT 15.725 31.040 16.860 31.180 ;
        RECT 17.065 31.180 17.355 31.225 ;
        RECT 18.255 31.180 18.545 31.225 ;
        RECT 20.775 31.180 21.065 31.225 ;
        RECT 17.065 31.040 21.065 31.180 ;
        RECT 15.725 30.995 16.015 31.040 ;
        RECT 17.065 30.995 17.355 31.040 ;
        RECT 18.255 30.995 18.545 31.040 ;
        RECT 20.775 30.995 21.065 31.040 ;
        RECT 33.190 31.180 33.510 31.240 ;
        RECT 34.200 31.180 34.340 31.335 ;
        RECT 33.190 31.040 34.340 31.180 ;
        RECT 47.540 31.180 47.680 31.335 ;
        RECT 48.370 31.320 48.690 31.580 ;
        RECT 48.830 31.320 49.150 31.580 ;
        RECT 49.305 31.520 49.595 31.565 ;
        RECT 49.750 31.520 50.070 31.580 ;
        RECT 49.305 31.380 50.070 31.520 ;
        RECT 49.305 31.335 49.595 31.380 ;
        RECT 49.750 31.320 50.070 31.380 ;
        RECT 48.920 31.180 49.060 31.320 ;
        RECT 47.540 31.040 49.060 31.180 ;
        RECT 33.190 30.980 33.510 31.040 ;
        RECT 50.210 30.980 50.530 31.240 ;
        RECT 53.060 31.180 53.200 31.720 ;
        RECT 53.445 31.675 53.735 31.905 ;
        RECT 64.470 31.860 64.790 31.920 ;
        RECT 62.030 31.720 64.790 31.860 ;
        RECT 53.520 31.520 53.660 31.675 ;
        RECT 53.905 31.520 54.195 31.565 ;
        RECT 55.730 31.520 56.050 31.580 ;
        RECT 57.585 31.520 57.875 31.565 ;
        RECT 62.030 31.520 62.170 31.720 ;
        RECT 64.470 31.660 64.790 31.720 ;
        RECT 65.020 31.720 71.600 31.860 ;
        RECT 65.020 31.565 65.160 31.720 ;
        RECT 53.520 31.380 62.170 31.520 ;
        RECT 63.105 31.520 63.395 31.565 ;
        RECT 63.105 31.380 64.700 31.520 ;
        RECT 53.905 31.335 54.195 31.380 ;
        RECT 55.730 31.320 56.050 31.380 ;
        RECT 57.585 31.335 57.875 31.380 ;
        RECT 63.105 31.335 63.395 31.380 ;
        RECT 55.270 31.180 55.590 31.240 ;
        RECT 56.190 31.180 56.510 31.240 ;
        RECT 53.060 31.040 56.510 31.180 ;
        RECT 55.270 30.980 55.590 31.040 ;
        RECT 56.190 30.980 56.510 31.040 ;
        RECT 58.965 30.995 59.255 31.225 ;
        RECT 64.560 31.180 64.700 31.380 ;
        RECT 64.945 31.335 65.235 31.565 ;
        RECT 66.325 31.335 66.615 31.565 ;
        RECT 67.245 31.520 67.535 31.565 ;
        RECT 67.690 31.520 68.010 31.580 ;
        RECT 67.245 31.380 68.010 31.520 ;
        RECT 67.245 31.335 67.535 31.380 ;
        RECT 66.400 31.180 66.540 31.335 ;
        RECT 67.690 31.320 68.010 31.380 ;
        RECT 68.625 31.335 68.915 31.565 ;
        RECT 68.150 31.180 68.470 31.240 ;
        RECT 64.560 31.040 68.470 31.180 ;
        RECT 68.700 31.180 68.840 31.335 ;
        RECT 69.530 31.320 69.850 31.580 ;
        RECT 71.460 31.565 71.600 31.720 ;
        RECT 72.290 31.660 72.610 31.920 ;
        RECT 73.210 31.860 73.530 31.920 ;
        RECT 79.740 31.905 79.880 32.060 ;
        RECT 80.110 32.000 80.430 32.060 ;
        RECT 73.210 31.720 79.420 31.860 ;
        RECT 73.210 31.660 73.530 31.720 ;
        RECT 71.385 31.520 71.675 31.565 ;
        RECT 71.830 31.520 72.150 31.580 ;
        RECT 71.385 31.380 72.150 31.520 ;
        RECT 71.385 31.335 71.675 31.380 ;
        RECT 71.830 31.320 72.150 31.380 ;
        RECT 72.750 31.320 73.070 31.580 ;
        RECT 74.605 31.550 74.895 31.565 ;
        RECT 75.050 31.550 75.370 31.570 ;
        RECT 74.605 31.410 75.370 31.550 ;
        RECT 74.605 31.335 74.895 31.410 ;
        RECT 75.050 31.310 75.370 31.410 ;
        RECT 75.525 31.350 75.815 31.580 ;
        RECT 76.015 31.565 76.335 31.580 ;
        RECT 76.000 31.520 76.335 31.565 ;
        RECT 76.675 31.520 76.965 31.565 ;
        RECT 78.730 31.520 79.050 31.580 ;
        RECT 79.280 31.565 79.420 31.720 ;
        RECT 79.665 31.675 79.955 31.905 ;
        RECT 76.000 31.380 76.500 31.520 ;
        RECT 76.675 31.380 79.050 31.520 ;
        RECT 69.990 31.180 70.310 31.240 ;
        RECT 68.700 31.040 70.310 31.180 ;
        RECT 16.670 30.840 16.960 30.885 ;
        RECT 18.770 30.840 19.060 30.885 ;
        RECT 20.340 30.840 20.630 30.885 ;
        RECT 16.670 30.700 20.630 30.840 ;
        RECT 16.670 30.655 16.960 30.700 ;
        RECT 18.770 30.655 19.060 30.700 ;
        RECT 20.340 30.655 20.630 30.700 ;
        RECT 28.145 30.840 28.435 30.885 ;
        RECT 30.890 30.840 31.210 30.900 ;
        RECT 59.040 30.840 59.180 30.995 ;
        RECT 68.150 30.980 68.470 31.040 ;
        RECT 69.990 30.980 70.310 31.040 ;
        RECT 70.450 31.180 70.770 31.240 ;
        RECT 70.450 31.140 73.900 31.180 ;
        RECT 75.600 31.140 75.740 31.350 ;
        RECT 76.000 31.335 76.335 31.380 ;
        RECT 76.675 31.335 76.965 31.380 ;
        RECT 76.015 31.320 76.335 31.335 ;
        RECT 78.730 31.320 79.050 31.380 ;
        RECT 79.205 31.335 79.495 31.565 ;
        RECT 80.110 31.320 80.430 31.580 ;
        RECT 81.030 31.320 81.350 31.580 ;
        RECT 70.450 31.040 75.740 31.140 ;
        RECT 70.450 30.980 70.770 31.040 ;
        RECT 73.760 31.000 75.740 31.040 ;
        RECT 28.145 30.700 31.210 30.840 ;
        RECT 28.145 30.655 28.435 30.700 ;
        RECT 30.890 30.640 31.210 30.700 ;
        RECT 55.820 30.700 59.180 30.840 ;
        RECT 17.090 30.500 17.410 30.560 ;
        RECT 23.085 30.500 23.375 30.545 ;
        RECT 17.090 30.360 23.375 30.500 ;
        RECT 17.090 30.300 17.410 30.360 ;
        RECT 23.085 30.315 23.375 30.360 ;
        RECT 23.530 30.300 23.850 30.560 ;
        RECT 23.990 30.500 24.310 30.560 ;
        RECT 24.465 30.500 24.755 30.545 ;
        RECT 23.990 30.360 24.755 30.500 ;
        RECT 23.990 30.300 24.310 30.360 ;
        RECT 24.465 30.315 24.755 30.360 ;
        RECT 27.210 30.300 27.530 30.560 ;
        RECT 49.750 30.300 50.070 30.560 ;
        RECT 52.525 30.500 52.815 30.545 ;
        RECT 54.350 30.500 54.670 30.560 ;
        RECT 55.820 30.545 55.960 30.700 ;
        RECT 55.745 30.500 56.035 30.545 ;
        RECT 52.525 30.360 56.035 30.500 ;
        RECT 52.525 30.315 52.815 30.360 ;
        RECT 54.350 30.300 54.670 30.360 ;
        RECT 55.745 30.315 56.035 30.360 ;
        RECT 58.490 30.300 58.810 30.560 ;
        RECT 59.040 30.500 59.180 30.700 ;
        RECT 62.185 30.840 62.475 30.885 ;
        RECT 75.970 30.840 76.290 30.900 ;
        RECT 62.185 30.700 76.290 30.840 ;
        RECT 62.185 30.655 62.475 30.700 ;
        RECT 75.970 30.640 76.290 30.700 ;
        RECT 63.550 30.500 63.870 30.560 ;
        RECT 59.040 30.360 63.870 30.500 ;
        RECT 63.550 30.300 63.870 30.360 ;
        RECT 64.010 30.300 64.330 30.560 ;
        RECT 65.405 30.500 65.695 30.545 ;
        RECT 68.610 30.500 68.930 30.560 ;
        RECT 65.405 30.360 68.930 30.500 ;
        RECT 65.405 30.315 65.695 30.360 ;
        RECT 68.610 30.300 68.930 30.360 ;
        RECT 69.070 30.500 69.390 30.560 ;
        RECT 75.050 30.500 75.370 30.560 ;
        RECT 69.070 30.360 75.370 30.500 ;
        RECT 69.070 30.300 69.390 30.360 ;
        RECT 75.050 30.300 75.370 30.360 ;
        RECT 5.520 29.680 83.260 30.160 ;
        RECT 18.945 29.480 19.235 29.525 ;
        RECT 19.390 29.480 19.710 29.540 ;
        RECT 18.945 29.340 19.710 29.480 ;
        RECT 18.945 29.295 19.235 29.340 ;
        RECT 19.390 29.280 19.710 29.340 ;
        RECT 33.205 29.480 33.495 29.525 ;
        RECT 34.570 29.480 34.890 29.540 ;
        RECT 33.205 29.340 34.890 29.480 ;
        RECT 33.205 29.295 33.495 29.340 ;
        RECT 34.570 29.280 34.890 29.340 ;
        RECT 52.970 29.280 53.290 29.540 ;
        RECT 59.885 29.480 60.175 29.525 ;
        RECT 60.330 29.480 60.650 29.540 ;
        RECT 59.885 29.340 60.650 29.480 ;
        RECT 59.885 29.295 60.175 29.340 ;
        RECT 60.330 29.280 60.650 29.340 ;
        RECT 63.105 29.480 63.395 29.525 ;
        RECT 70.450 29.480 70.770 29.540 ;
        RECT 80.110 29.480 80.430 29.540 ;
        RECT 63.105 29.340 70.770 29.480 ;
        RECT 63.105 29.295 63.395 29.340 ;
        RECT 70.450 29.280 70.770 29.340 ;
        RECT 75.600 29.340 80.430 29.480 ;
        RECT 13.410 29.140 13.730 29.200 ;
        RECT 20.310 29.140 20.630 29.200 ;
        RECT 13.410 29.000 20.630 29.140 ;
        RECT 13.410 28.940 13.730 29.000 ;
        RECT 20.310 28.940 20.630 29.000 ;
        RECT 21.690 29.140 21.980 29.185 ;
        RECT 23.260 29.140 23.550 29.185 ;
        RECT 25.360 29.140 25.650 29.185 ;
        RECT 21.690 29.000 25.650 29.140 ;
        RECT 21.690 28.955 21.980 29.000 ;
        RECT 23.260 28.955 23.550 29.000 ;
        RECT 25.360 28.955 25.650 29.000 ;
        RECT 26.790 29.140 27.080 29.185 ;
        RECT 28.890 29.140 29.180 29.185 ;
        RECT 30.460 29.140 30.750 29.185 ;
        RECT 26.790 29.000 30.750 29.140 ;
        RECT 26.790 28.955 27.080 29.000 ;
        RECT 28.890 28.955 29.180 29.000 ;
        RECT 30.460 28.955 30.750 29.000 ;
        RECT 70.910 28.940 71.230 29.200 ;
        RECT 73.670 28.940 73.990 29.200 ;
        RECT 21.255 28.800 21.545 28.845 ;
        RECT 23.775 28.800 24.065 28.845 ;
        RECT 24.965 28.800 25.255 28.845 ;
        RECT 21.255 28.660 25.255 28.800 ;
        RECT 21.255 28.615 21.545 28.660 ;
        RECT 23.775 28.615 24.065 28.660 ;
        RECT 24.965 28.615 25.255 28.660 ;
        RECT 27.185 28.800 27.475 28.845 ;
        RECT 28.375 28.800 28.665 28.845 ;
        RECT 30.895 28.800 31.185 28.845 ;
        RECT 69.530 28.800 69.850 28.860 ;
        RECT 27.185 28.660 31.185 28.800 ;
        RECT 27.185 28.615 27.475 28.660 ;
        RECT 28.375 28.615 28.665 28.660 ;
        RECT 30.895 28.615 31.185 28.660 ;
        RECT 53.520 28.660 56.880 28.800 ;
        RECT 25.845 28.460 26.135 28.505 ;
        RECT 26.305 28.460 26.595 28.505 ;
        RECT 25.845 28.320 26.980 28.460 ;
        RECT 25.845 28.275 26.135 28.320 ;
        RECT 26.305 28.275 26.595 28.320 ;
        RECT 23.530 28.120 23.850 28.180 ;
        RECT 24.510 28.120 24.800 28.165 ;
        RECT 23.530 27.980 24.800 28.120 ;
        RECT 23.530 27.920 23.850 27.980 ;
        RECT 24.510 27.935 24.800 27.980 ;
        RECT 26.840 27.780 26.980 28.320 ;
        RECT 27.640 28.275 27.930 28.505 ;
        RECT 49.750 28.460 50.070 28.520 ;
        RECT 53.520 28.505 53.660 28.660 ;
        RECT 52.525 28.460 52.815 28.505 ;
        RECT 49.750 28.320 52.815 28.460 ;
        RECT 27.210 28.120 27.530 28.180 ;
        RECT 27.760 28.120 27.900 28.275 ;
        RECT 49.750 28.260 50.070 28.320 ;
        RECT 52.525 28.275 52.815 28.320 ;
        RECT 53.445 28.275 53.735 28.505 ;
        RECT 53.890 28.260 54.210 28.520 ;
        RECT 54.350 28.460 54.670 28.520 ;
        RECT 56.740 28.505 56.880 28.660 ;
        RECT 65.480 28.660 69.850 28.800 ;
        RECT 71.000 28.800 71.140 28.940 ;
        RECT 75.600 28.800 75.740 29.340 ;
        RECT 80.110 29.280 80.430 29.340 ;
        RECT 76.430 28.940 76.750 29.200 ;
        RECT 71.000 28.660 75.740 28.800 ;
        RECT 76.520 28.800 76.660 28.940 ;
        RECT 76.520 28.660 79.420 28.800 ;
        RECT 54.825 28.460 55.115 28.505 ;
        RECT 54.350 28.320 55.115 28.460 ;
        RECT 54.350 28.260 54.670 28.320 ;
        RECT 54.825 28.275 55.115 28.320 ;
        RECT 56.665 28.460 56.955 28.505 ;
        RECT 58.490 28.460 58.810 28.520 ;
        RECT 56.665 28.320 58.810 28.460 ;
        RECT 56.665 28.275 56.955 28.320 ;
        RECT 58.490 28.260 58.810 28.320 ;
        RECT 60.805 28.460 61.095 28.505 ;
        RECT 61.250 28.460 61.570 28.520 ;
        RECT 60.805 28.320 61.570 28.460 ;
        RECT 60.805 28.275 61.095 28.320 ;
        RECT 61.250 28.260 61.570 28.320 ;
        RECT 62.645 28.460 62.935 28.505 ;
        RECT 64.010 28.460 64.330 28.520 ;
        RECT 62.645 28.320 64.330 28.460 ;
        RECT 62.645 28.275 62.935 28.320 ;
        RECT 64.010 28.260 64.330 28.320 ;
        RECT 65.480 28.180 65.620 28.660 ;
        RECT 69.530 28.600 69.850 28.660 ;
        RECT 66.325 28.460 66.615 28.505 ;
        RECT 70.465 28.460 70.755 28.505 ;
        RECT 70.910 28.460 71.230 28.520 ;
        RECT 71.460 28.505 71.600 28.660 ;
        RECT 66.325 28.320 71.230 28.460 ;
        RECT 66.325 28.275 66.615 28.320 ;
        RECT 70.465 28.275 70.755 28.320 ;
        RECT 70.910 28.260 71.230 28.320 ;
        RECT 71.385 28.275 71.675 28.505 ;
        RECT 71.845 28.275 72.135 28.505 ;
        RECT 72.305 28.460 72.595 28.505 ;
        RECT 73.210 28.460 73.530 28.520 ;
        RECT 75.600 28.505 75.740 28.660 ;
        RECT 79.280 28.520 79.420 28.660 ;
        RECT 74.605 28.460 74.895 28.505 ;
        RECT 72.305 28.320 74.895 28.460 ;
        RECT 72.305 28.275 72.595 28.320 ;
        RECT 27.210 27.980 27.900 28.120 ;
        RECT 64.945 28.120 65.235 28.165 ;
        RECT 65.390 28.120 65.710 28.180 ;
        RECT 64.945 27.980 65.710 28.120 ;
        RECT 27.210 27.920 27.530 27.980 ;
        RECT 64.945 27.935 65.235 27.980 ;
        RECT 65.390 27.920 65.710 27.980 ;
        RECT 67.690 27.920 68.010 28.180 ;
        RECT 68.625 27.935 68.915 28.165 ;
        RECT 69.070 28.120 69.390 28.180 ;
        RECT 69.545 28.120 69.835 28.165 ;
        RECT 69.070 27.980 69.835 28.120 ;
        RECT 71.920 28.120 72.060 28.275 ;
        RECT 73.210 28.260 73.530 28.320 ;
        RECT 74.605 28.275 74.895 28.320 ;
        RECT 75.525 28.275 75.815 28.505 ;
        RECT 76.445 28.275 76.735 28.505 ;
        RECT 78.270 28.460 78.590 28.520 ;
        RECT 78.745 28.460 79.035 28.505 ;
        RECT 78.270 28.320 79.035 28.460 ;
        RECT 72.750 28.120 73.070 28.180 ;
        RECT 73.670 28.120 73.990 28.180 ;
        RECT 71.920 27.980 73.070 28.120 ;
        RECT 27.670 27.780 27.990 27.840 ;
        RECT 26.840 27.640 27.990 27.780 ;
        RECT 27.670 27.580 27.990 27.640 ;
        RECT 54.365 27.780 54.655 27.825 ;
        RECT 54.810 27.780 55.130 27.840 ;
        RECT 54.365 27.640 55.130 27.780 ;
        RECT 54.365 27.595 54.655 27.640 ;
        RECT 54.810 27.580 55.130 27.640 ;
        RECT 57.125 27.780 57.415 27.825 ;
        RECT 57.570 27.780 57.890 27.840 ;
        RECT 57.125 27.640 57.890 27.780 ;
        RECT 57.125 27.595 57.415 27.640 ;
        RECT 57.570 27.580 57.890 27.640 ;
        RECT 61.710 27.580 62.030 27.840 ;
        RECT 67.245 27.780 67.535 27.825 ;
        RECT 68.150 27.780 68.470 27.840 ;
        RECT 67.245 27.640 68.470 27.780 ;
        RECT 68.700 27.780 68.840 27.935 ;
        RECT 69.070 27.920 69.390 27.980 ;
        RECT 69.545 27.935 69.835 27.980 ;
        RECT 70.910 27.780 71.230 27.840 ;
        RECT 68.700 27.640 71.230 27.780 ;
        RECT 67.245 27.595 67.535 27.640 ;
        RECT 68.150 27.580 68.470 27.640 ;
        RECT 70.910 27.580 71.230 27.640 ;
        RECT 71.830 27.780 72.150 27.840 ;
        RECT 72.380 27.780 72.520 27.980 ;
        RECT 72.750 27.920 73.070 27.980 ;
        RECT 73.300 27.980 73.990 28.120 ;
        RECT 73.300 27.825 73.440 27.980 ;
        RECT 73.670 27.920 73.990 27.980 ;
        RECT 75.050 27.920 75.370 28.180 ;
        RECT 76.520 28.120 76.660 28.275 ;
        RECT 78.270 28.260 78.590 28.320 ;
        RECT 78.745 28.275 79.035 28.320 ;
        RECT 79.190 28.260 79.510 28.520 ;
        RECT 79.650 28.260 79.970 28.520 ;
        RECT 80.570 28.260 80.890 28.520 ;
        RECT 75.600 27.980 76.660 28.120 ;
        RECT 71.830 27.640 72.520 27.780 ;
        RECT 71.830 27.580 72.150 27.640 ;
        RECT 73.225 27.595 73.515 27.825 ;
        RECT 74.130 27.780 74.450 27.840 ;
        RECT 75.600 27.780 75.740 27.980 ;
        RECT 74.130 27.640 75.740 27.780 ;
        RECT 76.430 27.780 76.750 27.840 ;
        RECT 77.365 27.780 77.655 27.825 ;
        RECT 76.430 27.640 77.655 27.780 ;
        RECT 74.130 27.580 74.450 27.640 ;
        RECT 76.430 27.580 76.750 27.640 ;
        RECT 77.365 27.595 77.655 27.640 ;
        RECT 5.520 26.960 83.260 27.440 ;
        RECT 46.990 26.760 47.310 26.820 ;
        RECT 50.225 26.760 50.515 26.805 ;
        RECT 53.890 26.760 54.210 26.820 ;
        RECT 46.990 26.620 54.210 26.760 ;
        RECT 46.990 26.560 47.310 26.620 ;
        RECT 50.225 26.575 50.515 26.620 ;
        RECT 53.890 26.560 54.210 26.620 ;
        RECT 59.870 26.760 60.190 26.820 ;
        RECT 63.550 26.760 63.870 26.820 ;
        RECT 59.870 26.620 63.870 26.760 ;
        RECT 59.870 26.560 60.190 26.620 ;
        RECT 63.550 26.560 63.870 26.620 ;
        RECT 64.025 26.760 64.315 26.805 ;
        RECT 70.005 26.760 70.295 26.805 ;
        RECT 64.025 26.620 70.295 26.760 ;
        RECT 64.025 26.575 64.315 26.620 ;
        RECT 70.005 26.575 70.295 26.620 ;
        RECT 76.890 26.760 77.210 26.820 ;
        RECT 76.890 26.620 80.340 26.760 ;
        RECT 76.890 26.560 77.210 26.620 ;
        RECT 46.070 26.420 46.390 26.480 ;
        RECT 47.450 26.420 47.770 26.480 ;
        RECT 52.985 26.420 53.275 26.465 ;
        RECT 55.270 26.420 55.590 26.480 ;
        RECT 46.070 26.280 47.770 26.420 ;
        RECT 46.070 26.220 46.390 26.280 ;
        RECT 47.450 26.220 47.770 26.280 ;
        RECT 50.760 26.280 55.590 26.420 ;
        RECT 63.640 26.420 63.780 26.560 ;
        RECT 66.770 26.420 67.090 26.480 ;
        RECT 69.070 26.420 69.390 26.480 ;
        RECT 63.640 26.280 65.620 26.420 ;
        RECT 50.760 26.125 50.900 26.280 ;
        RECT 52.985 26.235 53.275 26.280 ;
        RECT 55.270 26.220 55.590 26.280 ;
        RECT 49.765 25.895 50.055 26.125 ;
        RECT 50.685 25.895 50.975 26.125 ;
        RECT 52.065 25.895 52.355 26.125 ;
        RECT 53.905 26.080 54.195 26.125 ;
        RECT 54.350 26.080 54.670 26.140 ;
        RECT 53.905 25.940 54.670 26.080 ;
        RECT 53.905 25.895 54.195 25.940 ;
        RECT 49.840 25.740 49.980 25.895 ;
        RECT 52.140 25.740 52.280 25.895 ;
        RECT 54.350 25.880 54.670 25.940 ;
        RECT 55.745 26.080 56.035 26.125 ;
        RECT 58.490 26.080 58.810 26.140 ;
        RECT 55.745 25.940 58.810 26.080 ;
        RECT 55.745 25.895 56.035 25.940 ;
        RECT 58.490 25.880 58.810 25.940 ;
        RECT 64.470 25.880 64.790 26.140 ;
        RECT 65.480 26.080 65.620 26.280 ;
        RECT 66.770 26.280 68.380 26.420 ;
        RECT 66.770 26.220 67.090 26.280 ;
        RECT 68.240 26.125 68.380 26.280 ;
        RECT 69.070 26.280 79.880 26.420 ;
        RECT 69.070 26.220 69.390 26.280 ;
        RECT 67.705 26.080 67.995 26.125 ;
        RECT 65.480 25.940 67.995 26.080 ;
        RECT 67.705 25.895 67.995 25.940 ;
        RECT 68.165 25.895 68.455 26.125 ;
        RECT 68.625 26.080 68.915 26.125 ;
        RECT 68.625 25.940 69.300 26.080 ;
        RECT 68.625 25.895 68.915 25.940 ;
        RECT 49.840 25.600 55.960 25.740 ;
        RECT 47.450 25.400 47.770 25.460 ;
        RECT 51.145 25.400 51.435 25.445 ;
        RECT 47.450 25.260 51.435 25.400 ;
        RECT 47.450 25.200 47.770 25.260 ;
        RECT 51.145 25.215 51.435 25.260 ;
        RECT 55.820 25.120 55.960 25.600 ;
        RECT 60.330 25.540 60.650 25.800 ;
        RECT 60.790 25.540 61.110 25.800 ;
        RECT 64.930 25.540 65.250 25.800 ;
        RECT 56.665 25.400 56.955 25.445 ;
        RECT 64.470 25.400 64.790 25.460 ;
        RECT 56.665 25.260 64.790 25.400 ;
        RECT 56.665 25.215 56.955 25.260 ;
        RECT 64.470 25.200 64.790 25.260 ;
        RECT 55.730 24.860 56.050 25.120 ;
        RECT 58.045 25.060 58.335 25.105 ;
        RECT 58.490 25.060 58.810 25.120 ;
        RECT 58.045 24.920 58.810 25.060 ;
        RECT 58.045 24.875 58.335 24.920 ;
        RECT 58.490 24.860 58.810 24.920 ;
        RECT 62.170 24.860 62.490 25.120 ;
        RECT 66.325 25.060 66.615 25.105 ;
        RECT 66.770 25.060 67.090 25.120 ;
        RECT 66.325 24.920 67.090 25.060 ;
        RECT 67.780 25.060 67.920 25.895 ;
        RECT 68.150 25.400 68.470 25.460 ;
        RECT 69.160 25.400 69.300 25.940 ;
        RECT 69.530 25.880 69.850 26.140 ;
        RECT 71.830 26.080 72.150 26.140 ;
        RECT 75.065 26.080 75.355 26.125 ;
        RECT 71.830 25.940 75.355 26.080 ;
        RECT 71.830 25.880 72.150 25.940 ;
        RECT 75.065 25.895 75.355 25.940 ;
        RECT 75.510 25.880 75.830 26.140 ;
        RECT 75.970 25.880 76.290 26.140 ;
        RECT 76.890 25.880 77.210 26.140 ;
        RECT 79.740 26.125 79.880 26.280 ;
        RECT 78.745 25.895 79.035 26.125 ;
        RECT 79.205 25.895 79.495 26.125 ;
        RECT 79.665 25.895 79.955 26.125 ;
        RECT 80.200 26.080 80.340 26.620 ;
        RECT 80.570 26.080 80.890 26.140 ;
        RECT 80.200 25.940 80.890 26.080 ;
        RECT 70.910 25.740 71.230 25.800 ;
        RECT 72.765 25.740 73.055 25.785 ;
        RECT 70.910 25.600 73.055 25.740 ;
        RECT 70.910 25.540 71.230 25.600 ;
        RECT 72.765 25.555 73.055 25.600 ;
        RECT 73.210 25.740 73.530 25.800 ;
        RECT 78.820 25.740 78.960 25.895 ;
        RECT 73.210 25.600 78.960 25.740 ;
        RECT 73.210 25.540 73.530 25.600 ;
        RECT 68.150 25.260 69.300 25.400 ;
        RECT 69.530 25.400 69.850 25.460 ;
        RECT 75.510 25.400 75.830 25.460 ;
        RECT 79.280 25.400 79.420 25.895 ;
        RECT 80.570 25.880 80.890 25.940 ;
        RECT 69.530 25.260 75.280 25.400 ;
        RECT 68.150 25.200 68.470 25.260 ;
        RECT 69.530 25.200 69.850 25.260 ;
        RECT 71.830 25.060 72.150 25.120 ;
        RECT 67.780 24.920 72.150 25.060 ;
        RECT 66.325 24.875 66.615 24.920 ;
        RECT 66.770 24.860 67.090 24.920 ;
        RECT 71.830 24.860 72.150 24.920 ;
        RECT 73.670 24.860 73.990 25.120 ;
        RECT 75.140 25.060 75.280 25.260 ;
        RECT 75.510 25.260 79.420 25.400 ;
        RECT 75.510 25.200 75.830 25.260 ;
        RECT 76.890 25.060 77.210 25.120 ;
        RECT 75.140 24.920 77.210 25.060 ;
        RECT 76.890 24.860 77.210 24.920 ;
        RECT 77.350 24.860 77.670 25.120 ;
        RECT 5.520 24.240 83.260 24.720 ;
        RECT 44.690 24.040 45.010 24.100 ;
        RECT 45.165 24.040 45.455 24.085 ;
        RECT 44.690 23.900 45.455 24.040 ;
        RECT 44.690 23.840 45.010 23.900 ;
        RECT 45.165 23.855 45.455 23.900 ;
        RECT 55.730 23.840 56.050 24.100 ;
        RECT 63.550 24.040 63.870 24.100 ;
        RECT 64.025 24.040 64.315 24.085 ;
        RECT 63.550 23.900 64.315 24.040 ;
        RECT 63.550 23.840 63.870 23.900 ;
        RECT 64.025 23.855 64.315 23.900 ;
        RECT 70.465 24.040 70.755 24.085 ;
        RECT 71.370 24.040 71.690 24.100 ;
        RECT 70.465 23.900 71.690 24.040 ;
        RECT 70.465 23.855 70.755 23.900 ;
        RECT 71.370 23.840 71.690 23.900 ;
        RECT 49.330 23.700 49.620 23.745 ;
        RECT 51.430 23.700 51.720 23.745 ;
        RECT 53.000 23.700 53.290 23.745 ;
        RECT 49.330 23.560 53.290 23.700 ;
        RECT 49.330 23.515 49.620 23.560 ;
        RECT 51.430 23.515 51.720 23.560 ;
        RECT 53.000 23.515 53.290 23.560 ;
        RECT 57.610 23.700 57.900 23.745 ;
        RECT 59.710 23.700 60.000 23.745 ;
        RECT 61.280 23.700 61.570 23.745 ;
        RECT 57.610 23.560 61.570 23.700 ;
        RECT 57.610 23.515 57.900 23.560 ;
        RECT 59.710 23.515 60.000 23.560 ;
        RECT 61.280 23.515 61.570 23.560 ;
        RECT 73.210 23.700 73.500 23.745 ;
        RECT 74.780 23.700 75.070 23.745 ;
        RECT 76.880 23.700 77.170 23.745 ;
        RECT 73.210 23.560 77.170 23.700 ;
        RECT 73.210 23.515 73.500 23.560 ;
        RECT 74.780 23.515 75.070 23.560 ;
        RECT 76.880 23.515 77.170 23.560 ;
        RECT 79.190 23.500 79.510 23.760 ;
        RECT 45.610 23.360 45.930 23.420 ;
        RECT 46.085 23.360 46.375 23.405 ;
        RECT 45.610 23.220 46.375 23.360 ;
        RECT 45.610 23.160 45.930 23.220 ;
        RECT 46.085 23.175 46.375 23.220 ;
        RECT 49.725 23.360 50.015 23.405 ;
        RECT 50.915 23.360 51.205 23.405 ;
        RECT 53.435 23.360 53.725 23.405 ;
        RECT 49.725 23.220 53.725 23.360 ;
        RECT 49.725 23.175 50.015 23.220 ;
        RECT 50.915 23.175 51.205 23.220 ;
        RECT 53.435 23.175 53.725 23.220 ;
        RECT 58.005 23.360 58.295 23.405 ;
        RECT 59.195 23.360 59.485 23.405 ;
        RECT 61.715 23.360 62.005 23.405 ;
        RECT 58.005 23.220 62.005 23.360 ;
        RECT 58.005 23.175 58.295 23.220 ;
        RECT 59.195 23.175 59.485 23.220 ;
        RECT 61.715 23.175 62.005 23.220 ;
        RECT 64.470 23.360 64.790 23.420 ;
        RECT 67.705 23.360 67.995 23.405 ;
        RECT 64.470 23.220 67.995 23.360 ;
        RECT 64.470 23.160 64.790 23.220 ;
        RECT 67.705 23.175 67.995 23.220 ;
        RECT 72.775 23.360 73.065 23.405 ;
        RECT 75.295 23.360 75.585 23.405 ;
        RECT 76.485 23.360 76.775 23.405 ;
        RECT 72.775 23.220 76.775 23.360 ;
        RECT 79.280 23.360 79.420 23.500 ;
        RECT 79.280 23.220 79.880 23.360 ;
        RECT 72.775 23.175 73.065 23.220 ;
        RECT 75.295 23.175 75.585 23.220 ;
        RECT 76.485 23.175 76.775 23.220 ;
        RECT 44.230 23.020 44.550 23.080 ;
        RECT 44.705 23.020 44.995 23.065 ;
        RECT 46.530 23.020 46.850 23.080 ;
        RECT 44.230 22.880 46.850 23.020 ;
        RECT 44.230 22.820 44.550 22.880 ;
        RECT 44.705 22.835 44.995 22.880 ;
        RECT 46.530 22.820 46.850 22.880 ;
        RECT 46.990 22.820 47.310 23.080 ;
        RECT 47.450 22.820 47.770 23.080 ;
        RECT 48.845 23.020 49.135 23.065 ;
        RECT 49.290 23.020 49.610 23.080 ;
        RECT 48.845 22.880 49.610 23.020 ;
        RECT 48.845 22.835 49.135 22.880 ;
        RECT 49.290 22.820 49.610 22.880 ;
        RECT 57.110 22.820 57.430 23.080 ;
        RECT 58.490 23.065 58.810 23.080 ;
        RECT 58.460 23.020 58.810 23.065 ;
        RECT 67.245 23.020 67.535 23.065 ;
        RECT 71.830 23.020 72.150 23.080 ;
        RECT 73.210 23.020 73.530 23.080 ;
        RECT 58.295 22.880 58.810 23.020 ;
        RECT 58.460 22.835 58.810 22.880 ;
        RECT 58.490 22.820 58.810 22.835 ;
        RECT 59.040 22.880 73.530 23.020 ;
        RECT 48.385 22.680 48.675 22.725 ;
        RECT 50.070 22.680 50.360 22.725 ;
        RECT 48.385 22.540 50.360 22.680 ;
        RECT 48.385 22.495 48.675 22.540 ;
        RECT 50.070 22.495 50.360 22.540 ;
        RECT 58.030 22.680 58.350 22.740 ;
        RECT 59.040 22.680 59.180 22.880 ;
        RECT 67.245 22.835 67.535 22.880 ;
        RECT 71.830 22.820 72.150 22.880 ;
        RECT 73.210 22.820 73.530 22.880 ;
        RECT 74.590 23.020 74.910 23.080 ;
        RECT 79.740 23.065 79.880 23.220 ;
        RECT 77.365 23.020 77.655 23.065 ;
        RECT 74.590 22.880 77.655 23.020 ;
        RECT 74.590 22.820 74.910 22.880 ;
        RECT 77.365 22.835 77.655 22.880 ;
        RECT 79.205 22.835 79.495 23.065 ;
        RECT 79.665 22.835 79.955 23.065 ;
        RECT 66.785 22.680 67.075 22.725 ;
        RECT 58.030 22.540 59.180 22.680 ;
        RECT 62.030 22.540 67.075 22.680 ;
        RECT 58.030 22.480 58.350 22.540 ;
        RECT 46.085 22.340 46.375 22.385 ;
        RECT 47.910 22.340 48.230 22.400 ;
        RECT 46.085 22.200 48.230 22.340 ;
        RECT 46.085 22.155 46.375 22.200 ;
        RECT 47.910 22.140 48.230 22.200 ;
        RECT 53.890 22.340 54.210 22.400 ;
        RECT 60.330 22.340 60.650 22.400 ;
        RECT 62.030 22.340 62.170 22.540 ;
        RECT 66.785 22.495 67.075 22.540 ;
        RECT 73.670 22.680 73.990 22.740 ;
        RECT 76.030 22.680 76.320 22.725 ;
        RECT 73.670 22.540 76.320 22.680 ;
        RECT 79.280 22.680 79.420 22.835 ;
        RECT 80.110 22.820 80.430 23.080 ;
        RECT 80.570 23.020 80.890 23.080 ;
        RECT 81.045 23.020 81.335 23.065 ;
        RECT 80.570 22.880 81.335 23.020 ;
        RECT 80.570 22.820 80.890 22.880 ;
        RECT 81.045 22.835 81.335 22.880 ;
        RECT 81.490 22.680 81.810 22.740 ;
        RECT 79.280 22.540 81.810 22.680 ;
        RECT 73.670 22.480 73.990 22.540 ;
        RECT 76.030 22.495 76.320 22.540 ;
        RECT 81.490 22.480 81.810 22.540 ;
        RECT 53.890 22.200 62.170 22.340 ;
        RECT 64.470 22.340 64.790 22.400 ;
        RECT 64.945 22.340 65.235 22.385 ;
        RECT 64.470 22.200 65.235 22.340 ;
        RECT 53.890 22.140 54.210 22.200 ;
        RECT 60.330 22.140 60.650 22.200 ;
        RECT 64.470 22.140 64.790 22.200 ;
        RECT 64.945 22.155 65.235 22.200 ;
        RECT 77.810 22.140 78.130 22.400 ;
        RECT 5.520 21.520 83.260 22.000 ;
        RECT 54.810 21.320 55.130 21.380 ;
        RECT 41.100 21.180 55.130 21.320 ;
        RECT 41.100 21.025 41.240 21.180 ;
        RECT 54.810 21.120 55.130 21.180 ;
        RECT 58.030 21.120 58.350 21.380 ;
        RECT 41.025 20.795 41.315 21.025 ;
        RECT 44.230 20.980 44.550 21.040 ;
        RECT 46.085 20.980 46.375 21.025 ;
        RECT 44.230 20.840 46.375 20.980 ;
        RECT 44.230 20.780 44.550 20.840 ;
        RECT 46.085 20.795 46.375 20.840 ;
        RECT 46.530 20.780 46.850 21.040 ;
        RECT 47.235 20.980 47.525 21.025 ;
        RECT 48.830 20.980 49.150 21.040 ;
        RECT 47.235 20.840 49.150 20.980 ;
        RECT 47.235 20.795 47.525 20.840 ;
        RECT 48.830 20.780 49.150 20.840 ;
        RECT 63.720 20.980 64.010 21.025 ;
        RECT 64.470 20.980 64.790 21.040 ;
        RECT 69.070 20.980 69.390 21.040 ;
        RECT 74.590 20.980 74.910 21.040 ;
        RECT 63.720 20.840 64.790 20.980 ;
        RECT 63.720 20.795 64.010 20.840 ;
        RECT 64.470 20.780 64.790 20.840 ;
        RECT 66.400 20.840 80.340 20.980 ;
        RECT 41.945 20.640 42.235 20.685 ;
        RECT 42.405 20.640 42.695 20.685 ;
        RECT 41.945 20.500 42.695 20.640 ;
        RECT 41.945 20.455 42.235 20.500 ;
        RECT 42.405 20.455 42.695 20.500 ;
        RECT 43.325 20.640 43.615 20.685 ;
        RECT 43.325 20.500 45.380 20.640 ;
        RECT 43.325 20.455 43.615 20.500 ;
        RECT 44.245 20.115 44.535 20.345 ;
        RECT 45.240 20.300 45.380 20.500 ;
        RECT 45.610 20.440 45.930 20.700 ;
        RECT 47.910 20.440 48.230 20.700 ;
        RECT 50.640 20.640 50.930 20.685 ;
        RECT 52.050 20.640 52.370 20.700 ;
        RECT 50.640 20.500 52.370 20.640 ;
        RECT 50.640 20.455 50.930 20.500 ;
        RECT 52.050 20.440 52.370 20.500 ;
        RECT 64.945 20.640 65.235 20.685 ;
        RECT 65.405 20.640 65.695 20.685 ;
        RECT 66.400 20.640 66.540 20.840 ;
        RECT 69.070 20.780 69.390 20.840 ;
        RECT 74.590 20.780 74.910 20.840 ;
        RECT 66.770 20.685 67.090 20.700 ;
        RECT 64.945 20.500 66.540 20.640 ;
        RECT 66.740 20.640 67.090 20.685 ;
        RECT 77.350 20.640 77.670 20.700 ;
        RECT 80.200 20.685 80.340 20.840 ;
        RECT 78.790 20.640 79.080 20.685 ;
        RECT 66.740 20.500 67.240 20.640 ;
        RECT 77.350 20.500 79.080 20.640 ;
        RECT 64.945 20.455 65.235 20.500 ;
        RECT 65.405 20.455 65.695 20.500 ;
        RECT 66.740 20.455 67.090 20.500 ;
        RECT 66.770 20.440 67.090 20.455 ;
        RECT 77.350 20.440 77.670 20.500 ;
        RECT 78.790 20.455 79.080 20.500 ;
        RECT 80.125 20.455 80.415 20.685 ;
        RECT 46.990 20.300 47.310 20.360 ;
        RECT 45.240 20.160 47.310 20.300 ;
        RECT 44.320 19.960 44.460 20.115 ;
        RECT 46.990 20.100 47.310 20.160 ;
        RECT 49.290 20.100 49.610 20.360 ;
        RECT 50.185 20.300 50.475 20.345 ;
        RECT 51.375 20.300 51.665 20.345 ;
        RECT 53.895 20.300 54.185 20.345 ;
        RECT 50.185 20.160 54.185 20.300 ;
        RECT 50.185 20.115 50.475 20.160 ;
        RECT 51.375 20.115 51.665 20.160 ;
        RECT 53.895 20.115 54.185 20.160 ;
        RECT 60.355 20.300 60.645 20.345 ;
        RECT 62.875 20.300 63.165 20.345 ;
        RECT 64.065 20.300 64.355 20.345 ;
        RECT 60.355 20.160 64.355 20.300 ;
        RECT 60.355 20.115 60.645 20.160 ;
        RECT 62.875 20.115 63.165 20.160 ;
        RECT 64.065 20.115 64.355 20.160 ;
        RECT 66.285 20.300 66.575 20.345 ;
        RECT 67.475 20.300 67.765 20.345 ;
        RECT 69.995 20.300 70.285 20.345 ;
        RECT 66.285 20.160 70.285 20.300 ;
        RECT 66.285 20.115 66.575 20.160 ;
        RECT 67.475 20.115 67.765 20.160 ;
        RECT 69.995 20.115 70.285 20.160 ;
        RECT 75.535 20.300 75.825 20.345 ;
        RECT 78.055 20.300 78.345 20.345 ;
        RECT 79.245 20.300 79.535 20.345 ;
        RECT 75.535 20.160 79.535 20.300 ;
        RECT 75.535 20.115 75.825 20.160 ;
        RECT 78.055 20.115 78.345 20.160 ;
        RECT 79.245 20.115 79.535 20.160 ;
        RECT 49.790 19.960 50.080 20.005 ;
        RECT 51.890 19.960 52.180 20.005 ;
        RECT 53.460 19.960 53.750 20.005 ;
        RECT 44.320 19.820 49.520 19.960 ;
        RECT 40.090 19.420 40.410 19.680 ;
        RECT 44.690 19.420 45.010 19.680 ;
        RECT 49.380 19.620 49.520 19.820 ;
        RECT 49.790 19.820 53.750 19.960 ;
        RECT 49.790 19.775 50.080 19.820 ;
        RECT 51.890 19.775 52.180 19.820 ;
        RECT 53.460 19.775 53.750 19.820 ;
        RECT 56.190 19.760 56.510 20.020 ;
        RECT 60.790 19.960 61.080 20.005 ;
        RECT 62.360 19.960 62.650 20.005 ;
        RECT 64.460 19.960 64.750 20.005 ;
        RECT 60.790 19.820 64.750 19.960 ;
        RECT 60.790 19.775 61.080 19.820 ;
        RECT 62.360 19.775 62.650 19.820 ;
        RECT 64.460 19.775 64.750 19.820 ;
        RECT 65.890 19.960 66.180 20.005 ;
        RECT 67.990 19.960 68.280 20.005 ;
        RECT 69.560 19.960 69.850 20.005 ;
        RECT 65.890 19.820 69.850 19.960 ;
        RECT 65.890 19.775 66.180 19.820 ;
        RECT 67.990 19.775 68.280 19.820 ;
        RECT 69.560 19.775 69.850 19.820 ;
        RECT 73.225 19.960 73.515 20.005 ;
        RECT 75.050 19.960 75.370 20.020 ;
        RECT 73.225 19.820 75.370 19.960 ;
        RECT 73.225 19.775 73.515 19.820 ;
        RECT 75.050 19.760 75.370 19.820 ;
        RECT 75.970 19.960 76.260 20.005 ;
        RECT 77.540 19.960 77.830 20.005 ;
        RECT 79.640 19.960 79.930 20.005 ;
        RECT 75.970 19.820 79.930 19.960 ;
        RECT 75.970 19.775 76.260 19.820 ;
        RECT 77.540 19.775 77.830 19.820 ;
        RECT 79.640 19.775 79.930 19.820 ;
        RECT 54.350 19.620 54.670 19.680 ;
        RECT 49.380 19.480 54.670 19.620 ;
        RECT 54.350 19.420 54.670 19.480 ;
        RECT 72.290 19.420 72.610 19.680 ;
        RECT 5.520 18.800 83.260 19.280 ;
        RECT 48.830 18.400 49.150 18.660 ;
        RECT 54.350 18.600 54.670 18.660 ;
        RECT 56.205 18.600 56.495 18.645 ;
        RECT 57.585 18.600 57.875 18.645 ;
        RECT 54.350 18.460 57.875 18.600 ;
        RECT 54.350 18.400 54.670 18.460 ;
        RECT 56.205 18.415 56.495 18.460 ;
        RECT 57.585 18.415 57.875 18.460 ;
        RECT 58.505 18.600 58.795 18.645 ;
        RECT 60.790 18.600 61.110 18.660 ;
        RECT 58.505 18.460 61.110 18.600 ;
        RECT 58.505 18.415 58.795 18.460 ;
        RECT 60.790 18.400 61.110 18.460 ;
        RECT 66.785 18.600 67.075 18.645 ;
        RECT 70.910 18.600 71.230 18.660 ;
        RECT 78.270 18.600 78.590 18.660 ;
        RECT 81.505 18.600 81.795 18.645 ;
        RECT 66.785 18.460 71.230 18.600 ;
        RECT 66.785 18.415 67.075 18.460 ;
        RECT 70.910 18.400 71.230 18.460 ;
        RECT 71.460 18.460 73.440 18.600 ;
        RECT 49.790 18.260 50.080 18.305 ;
        RECT 51.890 18.260 52.180 18.305 ;
        RECT 53.460 18.260 53.750 18.305 ;
        RECT 49.790 18.120 53.750 18.260 ;
        RECT 49.790 18.075 50.080 18.120 ;
        RECT 51.890 18.075 52.180 18.120 ;
        RECT 53.460 18.075 53.750 18.120 ;
        RECT 60.370 18.260 60.660 18.305 ;
        RECT 62.470 18.260 62.760 18.305 ;
        RECT 64.040 18.260 64.330 18.305 ;
        RECT 69.530 18.260 69.850 18.320 ;
        RECT 71.460 18.260 71.600 18.460 ;
        RECT 60.370 18.120 64.330 18.260 ;
        RECT 60.370 18.075 60.660 18.120 ;
        RECT 62.470 18.075 62.760 18.120 ;
        RECT 64.040 18.075 64.330 18.120 ;
        RECT 65.020 18.120 71.600 18.260 ;
        RECT 71.920 18.120 72.980 18.260 ;
        RECT 40.090 17.920 40.410 17.980 ;
        RECT 40.090 17.780 46.760 17.920 ;
        RECT 40.090 17.720 40.410 17.780 ;
        RECT 43.770 17.380 44.090 17.640 ;
        RECT 46.070 17.380 46.390 17.640 ;
        RECT 46.620 17.580 46.760 17.780 ;
        RECT 49.290 17.720 49.610 17.980 ;
        RECT 50.185 17.920 50.475 17.965 ;
        RECT 51.375 17.920 51.665 17.965 ;
        RECT 53.895 17.920 54.185 17.965 ;
        RECT 50.185 17.780 54.185 17.920 ;
        RECT 50.185 17.735 50.475 17.780 ;
        RECT 51.375 17.735 51.665 17.780 ;
        RECT 53.895 17.735 54.185 17.780 ;
        RECT 57.110 17.920 57.430 17.980 ;
        RECT 59.870 17.920 60.190 17.980 ;
        RECT 57.110 17.780 60.190 17.920 ;
        RECT 57.110 17.720 57.430 17.780 ;
        RECT 59.870 17.720 60.190 17.780 ;
        RECT 60.765 17.920 61.055 17.965 ;
        RECT 61.955 17.920 62.245 17.965 ;
        RECT 64.475 17.920 64.765 17.965 ;
        RECT 60.765 17.780 64.765 17.920 ;
        RECT 60.765 17.735 61.055 17.780 ;
        RECT 61.955 17.735 62.245 17.780 ;
        RECT 64.475 17.735 64.765 17.780 ;
        RECT 50.585 17.580 50.875 17.625 ;
        RECT 65.020 17.580 65.160 18.120 ;
        RECT 69.530 18.060 69.850 18.120 ;
        RECT 69.085 17.920 69.375 17.965 ;
        RECT 71.920 17.920 72.060 18.120 ;
        RECT 69.085 17.780 72.060 17.920 ;
        RECT 69.085 17.735 69.375 17.780 ;
        RECT 46.620 17.440 50.875 17.580 ;
        RECT 50.585 17.395 50.875 17.440 ;
        RECT 55.360 17.440 65.160 17.580 ;
        RECT 65.390 17.580 65.710 17.640 ;
        RECT 67.245 17.580 67.535 17.625 ;
        RECT 71.370 17.580 71.690 17.640 ;
        RECT 65.390 17.440 71.690 17.580 ;
        RECT 45.610 17.240 45.930 17.300 ;
        RECT 55.360 17.240 55.500 17.440 ;
        RECT 65.390 17.380 65.710 17.440 ;
        RECT 67.245 17.395 67.535 17.440 ;
        RECT 71.370 17.380 71.690 17.440 ;
        RECT 71.830 17.380 72.150 17.640 ;
        RECT 72.840 17.625 72.980 18.120 ;
        RECT 72.305 17.395 72.595 17.625 ;
        RECT 72.765 17.395 73.055 17.625 ;
        RECT 73.300 17.580 73.440 18.460 ;
        RECT 78.270 18.460 81.795 18.600 ;
        RECT 78.270 18.400 78.590 18.460 ;
        RECT 81.505 18.415 81.795 18.460 ;
        RECT 75.090 18.260 75.380 18.305 ;
        RECT 77.190 18.260 77.480 18.305 ;
        RECT 78.760 18.260 79.050 18.305 ;
        RECT 75.090 18.120 79.050 18.260 ;
        RECT 75.090 18.075 75.380 18.120 ;
        RECT 77.190 18.075 77.480 18.120 ;
        RECT 78.760 18.075 79.050 18.120 ;
        RECT 74.590 17.720 74.910 17.980 ;
        RECT 75.485 17.920 75.775 17.965 ;
        RECT 76.675 17.920 76.965 17.965 ;
        RECT 79.195 17.920 79.485 17.965 ;
        RECT 75.485 17.780 79.485 17.920 ;
        RECT 75.485 17.735 75.775 17.780 ;
        RECT 76.675 17.735 76.965 17.780 ;
        RECT 79.195 17.735 79.485 17.780 ;
        RECT 73.685 17.580 73.975 17.625 ;
        RECT 73.300 17.440 73.975 17.580 ;
        RECT 73.685 17.395 73.975 17.440 ;
        RECT 75.940 17.580 76.230 17.625 ;
        RECT 77.810 17.580 78.130 17.640 ;
        RECT 75.940 17.440 78.130 17.580 ;
        RECT 75.940 17.395 76.230 17.440 ;
        RECT 45.610 17.100 55.500 17.240 ;
        RECT 55.730 17.240 56.050 17.300 ;
        RECT 57.570 17.285 57.890 17.300 ;
        RECT 56.665 17.240 56.955 17.285 ;
        RECT 55.730 17.100 56.955 17.240 ;
        RECT 45.610 17.040 45.930 17.100 ;
        RECT 55.730 17.040 56.050 17.100 ;
        RECT 56.665 17.055 56.955 17.100 ;
        RECT 57.570 17.055 57.955 17.285 ;
        RECT 61.220 17.240 61.510 17.285 ;
        RECT 62.170 17.240 62.490 17.300 ;
        RECT 61.220 17.100 62.490 17.240 ;
        RECT 61.220 17.055 61.510 17.100 ;
        RECT 57.570 17.040 57.890 17.055 ;
        RECT 62.170 17.040 62.490 17.100 ;
        RECT 68.165 17.240 68.455 17.285 ;
        RECT 69.530 17.240 69.850 17.300 ;
        RECT 68.165 17.100 69.850 17.240 ;
        RECT 72.380 17.240 72.520 17.395 ;
        RECT 77.810 17.380 78.130 17.440 ;
        RECT 79.190 17.240 79.510 17.300 ;
        RECT 72.380 17.100 79.510 17.240 ;
        RECT 68.165 17.055 68.455 17.100 ;
        RECT 69.530 17.040 69.850 17.100 ;
        RECT 79.190 17.040 79.510 17.100 ;
        RECT 42.865 16.900 43.155 16.945 ;
        RECT 43.770 16.900 44.090 16.960 ;
        RECT 42.865 16.760 44.090 16.900 ;
        RECT 42.865 16.715 43.155 16.760 ;
        RECT 43.770 16.700 44.090 16.760 ;
        RECT 70.450 16.700 70.770 16.960 ;
        RECT 5.520 16.080 83.260 16.560 ;
        RECT 46.070 15.880 46.390 15.940 ;
        RECT 47.005 15.880 47.295 15.925 ;
        RECT 46.070 15.740 47.295 15.880 ;
        RECT 46.070 15.680 46.390 15.740 ;
        RECT 47.005 15.695 47.295 15.740 ;
        RECT 52.050 15.680 52.370 15.940 ;
        RECT 53.905 15.880 54.195 15.925 ;
        RECT 56.190 15.880 56.510 15.940 ;
        RECT 53.905 15.740 56.510 15.880 ;
        RECT 53.905 15.695 54.195 15.740 ;
        RECT 56.190 15.680 56.510 15.740 ;
        RECT 69.530 15.880 69.850 15.940 ;
        RECT 70.465 15.880 70.755 15.925 ;
        RECT 72.750 15.880 73.070 15.940 ;
        RECT 69.530 15.740 73.070 15.880 ;
        RECT 69.530 15.680 69.850 15.740 ;
        RECT 70.465 15.695 70.755 15.740 ;
        RECT 72.750 15.680 73.070 15.740 ;
        RECT 74.145 15.880 74.435 15.925 ;
        RECT 79.650 15.880 79.970 15.940 ;
        RECT 74.145 15.740 79.970 15.880 ;
        RECT 74.145 15.695 74.435 15.740 ;
        RECT 79.650 15.680 79.970 15.740 ;
        RECT 41.440 15.540 41.730 15.585 ;
        RECT 44.690 15.540 45.010 15.600 ;
        RECT 41.440 15.400 45.010 15.540 ;
        RECT 41.440 15.355 41.730 15.400 ;
        RECT 44.690 15.340 45.010 15.400 ;
        RECT 59.870 15.540 60.190 15.600 ;
        RECT 69.070 15.540 69.390 15.600 ;
        RECT 59.870 15.400 69.390 15.540 ;
        RECT 59.870 15.340 60.190 15.400 ;
        RECT 27.670 15.200 27.990 15.260 ;
        RECT 63.640 15.245 63.780 15.400 ;
        RECT 69.070 15.340 69.390 15.400 ;
        RECT 73.225 15.540 73.515 15.585 ;
        RECT 73.670 15.540 73.990 15.600 ;
        RECT 73.225 15.400 73.990 15.540 ;
        RECT 73.225 15.355 73.515 15.400 ;
        RECT 73.670 15.340 73.990 15.400 ;
        RECT 75.940 15.540 76.230 15.585 ;
        RECT 76.430 15.540 76.750 15.600 ;
        RECT 75.940 15.400 76.750 15.540 ;
        RECT 75.940 15.355 76.230 15.400 ;
        RECT 76.430 15.340 76.750 15.400 ;
        RECT 40.105 15.200 40.395 15.245 ;
        RECT 27.670 15.060 40.395 15.200 ;
        RECT 27.670 15.000 27.990 15.060 ;
        RECT 40.105 15.015 40.395 15.060 ;
        RECT 63.565 15.200 63.855 15.245 ;
        RECT 64.900 15.200 65.190 15.245 ;
        RECT 70.450 15.200 70.770 15.260 ;
        RECT 63.565 15.060 63.965 15.200 ;
        RECT 64.900 15.060 70.770 15.200 ;
        RECT 63.565 15.015 63.855 15.060 ;
        RECT 64.900 15.015 65.190 15.060 ;
        RECT 70.450 15.000 70.770 15.060 ;
        RECT 70.910 15.000 71.230 15.260 ;
        RECT 71.370 15.200 71.690 15.260 ;
        RECT 72.305 15.200 72.595 15.245 ;
        RECT 72.750 15.200 73.070 15.260 ;
        RECT 71.370 15.060 73.070 15.200 ;
        RECT 71.370 15.000 71.690 15.060 ;
        RECT 72.305 15.015 72.595 15.060 ;
        RECT 72.750 15.000 73.070 15.060 ;
        RECT 74.590 15.000 74.910 15.260 ;
        RECT 40.985 14.860 41.275 14.905 ;
        RECT 42.175 14.860 42.465 14.905 ;
        RECT 44.695 14.860 44.985 14.905 ;
        RECT 40.985 14.720 44.985 14.860 ;
        RECT 40.985 14.675 41.275 14.720 ;
        RECT 42.175 14.675 42.465 14.720 ;
        RECT 44.695 14.675 44.985 14.720 ;
        RECT 54.350 14.660 54.670 14.920 ;
        RECT 54.810 14.660 55.130 14.920 ;
        RECT 64.445 14.860 64.735 14.905 ;
        RECT 65.635 14.860 65.925 14.905 ;
        RECT 68.155 14.860 68.445 14.905 ;
        RECT 64.445 14.720 68.445 14.860 ;
        RECT 64.445 14.675 64.735 14.720 ;
        RECT 65.635 14.675 65.925 14.720 ;
        RECT 68.155 14.675 68.445 14.720 ;
        RECT 75.485 14.860 75.775 14.905 ;
        RECT 76.675 14.860 76.965 14.905 ;
        RECT 79.195 14.860 79.485 14.905 ;
        RECT 75.485 14.720 79.485 14.860 ;
        RECT 75.485 14.675 75.775 14.720 ;
        RECT 76.675 14.675 76.965 14.720 ;
        RECT 79.195 14.675 79.485 14.720 ;
        RECT 40.590 14.520 40.880 14.565 ;
        RECT 42.690 14.520 42.980 14.565 ;
        RECT 44.260 14.520 44.550 14.565 ;
        RECT 40.590 14.380 44.550 14.520 ;
        RECT 40.590 14.335 40.880 14.380 ;
        RECT 42.690 14.335 42.980 14.380 ;
        RECT 44.260 14.335 44.550 14.380 ;
        RECT 64.050 14.520 64.340 14.565 ;
        RECT 66.150 14.520 66.440 14.565 ;
        RECT 67.720 14.520 68.010 14.565 ;
        RECT 64.050 14.380 68.010 14.520 ;
        RECT 64.050 14.335 64.340 14.380 ;
        RECT 66.150 14.335 66.440 14.380 ;
        RECT 67.720 14.335 68.010 14.380 ;
        RECT 69.070 14.520 69.390 14.580 ;
        RECT 72.290 14.520 72.610 14.580 ;
        RECT 69.070 14.380 72.610 14.520 ;
        RECT 69.070 14.320 69.390 14.380 ;
        RECT 72.290 14.320 72.610 14.380 ;
        RECT 75.090 14.520 75.380 14.565 ;
        RECT 77.190 14.520 77.480 14.565 ;
        RECT 78.760 14.520 79.050 14.565 ;
        RECT 75.090 14.380 79.050 14.520 ;
        RECT 75.090 14.335 75.380 14.380 ;
        RECT 77.190 14.335 77.480 14.380 ;
        RECT 78.760 14.335 79.050 14.380 ;
        RECT 71.845 14.180 72.135 14.225 ;
        RECT 73.210 14.180 73.530 14.240 ;
        RECT 71.845 14.040 73.530 14.180 ;
        RECT 71.845 13.995 72.135 14.040 ;
        RECT 73.210 13.980 73.530 14.040 ;
        RECT 73.670 14.180 73.990 14.240 ;
        RECT 81.505 14.180 81.795 14.225 ;
        RECT 73.670 14.040 81.795 14.180 ;
        RECT 73.670 13.980 73.990 14.040 ;
        RECT 81.505 13.995 81.795 14.040 ;
        RECT 5.520 13.360 83.260 13.840 ;
        RECT 74.130 12.960 74.450 13.220 ;
        RECT 75.970 12.960 76.290 13.220 ;
        RECT 78.745 13.160 79.035 13.205 ;
        RECT 80.110 13.160 80.430 13.220 ;
        RECT 78.745 13.020 80.430 13.160 ;
        RECT 78.745 12.975 79.035 13.020 ;
        RECT 80.110 12.960 80.430 13.020 ;
        RECT 81.030 12.960 81.350 13.220 ;
        RECT 41.945 12.820 42.235 12.865 ;
        RECT 44.230 12.820 44.550 12.880 ;
        RECT 41.945 12.680 44.550 12.820 ;
        RECT 41.945 12.635 42.235 12.680 ;
        RECT 44.230 12.620 44.550 12.680 ;
        RECT 50.225 12.820 50.515 12.865 ;
        RECT 54.350 12.820 54.670 12.880 ;
        RECT 50.225 12.680 54.670 12.820 ;
        RECT 50.225 12.635 50.515 12.680 ;
        RECT 54.350 12.620 54.670 12.680 ;
        RECT 72.750 12.820 73.070 12.880 ;
        RECT 72.750 12.680 77.120 12.820 ;
        RECT 72.750 12.620 73.070 12.680 ;
        RECT 37.345 12.480 37.635 12.525 ;
        RECT 46.530 12.480 46.850 12.540 ;
        RECT 37.345 12.340 46.850 12.480 ;
        RECT 37.345 12.295 37.635 12.340 ;
        RECT 46.530 12.280 46.850 12.340 ;
        RECT 35.490 12.140 35.810 12.200 ;
        RECT 35.965 12.140 36.255 12.185 ;
        RECT 35.490 12.000 36.255 12.140 ;
        RECT 35.490 11.940 35.810 12.000 ;
        RECT 35.965 11.955 36.255 12.000 ;
        RECT 43.770 11.940 44.090 12.200 ;
        RECT 46.070 12.140 46.390 12.200 ;
        RECT 47.005 12.140 47.295 12.185 ;
        RECT 46.070 12.000 47.295 12.140 ;
        RECT 46.070 11.940 46.390 12.000 ;
        RECT 47.005 11.955 47.295 12.000 ;
        RECT 66.325 12.140 66.615 12.185 ;
        RECT 69.070 12.140 69.390 12.200 ;
        RECT 66.325 12.000 69.390 12.140 ;
        RECT 66.325 11.955 66.615 12.000 ;
        RECT 69.070 11.940 69.390 12.000 ;
        RECT 69.530 11.940 69.850 12.200 ;
        RECT 69.990 12.140 70.310 12.200 ;
        RECT 72.765 12.140 73.055 12.185 ;
        RECT 69.990 12.000 73.055 12.140 ;
        RECT 69.990 11.940 70.310 12.000 ;
        RECT 72.765 11.955 73.055 12.000 ;
        RECT 73.210 11.940 73.530 12.200 ;
        RECT 73.670 12.140 73.990 12.200 ;
        RECT 76.980 12.185 77.120 12.680 ;
        RECT 75.065 12.140 75.355 12.185 ;
        RECT 73.670 12.000 75.355 12.140 ;
        RECT 73.670 11.940 73.990 12.000 ;
        RECT 75.065 11.955 75.355 12.000 ;
        RECT 76.905 11.955 77.195 12.185 ;
        RECT 77.825 12.140 78.115 12.185 ;
        RECT 78.270 12.140 78.590 12.200 ;
        RECT 80.125 12.140 80.415 12.185 ;
        RECT 77.825 12.000 80.415 12.140 ;
        RECT 77.825 11.955 78.115 12.000 ;
        RECT 78.270 11.940 78.590 12.000 ;
        RECT 80.125 11.955 80.415 12.000 ;
        RECT 38.710 11.800 39.030 11.860 ;
        RECT 41.025 11.800 41.315 11.845 ;
        RECT 38.710 11.660 41.315 11.800 ;
        RECT 38.710 11.600 39.030 11.660 ;
        RECT 41.025 11.615 41.315 11.660 ;
        RECT 48.370 11.800 48.690 11.860 ;
        RECT 49.305 11.800 49.595 11.845 ;
        RECT 48.370 11.660 49.595 11.800 ;
        RECT 48.370 11.600 48.690 11.660 ;
        RECT 49.305 11.615 49.595 11.660 ;
        RECT 41.930 11.460 42.250 11.520 ;
        RECT 42.865 11.460 43.155 11.505 ;
        RECT 41.930 11.320 43.155 11.460 ;
        RECT 41.930 11.260 42.250 11.320 ;
        RECT 42.865 11.275 43.155 11.320 ;
        RECT 45.150 11.460 45.470 11.520 ;
        RECT 46.085 11.460 46.375 11.505 ;
        RECT 45.150 11.320 46.375 11.460 ;
        RECT 45.150 11.260 45.470 11.320 ;
        RECT 46.085 11.275 46.375 11.320 ;
        RECT 64.470 11.460 64.790 11.520 ;
        RECT 65.405 11.460 65.695 11.505 ;
        RECT 64.470 11.320 65.695 11.460 ;
        RECT 64.470 11.260 64.790 11.320 ;
        RECT 65.405 11.275 65.695 11.320 ;
        RECT 67.690 11.460 68.010 11.520 ;
        RECT 68.625 11.460 68.915 11.505 ;
        RECT 67.690 11.320 68.915 11.460 ;
        RECT 67.690 11.260 68.010 11.320 ;
        RECT 68.625 11.275 68.915 11.320 ;
        RECT 70.910 11.460 71.230 11.520 ;
        RECT 71.845 11.460 72.135 11.505 ;
        RECT 70.910 11.320 72.135 11.460 ;
        RECT 70.910 11.260 71.230 11.320 ;
        RECT 71.845 11.275 72.135 11.320 ;
        RECT 5.520 10.640 83.260 11.120 ;
      LAYER met2 ;
        RECT 21.070 165.735 22.610 166.105 ;
        RECT 38.800 165.570 38.940 173.570 ;
        RECT 64.560 165.570 64.700 173.570 ;
        RECT 38.740 165.250 39.000 165.570 ;
        RECT 64.500 165.250 64.760 165.570 ;
        RECT 64.960 165.250 65.220 165.570 ;
        RECT 40.580 164.230 40.840 164.550 ;
        RECT 53.000 164.230 53.260 164.550 ;
        RECT 54.380 164.230 54.640 164.550 ;
        RECT 56.680 164.230 56.940 164.550 ;
        RECT 57.600 164.230 57.860 164.550 ;
        RECT 24.370 163.015 25.910 163.385 ;
        RECT 35.980 161.850 36.240 162.170 ;
        RECT 36.900 161.850 37.160 162.170 ;
        RECT 37.360 161.850 37.620 162.170 ;
        RECT 35.060 161.170 35.320 161.490 ;
        RECT 35.520 161.170 35.780 161.490 ;
        RECT 33.680 160.830 33.940 161.150 ;
        RECT 21.070 160.295 22.610 160.665 ;
        RECT 33.740 158.770 33.880 160.830 ;
        RECT 35.120 159.645 35.260 161.170 ;
        RECT 35.050 159.275 35.330 159.645 ;
        RECT 33.680 158.450 33.940 158.770 ;
        RECT 34.600 158.450 34.860 158.770 ;
        RECT 24.370 157.575 25.910 157.945 ;
        RECT 30.460 156.070 30.720 156.390 ;
        RECT 21.070 154.855 22.610 155.225 ;
        RECT 30.520 154.690 30.660 156.070 ;
        RECT 34.660 156.050 34.800 158.450 ;
        RECT 35.580 156.730 35.720 161.170 ;
        RECT 36.040 158.965 36.180 161.850 ;
        RECT 35.970 158.595 36.250 158.965 ;
        RECT 36.960 157.410 37.100 161.850 ;
        RECT 36.900 157.090 37.160 157.410 ;
        RECT 35.520 156.410 35.780 156.730 ;
        RECT 34.600 155.730 34.860 156.050 ;
        RECT 33.680 155.390 33.940 155.710 ;
        RECT 30.460 154.370 30.720 154.690 ;
        RECT 24.370 152.135 25.910 152.505 ;
        RECT 29.540 150.970 29.800 151.290 ;
        RECT 0.550 150.435 0.830 150.805 ;
        RECT 0.620 88.730 0.760 150.435 ;
        RECT 27.700 149.950 27.960 150.270 ;
        RECT 21.070 149.415 22.610 149.785 ;
        RECT 24.370 146.695 25.910 147.065 ;
        RECT 27.760 145.850 27.900 149.950 ;
        RECT 28.620 147.230 28.880 147.550 ;
        RECT 27.700 145.530 27.960 145.850 ;
        RECT 21.070 143.975 22.610 144.345 ;
        RECT 28.680 142.790 28.820 147.230 ;
        RECT 29.600 146.190 29.740 150.970 ;
        RECT 30.520 150.950 30.660 154.370 ;
        RECT 32.300 153.350 32.560 153.670 ;
        RECT 32.360 151.630 32.500 153.350 ;
        RECT 33.740 151.970 33.880 155.390 ;
        RECT 34.660 153.670 34.800 155.730 ;
        RECT 37.420 154.090 37.560 161.850 ;
        RECT 38.280 161.510 38.540 161.830 ;
        RECT 37.820 156.410 38.080 156.730 ;
        RECT 36.960 153.950 37.560 154.090 ;
        RECT 34.600 153.350 34.860 153.670 ;
        RECT 35.060 153.010 35.320 153.330 ;
        RECT 33.680 151.650 33.940 151.970 ;
        RECT 34.140 151.650 34.400 151.970 ;
        RECT 32.300 151.310 32.560 151.630 ;
        RECT 30.920 150.970 31.180 151.290 ;
        RECT 30.460 150.630 30.720 150.950 ;
        RECT 30.520 149.250 30.660 150.630 ;
        RECT 30.460 148.930 30.720 149.250 ;
        RECT 30.520 147.550 30.660 148.930 ;
        RECT 30.980 148.230 31.120 150.970 ;
        RECT 30.920 147.910 31.180 148.230 ;
        RECT 34.200 147.970 34.340 151.650 ;
        RECT 35.120 150.270 35.260 153.010 ;
        RECT 35.060 149.950 35.320 150.270 ;
        RECT 36.960 149.250 37.100 153.950 ;
        RECT 37.360 153.350 37.620 153.670 ;
        RECT 37.420 151.290 37.560 153.350 ;
        RECT 37.360 150.970 37.620 151.290 ;
        RECT 37.880 150.690 38.020 156.410 ;
        RECT 38.340 156.390 38.480 161.510 ;
        RECT 40.640 160.130 40.780 164.230 ;
        RECT 52.080 163.550 52.340 163.870 ;
        RECT 45.640 161.850 45.900 162.170 ;
        RECT 41.960 160.830 42.220 161.150 ;
        RECT 40.580 159.810 40.840 160.130 ;
        RECT 40.640 159.110 40.780 159.810 ;
        RECT 42.020 159.450 42.160 160.830 ;
        RECT 45.700 160.130 45.840 161.850 ;
        RECT 45.640 159.810 45.900 160.130 ;
        RECT 41.960 159.130 42.220 159.450 ;
        RECT 40.580 158.790 40.840 159.110 ;
        RECT 42.420 158.850 42.680 159.110 ;
        RECT 42.020 158.790 42.680 158.850 ;
        RECT 47.020 158.790 47.280 159.110 ;
        RECT 48.400 158.790 48.660 159.110 ;
        RECT 42.020 158.710 42.620 158.790 ;
        RECT 39.660 158.110 39.920 158.430 ;
        RECT 39.720 157.070 39.860 158.110 ;
        RECT 39.660 156.750 39.920 157.070 ;
        RECT 38.280 156.070 38.540 156.390 ;
        RECT 40.120 156.070 40.380 156.390 ;
        RECT 37.420 150.550 38.020 150.690 ;
        RECT 35.520 148.930 35.780 149.250 ;
        RECT 36.900 148.930 37.160 149.250 ;
        RECT 34.590 148.395 34.870 148.765 ;
        RECT 34.660 148.230 34.800 148.395 ;
        RECT 33.280 147.830 34.340 147.970 ;
        RECT 34.600 147.910 34.860 148.230 ;
        RECT 35.580 147.890 35.720 148.930 ;
        RECT 35.980 148.590 36.240 148.910 ;
        RECT 30.460 147.230 30.720 147.550 ;
        RECT 33.280 146.530 33.420 147.830 ;
        RECT 35.520 147.570 35.780 147.890 ;
        RECT 33.680 147.230 33.940 147.550 ;
        RECT 34.600 147.230 34.860 147.550 ;
        RECT 33.740 146.530 33.880 147.230 ;
        RECT 33.220 146.210 33.480 146.530 ;
        RECT 33.680 146.210 33.940 146.530 ;
        RECT 29.540 145.870 29.800 146.190 ;
        RECT 34.140 145.870 34.400 146.190 ;
        RECT 33.220 145.530 33.480 145.850 ;
        RECT 33.280 143.210 33.420 145.530 ;
        RECT 34.200 143.810 34.340 145.870 ;
        RECT 34.660 145.850 34.800 147.230 ;
        RECT 34.600 145.530 34.860 145.850 ;
        RECT 36.040 145.170 36.180 148.590 ;
        RECT 36.430 148.395 36.710 148.765 ;
        RECT 36.500 145.170 36.640 148.395 ;
        RECT 35.980 144.850 36.240 145.170 ;
        RECT 36.440 144.850 36.700 145.170 ;
        RECT 34.140 143.490 34.400 143.810 ;
        RECT 33.280 143.070 34.340 143.210 ;
        RECT 34.200 142.790 34.340 143.070 ;
        RECT 36.040 142.790 36.180 144.850 ;
        RECT 28.620 142.470 28.880 142.790 ;
        RECT 34.140 142.470 34.400 142.790 ;
        RECT 35.980 142.470 36.240 142.790 ;
        RECT 14.820 142.130 15.080 142.450 ;
        RECT 12.980 140.090 13.240 140.410 ;
        RECT 12.060 136.690 12.320 137.010 ;
        RECT 10.680 135.330 10.940 135.650 ;
        RECT 8.380 134.650 8.640 134.970 ;
        RECT 8.440 132.590 8.580 134.650 ;
        RECT 10.220 134.310 10.480 134.630 ;
        RECT 8.380 132.270 8.640 132.590 ;
        RECT 4.230 126.635 4.510 127.005 ;
        RECT 4.300 126.470 4.440 126.635 ;
        RECT 4.240 126.150 4.500 126.470 ;
        RECT 10.280 124.770 10.420 134.310 ;
        RECT 10.220 124.450 10.480 124.770 ;
        RECT 9.300 123.430 9.560 123.750 ;
        RECT 8.840 122.750 9.100 123.070 ;
        RECT 8.900 121.030 9.040 122.750 ;
        RECT 9.360 122.050 9.500 123.430 ;
        RECT 9.300 121.730 9.560 122.050 ;
        RECT 7.000 120.710 7.260 121.030 ;
        RECT 8.840 120.710 9.100 121.030 ;
        RECT 10.220 120.710 10.480 121.030 ;
        RECT 7.060 118.650 7.200 120.710 ;
        RECT 7.000 118.330 7.260 118.650 ;
        RECT 8.380 118.330 8.640 118.650 ;
        RECT 8.440 116.610 8.580 118.330 ;
        RECT 8.380 116.290 8.640 116.610 ;
        RECT 10.280 115.930 10.420 120.710 ;
        RECT 10.220 115.610 10.480 115.930 ;
        RECT 4.240 107.450 4.500 107.770 ;
        RECT 4.300 106.605 4.440 107.450 ;
        RECT 4.230 106.235 4.510 106.605 ;
        RECT 10.280 105.390 10.420 115.610 ;
        RECT 10.740 115.590 10.880 135.330 ;
        RECT 11.600 134.990 11.860 135.310 ;
        RECT 11.140 134.310 11.400 134.630 ;
        RECT 11.200 132.930 11.340 134.310 ;
        RECT 11.140 132.610 11.400 132.930 ;
        RECT 11.660 132.840 11.800 134.990 ;
        RECT 12.120 134.290 12.260 136.690 ;
        RECT 12.060 133.970 12.320 134.290 ;
        RECT 13.040 132.930 13.180 140.090 ;
        RECT 13.900 139.750 14.160 140.070 ;
        RECT 13.960 137.350 14.100 139.750 ;
        RECT 13.900 137.030 14.160 137.350 ;
        RECT 14.360 135.330 14.620 135.650 ;
        RECT 13.900 135.165 14.160 135.310 ;
        RECT 13.890 135.050 14.170 135.165 ;
        RECT 13.500 134.910 14.170 135.050 ;
        RECT 11.660 132.700 12.720 132.840 ;
        RECT 12.580 132.250 12.720 132.700 ;
        RECT 12.980 132.610 13.240 132.930 ;
        RECT 12.060 131.930 12.320 132.250 ;
        RECT 12.520 131.930 12.780 132.250 ;
        RECT 12.970 132.075 13.250 132.445 ;
        RECT 12.120 129.870 12.260 131.930 ;
        RECT 12.060 129.550 12.320 129.870 ;
        RECT 13.040 123.750 13.180 132.075 ;
        RECT 12.980 123.430 13.240 123.750 ;
        RECT 12.980 120.370 13.240 120.690 ;
        RECT 13.040 116.610 13.180 120.370 ;
        RECT 12.980 116.290 13.240 116.610 ;
        RECT 13.500 116.270 13.640 134.910 ;
        RECT 13.890 134.795 14.170 134.910 ;
        RECT 14.420 134.485 14.560 135.330 ;
        RECT 14.880 134.630 15.020 142.130 ;
        RECT 24.370 141.255 25.910 141.625 ;
        RECT 17.120 140.090 17.380 140.410 ;
        RECT 23.560 140.090 23.820 140.410 ;
        RECT 33.680 140.090 33.940 140.410 ;
        RECT 16.660 136.350 16.920 136.670 ;
        RECT 14.350 134.115 14.630 134.485 ;
        RECT 14.820 134.310 15.080 134.630 ;
        RECT 16.720 134.540 16.860 136.350 ;
        RECT 16.260 134.400 16.860 134.540 ;
        RECT 13.900 132.610 14.160 132.930 ;
        RECT 13.960 132.445 14.100 132.610 ;
        RECT 13.890 132.075 14.170 132.445 ;
        RECT 14.880 131.820 15.020 134.310 ;
        RECT 15.280 133.970 15.540 134.290 ;
        RECT 15.340 133.805 15.480 133.970 ;
        RECT 15.270 133.435 15.550 133.805 ;
        RECT 15.740 131.820 16.000 131.910 ;
        RECT 14.880 131.680 16.000 131.820 ;
        RECT 14.360 130.910 14.620 131.230 ;
        RECT 14.420 124.090 14.560 130.910 ;
        RECT 14.360 123.770 14.620 124.090 ;
        RECT 15.340 121.370 15.480 131.680 ;
        RECT 15.740 131.590 16.000 131.680 ;
        RECT 16.260 131.230 16.400 134.400 ;
        RECT 17.180 133.950 17.320 140.090 ;
        RECT 18.960 139.410 19.220 139.730 ;
        RECT 19.020 137.350 19.160 139.410 ;
        RECT 19.880 139.070 20.140 139.390 ;
        RECT 18.960 137.030 19.220 137.350 ;
        RECT 19.420 136.350 19.680 136.670 ;
        RECT 19.480 135.650 19.620 136.350 ;
        RECT 19.420 135.330 19.680 135.650 ;
        RECT 17.580 134.650 17.840 134.970 ;
        RECT 17.120 133.630 17.380 133.950 ;
        RECT 17.640 133.805 17.780 134.650 ;
        RECT 16.660 131.590 16.920 131.910 ;
        RECT 16.200 130.910 16.460 131.230 ;
        RECT 15.740 129.550 16.000 129.870 ;
        RECT 15.280 121.050 15.540 121.370 ;
        RECT 15.800 121.030 15.940 129.550 ;
        RECT 16.260 128.510 16.400 130.910 ;
        RECT 16.720 129.870 16.860 131.590 ;
        RECT 16.660 129.550 16.920 129.870 ;
        RECT 17.180 128.850 17.320 133.630 ;
        RECT 17.570 133.435 17.850 133.805 ;
        RECT 18.960 132.610 19.220 132.930 ;
        RECT 19.020 131.570 19.160 132.610 ;
        RECT 19.420 131.820 19.680 131.910 ;
        RECT 19.940 131.820 20.080 139.070 ;
        RECT 21.070 138.535 22.610 138.905 ;
        RECT 20.800 137.030 21.060 137.350 ;
        RECT 20.340 136.690 20.600 137.010 ;
        RECT 19.420 131.680 20.080 131.820 ;
        RECT 19.420 131.590 19.680 131.680 ;
        RECT 17.580 131.250 17.840 131.570 ;
        RECT 18.960 131.250 19.220 131.570 ;
        RECT 17.120 128.530 17.380 128.850 ;
        RECT 16.200 128.190 16.460 128.510 ;
        RECT 17.640 128.250 17.780 131.250 ;
        RECT 19.940 130.210 20.080 131.680 ;
        RECT 19.880 129.890 20.140 130.210 ;
        RECT 14.820 120.710 15.080 121.030 ;
        RECT 15.740 120.710 16.000 121.030 ;
        RECT 14.880 119.330 15.020 120.710 ;
        RECT 15.280 120.030 15.540 120.350 ;
        RECT 15.740 120.260 16.000 120.350 ;
        RECT 16.260 120.260 16.400 128.190 ;
        RECT 17.180 128.110 17.780 128.250 ;
        RECT 17.180 124.090 17.320 128.110 ;
        RECT 17.580 125.470 17.840 125.790 ;
        RECT 17.640 124.090 17.780 125.470 ;
        RECT 18.040 124.110 18.300 124.430 ;
        RECT 17.120 123.770 17.380 124.090 ;
        RECT 17.580 123.770 17.840 124.090 ;
        RECT 17.180 123.490 17.320 123.770 ;
        RECT 17.180 123.350 17.780 123.490 ;
        RECT 17.120 122.750 17.380 123.070 ;
        RECT 17.180 121.030 17.320 122.750 ;
        RECT 17.120 120.885 17.380 121.030 ;
        RECT 16.660 120.370 16.920 120.690 ;
        RECT 17.110 120.515 17.390 120.885 ;
        RECT 15.740 120.120 16.400 120.260 ;
        RECT 15.740 120.030 16.000 120.120 ;
        RECT 14.820 119.010 15.080 119.330 ;
        RECT 15.340 118.650 15.480 120.030 ;
        RECT 15.800 118.650 15.940 120.030 ;
        RECT 16.720 118.650 16.860 120.370 ;
        RECT 14.360 118.330 14.620 118.650 ;
        RECT 15.280 118.330 15.540 118.650 ;
        RECT 15.740 118.330 16.000 118.650 ;
        RECT 16.660 118.330 16.920 118.650 ;
        RECT 17.120 118.330 17.380 118.650 ;
        RECT 13.440 116.180 13.700 116.270 ;
        RECT 13.440 116.040 14.100 116.180 ;
        RECT 13.440 115.950 13.700 116.040 ;
        RECT 10.680 115.270 10.940 115.590 ;
        RECT 11.600 115.270 11.860 115.590 ;
        RECT 10.220 105.070 10.480 105.390 ;
        RECT 10.740 105.050 10.880 115.270 ;
        RECT 11.140 113.570 11.400 113.890 ;
        RECT 10.680 104.730 10.940 105.050 ;
        RECT 11.200 104.565 11.340 113.570 ;
        RECT 11.660 112.530 11.800 115.270 ;
        RECT 12.520 114.590 12.780 114.910 ;
        RECT 12.580 113.890 12.720 114.590 ;
        RECT 12.520 113.570 12.780 113.890 ;
        RECT 12.060 112.550 12.320 112.870 ;
        RECT 11.600 112.210 11.860 112.530 ;
        RECT 12.120 110.470 12.260 112.550 ;
        RECT 11.660 110.330 12.260 110.470 ;
        RECT 11.130 104.195 11.410 104.565 ;
        RECT 11.140 104.050 11.400 104.195 ;
        RECT 7.460 103.710 7.720 104.030 ;
        RECT 7.000 101.670 7.260 101.990 ;
        RECT 7.060 100.290 7.200 101.670 ;
        RECT 7.000 99.970 7.260 100.290 ;
        RECT 7.060 99.610 7.200 99.970 ;
        RECT 7.000 99.290 7.260 99.610 ;
        RECT 7.520 99.270 7.660 103.710 ;
        RECT 7.460 98.950 7.720 99.270 ;
        RECT 11.660 95.870 11.800 110.330 ;
        RECT 13.960 105.050 14.100 116.040 ;
        RECT 14.420 115.590 14.560 118.330 ;
        RECT 14.820 117.310 15.080 117.630 ;
        RECT 14.880 116.610 15.020 117.310 ;
        RECT 14.820 116.290 15.080 116.610 ;
        RECT 14.880 115.590 15.020 116.290 ;
        RECT 15.340 116.270 15.480 118.330 ;
        RECT 15.280 115.950 15.540 116.270 ;
        RECT 16.660 115.610 16.920 115.930 ;
        RECT 14.360 115.270 14.620 115.590 ;
        RECT 14.820 115.270 15.080 115.590 ;
        RECT 16.200 115.270 16.460 115.590 ;
        RECT 14.420 113.890 14.560 115.270 ;
        RECT 14.880 114.650 15.020 115.270 ;
        RECT 15.280 115.160 15.540 115.250 ;
        RECT 15.280 115.020 15.940 115.160 ;
        RECT 15.280 114.930 15.540 115.020 ;
        RECT 14.880 114.510 15.480 114.650 ;
        RECT 14.360 113.570 14.620 113.890 ;
        RECT 15.340 113.210 15.480 114.510 ;
        RECT 15.280 112.890 15.540 113.210 ;
        RECT 15.800 112.190 15.940 115.020 ;
        RECT 16.260 112.870 16.400 115.270 ;
        RECT 16.200 112.550 16.460 112.870 ;
        RECT 15.740 111.870 16.000 112.190 ;
        RECT 15.800 107.770 15.940 111.870 ;
        RECT 16.720 111.170 16.860 115.610 ;
        RECT 16.660 110.850 16.920 111.170 ;
        RECT 16.660 110.470 16.920 110.490 ;
        RECT 17.180 110.470 17.320 118.330 ;
        RECT 17.640 113.890 17.780 123.350 ;
        RECT 18.100 121.030 18.240 124.110 ;
        RECT 19.940 124.090 20.080 129.890 ;
        RECT 20.400 128.850 20.540 136.690 ;
        RECT 20.860 135.310 21.000 137.030 ;
        RECT 23.100 136.690 23.360 137.010 ;
        RECT 20.800 134.990 21.060 135.310 ;
        RECT 20.860 133.950 21.000 134.990 ;
        RECT 20.800 133.630 21.060 133.950 ;
        RECT 21.070 133.095 22.610 133.465 ;
        RECT 23.160 132.590 23.300 136.690 ;
        RECT 23.620 135.650 23.760 140.090 ;
        RECT 29.080 139.410 29.340 139.730 ;
        RECT 28.160 137.030 28.420 137.350 ;
        RECT 26.320 136.350 26.580 136.670 ;
        RECT 24.370 135.815 25.910 136.185 ;
        RECT 23.560 135.330 23.820 135.650 ;
        RECT 23.100 132.270 23.360 132.590 ;
        RECT 21.260 131.930 21.520 132.250 ;
        RECT 21.320 131.230 21.460 131.930 ;
        RECT 22.180 131.250 22.440 131.570 ;
        RECT 21.260 130.910 21.520 131.230 ;
        RECT 22.240 129.190 22.380 131.250 ;
        RECT 23.100 130.910 23.360 131.230 ;
        RECT 22.180 128.870 22.440 129.190 ;
        RECT 20.340 128.530 20.600 128.850 ;
        RECT 21.070 127.655 22.610 128.025 ;
        RECT 23.160 126.810 23.300 130.910 ;
        RECT 23.620 129.870 23.760 135.330 ;
        RECT 24.010 134.795 24.290 135.165 ;
        RECT 24.080 132.250 24.220 134.795 ;
        RECT 24.940 134.650 25.200 134.970 ;
        RECT 24.020 131.930 24.280 132.250 ;
        RECT 24.020 131.250 24.280 131.570 ;
        RECT 23.560 129.550 23.820 129.870 ;
        RECT 23.100 126.490 23.360 126.810 ;
        RECT 23.160 124.770 23.300 126.490 ;
        RECT 23.100 124.450 23.360 124.770 ;
        RECT 23.620 124.430 23.760 129.550 ;
        RECT 24.080 129.530 24.220 131.250 ;
        RECT 25.000 131.230 25.140 134.650 ;
        RECT 25.390 134.115 25.670 134.485 ;
        RECT 25.460 132.250 25.600 134.115 ;
        RECT 25.400 131.930 25.660 132.250 ;
        RECT 24.940 130.910 25.200 131.230 ;
        RECT 25.460 131.140 25.600 131.930 ;
        RECT 26.380 131.570 26.520 136.350 ;
        RECT 28.220 133.950 28.360 137.030 ;
        RECT 28.160 133.630 28.420 133.950 ;
        RECT 27.700 131.930 27.960 132.250 ;
        RECT 26.780 131.590 27.040 131.910 ;
        RECT 26.320 131.250 26.580 131.570 ;
        RECT 25.460 131.000 26.185 131.140 ;
        RECT 26.045 130.970 26.185 131.000 ;
        RECT 26.045 130.830 26.520 130.970 ;
        RECT 24.370 130.375 25.910 130.745 ;
        RECT 24.020 129.210 24.280 129.530 ;
        RECT 24.080 128.510 24.220 129.210 ;
        RECT 24.020 128.190 24.280 128.510 ;
        RECT 24.080 124.680 24.220 128.190 ;
        RECT 24.370 124.935 25.910 125.305 ;
        RECT 24.080 124.540 24.680 124.680 ;
        RECT 23.560 124.110 23.820 124.430 ;
        RECT 19.880 123.770 20.140 124.090 ;
        RECT 19.420 123.430 19.680 123.750 ;
        RECT 23.620 123.490 23.760 124.110 ;
        RECT 24.540 123.750 24.680 124.540 ;
        RECT 18.960 123.090 19.220 123.410 ;
        RECT 18.040 120.710 18.300 121.030 ;
        RECT 18.500 118.560 18.760 118.650 ;
        RECT 19.020 118.560 19.160 123.090 ;
        RECT 19.480 120.770 19.620 123.430 ;
        RECT 23.100 123.090 23.360 123.410 ;
        RECT 23.620 123.350 24.220 123.490 ;
        RECT 24.480 123.430 24.740 123.750 ;
        RECT 20.340 122.750 20.600 123.070 ;
        RECT 19.880 121.565 20.140 121.710 ;
        RECT 19.870 121.195 20.150 121.565 ;
        RECT 20.400 121.030 20.540 122.750 ;
        RECT 21.070 122.215 22.610 122.585 ;
        RECT 21.260 121.730 21.520 122.050 ;
        RECT 19.480 120.630 20.080 120.770 ;
        RECT 20.340 120.710 20.600 121.030 ;
        RECT 19.940 120.090 20.080 120.630 ;
        RECT 20.340 120.090 20.600 120.350 ;
        RECT 19.940 120.030 20.600 120.090 ;
        RECT 19.940 119.950 20.540 120.030 ;
        RECT 18.500 118.420 19.160 118.560 ;
        RECT 18.500 118.330 18.760 118.420 ;
        RECT 18.040 117.990 18.300 118.310 ;
        RECT 17.580 113.570 17.840 113.890 ;
        RECT 16.660 110.400 17.320 110.470 ;
        RECT 16.260 110.330 17.320 110.400 ;
        RECT 16.260 110.260 16.920 110.330 ;
        RECT 15.740 107.450 16.000 107.770 ;
        RECT 13.900 104.960 14.160 105.050 ;
        RECT 13.040 104.820 14.160 104.960 ;
        RECT 12.060 104.620 12.320 104.710 ;
        RECT 13.040 104.620 13.180 104.820 ;
        RECT 13.900 104.730 14.160 104.820 ;
        RECT 12.060 104.480 13.180 104.620 ;
        RECT 14.360 104.565 14.620 104.710 ;
        RECT 12.060 104.390 12.320 104.480 ;
        RECT 14.350 104.195 14.630 104.565 ;
        RECT 12.060 103.710 12.320 104.030 ;
        RECT 12.120 102.670 12.260 103.710 ;
        RECT 12.060 102.350 12.320 102.670 ;
        RECT 14.420 102.330 14.560 104.195 ;
        RECT 14.820 104.050 15.080 104.370 ;
        RECT 14.360 102.010 14.620 102.330 ;
        RECT 14.420 99.950 14.560 102.010 ;
        RECT 14.880 101.990 15.020 104.050 ;
        RECT 15.800 103.010 15.940 107.450 ;
        RECT 15.740 102.690 16.000 103.010 ;
        RECT 15.800 102.330 15.940 102.690 ;
        RECT 15.740 102.010 16.000 102.330 ;
        RECT 14.820 101.670 15.080 101.990 ;
        RECT 14.360 99.630 14.620 99.950 ;
        RECT 11.600 95.550 11.860 95.870 ;
        RECT 13.440 95.550 13.700 95.870 ;
        RECT 15.740 95.780 16.000 95.870 ;
        RECT 16.260 95.780 16.400 110.260 ;
        RECT 16.660 110.170 16.920 110.260 ;
        RECT 18.100 108.450 18.240 117.990 ;
        RECT 18.040 108.130 18.300 108.450 ;
        RECT 16.660 107.450 16.920 107.770 ;
        RECT 16.720 105.730 16.860 107.450 ;
        RECT 17.120 106.430 17.380 106.750 ;
        RECT 16.660 105.410 16.920 105.730 ;
        RECT 17.180 104.710 17.320 106.430 ;
        RECT 17.120 104.390 17.380 104.710 ;
        RECT 17.180 98.590 17.320 104.390 ;
        RECT 18.100 103.090 18.240 108.130 ;
        RECT 18.560 103.770 18.700 118.330 ;
        RECT 20.400 118.310 20.540 119.950 ;
        RECT 21.320 118.650 21.460 121.730 ;
        RECT 21.260 118.330 21.520 118.650 ;
        RECT 20.340 117.990 20.600 118.310 ;
        RECT 18.960 117.310 19.220 117.630 ;
        RECT 20.340 117.310 20.600 117.630 ;
        RECT 19.020 115.590 19.160 117.310 ;
        RECT 18.960 115.270 19.220 115.590 ;
        RECT 20.400 115.500 20.540 117.310 ;
        RECT 21.070 116.775 22.610 117.145 ;
        RECT 20.800 115.500 21.060 115.590 ;
        RECT 20.400 115.360 21.060 115.500 ;
        RECT 18.960 113.570 19.220 113.890 ;
        RECT 19.020 105.730 19.160 113.570 ;
        RECT 20.400 113.210 20.540 115.360 ;
        RECT 20.800 115.270 21.060 115.360 ;
        RECT 23.160 115.330 23.300 123.090 ;
        RECT 23.560 122.750 23.820 123.070 ;
        RECT 21.260 114.930 21.520 115.250 ;
        RECT 22.240 115.190 23.300 115.330 ;
        RECT 20.340 112.890 20.600 113.210 ;
        RECT 21.320 112.530 21.460 114.930 ;
        RECT 22.240 113.210 22.380 115.190 ;
        RECT 23.620 114.910 23.760 122.750 ;
        RECT 24.080 117.970 24.220 123.350 ;
        RECT 24.540 122.050 24.680 123.430 ;
        RECT 24.480 121.730 24.740 122.050 ;
        RECT 24.940 121.280 25.200 121.370 ;
        RECT 26.380 121.280 26.520 130.830 ;
        RECT 26.840 130.210 26.980 131.590 ;
        RECT 27.760 130.210 27.900 131.930 ;
        RECT 26.780 129.890 27.040 130.210 ;
        RECT 27.700 129.890 27.960 130.210 ;
        RECT 26.840 129.190 26.980 129.890 ;
        RECT 26.780 128.870 27.040 129.190 ;
        RECT 26.840 122.050 26.980 128.870 ;
        RECT 28.220 126.130 28.360 133.630 ;
        RECT 29.140 131.570 29.280 139.410 ;
        RECT 30.000 136.690 30.260 137.010 ;
        RECT 29.530 134.795 29.810 135.165 ;
        RECT 29.080 131.250 29.340 131.570 ;
        RECT 29.600 131.230 29.740 134.795 ;
        RECT 30.060 132.590 30.200 136.690 ;
        RECT 33.740 136.670 33.880 140.090 ;
        RECT 31.380 136.350 31.640 136.670 ;
        RECT 33.680 136.350 33.940 136.670 ;
        RECT 30.460 133.630 30.720 133.950 ;
        RECT 30.000 132.270 30.260 132.590 ;
        RECT 30.000 131.820 30.260 131.910 ;
        RECT 30.520 131.820 30.660 133.630 ;
        RECT 31.440 131.910 31.580 136.350 ;
        RECT 30.000 131.680 30.660 131.820 ;
        RECT 30.000 131.590 30.260 131.680 ;
        RECT 28.620 130.910 28.880 131.230 ;
        RECT 29.540 130.910 29.800 131.230 ;
        RECT 28.680 129.530 28.820 130.910 ;
        RECT 28.620 129.210 28.880 129.530 ;
        RECT 29.080 129.210 29.340 129.530 ;
        RECT 29.140 128.510 29.280 129.210 ;
        RECT 29.080 128.190 29.340 128.510 ;
        RECT 28.160 125.810 28.420 126.130 ;
        RECT 28.220 124.090 28.360 125.810 ;
        RECT 29.140 124.090 29.280 128.190 ;
        RECT 28.160 123.770 28.420 124.090 ;
        RECT 29.080 123.770 29.340 124.090 ;
        RECT 27.240 122.750 27.500 123.070 ;
        RECT 26.780 121.730 27.040 122.050 ;
        RECT 27.300 121.370 27.440 122.750 ;
        RECT 24.940 121.140 26.980 121.280 ;
        RECT 24.940 121.050 25.200 121.140 ;
        RECT 26.840 120.770 26.980 121.140 ;
        RECT 27.240 121.050 27.500 121.370 ;
        RECT 25.860 120.600 26.120 120.690 ;
        RECT 26.840 120.630 27.440 120.770 ;
        RECT 25.860 120.460 26.520 120.600 ;
        RECT 25.860 120.370 26.120 120.460 ;
        RECT 24.370 119.495 25.910 119.865 ;
        RECT 24.020 117.650 24.280 117.970 ;
        RECT 23.100 114.590 23.360 114.910 ;
        RECT 23.560 114.590 23.820 114.910 ;
        RECT 24.020 114.590 24.280 114.910 ;
        RECT 22.180 112.890 22.440 113.210 ;
        RECT 21.260 112.210 21.520 112.530 ;
        RECT 21.070 111.335 22.610 111.705 ;
        RECT 22.180 110.850 22.440 111.170 ;
        RECT 21.720 110.510 21.980 110.830 ;
        RECT 19.880 109.830 20.140 110.150 ;
        RECT 19.420 109.490 19.680 109.810 ;
        RECT 19.480 108.450 19.620 109.490 ;
        RECT 19.420 108.130 19.680 108.450 ;
        RECT 19.420 107.450 19.680 107.770 ;
        RECT 19.480 106.750 19.620 107.450 ;
        RECT 19.420 106.430 19.680 106.750 ;
        RECT 18.960 105.410 19.220 105.730 ;
        RECT 18.560 103.630 19.160 103.770 ;
        RECT 18.100 102.950 18.700 103.090 ;
        RECT 18.040 102.010 18.300 102.330 ;
        RECT 18.100 100.290 18.240 102.010 ;
        RECT 18.040 99.970 18.300 100.290 ;
        RECT 17.120 98.270 17.380 98.590 ;
        RECT 17.180 97.570 17.320 98.270 ;
        RECT 17.120 97.250 17.380 97.570 ;
        RECT 18.560 97.230 18.700 102.950 ;
        RECT 18.500 96.910 18.760 97.230 ;
        RECT 15.740 95.640 16.400 95.780 ;
        RECT 15.740 95.550 16.000 95.640 ;
        RECT 12.060 91.360 12.320 91.450 ;
        RECT 12.060 91.220 12.720 91.360 ;
        RECT 12.060 91.130 12.320 91.220 ;
        RECT 10.680 90.110 10.940 90.430 ;
        RECT 9.760 89.090 10.020 89.410 ;
        RECT 0.560 88.410 0.820 88.730 ;
        RECT 8.840 87.730 9.100 88.050 ;
        RECT 7.000 87.620 7.260 87.710 ;
        RECT 7.000 87.480 7.660 87.620 ;
        RECT 7.000 87.390 7.260 87.480 ;
        RECT 7.000 85.690 7.260 86.010 ;
        RECT 7.060 83.290 7.200 85.690 ;
        RECT 7.000 82.970 7.260 83.290 ;
        RECT 7.060 80.570 7.200 82.970 ;
        RECT 7.520 82.950 7.660 87.480 ;
        RECT 7.920 87.390 8.180 87.710 ;
        RECT 7.460 82.630 7.720 82.950 ;
        RECT 7.000 80.250 7.260 80.570 ;
        RECT 7.980 75.810 8.120 87.390 ;
        RECT 8.380 80.250 8.640 80.570 ;
        RECT 8.440 78.530 8.580 80.250 ;
        RECT 8.900 78.530 9.040 87.730 ;
        RECT 9.300 87.390 9.560 87.710 ;
        RECT 9.360 86.010 9.500 87.390 ;
        RECT 9.300 85.690 9.560 86.010 ;
        RECT 8.380 78.210 8.640 78.530 ;
        RECT 8.840 78.210 9.100 78.530 ;
        RECT 9.820 77.170 9.960 89.090 ;
        RECT 10.220 80.250 10.480 80.570 ;
        RECT 9.760 77.080 10.020 77.170 ;
        RECT 9.360 76.940 10.020 77.080 ;
        RECT 7.920 75.490 8.180 75.810 ;
        RECT 8.380 65.970 8.640 66.290 ;
        RECT 8.440 64.930 8.580 65.970 ;
        RECT 8.380 64.610 8.640 64.930 ;
        RECT 9.360 64.250 9.500 76.940 ;
        RECT 9.760 76.850 10.020 76.940 ;
        RECT 10.280 75.130 10.420 80.250 ;
        RECT 10.740 75.130 10.880 90.110 ;
        RECT 12.060 88.245 12.320 88.390 ;
        RECT 11.600 87.730 11.860 88.050 ;
        RECT 12.050 87.875 12.330 88.245 ;
        RECT 11.660 83.970 11.800 87.730 ;
        RECT 12.580 87.710 12.720 91.220 ;
        RECT 13.500 88.390 13.640 95.550 ;
        RECT 15.280 91.130 15.540 91.450 ;
        RECT 13.960 89.410 14.560 89.490 ;
        RECT 13.960 89.350 14.620 89.410 ;
        RECT 13.440 88.070 13.700 88.390 ;
        RECT 12.060 87.390 12.320 87.710 ;
        RECT 12.520 87.390 12.780 87.710 ;
        RECT 11.600 83.650 11.860 83.970 ;
        RECT 10.220 74.810 10.480 75.130 ;
        RECT 10.680 74.810 10.940 75.130 ;
        RECT 10.280 69.690 10.420 74.810 ;
        RECT 10.220 69.370 10.480 69.690 ;
        RECT 9.760 68.350 10.020 68.670 ;
        RECT 9.820 64.930 9.960 68.350 ;
        RECT 9.760 64.610 10.020 64.930 ;
        RECT 10.280 64.250 10.420 69.370 ;
        RECT 9.300 63.930 9.560 64.250 ;
        RECT 10.220 63.930 10.480 64.250 ;
        RECT 7.460 60.530 7.720 60.850 ;
        RECT 7.520 59.490 7.660 60.530 ;
        RECT 8.840 60.190 9.100 60.510 ;
        RECT 7.460 59.170 7.720 59.490 ;
        RECT 8.900 56.770 9.040 60.190 ;
        RECT 9.360 59.150 9.500 63.930 ;
        RECT 11.660 63.910 11.800 83.650 ;
        RECT 12.120 75.810 12.260 87.390 ;
        RECT 12.060 75.490 12.320 75.810 ;
        RECT 12.580 75.130 12.720 87.390 ;
        RECT 13.960 85.410 14.100 89.350 ;
        RECT 14.360 89.090 14.620 89.350 ;
        RECT 14.820 88.750 15.080 89.070 ;
        RECT 14.880 86.690 15.020 88.750 ;
        RECT 15.340 88.390 15.480 91.130 ;
        RECT 15.280 88.070 15.540 88.390 ;
        RECT 14.820 86.370 15.080 86.690 ;
        RECT 13.960 85.270 14.560 85.410 ;
        RECT 14.420 82.610 14.560 85.270 ;
        RECT 14.360 82.290 14.620 82.610 ;
        RECT 14.420 80.650 14.560 82.290 ;
        RECT 14.880 81.250 15.020 86.370 ;
        RECT 15.340 82.270 15.480 88.070 ;
        RECT 15.800 87.710 15.940 95.550 ;
        RECT 19.020 91.790 19.160 103.630 ;
        RECT 19.480 101.310 19.620 106.430 ;
        RECT 19.940 102.670 20.080 109.830 ;
        RECT 21.780 107.770 21.920 110.510 ;
        RECT 22.240 107.770 22.380 110.850 ;
        RECT 23.160 110.490 23.300 114.590 ;
        RECT 23.560 112.890 23.820 113.210 ;
        RECT 23.620 112.530 23.760 112.890 ;
        RECT 23.560 112.210 23.820 112.530 ;
        RECT 23.100 110.170 23.360 110.490 ;
        RECT 23.620 109.810 23.760 112.210 ;
        RECT 24.080 110.150 24.220 114.590 ;
        RECT 24.370 114.055 25.910 114.425 ;
        RECT 24.940 112.550 25.200 112.870 ;
        RECT 24.480 111.870 24.740 112.190 ;
        RECT 24.020 109.830 24.280 110.150 ;
        RECT 23.560 109.490 23.820 109.810 ;
        RECT 23.100 109.150 23.360 109.470 ;
        RECT 24.540 109.380 24.680 111.870 ;
        RECT 25.000 111.170 25.140 112.550 ;
        RECT 25.400 112.210 25.660 112.530 ;
        RECT 24.940 110.850 25.200 111.170 ;
        RECT 25.460 110.830 25.600 112.210 ;
        RECT 25.400 110.510 25.660 110.830 ;
        RECT 24.080 109.240 24.680 109.380 ;
        RECT 21.720 107.450 21.980 107.770 ;
        RECT 22.180 107.450 22.440 107.770 ;
        RECT 21.070 105.895 22.610 106.265 ;
        RECT 21.720 104.390 21.980 104.710 ;
        RECT 22.640 104.390 22.900 104.710 ;
        RECT 20.790 102.835 21.070 103.205 ;
        RECT 21.780 103.010 21.920 104.390 ;
        RECT 19.880 102.350 20.140 102.670 ;
        RECT 19.420 100.990 19.680 101.310 ;
        RECT 19.940 97.230 20.080 102.350 ;
        RECT 20.860 102.330 21.000 102.835 ;
        RECT 21.720 102.690 21.980 103.010 ;
        RECT 20.800 102.010 21.060 102.330 ;
        RECT 20.340 101.670 20.600 101.990 ;
        RECT 22.700 101.730 22.840 104.390 ;
        RECT 23.160 102.330 23.300 109.150 ;
        RECT 23.560 106.430 23.820 106.750 ;
        RECT 23.100 102.010 23.360 102.330 ;
        RECT 20.400 100.200 20.540 101.670 ;
        RECT 22.700 101.590 23.300 101.730 ;
        RECT 21.070 100.455 22.610 100.825 ;
        RECT 20.800 100.200 21.060 100.290 ;
        RECT 20.400 100.060 21.060 100.200 ;
        RECT 20.800 99.970 21.060 100.060 ;
        RECT 21.720 99.970 21.980 100.290 ;
        RECT 22.640 99.970 22.900 100.290 ;
        RECT 21.260 98.950 21.520 99.270 ;
        RECT 20.800 98.610 21.060 98.930 ;
        RECT 20.860 97.570 21.000 98.610 ;
        RECT 20.800 97.250 21.060 97.570 ;
        RECT 19.880 96.910 20.140 97.230 ;
        RECT 21.320 96.890 21.460 98.950 ;
        RECT 21.780 98.590 21.920 99.970 ;
        RECT 22.180 98.950 22.440 99.270 ;
        RECT 21.720 98.270 21.980 98.590 ;
        RECT 20.340 96.570 20.600 96.890 ;
        RECT 21.260 96.570 21.520 96.890 ;
        RECT 19.880 95.890 20.140 96.210 ;
        RECT 19.940 92.130 20.080 95.890 ;
        RECT 20.400 94.760 20.540 96.570 ;
        RECT 21.320 96.405 21.460 96.570 ;
        RECT 21.250 96.035 21.530 96.405 ;
        RECT 21.780 95.870 21.920 98.270 ;
        RECT 22.240 96.550 22.380 98.950 ;
        RECT 22.180 96.230 22.440 96.550 ;
        RECT 22.700 96.210 22.840 99.970 ;
        RECT 22.640 95.890 22.900 96.210 ;
        RECT 21.720 95.550 21.980 95.870 ;
        RECT 21.070 95.015 22.610 95.385 ;
        RECT 20.400 94.620 21.000 94.760 ;
        RECT 19.880 91.810 20.140 92.130 ;
        RECT 20.860 91.790 21.000 94.620 ;
        RECT 16.200 91.470 16.460 91.790 ;
        RECT 18.960 91.470 19.220 91.790 ;
        RECT 20.800 91.470 21.060 91.790 ;
        RECT 15.740 87.390 16.000 87.710 ;
        RECT 15.730 85.835 16.010 86.205 ;
        RECT 15.740 85.690 16.000 85.835 ;
        RECT 15.280 81.950 15.540 82.270 ;
        RECT 14.820 80.930 15.080 81.250 ;
        RECT 14.420 80.510 15.020 80.650 ;
        RECT 13.900 79.570 14.160 79.890 ;
        RECT 13.440 78.210 13.700 78.530 ;
        RECT 13.500 78.045 13.640 78.210 ;
        RECT 13.430 77.675 13.710 78.045 ;
        RECT 13.960 77.850 14.100 79.570 ;
        RECT 14.880 79.550 15.020 80.510 ;
        RECT 15.340 80.480 15.480 81.950 ;
        RECT 15.740 80.480 16.000 80.570 ;
        RECT 15.340 80.340 16.000 80.480 ;
        RECT 14.820 79.230 15.080 79.550 ;
        RECT 14.350 78.355 14.630 78.725 ;
        RECT 13.900 77.530 14.160 77.850 ;
        RECT 14.420 77.510 14.560 78.355 ;
        RECT 14.360 77.190 14.620 77.510 ;
        RECT 12.520 74.810 12.780 75.130 ;
        RECT 14.360 70.050 14.620 70.370 ;
        RECT 12.060 69.030 12.320 69.350 ;
        RECT 12.120 67.310 12.260 69.030 ;
        RECT 12.060 66.990 12.320 67.310 ;
        RECT 12.120 64.590 12.260 66.990 ;
        RECT 14.420 66.630 14.560 70.050 ;
        RECT 14.360 66.540 14.620 66.630 ;
        RECT 13.960 66.400 14.620 66.540 ;
        RECT 12.060 64.330 12.320 64.590 ;
        RECT 12.060 64.270 13.640 64.330 ;
        RECT 12.120 64.190 13.640 64.270 ;
        RECT 11.600 63.590 11.860 63.910 ;
        RECT 12.520 63.590 12.780 63.910 ;
        RECT 12.580 61.190 12.720 63.590 ;
        RECT 12.980 63.250 13.240 63.570 ;
        RECT 12.520 60.870 12.780 61.190 ;
        RECT 11.140 60.190 11.400 60.510 ;
        RECT 11.600 60.190 11.860 60.510 ;
        RECT 11.200 59.490 11.340 60.190 ;
        RECT 11.140 59.170 11.400 59.490 ;
        RECT 9.300 58.830 9.560 59.150 ;
        RECT 8.840 56.450 9.100 56.770 ;
        RECT 8.380 55.090 8.640 55.410 ;
        RECT 8.440 54.050 8.580 55.090 ;
        RECT 8.380 53.730 8.640 54.050 ;
        RECT 9.360 52.350 9.500 58.830 ;
        RECT 11.200 55.410 11.340 59.170 ;
        RECT 11.140 55.090 11.400 55.410 ;
        RECT 10.220 54.750 10.480 55.070 ;
        RECT 10.280 53.710 10.420 54.750 ;
        RECT 10.220 53.390 10.480 53.710 ;
        RECT 9.300 52.030 9.560 52.350 ;
        RECT 9.360 45.890 9.500 52.030 ;
        RECT 9.300 45.570 9.560 45.890 ;
        RECT 7.920 45.230 8.180 45.550 ;
        RECT 7.460 44.210 7.720 44.530 ;
        RECT 7.520 37.390 7.660 44.210 ;
        RECT 7.460 37.070 7.720 37.390 ;
        RECT 7.980 37.050 8.120 45.230 ;
        RECT 8.840 43.870 9.100 44.190 ;
        RECT 8.380 39.110 8.640 39.430 ;
        RECT 8.900 39.340 9.040 43.870 ;
        RECT 9.360 39.850 9.500 45.570 ;
        RECT 10.280 44.530 10.420 53.390 ;
        RECT 11.660 53.370 11.800 60.190 ;
        RECT 13.040 55.070 13.180 63.250 ;
        RECT 13.500 61.530 13.640 64.190 ;
        RECT 13.960 63.910 14.100 66.400 ;
        RECT 14.360 66.310 14.620 66.400 ;
        RECT 14.360 65.630 14.620 65.950 ;
        RECT 14.420 64.590 14.560 65.630 ;
        RECT 14.360 64.270 14.620 64.590 ;
        RECT 13.900 63.820 14.160 63.910 ;
        RECT 13.900 63.680 14.560 63.820 ;
        RECT 13.900 63.590 14.160 63.680 ;
        RECT 13.440 61.210 13.700 61.530 ;
        RECT 13.900 60.530 14.160 60.850 ;
        RECT 13.960 56.770 14.100 60.530 ;
        RECT 14.420 60.365 14.560 63.680 ;
        RECT 14.350 59.995 14.630 60.365 ;
        RECT 14.360 59.170 14.620 59.490 ;
        RECT 14.420 57.530 14.560 59.170 ;
        RECT 14.880 58.210 15.020 79.230 ;
        RECT 15.340 78.190 15.480 80.340 ;
        RECT 15.740 80.250 16.000 80.340 ;
        RECT 16.260 78.440 16.400 91.470 ;
        RECT 21.070 89.575 22.610 89.945 ;
        RECT 23.160 89.410 23.300 101.590 ;
        RECT 23.620 99.610 23.760 106.430 ;
        RECT 24.080 105.390 24.220 109.240 ;
        RECT 24.370 108.615 25.910 108.985 ;
        RECT 26.380 108.450 26.520 120.460 ;
        RECT 27.300 120.350 27.440 120.630 ;
        RECT 27.700 120.370 27.960 120.690 ;
        RECT 26.780 120.030 27.040 120.350 ;
        RECT 27.240 120.030 27.500 120.350 ;
        RECT 26.840 118.650 26.980 120.030 ;
        RECT 26.780 118.330 27.040 118.650 ;
        RECT 26.780 114.590 27.040 114.910 ;
        RECT 26.840 112.530 26.980 114.590 ;
        RECT 27.300 113.550 27.440 120.030 ;
        RECT 27.240 113.230 27.500 113.550 ;
        RECT 26.780 112.210 27.040 112.530 ;
        RECT 27.300 111.930 27.440 113.230 ;
        RECT 27.760 112.870 27.900 120.370 ;
        RECT 28.220 118.990 28.360 123.770 ;
        RECT 29.080 123.090 29.340 123.410 ;
        RECT 28.160 118.670 28.420 118.990 ;
        RECT 29.140 113.210 29.280 123.090 ;
        RECT 29.600 121.370 29.740 130.910 ;
        RECT 30.520 129.870 30.660 131.680 ;
        RECT 31.380 131.590 31.640 131.910 ;
        RECT 30.460 129.550 30.720 129.870 ;
        RECT 29.540 121.050 29.800 121.370 ;
        RECT 30.520 120.690 30.660 129.550 ;
        RECT 32.760 128.870 33.020 129.190 ;
        RECT 32.820 127.490 32.960 128.870 ;
        RECT 32.760 127.170 33.020 127.490 ;
        RECT 34.200 127.150 34.340 142.470 ;
        RECT 35.060 140.430 35.320 140.750 ;
        RECT 37.420 140.490 37.560 150.550 ;
        RECT 38.340 143.130 38.480 156.070 ;
        RECT 40.180 154.690 40.320 156.070 ;
        RECT 40.120 154.370 40.380 154.690 ;
        RECT 42.020 153.670 42.160 158.710 ;
        RECT 44.260 158.450 44.520 158.770 ;
        RECT 42.420 158.110 42.680 158.430 ;
        RECT 42.480 156.730 42.620 158.110 ;
        RECT 42.420 156.410 42.680 156.730 ;
        RECT 42.420 154.030 42.680 154.350 ;
        RECT 42.480 153.670 42.620 154.030 ;
        RECT 44.320 153.670 44.460 158.450 ;
        RECT 47.080 155.710 47.220 158.790 ;
        RECT 48.460 156.730 48.600 158.790 ;
        RECT 52.140 158.770 52.280 163.550 ;
        RECT 52.140 158.630 52.740 158.770 ;
        RECT 48.400 156.410 48.660 156.730 ;
        RECT 49.780 156.410 50.040 156.730 ;
        RECT 47.020 155.390 47.280 155.710 ;
        RECT 41.960 153.350 42.220 153.670 ;
        RECT 42.420 153.350 42.680 153.670 ;
        RECT 44.260 153.350 44.520 153.670 ;
        RECT 45.640 153.350 45.900 153.670 ;
        RECT 46.100 153.350 46.360 153.670 ;
        RECT 40.120 152.670 40.380 152.990 ;
        RECT 40.180 151.630 40.320 152.670 ;
        RECT 40.120 151.310 40.380 151.630 ;
        RECT 39.660 150.970 39.920 151.290 ;
        RECT 38.740 149.950 39.000 150.270 ;
        RECT 38.800 148.570 38.940 149.950 ;
        RECT 39.200 148.930 39.460 149.250 ;
        RECT 38.740 148.250 39.000 148.570 ;
        RECT 38.280 142.810 38.540 143.130 ;
        RECT 37.820 141.790 38.080 142.110 ;
        RECT 34.600 139.070 34.860 139.390 ;
        RECT 34.660 134.970 34.800 139.070 ;
        RECT 35.120 138.370 35.260 140.430 ;
        RECT 35.520 140.090 35.780 140.410 ;
        RECT 36.440 140.090 36.700 140.410 ;
        RECT 36.960 140.350 37.560 140.490 ;
        RECT 35.060 138.050 35.320 138.370 ;
        RECT 35.580 138.030 35.720 140.090 ;
        RECT 35.980 139.750 36.240 140.070 ;
        RECT 35.520 137.710 35.780 138.030 ;
        RECT 35.060 136.350 35.320 136.670 ;
        RECT 34.600 134.650 34.860 134.970 ;
        RECT 34.600 131.250 34.860 131.570 ;
        RECT 34.660 130.210 34.800 131.250 ;
        RECT 34.600 129.890 34.860 130.210 ;
        RECT 35.120 127.490 35.260 136.350 ;
        RECT 35.520 134.990 35.780 135.310 ;
        RECT 35.580 131.910 35.720 134.990 ;
        RECT 35.520 131.590 35.780 131.910 ;
        RECT 36.040 128.850 36.180 139.750 ;
        RECT 36.500 137.010 36.640 140.090 ;
        RECT 36.960 138.370 37.100 140.350 ;
        RECT 36.900 138.050 37.160 138.370 ;
        RECT 36.440 136.690 36.700 137.010 ;
        RECT 36.500 132.930 36.640 136.690 ;
        RECT 36.440 132.610 36.700 132.930 ;
        RECT 35.980 128.530 36.240 128.850 ;
        RECT 35.060 127.170 35.320 127.490 ;
        RECT 34.140 126.830 34.400 127.150 ;
        RECT 33.220 126.490 33.480 126.810 ;
        RECT 30.920 123.090 31.180 123.410 ;
        RECT 31.380 123.090 31.640 123.410 ;
        RECT 30.980 122.050 31.120 123.090 ;
        RECT 30.920 121.730 31.180 122.050 ;
        RECT 30.460 120.370 30.720 120.690 ;
        RECT 29.540 117.310 29.800 117.630 ;
        RECT 29.080 112.890 29.340 113.210 ;
        RECT 27.700 112.550 27.960 112.870 ;
        RECT 26.840 111.790 27.440 111.930 ;
        RECT 28.160 111.870 28.420 112.190 ;
        RECT 26.840 108.450 26.980 111.790 ;
        RECT 27.240 109.830 27.500 110.150 ;
        RECT 26.320 108.130 26.580 108.450 ;
        RECT 26.780 108.130 27.040 108.450 ;
        RECT 24.940 107.790 25.200 108.110 ;
        RECT 24.480 107.450 24.740 107.770 ;
        RECT 24.020 105.070 24.280 105.390 ;
        RECT 24.540 104.710 24.680 107.450 ;
        RECT 25.000 105.390 25.140 107.790 ;
        RECT 25.400 107.110 25.660 107.430 ;
        RECT 24.940 105.070 25.200 105.390 ;
        RECT 25.460 105.050 25.600 107.110 ;
        RECT 26.380 107.090 26.520 108.130 ;
        RECT 26.320 106.770 26.580 107.090 ;
        RECT 25.400 104.730 25.660 105.050 ;
        RECT 26.380 104.710 26.520 106.770 ;
        RECT 24.480 104.390 24.740 104.710 ;
        RECT 26.320 104.390 26.580 104.710 ;
        RECT 26.840 104.370 26.980 108.130 ;
        RECT 26.780 104.050 27.040 104.370 ;
        RECT 24.020 103.710 24.280 104.030 ;
        RECT 24.080 100.290 24.220 103.710 ;
        RECT 24.370 103.175 25.910 103.545 ;
        RECT 26.320 101.670 26.580 101.990 ;
        RECT 24.480 101.330 24.740 101.650 ;
        RECT 24.020 99.970 24.280 100.290 ;
        RECT 23.560 99.290 23.820 99.610 ;
        RECT 23.620 96.890 23.760 99.290 ;
        RECT 24.540 99.270 24.680 101.330 ;
        RECT 25.860 99.290 26.120 99.610 ;
        RECT 24.480 98.950 24.740 99.270 ;
        RECT 25.920 99.125 26.060 99.290 ;
        RECT 25.850 98.755 26.130 99.125 ;
        RECT 24.370 97.735 25.910 98.105 ;
        RECT 26.380 97.570 26.520 101.670 ;
        RECT 27.300 99.270 27.440 109.830 ;
        RECT 28.220 108.110 28.360 111.870 ;
        RECT 29.140 110.490 29.280 112.890 ;
        RECT 29.080 110.170 29.340 110.490 ;
        RECT 28.160 107.790 28.420 108.110 ;
        RECT 29.080 107.790 29.340 108.110 ;
        RECT 29.140 107.170 29.280 107.790 ;
        RECT 29.600 107.770 29.740 117.310 ;
        RECT 29.540 107.450 29.800 107.770 ;
        RECT 29.140 107.030 29.740 107.170 ;
        RECT 28.160 106.430 28.420 106.750 ;
        RECT 29.080 106.430 29.340 106.750 ;
        RECT 28.220 99.270 28.360 106.430 ;
        RECT 26.770 98.755 27.050 99.125 ;
        RECT 27.240 98.950 27.500 99.270 ;
        RECT 28.160 98.950 28.420 99.270 ;
        RECT 29.140 98.930 29.280 106.430 ;
        RECT 29.600 105.810 29.740 107.030 ;
        RECT 29.600 105.670 30.200 105.810 ;
        RECT 24.020 97.250 24.280 97.570 ;
        RECT 26.320 97.250 26.580 97.570 ;
        RECT 23.560 96.570 23.820 96.890 ;
        RECT 23.560 95.550 23.820 95.870 ;
        RECT 16.660 89.090 16.920 89.410 ;
        RECT 23.100 89.090 23.360 89.410 ;
        RECT 16.720 88.390 16.860 89.090 ;
        RECT 17.180 88.670 18.240 88.810 ;
        RECT 18.960 88.750 19.220 89.070 ;
        RECT 17.180 88.390 17.320 88.670 ;
        RECT 16.660 88.070 16.920 88.390 ;
        RECT 17.120 88.070 17.380 88.390 ;
        RECT 16.720 82.270 16.860 88.070 ;
        RECT 17.580 87.730 17.840 88.050 ;
        RECT 17.120 87.390 17.380 87.710 ;
        RECT 16.660 81.950 16.920 82.270 ;
        RECT 16.720 80.910 16.860 81.950 ;
        RECT 16.660 80.590 16.920 80.910 ;
        RECT 15.800 78.300 16.400 78.440 ;
        RECT 15.280 77.870 15.540 78.190 ;
        RECT 15.800 77.365 15.940 78.300 ;
        RECT 16.190 77.675 16.470 78.045 ;
        RECT 15.730 76.995 16.010 77.365 ;
        RECT 15.800 76.830 15.940 76.995 ;
        RECT 15.740 76.510 16.000 76.830 ;
        RECT 15.800 70.370 15.940 76.510 ;
        RECT 16.260 71.300 16.400 77.675 ;
        RECT 16.660 77.530 16.920 77.850 ;
        RECT 16.720 72.070 16.860 77.530 ;
        RECT 17.180 77.510 17.320 87.390 ;
        RECT 17.640 86.010 17.780 87.730 ;
        RECT 17.580 85.690 17.840 86.010 ;
        RECT 17.580 81.950 17.840 82.270 ;
        RECT 17.640 81.250 17.780 81.950 ;
        RECT 17.580 80.930 17.840 81.250 ;
        RECT 18.100 80.570 18.240 88.670 ;
        RECT 19.020 88.390 19.160 88.750 ;
        RECT 18.960 88.070 19.220 88.390 ;
        RECT 19.420 88.245 19.680 88.390 ;
        RECT 19.410 87.875 19.690 88.245 ;
        RECT 18.500 85.690 18.760 86.010 ;
        RECT 18.560 83.970 18.700 85.690 ;
        RECT 18.960 84.670 19.220 84.990 ;
        RECT 18.500 83.650 18.760 83.970 ;
        RECT 19.020 82.950 19.160 84.670 ;
        RECT 18.960 82.630 19.220 82.950 ;
        RECT 18.040 80.250 18.300 80.570 ;
        RECT 18.100 79.890 18.240 80.250 ;
        RECT 19.480 80.140 19.620 87.875 ;
        RECT 20.340 87.730 20.600 88.050 ;
        RECT 20.400 84.990 20.540 87.730 ;
        RECT 20.340 84.670 20.600 84.990 ;
        RECT 20.400 82.950 20.540 84.670 ;
        RECT 21.070 84.135 22.610 84.505 ;
        RECT 23.160 82.950 23.300 89.090 ;
        RECT 23.620 83.290 23.760 95.550 ;
        RECT 23.560 82.970 23.820 83.290 ;
        RECT 20.340 82.630 20.600 82.950 ;
        RECT 21.260 82.630 21.520 82.950 ;
        RECT 23.100 82.630 23.360 82.950 ;
        RECT 19.880 82.290 20.140 82.610 ;
        RECT 19.940 81.250 20.080 82.290 ;
        RECT 19.880 80.930 20.140 81.250 ;
        RECT 20.400 80.570 20.540 82.630 ;
        RECT 20.800 81.950 21.060 82.270 ;
        RECT 20.340 80.250 20.600 80.570 ;
        RECT 19.880 80.140 20.140 80.230 ;
        RECT 19.480 80.000 20.140 80.140 ;
        RECT 18.040 79.570 18.300 79.890 ;
        RECT 18.100 78.190 18.240 79.570 ;
        RECT 19.480 78.530 19.620 80.000 ;
        RECT 19.880 79.910 20.140 80.000 ;
        RECT 20.860 79.970 21.000 81.950 ;
        RECT 21.320 80.570 21.460 82.630 ;
        RECT 23.560 82.290 23.820 82.610 ;
        RECT 22.640 81.950 22.900 82.270 ;
        RECT 21.260 80.250 21.520 80.570 ;
        RECT 21.720 80.250 21.980 80.570 ;
        RECT 20.400 79.830 21.000 79.970 ;
        RECT 21.780 79.890 21.920 80.250 ;
        RECT 19.420 78.210 19.680 78.530 ;
        RECT 20.400 78.440 20.540 79.830 ;
        RECT 21.720 79.570 21.980 79.890 ;
        RECT 22.700 79.550 22.840 81.950 ;
        RECT 23.100 80.930 23.360 81.250 ;
        RECT 22.640 79.230 22.900 79.550 ;
        RECT 23.160 79.290 23.300 80.930 ;
        RECT 23.620 80.570 23.760 82.290 ;
        RECT 23.560 80.250 23.820 80.570 ;
        RECT 23.160 79.150 23.760 79.290 ;
        RECT 21.070 78.695 22.610 79.065 ;
        RECT 20.400 78.300 21.000 78.440 ;
        RECT 18.040 77.870 18.300 78.190 ;
        RECT 19.480 77.510 19.620 78.210 ;
        RECT 17.120 77.190 17.380 77.510 ;
        RECT 19.420 77.190 19.680 77.510 ;
        RECT 20.340 77.365 20.600 77.510 ;
        RECT 18.500 76.850 18.760 77.170 ;
        RECT 20.330 76.995 20.610 77.365 ;
        RECT 18.560 75.810 18.700 76.850 ;
        RECT 19.420 76.510 19.680 76.830 ;
        RECT 19.880 76.510 20.140 76.830 ;
        RECT 18.500 75.490 18.760 75.810 ;
        RECT 16.660 71.750 16.920 72.070 ;
        RECT 16.260 71.160 16.860 71.300 ;
        RECT 15.740 70.050 16.000 70.370 ;
        RECT 15.740 66.990 16.000 67.310 ;
        RECT 15.280 66.310 15.540 66.630 ;
        RECT 15.340 61.870 15.480 66.310 ;
        RECT 15.800 64.250 15.940 66.990 ;
        RECT 16.200 65.970 16.460 66.290 ;
        RECT 15.740 63.930 16.000 64.250 ;
        RECT 15.740 62.910 16.000 63.230 ;
        RECT 15.280 61.550 15.540 61.870 ;
        RECT 15.800 60.510 15.940 62.910 ;
        RECT 16.260 62.210 16.400 65.970 ;
        RECT 16.200 61.890 16.460 62.210 ;
        RECT 15.740 60.190 16.000 60.510 ;
        RECT 16.720 59.570 16.860 71.160 ;
        RECT 17.120 71.070 17.380 71.390 ;
        RECT 17.180 67.165 17.320 71.070 ;
        RECT 18.030 69.515 18.310 69.885 ;
        RECT 18.960 69.710 19.220 70.030 ;
        RECT 18.040 69.370 18.300 69.515 ;
        RECT 18.040 68.920 18.300 69.010 ;
        RECT 17.640 68.780 18.300 68.920 ;
        RECT 17.110 66.795 17.390 67.165 ;
        RECT 17.640 66.370 17.780 68.780 ;
        RECT 18.040 68.690 18.300 68.780 ;
        RECT 18.030 68.155 18.310 68.525 ;
        RECT 18.500 68.350 18.760 68.670 ;
        RECT 18.100 66.630 18.240 68.155 ;
        RECT 17.180 66.290 17.780 66.370 ;
        RECT 18.040 66.310 18.300 66.630 ;
        RECT 17.120 66.230 17.780 66.290 ;
        RECT 17.120 65.970 17.380 66.230 ;
        RECT 17.580 65.630 17.840 65.950 ;
        RECT 17.120 63.140 17.380 63.230 ;
        RECT 17.640 63.140 17.780 65.630 ;
        RECT 18.100 63.650 18.240 66.310 ;
        RECT 18.560 64.250 18.700 68.350 ;
        RECT 19.020 64.930 19.160 69.710 ;
        RECT 19.480 67.165 19.620 76.510 ;
        RECT 19.940 68.670 20.080 76.510 ;
        RECT 20.860 74.360 21.000 78.300 ;
        RECT 23.100 78.210 23.360 78.530 ;
        RECT 20.400 74.220 21.000 74.360 ;
        RECT 20.400 72.410 20.540 74.220 ;
        RECT 21.070 73.255 22.610 73.625 ;
        RECT 20.340 72.090 20.600 72.410 ;
        RECT 20.400 69.350 20.540 72.090 ;
        RECT 23.160 72.070 23.300 78.210 ;
        RECT 23.620 75.130 23.760 79.150 ;
        RECT 24.080 78.530 24.220 97.250 ;
        RECT 25.850 96.715 26.130 97.085 ;
        RECT 25.860 96.570 26.120 96.715 ;
        RECT 24.370 92.295 25.910 92.665 ;
        RECT 24.940 91.130 25.200 91.450 ;
        RECT 25.860 91.130 26.120 91.450 ;
        RECT 25.000 88.390 25.140 91.130 ;
        RECT 25.920 88.390 26.060 91.130 ;
        RECT 26.840 89.410 26.980 98.755 ;
        RECT 29.080 98.610 29.340 98.930 ;
        RECT 29.140 96.890 29.280 98.610 ;
        RECT 29.540 98.270 29.800 98.590 ;
        RECT 29.600 97.230 29.740 98.270 ;
        RECT 29.540 96.910 29.800 97.230 ;
        RECT 30.060 97.085 30.200 105.670 ;
        RECT 30.520 101.990 30.660 120.370 ;
        RECT 31.440 120.350 31.580 123.090 ;
        RECT 30.920 120.030 31.180 120.350 ;
        RECT 31.380 120.030 31.640 120.350 ;
        RECT 30.980 115.590 31.120 120.030 ;
        RECT 31.440 117.630 31.580 120.030 ;
        RECT 31.380 117.310 31.640 117.630 ;
        RECT 30.920 115.270 31.180 115.590 ;
        RECT 31.840 115.270 32.100 115.590 ;
        RECT 31.380 112.550 31.640 112.870 ;
        RECT 30.920 112.210 31.180 112.530 ;
        RECT 30.980 108.110 31.120 112.210 ;
        RECT 30.920 107.790 31.180 108.110 ;
        RECT 31.440 105.390 31.580 112.550 ;
        RECT 31.900 110.830 32.040 115.270 ;
        RECT 32.300 112.890 32.560 113.210 ;
        RECT 31.840 110.510 32.100 110.830 ;
        RECT 31.900 110.150 32.040 110.510 ;
        RECT 31.840 109.830 32.100 110.150 ;
        RECT 31.900 105.390 32.040 109.830 ;
        RECT 31.380 105.070 31.640 105.390 ;
        RECT 31.840 105.070 32.100 105.390 ;
        RECT 30.460 101.670 30.720 101.990 ;
        RECT 31.440 100.290 31.580 105.070 ;
        RECT 32.360 104.710 32.500 112.890 ;
        RECT 33.280 107.770 33.420 126.490 ;
        RECT 36.040 126.470 36.180 128.530 ;
        RECT 35.980 126.150 36.240 126.470 ;
        RECT 35.520 123.770 35.780 124.090 ;
        RECT 35.580 122.050 35.720 123.770 ;
        RECT 35.520 121.730 35.780 122.050 ;
        RECT 36.960 121.370 37.100 138.050 ;
        RECT 37.360 133.630 37.620 133.950 ;
        RECT 36.900 121.050 37.160 121.370 ;
        RECT 34.600 114.590 34.860 114.910 ;
        RECT 34.140 109.830 34.400 110.150 ;
        RECT 33.680 109.150 33.940 109.470 ;
        RECT 33.220 107.450 33.480 107.770 ;
        RECT 32.760 106.430 33.020 106.750 ;
        RECT 32.300 104.390 32.560 104.710 ;
        RECT 32.360 103.010 32.500 104.390 ;
        RECT 32.300 102.690 32.560 103.010 ;
        RECT 31.380 99.970 31.640 100.290 ;
        RECT 32.360 97.570 32.500 102.690 ;
        RECT 32.300 97.250 32.560 97.570 ;
        RECT 29.080 96.570 29.340 96.890 ;
        RECT 29.990 96.715 30.270 97.085 ;
        RECT 32.820 95.870 32.960 106.430 ;
        RECT 33.280 101.650 33.420 107.450 ;
        RECT 33.740 105.050 33.880 109.150 ;
        RECT 34.200 108.110 34.340 109.830 ;
        RECT 34.140 107.790 34.400 108.110 ;
        RECT 34.660 107.770 34.800 114.590 ;
        RECT 35.060 109.490 35.320 109.810 ;
        RECT 35.120 108.110 35.260 109.490 ;
        RECT 35.060 107.790 35.320 108.110 ;
        RECT 34.600 107.450 34.860 107.770 ;
        RECT 36.440 105.410 36.700 105.730 ;
        RECT 33.680 104.730 33.940 105.050 ;
        RECT 36.500 102.670 36.640 105.410 ;
        RECT 36.440 102.350 36.700 102.670 ;
        RECT 33.220 101.330 33.480 101.650 ;
        RECT 34.600 96.230 34.860 96.550 ;
        RECT 32.760 95.550 33.020 95.870 ;
        RECT 33.220 95.550 33.480 95.870 ;
        RECT 30.000 92.830 30.260 93.150 ;
        RECT 30.060 91.450 30.200 92.830 ;
        RECT 33.280 91.450 33.420 95.550 ;
        RECT 34.660 93.830 34.800 96.230 ;
        RECT 34.600 93.510 34.860 93.830 ;
        RECT 34.660 91.450 34.800 93.510 ;
        RECT 35.060 93.170 35.320 93.490 ;
        RECT 35.120 91.790 35.260 93.170 ;
        RECT 35.520 92.830 35.780 93.150 ;
        RECT 35.060 91.470 35.320 91.790 ;
        RECT 30.000 91.130 30.260 91.450 ;
        RECT 33.220 91.130 33.480 91.450 ;
        RECT 34.600 91.130 34.860 91.450 ;
        RECT 26.780 89.090 27.040 89.410 ;
        RECT 24.940 88.070 25.200 88.390 ;
        RECT 25.860 88.070 26.120 88.390 ;
        RECT 25.920 87.710 26.060 88.070 ;
        RECT 25.860 87.390 26.120 87.710 ;
        RECT 24.370 86.855 25.910 87.225 ;
        RECT 26.840 86.770 26.980 89.090 ;
        RECT 30.460 87.390 30.720 87.710 ;
        RECT 26.840 86.630 27.440 86.770 ;
        RECT 25.400 86.030 25.660 86.350 ;
        RECT 26.780 86.030 27.040 86.350 ;
        RECT 25.460 83.290 25.600 86.030 ;
        RECT 26.320 84.670 26.580 84.990 ;
        RECT 26.380 83.970 26.520 84.670 ;
        RECT 26.320 83.650 26.580 83.970 ;
        RECT 25.400 82.970 25.660 83.290 ;
        RECT 26.320 82.970 26.580 83.290 ;
        RECT 24.370 81.415 25.910 81.785 ;
        RECT 25.400 80.590 25.660 80.910 ;
        RECT 24.940 79.570 25.200 79.890 ;
        RECT 24.480 79.230 24.740 79.550 ;
        RECT 24.020 78.210 24.280 78.530 ;
        RECT 24.540 77.930 24.680 79.230 ;
        RECT 24.080 77.850 24.680 77.930 ;
        RECT 24.020 77.790 24.680 77.850 ;
        RECT 24.020 77.530 24.280 77.790 ;
        RECT 23.560 74.810 23.820 75.130 ;
        RECT 23.560 73.790 23.820 74.110 ;
        RECT 21.720 71.750 21.980 72.070 ;
        RECT 23.100 71.750 23.360 72.070 ;
        RECT 21.260 71.070 21.520 71.390 ;
        RECT 21.320 69.690 21.460 71.070 ;
        RECT 21.260 69.370 21.520 69.690 ;
        RECT 20.340 69.030 20.600 69.350 ;
        RECT 21.780 69.010 21.920 71.750 ;
        RECT 23.100 71.070 23.360 71.390 ;
        RECT 22.180 69.370 22.440 69.690 ;
        RECT 21.720 68.690 21.980 69.010 ;
        RECT 22.240 68.670 22.380 69.370 ;
        RECT 19.880 68.350 20.140 68.670 ;
        RECT 20.340 68.350 20.600 68.670 ;
        RECT 22.180 68.350 22.440 68.670 ;
        RECT 19.410 66.795 19.690 67.165 ;
        RECT 18.960 64.610 19.220 64.930 ;
        RECT 19.940 64.250 20.080 68.350 ;
        RECT 18.500 63.930 18.760 64.250 ;
        RECT 19.880 63.930 20.140 64.250 ;
        RECT 18.100 63.510 18.700 63.650 ;
        RECT 19.420 63.590 19.680 63.910 ;
        RECT 17.120 63.000 17.780 63.140 ;
        RECT 17.120 62.910 17.380 63.000 ;
        RECT 18.040 62.910 18.300 63.230 ;
        RECT 17.110 61.440 17.390 61.725 ;
        RECT 17.110 61.355 17.780 61.440 ;
        RECT 17.120 61.300 17.780 61.355 ;
        RECT 17.120 61.210 17.380 61.300 ;
        RECT 16.260 59.430 16.860 59.570 ;
        RECT 16.260 59.150 16.400 59.430 ;
        RECT 15.740 58.830 16.000 59.150 ;
        RECT 16.200 58.830 16.460 59.150 ;
        RECT 14.880 58.070 15.480 58.210 ;
        RECT 15.340 57.790 15.480 58.070 ;
        RECT 14.820 57.530 15.080 57.790 ;
        RECT 14.420 57.470 15.080 57.530 ;
        RECT 15.280 57.470 15.540 57.790 ;
        RECT 14.420 57.390 15.020 57.470 ;
        RECT 15.800 56.770 15.940 58.830 ;
        RECT 13.900 56.450 14.160 56.770 ;
        RECT 15.740 56.450 16.000 56.770 ;
        RECT 13.900 55.430 14.160 55.750 ;
        RECT 12.980 54.750 13.240 55.070 ;
        RECT 13.040 53.710 13.180 54.750 ;
        RECT 12.980 53.390 13.240 53.710 ;
        RECT 11.600 53.050 11.860 53.370 ;
        RECT 11.660 45.210 11.800 53.050 ;
        RECT 13.960 50.650 14.100 55.430 ;
        RECT 15.740 55.090 16.000 55.410 ;
        RECT 13.900 50.330 14.160 50.650 ;
        RECT 11.600 44.890 11.860 45.210 ;
        RECT 11.660 44.610 11.800 44.890 ;
        RECT 10.220 44.440 10.480 44.530 ;
        RECT 11.660 44.470 12.260 44.610 ;
        RECT 10.220 44.300 11.340 44.440 ;
        RECT 10.220 44.210 10.480 44.300 ;
        RECT 9.360 39.710 9.960 39.850 ;
        RECT 9.300 39.340 9.560 39.430 ;
        RECT 8.900 39.200 9.560 39.340 ;
        RECT 9.300 39.110 9.560 39.200 ;
        RECT 8.440 37.050 8.580 39.110 ;
        RECT 7.920 36.730 8.180 37.050 ;
        RECT 8.380 36.730 8.640 37.050 ;
        RECT 9.820 36.030 9.960 39.710 ;
        RECT 11.200 37.050 11.340 44.300 ;
        RECT 11.600 43.870 11.860 44.190 ;
        RECT 11.660 43.170 11.800 43.870 ;
        RECT 11.600 42.850 11.860 43.170 ;
        RECT 12.120 42.830 12.260 44.470 ;
        RECT 12.060 42.510 12.320 42.830 ;
        RECT 12.120 39.090 12.260 42.510 ;
        RECT 13.960 42.490 14.100 50.330 ;
        RECT 14.820 47.270 15.080 47.590 ;
        RECT 14.880 44.530 15.020 47.270 ;
        RECT 15.800 44.870 15.940 55.090 ;
        RECT 16.260 54.050 16.400 58.830 ;
        RECT 17.640 58.810 17.780 61.300 ;
        RECT 17.120 58.490 17.380 58.810 ;
        RECT 17.580 58.490 17.840 58.810 ;
        RECT 17.180 57.790 17.320 58.490 ;
        RECT 17.120 57.470 17.380 57.790 ;
        RECT 17.580 57.470 17.840 57.790 ;
        RECT 16.200 53.730 16.460 54.050 ;
        RECT 16.260 51.330 16.400 53.730 ;
        RECT 17.180 52.690 17.320 57.470 ;
        RECT 17.640 53.370 17.780 57.470 ;
        RECT 17.580 53.050 17.840 53.370 ;
        RECT 17.120 52.370 17.380 52.690 ;
        RECT 16.200 51.010 16.460 51.330 ;
        RECT 18.100 50.310 18.240 62.910 ;
        RECT 16.660 49.990 16.920 50.310 ;
        RECT 18.040 49.990 18.300 50.310 ;
        RECT 16.720 48.610 16.860 49.990 ;
        RECT 16.660 48.290 16.920 48.610 ;
        RECT 16.660 47.610 16.920 47.930 ;
        RECT 15.740 44.550 16.000 44.870 ;
        RECT 14.820 44.210 15.080 44.530 ;
        RECT 14.360 43.870 14.620 44.190 ;
        RECT 14.420 42.830 14.560 43.870 ;
        RECT 14.360 42.510 14.620 42.830 ;
        RECT 12.520 42.170 12.780 42.490 ;
        RECT 13.900 42.170 14.160 42.490 ;
        RECT 12.060 38.770 12.320 39.090 ;
        RECT 11.140 36.730 11.400 37.050 ;
        RECT 9.760 35.710 10.020 36.030 ;
        RECT 11.200 33.650 11.340 36.730 ;
        RECT 11.600 35.710 11.860 36.030 ;
        RECT 11.660 35.010 11.800 35.710 ;
        RECT 11.600 34.690 11.860 35.010 ;
        RECT 12.120 34.670 12.260 38.770 ;
        RECT 12.060 34.350 12.320 34.670 ;
        RECT 11.600 34.010 11.860 34.330 ;
        RECT 11.660 33.650 11.800 34.010 ;
        RECT 11.140 33.330 11.400 33.650 ;
        RECT 11.600 33.330 11.860 33.650 ;
        RECT 12.580 33.310 12.720 42.170 ;
        RECT 13.960 40.450 14.100 42.170 ;
        RECT 14.420 40.450 14.560 42.510 ;
        RECT 14.820 41.490 15.080 41.810 ;
        RECT 13.900 40.130 14.160 40.450 ;
        RECT 14.360 40.130 14.620 40.450 ;
        RECT 12.980 39.790 13.240 40.110 ;
        RECT 13.040 33.310 13.180 39.790 ;
        RECT 13.960 34.330 14.100 40.130 ;
        RECT 14.360 38.430 14.620 38.750 ;
        RECT 13.900 34.010 14.160 34.330 ;
        RECT 14.420 33.990 14.560 38.430 ;
        RECT 14.880 37.730 15.020 41.490 ;
        RECT 15.800 41.470 15.940 44.550 ;
        RECT 16.720 44.190 16.860 47.610 ;
        RECT 18.040 47.270 18.300 47.590 ;
        RECT 18.100 45.890 18.240 47.270 ;
        RECT 18.040 45.570 18.300 45.890 ;
        RECT 18.560 45.210 18.700 63.510 ;
        RECT 19.480 62.170 19.620 63.590 ;
        RECT 19.020 62.030 19.620 62.170 ;
        RECT 19.020 57.530 19.160 62.030 ;
        RECT 19.420 60.530 19.680 60.850 ;
        RECT 19.480 58.130 19.620 60.530 ;
        RECT 19.880 60.190 20.140 60.510 ;
        RECT 19.940 59.490 20.080 60.190 ;
        RECT 19.880 59.170 20.140 59.490 ;
        RECT 19.880 58.490 20.140 58.810 ;
        RECT 19.420 57.810 19.680 58.130 ;
        RECT 19.940 57.530 20.080 58.490 ;
        RECT 19.020 57.390 20.080 57.530 ;
        RECT 19.020 55.410 19.160 57.390 ;
        RECT 18.960 55.090 19.220 55.410 ;
        RECT 20.400 53.370 20.540 68.350 ;
        RECT 21.070 67.815 22.610 68.185 ;
        RECT 21.260 67.165 21.520 67.310 ;
        RECT 21.250 66.795 21.530 67.165 ;
        RECT 21.260 66.485 21.520 66.630 ;
        RECT 21.250 66.115 21.530 66.485 ;
        RECT 20.800 65.630 21.060 65.950 ;
        RECT 20.860 64.250 21.000 65.630 ;
        RECT 20.800 63.930 21.060 64.250 ;
        RECT 21.070 62.375 22.610 62.745 ;
        RECT 23.160 62.170 23.300 71.070 ;
        RECT 23.620 63.230 23.760 73.790 ;
        RECT 24.080 71.730 24.220 77.530 ;
        RECT 25.000 77.510 25.140 79.570 ;
        RECT 24.480 77.365 24.740 77.510 ;
        RECT 24.470 76.995 24.750 77.365 ;
        RECT 24.940 77.190 25.200 77.510 ;
        RECT 25.460 77.365 25.600 80.590 ;
        RECT 25.850 77.675 26.130 78.045 ;
        RECT 25.920 77.510 26.060 77.675 ;
        RECT 25.390 76.995 25.670 77.365 ;
        RECT 25.860 77.190 26.120 77.510 ;
        RECT 24.370 75.975 25.910 76.345 ;
        RECT 24.480 75.490 24.740 75.810 ;
        RECT 24.540 72.410 24.680 75.490 ;
        RECT 25.860 74.810 26.120 75.130 ;
        RECT 24.480 72.090 24.740 72.410 ;
        RECT 24.020 71.410 24.280 71.730 ;
        RECT 24.080 69.885 24.220 71.410 ;
        RECT 25.920 71.390 26.060 74.810 ;
        RECT 26.380 72.070 26.520 82.970 ;
        RECT 26.840 78.530 26.980 86.030 ;
        RECT 26.780 78.210 27.040 78.530 ;
        RECT 27.300 77.850 27.440 86.630 ;
        RECT 28.160 85.690 28.420 86.010 ;
        RECT 29.540 85.690 29.800 86.010 ;
        RECT 27.700 84.670 27.960 84.990 ;
        RECT 27.760 82.950 27.900 84.670 ;
        RECT 27.700 82.630 27.960 82.950 ;
        RECT 28.220 80.910 28.360 85.690 ;
        RECT 28.620 85.350 28.880 85.670 ;
        RECT 28.680 80.910 28.820 85.350 ;
        RECT 29.080 84.670 29.340 84.990 ;
        RECT 28.160 80.590 28.420 80.910 ;
        RECT 28.620 80.590 28.880 80.910 ;
        RECT 27.700 79.570 27.960 79.890 ;
        RECT 28.620 79.570 28.880 79.890 ;
        RECT 27.240 77.530 27.500 77.850 ;
        RECT 27.240 75.150 27.500 75.470 ;
        RECT 27.300 72.070 27.440 75.150 ;
        RECT 27.760 75.130 27.900 79.570 ;
        RECT 28.160 79.230 28.420 79.550 ;
        RECT 28.220 78.530 28.360 79.230 ;
        RECT 28.160 78.210 28.420 78.530 ;
        RECT 28.220 77.510 28.360 78.210 ;
        RECT 28.160 77.190 28.420 77.510 ;
        RECT 27.700 74.810 27.960 75.130 ;
        RECT 28.220 73.090 28.360 77.190 ;
        RECT 28.680 75.810 28.820 79.570 ;
        RECT 29.140 79.550 29.280 84.670 ;
        RECT 29.600 83.970 29.740 85.690 ;
        RECT 29.540 83.650 29.800 83.970 ;
        RECT 29.600 81.250 29.740 83.650 ;
        RECT 30.000 82.290 30.260 82.610 ;
        RECT 30.060 81.250 30.200 82.290 ;
        RECT 29.540 80.930 29.800 81.250 ;
        RECT 30.000 80.930 30.260 81.250 ;
        RECT 29.080 79.230 29.340 79.550 ;
        RECT 29.600 77.510 29.740 80.930 ;
        RECT 29.540 77.190 29.800 77.510 ;
        RECT 29.080 76.850 29.340 77.170 ;
        RECT 29.140 76.685 29.280 76.850 ;
        RECT 29.070 76.315 29.350 76.685 ;
        RECT 28.620 75.720 28.880 75.810 ;
        RECT 28.620 75.580 29.740 75.720 ;
        RECT 28.620 75.490 28.880 75.580 ;
        RECT 28.160 72.770 28.420 73.090 ;
        RECT 26.320 71.750 26.580 72.070 ;
        RECT 27.240 71.750 27.500 72.070 ;
        RECT 25.860 71.070 26.120 71.390 ;
        RECT 24.370 70.535 25.910 70.905 ;
        RECT 25.860 70.050 26.120 70.370 ;
        RECT 24.010 69.515 24.290 69.885 ;
        RECT 25.920 69.690 26.060 70.050 ;
        RECT 25.860 69.370 26.120 69.690 ;
        RECT 24.480 68.690 24.740 69.010 ;
        RECT 24.020 67.330 24.280 67.650 ;
        RECT 23.560 62.910 23.820 63.230 ;
        RECT 23.160 62.030 23.760 62.170 ;
        RECT 23.100 60.870 23.360 61.190 ;
        RECT 20.790 59.995 21.070 60.365 ;
        RECT 22.180 60.190 22.440 60.510 ;
        RECT 20.860 58.810 21.000 59.995 ;
        RECT 22.240 59.490 22.380 60.190 ;
        RECT 22.180 59.170 22.440 59.490 ;
        RECT 20.800 58.490 21.060 58.810 ;
        RECT 23.160 58.210 23.300 60.870 ;
        RECT 23.620 58.810 23.760 62.030 ;
        RECT 24.080 61.190 24.220 67.330 ;
        RECT 24.540 66.970 24.680 68.690 ;
        RECT 24.480 66.650 24.740 66.970 ;
        RECT 25.920 66.370 26.060 69.370 ;
        RECT 26.380 67.650 26.520 71.750 ;
        RECT 27.300 70.370 27.440 71.750 ;
        RECT 27.700 71.070 27.960 71.390 ;
        RECT 28.160 71.070 28.420 71.390 ;
        RECT 27.240 70.050 27.500 70.370 ;
        RECT 26.780 68.350 27.040 68.670 ;
        RECT 26.320 67.330 26.580 67.650 ;
        RECT 26.380 66.970 26.520 67.330 ;
        RECT 26.320 66.650 26.580 66.970 ;
        RECT 25.920 66.230 26.520 66.370 ;
        RECT 24.370 65.095 25.910 65.465 ;
        RECT 24.470 64.075 24.750 64.445 ;
        RECT 24.540 63.570 24.680 64.075 ;
        RECT 24.940 63.930 25.200 64.250 ;
        RECT 24.480 63.250 24.740 63.570 ;
        RECT 24.020 60.870 24.280 61.190 ;
        RECT 24.080 59.150 24.220 60.870 ;
        RECT 24.540 60.850 24.680 63.250 ;
        RECT 25.000 62.405 25.140 63.930 ;
        RECT 24.930 62.035 25.210 62.405 ;
        RECT 25.860 62.120 26.120 62.210 ;
        RECT 26.380 62.120 26.520 66.230 ;
        RECT 26.840 63.910 26.980 68.350 ;
        RECT 27.760 64.250 27.900 71.070 ;
        RECT 28.220 64.250 28.360 71.070 ;
        RECT 28.620 69.370 28.880 69.690 ;
        RECT 28.680 64.930 28.820 69.370 ;
        RECT 29.080 68.350 29.340 68.670 ;
        RECT 29.140 64.930 29.280 68.350 ;
        RECT 28.620 64.610 28.880 64.930 ;
        RECT 29.080 64.610 29.340 64.930 ;
        RECT 29.600 64.250 29.740 75.580 ;
        RECT 30.520 75.210 30.660 87.390 ;
        RECT 31.380 86.030 31.640 86.350 ;
        RECT 31.440 82.270 31.580 86.030 ;
        RECT 35.580 84.990 35.720 92.830 ;
        RECT 36.900 91.470 37.160 91.790 ;
        RECT 36.960 89.410 37.100 91.470 ;
        RECT 36.900 89.090 37.160 89.410 ;
        RECT 35.520 84.670 35.780 84.990 ;
        RECT 31.380 81.950 31.640 82.270 ;
        RECT 31.440 78.530 31.580 81.950 ;
        RECT 32.300 80.590 32.560 80.910 ;
        RECT 31.380 78.210 31.640 78.530 ;
        RECT 31.440 77.510 31.580 78.210 ;
        RECT 31.380 77.190 31.640 77.510 ;
        RECT 30.920 76.850 31.180 77.170 ;
        RECT 30.980 75.810 31.120 76.850 ;
        RECT 31.840 76.510 32.100 76.830 ;
        RECT 30.920 75.490 31.180 75.810 ;
        RECT 30.000 74.810 30.260 75.130 ;
        RECT 30.520 75.070 31.580 75.210 ;
        RECT 30.060 71.390 30.200 74.810 ;
        RECT 31.440 72.750 31.580 75.070 ;
        RECT 31.900 74.790 32.040 76.510 ;
        RECT 31.840 74.470 32.100 74.790 ;
        RECT 31.380 72.430 31.640 72.750 ;
        RECT 30.460 71.750 30.720 72.070 ;
        RECT 30.920 71.750 31.180 72.070 ;
        RECT 30.000 71.070 30.260 71.390 ;
        RECT 30.060 66.970 30.200 71.070 ;
        RECT 30.000 66.650 30.260 66.970 ;
        RECT 27.700 63.930 27.960 64.250 ;
        RECT 28.160 63.930 28.420 64.250 ;
        RECT 28.620 63.930 28.880 64.250 ;
        RECT 29.540 63.930 29.800 64.250 ;
        RECT 26.780 63.590 27.040 63.910 ;
        RECT 26.780 62.910 27.040 63.230 ;
        RECT 27.700 62.970 27.960 63.230 ;
        RECT 27.300 62.910 27.960 62.970 ;
        RECT 25.860 61.980 26.520 62.120 ;
        RECT 25.860 61.890 26.120 61.980 ;
        RECT 24.480 60.530 24.740 60.850 ;
        RECT 26.320 60.530 26.580 60.850 ;
        RECT 24.370 59.655 25.910 60.025 ;
        RECT 26.380 59.490 26.520 60.530 ;
        RECT 24.480 59.170 24.740 59.490 ;
        RECT 26.320 59.170 26.580 59.490 ;
        RECT 24.020 58.830 24.280 59.150 ;
        RECT 23.560 58.490 23.820 58.810 ;
        RECT 23.160 58.070 23.760 58.210 ;
        RECT 21.070 56.935 22.610 57.305 ;
        RECT 22.630 55.915 22.910 56.285 ;
        RECT 23.100 56.110 23.360 56.430 ;
        RECT 22.700 55.750 22.840 55.915 ;
        RECT 20.800 55.430 21.060 55.750 ;
        RECT 22.640 55.430 22.900 55.750 ;
        RECT 20.340 53.050 20.600 53.370 ;
        RECT 20.860 52.770 21.000 55.430 ;
        RECT 20.400 52.630 21.000 52.770 ;
        RECT 22.700 52.690 22.840 55.430 ;
        RECT 19.880 50.330 20.140 50.650 ;
        RECT 19.420 47.950 19.680 48.270 ;
        RECT 18.500 44.890 18.760 45.210 ;
        RECT 17.580 44.550 17.840 44.870 ;
        RECT 17.120 44.210 17.380 44.530 ;
        RECT 16.660 43.870 16.920 44.190 ;
        RECT 15.740 41.150 16.000 41.470 ;
        RECT 15.280 39.110 15.540 39.430 ;
        RECT 15.340 37.730 15.480 39.110 ;
        RECT 15.800 38.750 15.940 41.150 ;
        RECT 17.180 38.750 17.320 44.210 ;
        RECT 17.640 42.490 17.780 44.550 ;
        RECT 19.480 43.170 19.620 47.950 ;
        RECT 19.940 47.930 20.080 50.330 ;
        RECT 19.880 47.610 20.140 47.930 ;
        RECT 20.400 47.330 20.540 52.630 ;
        RECT 22.640 52.370 22.900 52.690 ;
        RECT 21.070 51.495 22.610 51.865 ;
        RECT 22.640 49.310 22.900 49.630 ;
        RECT 19.940 47.190 20.540 47.330 ;
        RECT 22.700 47.330 22.840 49.310 ;
        RECT 23.160 48.270 23.300 56.110 ;
        RECT 23.620 55.410 23.760 58.070 ;
        RECT 24.540 55.750 24.680 59.170 ;
        RECT 25.400 58.830 25.660 59.150 ;
        RECT 24.480 55.430 24.740 55.750 ;
        RECT 23.560 55.090 23.820 55.410 ;
        RECT 25.460 55.070 25.600 58.830 ;
        RECT 26.320 57.810 26.580 58.130 ;
        RECT 26.380 56.770 26.520 57.810 ;
        RECT 26.320 56.450 26.580 56.770 ;
        RECT 24.020 54.750 24.280 55.070 ;
        RECT 25.400 54.750 25.660 55.070 ;
        RECT 24.080 53.450 24.220 54.750 ;
        RECT 24.370 54.215 25.910 54.585 ;
        RECT 23.560 53.050 23.820 53.370 ;
        RECT 24.080 53.310 24.680 53.450 ;
        RECT 23.620 50.310 23.760 53.050 ;
        RECT 24.020 52.370 24.280 52.690 ;
        RECT 23.560 49.990 23.820 50.310 ;
        RECT 23.620 48.610 23.760 49.990 ;
        RECT 23.560 48.290 23.820 48.610 ;
        RECT 23.100 47.950 23.360 48.270 ;
        RECT 22.700 47.190 23.300 47.330 ;
        RECT 19.940 45.210 20.080 47.190 ;
        RECT 20.340 46.590 20.600 46.910 ;
        RECT 20.400 45.890 20.540 46.590 ;
        RECT 21.070 46.055 22.610 46.425 ;
        RECT 20.340 45.570 20.600 45.890 ;
        RECT 19.880 44.890 20.140 45.210 ;
        RECT 19.420 42.850 19.680 43.170 ;
        RECT 19.940 42.830 20.080 44.890 ;
        RECT 19.880 42.510 20.140 42.830 ;
        RECT 17.580 42.170 17.840 42.490 ;
        RECT 17.640 39.430 17.780 42.170 ;
        RECT 19.940 39.430 20.080 42.510 ;
        RECT 20.340 41.490 20.600 41.810 ;
        RECT 20.400 40.360 20.540 41.490 ;
        RECT 23.160 41.470 23.300 47.190 ;
        RECT 24.080 45.890 24.220 52.370 ;
        RECT 24.540 49.970 24.680 53.310 ;
        RECT 24.930 53.195 25.210 53.565 ;
        RECT 24.940 53.050 25.200 53.195 ;
        RECT 26.320 52.710 26.580 53.030 ;
        RECT 24.480 49.650 24.740 49.970 ;
        RECT 24.370 48.775 25.910 49.145 ;
        RECT 24.020 45.570 24.280 45.890 ;
        RECT 23.560 42.850 23.820 43.170 ;
        RECT 23.100 41.150 23.360 41.470 ;
        RECT 21.070 40.615 22.610 40.985 ;
        RECT 20.400 40.220 21.000 40.360 ;
        RECT 20.860 39.430 21.000 40.220 ;
        RECT 17.580 39.110 17.840 39.430 ;
        RECT 19.880 39.340 20.140 39.430 ;
        RECT 19.480 39.200 20.140 39.340 ;
        RECT 15.740 38.430 16.000 38.750 ;
        RECT 17.120 38.430 17.380 38.750 ;
        RECT 14.820 37.410 15.080 37.730 ;
        RECT 15.280 37.410 15.540 37.730 ;
        RECT 17.180 35.010 17.320 38.430 ;
        RECT 15.740 34.690 16.000 35.010 ;
        RECT 17.120 34.690 17.380 35.010 ;
        RECT 14.360 33.670 14.620 33.990 ;
        RECT 13.440 33.330 13.700 33.650 ;
        RECT 14.810 33.475 15.090 33.845 ;
        RECT 14.820 33.330 15.080 33.475 ;
        RECT 12.520 32.990 12.780 33.310 ;
        RECT 12.980 32.990 13.240 33.310 ;
        RECT 13.500 29.230 13.640 33.330 ;
        RECT 14.360 32.990 14.620 33.310 ;
        RECT 14.420 31.270 14.560 32.990 ;
        RECT 15.800 31.950 15.940 34.690 ;
        RECT 16.200 34.010 16.460 34.330 ;
        RECT 15.740 31.630 16.000 31.950 ;
        RECT 16.260 31.610 16.400 34.010 ;
        RECT 16.200 31.290 16.460 31.610 ;
        RECT 14.360 30.950 14.620 31.270 ;
        RECT 17.180 30.590 17.320 34.690 ;
        RECT 19.480 33.990 19.620 39.200 ;
        RECT 19.880 39.110 20.140 39.200 ;
        RECT 20.800 39.110 21.060 39.430 ;
        RECT 21.260 38.430 21.520 38.750 ;
        RECT 21.320 37.730 21.460 38.430 ;
        RECT 23.620 37.730 23.760 42.850 ;
        RECT 24.080 42.150 24.220 45.570 ;
        RECT 26.380 44.870 26.520 52.710 ;
        RECT 26.320 44.550 26.580 44.870 ;
        RECT 24.370 43.335 25.910 43.705 ;
        RECT 24.020 41.830 24.280 42.150 ;
        RECT 26.380 39.285 26.520 44.550 ;
        RECT 26.840 43.170 26.980 62.910 ;
        RECT 27.300 62.830 27.900 62.910 ;
        RECT 27.300 50.310 27.440 62.830 ;
        RECT 28.680 62.210 28.820 63.930 ;
        RECT 29.600 62.970 29.740 63.930 ;
        RECT 30.060 63.570 30.200 66.650 ;
        RECT 30.000 63.250 30.260 63.570 ;
        RECT 29.600 62.830 30.200 62.970 ;
        RECT 28.620 61.890 28.880 62.210 ;
        RECT 30.060 60.850 30.200 62.830 ;
        RECT 30.520 61.190 30.660 71.750 ;
        RECT 30.980 61.530 31.120 71.750 ;
        RECT 30.920 61.210 31.180 61.530 ;
        RECT 30.460 60.870 30.720 61.190 ;
        RECT 30.000 60.530 30.260 60.850 ;
        RECT 29.080 60.190 29.340 60.510 ;
        RECT 29.140 58.810 29.280 60.190 ;
        RECT 30.980 59.490 31.120 61.210 ;
        RECT 30.920 59.170 31.180 59.490 ;
        RECT 29.080 58.490 29.340 58.810 ;
        RECT 28.160 58.150 28.420 58.470 ;
        RECT 27.700 55.320 27.960 55.410 ;
        RECT 28.220 55.320 28.360 58.150 ;
        RECT 28.620 56.450 28.880 56.770 ;
        RECT 28.680 55.750 28.820 56.450 ;
        RECT 28.620 55.430 28.880 55.750 ;
        RECT 27.700 55.180 28.360 55.320 ;
        RECT 27.700 55.090 27.960 55.180 ;
        RECT 28.220 53.370 28.360 55.180 ;
        RECT 28.680 53.710 28.820 55.430 ;
        RECT 29.140 55.410 29.280 58.490 ;
        RECT 30.980 56.770 31.120 59.170 ;
        RECT 30.920 56.450 31.180 56.770 ;
        RECT 29.080 55.090 29.340 55.410 ;
        RECT 28.620 53.390 28.880 53.710 ;
        RECT 28.160 53.050 28.420 53.370 ;
        RECT 27.240 49.990 27.500 50.310 ;
        RECT 27.300 48.690 27.440 49.990 ;
        RECT 27.300 48.550 27.900 48.690 ;
        RECT 27.240 47.270 27.500 47.590 ;
        RECT 26.780 42.850 27.040 43.170 ;
        RECT 27.300 42.490 27.440 47.270 ;
        RECT 27.760 44.870 27.900 48.550 ;
        RECT 27.700 44.550 27.960 44.870 ;
        RECT 27.700 42.510 27.960 42.830 ;
        RECT 27.240 42.170 27.500 42.490 ;
        RECT 27.760 41.810 27.900 42.510 ;
        RECT 27.700 41.490 27.960 41.810 ;
        RECT 26.780 41.150 27.040 41.470 ;
        RECT 24.020 38.770 24.280 39.090 ;
        RECT 26.310 38.915 26.590 39.285 ;
        RECT 21.260 37.410 21.520 37.730 ;
        RECT 23.560 37.410 23.820 37.730 ;
        RECT 19.880 36.730 20.140 37.050 ;
        RECT 20.330 36.875 20.610 37.245 ;
        RECT 24.080 37.130 24.220 38.770 ;
        RECT 26.840 38.750 26.980 41.150 ;
        RECT 27.240 39.790 27.500 40.110 ;
        RECT 26.320 38.430 26.580 38.750 ;
        RECT 26.780 38.430 27.040 38.750 ;
        RECT 24.370 37.895 25.910 38.265 ;
        RECT 23.620 37.050 24.220 37.130 ;
        RECT 23.560 36.990 24.220 37.050 ;
        RECT 20.340 36.730 20.600 36.875 ;
        RECT 23.560 36.730 23.820 36.990 ;
        RECT 25.850 36.875 26.130 37.245 ;
        RECT 26.380 37.130 26.520 38.430 ;
        RECT 26.380 37.050 26.980 37.130 ;
        RECT 26.380 36.990 27.040 37.050 ;
        RECT 19.420 33.670 19.680 33.990 ;
        RECT 19.480 32.290 19.620 33.670 ;
        RECT 19.940 33.310 20.080 36.730 ;
        RECT 23.100 36.050 23.360 36.370 ;
        RECT 21.070 35.175 22.610 35.545 ;
        RECT 23.160 33.990 23.300 36.050 ;
        RECT 25.920 35.010 26.060 36.875 ;
        RECT 26.780 36.730 27.040 36.990 ;
        RECT 24.020 34.690 24.280 35.010 ;
        RECT 25.860 34.690 26.120 35.010 ;
        RECT 23.100 33.670 23.360 33.990 ;
        RECT 19.880 32.990 20.140 33.310 ;
        RECT 19.420 31.970 19.680 32.290 ;
        RECT 17.120 30.270 17.380 30.590 ;
        RECT 19.480 29.570 19.620 31.970 ;
        RECT 20.340 31.290 20.600 31.610 ;
        RECT 19.420 29.250 19.680 29.570 ;
        RECT 20.400 29.230 20.540 31.290 ;
        RECT 24.080 30.590 24.220 34.690 ;
        RECT 27.300 33.990 27.440 39.790 ;
        RECT 26.770 33.475 27.050 33.845 ;
        RECT 27.240 33.670 27.500 33.990 ;
        RECT 26.780 33.330 27.040 33.475 ;
        RECT 24.370 32.455 25.910 32.825 ;
        RECT 27.760 32.290 27.900 41.490 ;
        RECT 28.220 40.110 28.360 53.050 ;
        RECT 28.680 51.330 28.820 53.390 ;
        RECT 29.540 52.030 29.800 52.350 ;
        RECT 28.620 51.010 28.880 51.330 ;
        RECT 29.600 48.270 29.740 52.030 ;
        RECT 29.540 47.950 29.800 48.270 ;
        RECT 31.440 47.930 31.580 72.430 ;
        RECT 31.840 71.925 32.100 72.070 ;
        RECT 31.830 71.555 32.110 71.925 ;
        RECT 32.360 62.405 32.500 80.590 ;
        RECT 36.900 80.250 37.160 80.570 ;
        RECT 35.980 79.230 36.240 79.550 ;
        RECT 34.600 78.210 34.860 78.530 ;
        RECT 32.760 76.510 33.020 76.830 ;
        RECT 32.820 69.090 32.960 76.510 ;
        RECT 34.660 75.810 34.800 78.210 ;
        RECT 36.040 77.510 36.180 79.230 ;
        RECT 36.960 78.530 37.100 80.250 ;
        RECT 36.900 78.210 37.160 78.530 ;
        RECT 35.980 77.190 36.240 77.510 ;
        RECT 34.600 75.490 34.860 75.810 ;
        RECT 34.660 72.410 34.800 75.490 ;
        RECT 34.600 72.090 34.860 72.410 ;
        RECT 35.980 72.090 36.240 72.410 ;
        RECT 33.670 71.555 33.950 71.925 ;
        RECT 32.820 69.010 33.420 69.090 ;
        RECT 32.820 68.950 33.480 69.010 ;
        RECT 33.220 68.690 33.480 68.950 ;
        RECT 32.760 65.630 33.020 65.950 ;
        RECT 32.820 64.250 32.960 65.630 ;
        RECT 32.760 63.930 33.020 64.250 ;
        RECT 32.290 62.035 32.570 62.405 ;
        RECT 32.360 59.150 32.500 62.035 ;
        RECT 33.220 60.420 33.480 60.510 ;
        RECT 33.740 60.420 33.880 71.555 ;
        RECT 34.600 71.070 34.860 71.390 ;
        RECT 34.660 69.690 34.800 71.070 ;
        RECT 35.520 70.050 35.780 70.370 ;
        RECT 34.140 69.370 34.400 69.690 ;
        RECT 34.600 69.370 34.860 69.690 ;
        RECT 35.060 69.370 35.320 69.690 ;
        RECT 34.200 66.290 34.340 69.370 ;
        RECT 35.120 66.630 35.260 69.370 ;
        RECT 35.060 66.310 35.320 66.630 ;
        RECT 34.140 65.970 34.400 66.290 ;
        RECT 34.200 64.590 34.340 65.970 ;
        RECT 34.140 64.270 34.400 64.590 ;
        RECT 34.200 62.210 34.340 64.270 ;
        RECT 34.600 63.590 34.860 63.910 ;
        RECT 34.140 61.890 34.400 62.210 ;
        RECT 33.220 60.280 33.880 60.420 ;
        RECT 33.220 60.190 33.480 60.280 ;
        RECT 32.300 58.830 32.560 59.150 ;
        RECT 31.840 49.650 32.100 49.970 ;
        RECT 31.900 48.610 32.040 49.650 ;
        RECT 32.360 49.630 32.500 58.830 ;
        RECT 32.760 55.770 33.020 56.090 ;
        RECT 32.300 49.310 32.560 49.630 ;
        RECT 31.840 48.290 32.100 48.610 ;
        RECT 31.380 47.610 31.640 47.930 ;
        RECT 31.440 45.550 31.580 47.610 ;
        RECT 32.360 47.590 32.500 49.310 ;
        RECT 32.300 47.270 32.560 47.590 ;
        RECT 32.820 46.910 32.960 55.770 ;
        RECT 33.220 49.990 33.480 50.310 ;
        RECT 32.760 46.590 33.020 46.910 ;
        RECT 31.380 45.230 31.640 45.550 ;
        RECT 33.280 44.530 33.420 49.990 ;
        RECT 33.740 47.250 33.880 60.280 ;
        RECT 34.660 57.790 34.800 63.590 ;
        RECT 35.120 63.230 35.260 66.310 ;
        RECT 35.060 62.910 35.320 63.230 ;
        RECT 35.580 58.810 35.720 70.050 ;
        RECT 36.040 67.650 36.180 72.090 ;
        RECT 36.440 71.410 36.700 71.730 ;
        RECT 35.980 67.330 36.240 67.650 ;
        RECT 36.500 67.310 36.640 71.410 ;
        RECT 36.440 66.990 36.700 67.310 ;
        RECT 37.420 66.630 37.560 133.630 ;
        RECT 37.880 121.030 38.020 141.790 ;
        RECT 38.340 131.230 38.480 142.810 ;
        RECT 39.260 141.090 39.400 148.930 ;
        RECT 39.720 146.190 39.860 150.970 ;
        RECT 40.570 148.395 40.850 148.765 ;
        RECT 40.580 148.250 40.840 148.395 ;
        RECT 42.020 146.530 42.160 153.350 ;
        RECT 42.480 151.970 42.620 153.350 ;
        RECT 42.420 151.650 42.680 151.970 ;
        RECT 44.320 150.270 44.460 153.350 ;
        RECT 44.260 149.950 44.520 150.270 ;
        RECT 44.320 148.230 44.460 149.950 ;
        RECT 44.260 147.910 44.520 148.230 ;
        RECT 43.340 147.230 43.600 147.550 ;
        RECT 43.400 146.530 43.540 147.230 ;
        RECT 41.960 146.210 42.220 146.530 ;
        RECT 43.340 146.210 43.600 146.530 ;
        RECT 39.660 145.870 39.920 146.190 ;
        RECT 39.200 140.770 39.460 141.090 ;
        RECT 39.200 140.090 39.460 140.410 ;
        RECT 39.260 138.030 39.400 140.090 ;
        RECT 39.200 137.710 39.460 138.030 ;
        RECT 39.260 131.230 39.400 137.710 ;
        RECT 39.720 135.310 39.860 145.870 ;
        RECT 44.320 143.210 44.460 147.910 ;
        RECT 45.180 147.230 45.440 147.550 ;
        RECT 45.240 146.190 45.380 147.230 ;
        RECT 45.180 145.870 45.440 146.190 ;
        RECT 44.720 145.530 44.980 145.850 ;
        RECT 44.780 143.810 44.920 145.530 ;
        RECT 45.180 144.510 45.440 144.830 ;
        RECT 45.240 143.810 45.380 144.510 ;
        RECT 44.720 143.490 44.980 143.810 ;
        RECT 45.180 143.490 45.440 143.810 ;
        RECT 44.320 143.070 44.920 143.210 ;
        RECT 41.040 142.130 41.300 142.450 ;
        RECT 41.100 140.410 41.240 142.130 ;
        RECT 44.260 141.790 44.520 142.110 ;
        RECT 41.040 140.090 41.300 140.410 ;
        RECT 43.800 140.090 44.060 140.410 ;
        RECT 41.100 135.650 41.240 140.090 ;
        RECT 43.860 137.350 44.000 140.090 ;
        RECT 43.800 137.030 44.060 137.350 ;
        RECT 42.420 136.350 42.680 136.670 ;
        RECT 41.040 135.330 41.300 135.650 ;
        RECT 39.660 134.990 39.920 135.310 ;
        RECT 40.580 134.650 40.840 134.970 ;
        RECT 40.640 132.930 40.780 134.650 ;
        RECT 40.580 132.610 40.840 132.930 ;
        RECT 42.480 132.250 42.620 136.350 ;
        RECT 43.860 135.650 44.000 137.030 ;
        RECT 43.800 135.330 44.060 135.650 ;
        RECT 42.420 131.930 42.680 132.250 ;
        RECT 39.660 131.590 39.920 131.910 ;
        RECT 38.280 130.910 38.540 131.230 ;
        RECT 39.200 130.910 39.460 131.230 ;
        RECT 38.340 128.250 38.480 130.910 ;
        RECT 39.260 129.530 39.400 130.910 ;
        RECT 39.720 129.530 39.860 131.590 ;
        RECT 41.040 129.550 41.300 129.870 ;
        RECT 39.200 129.210 39.460 129.530 ;
        RECT 39.660 129.210 39.920 129.530 ;
        RECT 38.340 128.110 38.940 128.250 ;
        RECT 38.270 127.315 38.550 127.685 ;
        RECT 38.280 127.170 38.540 127.315 ;
        RECT 38.340 124.770 38.480 127.170 ;
        RECT 38.800 126.810 38.940 128.110 ;
        RECT 39.260 127.490 39.400 129.210 ;
        RECT 39.200 127.170 39.460 127.490 ;
        RECT 39.720 126.890 39.860 129.210 ;
        RECT 40.570 127.315 40.850 127.685 ;
        RECT 40.580 127.170 40.840 127.315 ;
        RECT 38.740 126.490 39.000 126.810 ;
        RECT 39.260 126.750 39.860 126.890 ;
        RECT 38.280 124.450 38.540 124.770 ;
        RECT 38.800 123.070 38.940 126.490 ;
        RECT 39.260 126.470 39.400 126.750 ;
        RECT 39.200 126.150 39.460 126.470 ;
        RECT 40.120 126.150 40.380 126.470 ;
        RECT 39.260 124.430 39.400 126.150 ;
        RECT 39.660 125.470 39.920 125.790 ;
        RECT 39.200 124.110 39.460 124.430 ;
        RECT 38.740 122.750 39.000 123.070 ;
        RECT 37.820 120.710 38.080 121.030 ;
        RECT 39.720 110.470 39.860 125.470 ;
        RECT 40.180 116.610 40.320 126.150 ;
        RECT 40.640 124.770 40.780 127.170 ;
        RECT 41.100 126.130 41.240 129.550 ;
        RECT 41.500 126.830 41.760 127.150 ;
        RECT 41.040 125.810 41.300 126.130 ;
        RECT 40.580 124.450 40.840 124.770 ;
        RECT 40.120 116.290 40.380 116.610 ;
        RECT 38.340 110.330 39.860 110.470 ;
        RECT 37.820 109.490 38.080 109.810 ;
        RECT 37.880 108.450 38.020 109.490 ;
        RECT 37.820 108.130 38.080 108.450 ;
        RECT 37.820 96.570 38.080 96.890 ;
        RECT 37.880 89.410 38.020 96.570 ;
        RECT 37.820 89.090 38.080 89.410 ;
        RECT 36.440 66.310 36.700 66.630 ;
        RECT 37.360 66.310 37.620 66.630 ;
        RECT 36.500 64.930 36.640 66.310 ;
        RECT 36.900 65.630 37.160 65.950 ;
        RECT 36.440 64.610 36.700 64.930 ;
        RECT 36.440 60.530 36.700 60.850 ;
        RECT 35.520 58.490 35.780 58.810 ;
        RECT 36.500 58.130 36.640 60.530 ;
        RECT 35.980 57.810 36.240 58.130 ;
        RECT 36.440 57.810 36.700 58.130 ;
        RECT 34.600 57.470 34.860 57.790 ;
        RECT 36.040 54.050 36.180 57.810 ;
        RECT 35.980 53.730 36.240 54.050 ;
        RECT 36.040 51.330 36.180 53.730 ;
        RECT 36.960 53.370 37.100 65.630 ;
        RECT 38.340 62.170 38.480 110.330 ;
        RECT 39.200 109.490 39.460 109.810 ;
        RECT 39.260 107.770 39.400 109.490 ;
        RECT 41.100 108.110 41.240 125.810 ;
        RECT 41.560 123.750 41.700 126.830 ;
        RECT 44.320 126.810 44.460 141.790 ;
        RECT 44.780 138.030 44.920 143.070 ;
        RECT 45.240 142.790 45.380 143.490 ;
        RECT 45.180 142.470 45.440 142.790 ;
        RECT 45.700 141.090 45.840 153.350 ;
        RECT 46.160 148.230 46.300 153.350 ;
        RECT 47.080 152.990 47.220 155.390 ;
        RECT 48.460 154.350 48.600 156.410 ;
        RECT 49.840 154.690 49.980 156.410 ;
        RECT 49.320 154.370 49.580 154.690 ;
        RECT 49.780 154.370 50.040 154.690 ;
        RECT 48.400 154.030 48.660 154.350 ;
        RECT 47.480 153.350 47.740 153.670 ;
        RECT 47.020 152.670 47.280 152.990 ;
        RECT 47.080 148.230 47.220 152.670 ;
        RECT 47.540 149.250 47.680 153.350 ;
        RECT 47.940 151.650 48.200 151.970 ;
        RECT 47.480 148.930 47.740 149.250 ;
        RECT 48.000 148.910 48.140 151.650 ;
        RECT 47.940 148.590 48.200 148.910 ;
        RECT 48.000 148.230 48.140 148.590 ;
        RECT 46.100 147.910 46.360 148.230 ;
        RECT 47.020 147.910 47.280 148.230 ;
        RECT 47.940 147.910 48.200 148.230 ;
        RECT 46.160 143.470 46.300 147.910 ;
        RECT 46.100 143.150 46.360 143.470 ;
        RECT 47.080 142.450 47.220 147.910 ;
        RECT 48.000 146.610 48.140 147.910 ;
        RECT 47.540 146.470 48.140 146.610 ;
        RECT 47.540 144.830 47.680 146.470 ;
        RECT 48.460 145.930 48.600 154.030 ;
        RECT 48.860 152.670 49.120 152.990 ;
        RECT 48.920 148.230 49.060 152.670 ;
        RECT 49.380 151.970 49.520 154.370 ;
        RECT 49.780 153.690 50.040 154.010 ;
        RECT 51.160 153.690 51.420 154.010 ;
        RECT 49.320 151.650 49.580 151.970 ;
        RECT 49.320 149.950 49.580 150.270 ;
        RECT 49.380 148.230 49.520 149.950 ;
        RECT 49.840 149.250 49.980 153.690 ;
        RECT 50.700 153.350 50.960 153.670 ;
        RECT 50.760 151.630 50.900 153.350 ;
        RECT 50.700 151.310 50.960 151.630 ;
        RECT 50.240 150.970 50.500 151.290 ;
        RECT 49.780 148.930 50.040 149.250 ;
        RECT 49.780 148.250 50.040 148.570 ;
        RECT 48.860 147.910 49.120 148.230 ;
        RECT 49.320 147.910 49.580 148.230 ;
        RECT 48.000 145.850 48.600 145.930 ;
        RECT 47.940 145.790 48.600 145.850 ;
        RECT 47.940 145.530 48.200 145.790 ;
        RECT 47.480 144.510 47.740 144.830 ;
        RECT 48.460 142.450 48.600 145.790 ;
        RECT 47.020 142.130 47.280 142.450 ;
        RECT 48.400 142.130 48.660 142.450 ;
        RECT 45.640 140.770 45.900 141.090 ;
        RECT 46.100 139.750 46.360 140.070 ;
        RECT 44.720 137.710 44.980 138.030 ;
        RECT 46.160 130.210 46.300 139.750 ;
        RECT 48.460 137.350 48.600 142.130 ;
        RECT 49.840 140.070 49.980 148.250 ;
        RECT 50.300 143.810 50.440 150.970 ;
        RECT 50.760 148.570 50.900 151.310 ;
        RECT 50.700 148.250 50.960 148.570 ;
        RECT 50.700 145.530 50.960 145.850 ;
        RECT 50.760 143.810 50.900 145.530 ;
        RECT 50.240 143.490 50.500 143.810 ;
        RECT 50.700 143.490 50.960 143.810 ;
        RECT 51.220 143.130 51.360 153.690 ;
        RECT 52.600 153.525 52.740 158.630 ;
        RECT 52.080 153.010 52.340 153.330 ;
        RECT 52.530 153.155 52.810 153.525 ;
        RECT 51.620 149.950 51.880 150.270 ;
        RECT 51.680 149.250 51.820 149.950 ;
        RECT 52.140 149.250 52.280 153.010 ;
        RECT 53.060 151.290 53.200 164.230 ;
        RECT 53.920 163.550 54.180 163.870 ;
        RECT 53.980 162.510 54.120 163.550 ;
        RECT 53.920 162.190 54.180 162.510 ;
        RECT 53.920 161.510 54.180 161.830 ;
        RECT 53.980 159.790 54.120 161.510 ;
        RECT 53.920 159.470 54.180 159.790 ;
        RECT 54.440 158.770 54.580 164.230 ;
        RECT 56.740 162.850 56.880 164.230 ;
        RECT 56.680 162.530 56.940 162.850 ;
        RECT 55.300 161.170 55.560 161.490 ;
        RECT 54.840 159.470 55.100 159.790 ;
        RECT 53.460 158.450 53.720 158.770 ;
        RECT 53.980 158.630 54.580 158.770 ;
        RECT 53.520 154.010 53.660 158.450 ;
        RECT 53.460 153.690 53.720 154.010 ;
        RECT 53.980 152.165 54.120 158.630 ;
        RECT 53.910 151.795 54.190 152.165 ;
        RECT 54.380 151.650 54.640 151.970 ;
        RECT 53.920 151.310 54.180 151.630 ;
        RECT 53.000 150.970 53.260 151.290 ;
        RECT 53.460 150.290 53.720 150.610 ;
        RECT 51.620 148.930 51.880 149.250 ;
        RECT 52.080 148.930 52.340 149.250 ;
        RECT 53.520 148.230 53.660 150.290 ;
        RECT 53.460 147.910 53.720 148.230 ;
        RECT 51.620 147.230 51.880 147.550 ;
        RECT 52.540 147.230 52.800 147.550 ;
        RECT 51.160 142.810 51.420 143.130 ;
        RECT 49.780 139.750 50.040 140.070 ;
        RECT 51.220 139.390 51.360 142.810 ;
        RECT 51.160 139.070 51.420 139.390 ;
        RECT 48.400 137.030 48.660 137.350 ;
        RECT 48.460 135.310 48.600 137.030 ;
        RECT 51.220 135.650 51.360 139.070 ;
        RECT 51.160 135.330 51.420 135.650 ;
        RECT 48.400 134.990 48.660 135.310 ;
        RECT 47.940 133.630 48.200 133.950 ;
        RECT 46.560 132.610 46.820 132.930 ;
        RECT 46.100 129.890 46.360 130.210 ;
        RECT 45.180 129.210 45.440 129.530 ;
        RECT 45.240 127.490 45.380 129.210 ;
        RECT 45.180 127.170 45.440 127.490 ;
        RECT 44.260 126.490 44.520 126.810 ;
        RECT 43.340 124.110 43.600 124.430 ;
        RECT 41.500 123.430 41.760 123.750 ;
        RECT 42.420 122.750 42.680 123.070 ;
        RECT 42.480 121.030 42.620 122.750 ;
        RECT 42.420 120.710 42.680 121.030 ;
        RECT 43.400 116.610 43.540 124.110 ;
        RECT 44.320 122.050 44.460 126.490 ;
        RECT 46.160 126.470 46.300 129.890 ;
        RECT 46.620 126.810 46.760 132.610 ;
        RECT 48.000 131.910 48.140 133.630 ;
        RECT 48.460 131.910 48.600 134.990 ;
        RECT 51.220 134.630 51.360 135.330 ;
        RECT 51.680 134.630 51.820 147.230 ;
        RECT 52.600 142.790 52.740 147.230 ;
        RECT 53.520 146.190 53.660 147.910 ;
        RECT 53.460 145.870 53.720 146.190 ;
        RECT 53.980 145.170 54.120 151.310 ;
        RECT 54.440 146.530 54.580 151.650 ;
        RECT 54.900 150.610 55.040 159.470 ;
        RECT 55.360 153.330 55.500 161.170 ;
        RECT 56.680 160.830 56.940 161.150 ;
        RECT 56.740 159.450 56.880 160.830 ;
        RECT 57.660 160.130 57.800 164.230 ;
        RECT 62.660 163.890 62.920 164.210 ;
        RECT 64.030 164.035 64.310 164.405 ;
        RECT 65.020 164.210 65.160 165.250 ;
        RECT 67.780 165.230 67.920 173.570 ;
        RECT 74.220 165.570 74.360 173.570 ;
        RECT 74.160 165.250 74.420 165.570 ;
        RECT 76.460 165.250 76.720 165.570 ;
        RECT 67.720 164.910 67.980 165.230 ;
        RECT 69.620 164.830 71.600 164.970 ;
        RECT 69.620 164.550 69.760 164.830 ;
        RECT 69.560 164.230 69.820 164.550 ;
        RECT 71.460 164.210 71.600 164.830 ;
        RECT 76.520 164.550 76.660 165.250 ;
        RECT 77.440 164.890 77.580 173.570 ;
        RECT 82.440 165.250 82.700 165.570 ;
        RECT 77.380 164.570 77.640 164.890 ;
        RECT 74.620 164.230 74.880 164.550 ;
        RECT 76.460 164.405 76.720 164.550 ;
        RECT 64.040 163.890 64.300 164.035 ;
        RECT 64.960 163.890 65.220 164.210 ;
        RECT 66.800 163.890 67.060 164.210 ;
        RECT 67.260 163.890 67.520 164.210 ;
        RECT 70.940 163.890 71.200 164.210 ;
        RECT 71.400 163.890 71.660 164.210 ;
        RECT 71.860 163.890 72.120 164.210 ;
        RECT 73.240 163.890 73.500 164.210 ;
        RECT 61.280 163.550 61.540 163.870 ;
        RECT 62.720 163.725 62.860 163.890 ;
        RECT 60.360 161.510 60.620 161.830 ;
        RECT 59.890 160.635 60.170 161.005 ;
        RECT 57.600 159.810 57.860 160.130 ;
        RECT 56.680 159.130 56.940 159.450 ;
        RECT 57.660 158.850 57.800 159.810 ;
        RECT 58.510 159.275 58.790 159.645 ;
        RECT 57.200 158.710 57.800 158.850 ;
        RECT 56.220 157.090 56.480 157.410 ;
        RECT 55.300 153.010 55.560 153.330 ;
        RECT 54.840 150.290 55.100 150.610 ;
        RECT 55.300 150.290 55.560 150.610 ;
        RECT 54.380 146.210 54.640 146.530 ;
        RECT 53.920 144.850 54.180 145.170 ;
        RECT 55.360 143.890 55.500 150.290 ;
        RECT 56.280 148.910 56.420 157.090 ;
        RECT 56.680 150.630 56.940 150.950 ;
        RECT 56.220 148.590 56.480 148.910 ;
        RECT 55.760 148.250 56.020 148.570 ;
        RECT 55.820 144.830 55.960 148.250 ;
        RECT 55.760 144.510 56.020 144.830 ;
        RECT 55.360 143.750 55.960 143.890 ;
        RECT 52.540 142.470 52.800 142.790 ;
        RECT 52.540 141.790 52.800 142.110 ;
        RECT 52.600 141.090 52.740 141.790 ;
        RECT 52.540 140.770 52.800 141.090 ;
        RECT 55.820 140.070 55.960 143.750 ;
        RECT 56.210 142.955 56.490 143.325 ;
        RECT 54.380 139.750 54.640 140.070 ;
        RECT 55.760 139.750 56.020 140.070 ;
        RECT 53.000 136.690 53.260 137.010 ;
        RECT 51.160 134.310 51.420 134.630 ;
        RECT 51.620 134.310 51.880 134.630 ;
        RECT 51.220 132.930 51.360 134.310 ;
        RECT 51.680 132.930 51.820 134.310 ;
        RECT 51.160 132.610 51.420 132.930 ;
        RECT 51.620 132.610 51.880 132.930 ;
        RECT 47.940 131.590 48.200 131.910 ;
        RECT 48.400 131.590 48.660 131.910 ;
        RECT 46.560 126.490 46.820 126.810 ;
        RECT 46.100 126.150 46.360 126.470 ;
        RECT 46.620 124.770 46.760 126.490 ;
        RECT 46.560 124.450 46.820 124.770 ;
        RECT 46.620 123.750 46.760 124.450 ;
        RECT 48.460 124.090 48.600 131.590 ;
        RECT 48.860 131.250 49.120 131.570 ;
        RECT 48.920 130.210 49.060 131.250 ;
        RECT 48.860 129.890 49.120 130.210 ;
        RECT 52.080 129.210 52.340 129.530 ;
        RECT 51.160 128.870 51.420 129.190 ;
        RECT 50.700 125.810 50.960 126.130 ;
        RECT 48.400 123.770 48.660 124.090 ;
        RECT 46.560 123.430 46.820 123.750 ;
        RECT 50.760 122.050 50.900 125.810 ;
        RECT 51.220 122.050 51.360 128.870 ;
        RECT 44.260 121.730 44.520 122.050 ;
        RECT 50.700 121.730 50.960 122.050 ;
        RECT 51.160 121.730 51.420 122.050 ;
        RECT 46.100 120.710 46.360 121.030 ;
        RECT 49.320 120.710 49.580 121.030 ;
        RECT 46.160 118.990 46.300 120.710 ;
        RECT 48.400 120.030 48.660 120.350 ;
        RECT 46.100 118.670 46.360 118.990 ;
        RECT 46.160 118.310 46.300 118.670 ;
        RECT 46.100 117.990 46.360 118.310 ;
        RECT 43.340 116.290 43.600 116.610 ;
        RECT 41.500 115.610 41.760 115.930 ;
        RECT 41.560 113.550 41.700 115.610 ;
        RECT 42.880 115.270 43.140 115.590 ;
        RECT 41.960 114.930 42.220 115.250 ;
        RECT 41.500 113.230 41.760 113.550 ;
        RECT 41.560 112.870 41.700 113.230 ;
        RECT 41.500 112.550 41.760 112.870 ;
        RECT 41.040 107.790 41.300 108.110 ;
        RECT 39.200 107.450 39.460 107.770 ;
        RECT 41.560 104.710 41.700 112.550 ;
        RECT 42.020 111.170 42.160 114.930 ;
        RECT 42.420 112.890 42.680 113.210 ;
        RECT 42.480 111.170 42.620 112.890 ;
        RECT 41.960 110.850 42.220 111.170 ;
        RECT 42.420 110.850 42.680 111.170 ;
        RECT 42.940 110.470 43.080 115.270 ;
        RECT 42.480 110.330 43.080 110.470 ;
        RECT 42.480 105.730 42.620 110.330 ;
        RECT 45.640 109.150 45.900 109.470 ;
        RECT 44.720 107.110 44.980 107.430 ;
        RECT 43.340 106.430 43.600 106.750 ;
        RECT 42.420 105.410 42.680 105.730 ;
        RECT 41.500 104.390 41.760 104.710 ;
        RECT 41.560 101.990 41.700 104.390 ;
        RECT 42.480 102.330 42.620 105.410 ;
        RECT 42.420 102.010 42.680 102.330 ;
        RECT 41.500 101.670 41.760 101.990 ;
        RECT 41.960 101.670 42.220 101.990 ;
        RECT 39.660 100.990 39.920 101.310 ;
        RECT 39.720 99.270 39.860 100.990 ;
        RECT 41.040 99.970 41.300 100.290 ;
        RECT 39.200 98.950 39.460 99.270 ;
        RECT 39.660 98.950 39.920 99.270 ;
        RECT 39.260 93.570 39.400 98.950 ;
        RECT 40.580 98.610 40.840 98.930 ;
        RECT 40.640 95.870 40.780 98.610 ;
        RECT 40.580 95.550 40.840 95.870 ;
        RECT 38.800 93.430 39.400 93.570 ;
        RECT 38.800 91.450 38.940 93.430 ;
        RECT 39.200 92.830 39.460 93.150 ;
        RECT 40.640 92.890 40.780 95.550 ;
        RECT 41.100 93.490 41.240 99.970 ;
        RECT 41.560 96.550 41.700 101.670 ;
        RECT 42.020 99.610 42.160 101.670 ;
        RECT 41.960 99.290 42.220 99.610 ;
        RECT 43.400 99.270 43.540 106.430 ;
        RECT 44.780 104.710 44.920 107.110 ;
        RECT 44.720 104.390 44.980 104.710 ;
        RECT 44.260 104.050 44.520 104.370 ;
        RECT 44.320 103.010 44.460 104.050 ;
        RECT 44.260 102.690 44.520 103.010 ;
        RECT 43.800 99.630 44.060 99.950 ;
        RECT 43.340 98.950 43.600 99.270 ;
        RECT 41.960 98.270 42.220 98.590 ;
        RECT 42.020 97.570 42.160 98.270 ;
        RECT 43.400 97.650 43.540 98.950 ;
        RECT 41.960 97.250 42.220 97.570 ;
        RECT 42.940 97.510 43.540 97.650 ;
        RECT 41.500 96.230 41.760 96.550 ;
        RECT 41.560 93.830 41.700 96.230 ;
        RECT 41.500 93.510 41.760 93.830 ;
        RECT 41.040 93.170 41.300 93.490 ;
        RECT 41.500 92.890 41.760 93.150 ;
        RECT 40.640 92.830 41.760 92.890 ;
        RECT 38.740 91.130 39.000 91.450 ;
        RECT 39.260 88.390 39.400 92.830 ;
        RECT 40.640 92.750 41.700 92.830 ;
        RECT 39.660 91.810 39.920 92.130 ;
        RECT 39.720 88.390 39.860 91.810 ;
        RECT 39.200 88.070 39.460 88.390 ;
        RECT 39.660 88.070 39.920 88.390 ;
        RECT 40.580 82.630 40.840 82.950 ;
        RECT 40.640 77.850 40.780 82.630 ;
        RECT 41.100 78.530 41.240 92.750 ;
        RECT 42.020 91.790 42.160 97.250 ;
        RECT 42.940 94.510 43.080 97.510 ;
        RECT 43.340 96.910 43.600 97.230 ;
        RECT 42.880 94.190 43.140 94.510 ;
        RECT 42.420 93.510 42.680 93.830 ;
        RECT 42.480 92.130 42.620 93.510 ;
        RECT 43.400 93.150 43.540 96.910 ;
        RECT 43.860 95.870 44.000 99.630 ;
        RECT 44.720 98.950 44.980 99.270 ;
        RECT 44.260 98.610 44.520 98.930 ;
        RECT 43.800 95.550 44.060 95.870 ;
        RECT 43.340 92.830 43.600 93.150 ;
        RECT 42.420 91.810 42.680 92.130 ;
        RECT 41.960 91.470 42.220 91.790 ;
        RECT 42.020 88.810 42.160 91.470 ;
        RECT 43.860 90.770 44.000 95.550 ;
        RECT 44.320 94.850 44.460 98.610 ;
        RECT 44.260 94.530 44.520 94.850 ;
        RECT 43.800 90.450 44.060 90.770 ;
        RECT 41.560 88.670 43.540 88.810 ;
        RECT 43.800 88.750 44.060 89.070 ;
        RECT 41.560 88.390 41.700 88.670 ;
        RECT 43.400 88.390 43.540 88.670 ;
        RECT 41.500 88.070 41.760 88.390 ;
        RECT 41.960 88.070 42.220 88.390 ;
        RECT 43.340 88.070 43.600 88.390 ;
        RECT 42.020 86.690 42.160 88.070 ;
        RECT 41.960 86.370 42.220 86.690 ;
        RECT 43.400 85.670 43.540 88.070 ;
        RECT 43.860 86.350 44.000 88.750 ;
        RECT 44.320 88.050 44.460 94.530 ;
        RECT 44.260 87.730 44.520 88.050 ;
        RECT 44.780 86.690 44.920 98.950 ;
        RECT 45.180 94.530 45.440 94.850 ;
        RECT 44.720 86.370 44.980 86.690 ;
        RECT 43.800 86.030 44.060 86.350 ;
        RECT 43.340 85.350 43.600 85.670 ;
        RECT 43.860 80.570 44.000 86.030 ;
        RECT 45.240 85.410 45.380 94.530 ;
        RECT 45.700 93.490 45.840 109.150 ;
        RECT 46.160 107.770 46.300 117.990 ;
        RECT 47.480 115.610 47.740 115.930 ;
        RECT 47.540 115.445 47.680 115.610 ;
        RECT 47.470 115.075 47.750 115.445 ;
        RECT 47.480 114.590 47.740 114.910 ;
        RECT 47.540 112.530 47.680 114.590 ;
        RECT 47.480 112.210 47.740 112.530 ;
        RECT 48.460 111.365 48.600 120.030 ;
        RECT 49.380 117.630 49.520 120.710 ;
        RECT 49.320 117.310 49.580 117.630 ;
        RECT 51.220 116.610 51.360 121.730 ;
        RECT 51.160 116.290 51.420 116.610 ;
        RECT 51.610 116.435 51.890 116.805 ;
        RECT 50.700 115.610 50.960 115.930 ;
        RECT 48.860 115.270 49.120 115.590 ;
        RECT 48.920 113.890 49.060 115.270 ;
        RECT 48.860 113.570 49.120 113.890 ;
        RECT 49.320 111.870 49.580 112.190 ;
        RECT 50.240 111.870 50.500 112.190 ;
        RECT 48.390 110.995 48.670 111.365 ;
        RECT 47.020 110.170 47.280 110.490 ;
        RECT 46.560 109.830 46.820 110.150 ;
        RECT 46.100 107.450 46.360 107.770 ;
        RECT 46.620 105.050 46.760 109.830 ;
        RECT 46.560 104.730 46.820 105.050 ;
        RECT 46.620 99.950 46.760 104.730 ;
        RECT 47.080 103.885 47.220 110.170 ;
        RECT 47.480 109.490 47.740 109.810 ;
        RECT 47.540 106.750 47.680 109.490 ;
        RECT 49.380 109.470 49.520 111.870 ;
        RECT 49.780 109.830 50.040 110.150 ;
        RECT 49.320 109.150 49.580 109.470 ;
        RECT 48.860 107.450 49.120 107.770 ;
        RECT 47.480 106.430 47.740 106.750 ;
        RECT 48.920 105.730 49.060 107.450 ;
        RECT 48.860 105.410 49.120 105.730 ;
        RECT 49.840 104.710 49.980 109.830 ;
        RECT 49.780 104.390 50.040 104.710 ;
        RECT 47.010 103.515 47.290 103.885 ;
        RECT 49.840 102.670 49.980 104.390 ;
        RECT 49.780 102.350 50.040 102.670 ;
        RECT 46.560 99.630 46.820 99.950 ;
        RECT 46.100 98.610 46.360 98.930 ;
        RECT 45.640 93.170 45.900 93.490 ;
        RECT 45.640 91.810 45.900 92.130 ;
        RECT 45.700 86.010 45.840 91.810 ;
        RECT 45.640 85.690 45.900 86.010 ;
        RECT 45.240 85.270 45.840 85.410 ;
        RECT 44.720 83.650 44.980 83.970 ;
        RECT 44.780 80.570 44.920 83.650 ;
        RECT 45.180 82.290 45.440 82.610 ;
        RECT 45.240 81.250 45.380 82.290 ;
        RECT 45.180 80.930 45.440 81.250 ;
        RECT 43.800 80.250 44.060 80.570 ;
        RECT 44.720 80.250 44.980 80.570 ;
        RECT 41.040 78.210 41.300 78.530 ;
        RECT 42.880 78.210 43.140 78.530 ;
        RECT 40.580 77.530 40.840 77.850 ;
        RECT 40.640 75.130 40.780 77.530 ;
        RECT 41.960 77.190 42.220 77.510 ;
        RECT 41.500 76.510 41.760 76.830 ;
        RECT 41.560 75.810 41.700 76.510 ;
        RECT 41.500 75.490 41.760 75.810 ;
        RECT 40.580 74.810 40.840 75.130 ;
        RECT 40.120 71.980 40.380 72.070 ;
        RECT 40.640 71.980 40.780 74.810 ;
        RECT 41.560 72.070 41.700 75.490 ;
        RECT 40.120 71.840 40.780 71.980 ;
        RECT 40.120 71.750 40.380 71.840 ;
        RECT 41.500 71.750 41.760 72.070 ;
        RECT 40.180 69.690 40.320 71.750 ;
        RECT 42.020 71.730 42.160 77.190 ;
        RECT 42.940 72.070 43.080 78.210 ;
        RECT 43.860 76.685 44.000 80.250 ;
        RECT 44.720 79.230 44.980 79.550 ;
        RECT 44.250 77.675 44.530 78.045 ;
        RECT 44.260 77.530 44.520 77.675 ;
        RECT 43.790 76.315 44.070 76.685 ;
        RECT 43.860 72.750 44.000 76.315 ;
        RECT 44.780 75.470 44.920 79.230 ;
        RECT 44.720 75.150 44.980 75.470 ;
        RECT 43.800 72.430 44.060 72.750 ;
        RECT 44.780 72.070 44.920 75.150 ;
        RECT 45.240 72.750 45.380 80.930 ;
        RECT 45.700 80.570 45.840 85.270 ;
        RECT 45.640 80.250 45.900 80.570 ;
        RECT 45.180 72.430 45.440 72.750 ;
        RECT 42.880 71.750 43.140 72.070 ;
        RECT 44.720 71.750 44.980 72.070 ;
        RECT 41.960 71.410 42.220 71.730 ;
        RECT 41.500 71.070 41.760 71.390 ;
        RECT 40.580 69.710 40.840 70.030 ;
        RECT 40.120 69.370 40.380 69.690 ;
        RECT 38.740 65.630 39.000 65.950 ;
        RECT 38.800 64.250 38.940 65.630 ;
        RECT 40.180 64.250 40.320 69.370 ;
        RECT 38.740 63.930 39.000 64.250 ;
        RECT 40.120 63.930 40.380 64.250 ;
        RECT 38.340 62.030 38.940 62.170 ;
        RECT 36.900 53.050 37.160 53.370 ;
        RECT 35.980 51.010 36.240 51.330 ;
        RECT 34.600 49.990 34.860 50.310 ;
        RECT 34.660 48.610 34.800 49.990 ;
        RECT 36.960 49.630 37.100 53.050 ;
        RECT 38.280 52.030 38.540 52.350 ;
        RECT 36.900 49.310 37.160 49.630 ;
        RECT 34.600 48.290 34.860 48.610 ;
        RECT 33.680 46.930 33.940 47.250 ;
        RECT 31.840 44.210 32.100 44.530 ;
        RECT 33.220 44.210 33.480 44.530 ;
        RECT 28.620 42.170 28.880 42.490 ;
        RECT 31.380 42.170 31.640 42.490 ;
        RECT 28.160 39.790 28.420 40.110 ;
        RECT 28.680 39.430 28.820 42.170 ;
        RECT 29.540 41.830 29.800 42.150 ;
        RECT 28.620 39.110 28.880 39.430 ;
        RECT 28.620 38.430 28.880 38.750 ;
        RECT 28.160 36.730 28.420 37.050 ;
        RECT 28.220 33.990 28.360 36.730 ;
        RECT 28.680 35.010 28.820 38.430 ;
        RECT 28.620 34.690 28.880 35.010 ;
        RECT 28.160 33.670 28.420 33.990 ;
        RECT 27.700 31.970 27.960 32.290 ;
        RECT 28.220 31.690 28.360 33.670 ;
        RECT 29.600 33.650 29.740 41.830 ;
        RECT 31.440 40.110 31.580 42.170 ;
        RECT 31.900 41.810 32.040 44.210 ;
        RECT 33.740 42.150 33.880 46.930 ;
        RECT 38.340 44.870 38.480 52.030 ;
        RECT 38.280 44.550 38.540 44.870 ;
        RECT 33.680 41.830 33.940 42.150 ;
        RECT 31.840 41.490 32.100 41.810 ;
        RECT 31.380 39.790 31.640 40.110 ;
        RECT 31.440 39.430 31.580 39.790 ;
        RECT 30.460 39.340 30.720 39.430 ;
        RECT 30.460 39.200 31.120 39.340 ;
        RECT 30.460 39.110 30.720 39.200 ;
        RECT 30.000 38.430 30.260 38.750 ;
        RECT 30.460 38.430 30.720 38.750 ;
        RECT 30.060 37.130 30.200 38.430 ;
        RECT 30.520 37.730 30.660 38.430 ;
        RECT 30.980 37.730 31.120 39.200 ;
        RECT 31.380 39.110 31.640 39.430 ;
        RECT 30.460 37.410 30.720 37.730 ;
        RECT 30.920 37.410 31.180 37.730 ;
        RECT 31.440 37.130 31.580 39.110 ;
        RECT 30.060 36.990 31.580 37.130 ;
        RECT 31.900 37.050 32.040 41.490 ;
        RECT 33.680 39.110 33.940 39.430 ;
        RECT 33.740 38.750 33.880 39.110 ;
        RECT 34.600 38.770 34.860 39.090 ;
        RECT 33.680 38.430 33.940 38.750 ;
        RECT 30.060 36.030 30.200 36.990 ;
        RECT 31.840 36.730 32.100 37.050 ;
        RECT 30.000 35.710 30.260 36.030 ;
        RECT 33.220 35.710 33.480 36.030 ;
        RECT 30.920 34.690 31.180 35.010 ;
        RECT 29.540 33.330 29.800 33.650 ;
        RECT 27.760 31.550 28.360 31.690 ;
        RECT 23.560 30.270 23.820 30.590 ;
        RECT 24.020 30.270 24.280 30.590 ;
        RECT 27.240 30.270 27.500 30.590 ;
        RECT 21.070 29.735 22.610 30.105 ;
        RECT 13.440 28.910 13.700 29.230 ;
        RECT 20.340 28.910 20.600 29.230 ;
        RECT 23.620 28.210 23.760 30.270 ;
        RECT 27.300 28.210 27.440 30.270 ;
        RECT 23.560 27.890 23.820 28.210 ;
        RECT 27.240 27.890 27.500 28.210 ;
        RECT 27.760 27.870 27.900 31.550 ;
        RECT 30.980 30.930 31.120 34.690 ;
        RECT 33.280 31.270 33.420 35.710 ;
        RECT 33.740 35.010 33.880 38.430 ;
        RECT 33.680 34.690 33.940 35.010 ;
        RECT 33.740 31.610 33.880 34.690 ;
        RECT 34.660 33.990 34.800 38.770 ;
        RECT 35.520 38.430 35.780 38.750 ;
        RECT 35.060 36.730 35.320 37.050 ;
        RECT 35.120 35.010 35.260 36.730 ;
        RECT 35.060 34.690 35.320 35.010 ;
        RECT 34.600 33.670 34.860 33.990 ;
        RECT 34.660 32.290 34.800 33.670 ;
        RECT 35.580 33.650 35.720 38.430 ;
        RECT 35.520 33.330 35.780 33.650 ;
        RECT 34.600 31.970 34.860 32.290 ;
        RECT 33.680 31.290 33.940 31.610 ;
        RECT 33.220 30.950 33.480 31.270 ;
        RECT 30.920 30.610 31.180 30.930 ;
        RECT 34.660 29.570 34.800 31.970 ;
        RECT 38.800 30.445 38.940 62.030 ;
        RECT 40.180 61.190 40.320 63.930 ;
        RECT 40.640 63.230 40.780 69.710 ;
        RECT 41.560 69.690 41.700 71.070 ;
        RECT 41.500 69.370 41.760 69.690 ;
        RECT 41.040 66.310 41.300 66.630 ;
        RECT 41.500 66.310 41.760 66.630 ;
        RECT 41.100 64.250 41.240 66.310 ;
        RECT 41.560 64.930 41.700 66.310 ;
        RECT 41.500 64.610 41.760 64.930 ;
        RECT 41.040 63.930 41.300 64.250 ;
        RECT 41.040 63.250 41.300 63.570 ;
        RECT 40.580 62.910 40.840 63.230 ;
        RECT 41.100 62.170 41.240 63.250 ;
        RECT 41.500 62.910 41.760 63.230 ;
        RECT 40.640 62.030 41.240 62.170 ;
        RECT 40.120 60.870 40.380 61.190 ;
        RECT 39.660 58.720 39.920 58.810 ;
        RECT 40.180 58.720 40.320 60.870 ;
        RECT 39.660 58.580 40.320 58.720 ;
        RECT 39.660 58.490 39.920 58.580 ;
        RECT 40.640 55.070 40.780 62.030 ;
        RECT 41.560 59.150 41.700 62.910 ;
        RECT 41.500 58.830 41.760 59.150 ;
        RECT 42.020 58.810 42.160 71.410 ;
        RECT 41.960 58.490 42.220 58.810 ;
        RECT 42.940 56.770 43.080 71.750 ;
        RECT 45.700 70.370 45.840 80.250 ;
        RECT 46.160 74.790 46.300 98.610 ;
        RECT 46.620 94.930 46.760 99.630 ;
        RECT 47.020 99.290 47.280 99.610 ;
        RECT 47.080 95.870 47.220 99.290 ;
        RECT 50.300 99.270 50.440 111.870 ;
        RECT 50.760 105.390 50.900 115.610 ;
        RECT 51.680 110.470 51.820 116.435 ;
        RECT 52.140 113.210 52.280 129.210 ;
        RECT 53.060 129.190 53.200 136.690 ;
        RECT 53.920 132.610 54.180 132.930 ;
        RECT 53.460 131.250 53.720 131.570 ;
        RECT 53.520 130.210 53.660 131.250 ;
        RECT 53.980 130.210 54.120 132.610 ;
        RECT 53.460 129.890 53.720 130.210 ;
        RECT 53.920 129.890 54.180 130.210 ;
        RECT 53.000 128.870 53.260 129.190 ;
        RECT 53.460 121.730 53.720 122.050 ;
        RECT 53.520 121.370 53.660 121.730 ;
        RECT 53.000 121.050 53.260 121.370 ;
        RECT 53.460 121.050 53.720 121.370 ;
        RECT 53.060 119.330 53.200 121.050 ;
        RECT 53.000 119.010 53.260 119.330 ;
        RECT 53.060 118.650 53.200 119.010 ;
        RECT 52.540 118.330 52.800 118.650 ;
        RECT 53.000 118.330 53.260 118.650 ;
        RECT 52.600 116.610 52.740 118.330 ;
        RECT 52.540 116.290 52.800 116.610 ;
        RECT 53.460 115.270 53.720 115.590 ;
        RECT 53.000 114.590 53.260 114.910 ;
        RECT 53.060 113.210 53.200 114.590 ;
        RECT 52.080 112.890 52.340 113.210 ;
        RECT 53.000 112.890 53.260 113.210 ;
        RECT 52.540 112.550 52.800 112.870 ;
        RECT 52.600 110.740 52.740 112.550 ;
        RECT 53.000 110.740 53.260 110.830 ;
        RECT 52.600 110.600 53.260 110.740 ;
        RECT 52.080 110.470 52.340 110.490 ;
        RECT 51.680 110.330 52.340 110.470 ;
        RECT 52.080 110.170 52.340 110.330 ;
        RECT 51.620 109.830 51.880 110.150 ;
        RECT 51.160 109.490 51.420 109.810 ;
        RECT 51.220 108.110 51.360 109.490 ;
        RECT 51.160 107.790 51.420 108.110 ;
        RECT 50.700 105.070 50.960 105.390 ;
        RECT 49.320 98.950 49.580 99.270 ;
        RECT 50.240 98.950 50.500 99.270 ;
        RECT 47.480 98.270 47.740 98.590 ;
        RECT 47.540 97.230 47.680 98.270 ;
        RECT 47.480 96.910 47.740 97.230 ;
        RECT 49.380 96.670 49.520 98.950 ;
        RECT 50.300 96.670 50.440 98.950 ;
        RECT 49.380 96.530 49.980 96.670 ;
        RECT 50.300 96.530 50.900 96.670 ;
        RECT 49.840 95.870 49.980 96.530 ;
        RECT 50.240 95.890 50.500 96.210 ;
        RECT 47.020 95.780 47.280 95.870 ;
        RECT 47.020 95.640 47.680 95.780 ;
        RECT 47.020 95.550 47.280 95.640 ;
        RECT 46.620 94.790 47.220 94.930 ;
        RECT 46.560 93.170 46.820 93.490 ;
        RECT 46.620 86.690 46.760 93.170 ;
        RECT 47.080 90.430 47.220 94.790 ;
        RECT 47.540 93.830 47.680 95.640 ;
        RECT 49.780 95.550 50.040 95.870 ;
        RECT 49.840 94.510 49.980 95.550 ;
        RECT 50.300 94.850 50.440 95.890 ;
        RECT 50.240 94.530 50.500 94.850 ;
        RECT 48.860 94.190 49.120 94.510 ;
        RECT 49.780 94.190 50.040 94.510 ;
        RECT 48.400 93.850 48.660 94.170 ;
        RECT 47.480 93.510 47.740 93.830 ;
        RECT 47.940 93.510 48.200 93.830 ;
        RECT 47.540 90.850 47.680 93.510 ;
        RECT 48.000 91.790 48.140 93.510 ;
        RECT 47.940 91.470 48.200 91.790 ;
        RECT 48.460 91.450 48.600 93.850 ;
        RECT 48.920 93.150 49.060 94.190 ;
        RECT 49.840 93.490 49.980 94.190 ;
        RECT 49.780 93.170 50.040 93.490 ;
        RECT 48.860 92.830 49.120 93.150 ;
        RECT 48.400 91.360 48.660 91.450 ;
        RECT 49.320 91.360 49.580 91.450 ;
        RECT 49.840 91.360 49.980 93.170 ;
        RECT 50.760 92.130 50.900 96.530 ;
        RECT 50.700 91.810 50.960 92.130 ;
        RECT 48.400 91.220 49.060 91.360 ;
        RECT 48.400 91.130 48.660 91.220 ;
        RECT 47.540 90.710 48.140 90.850 ;
        RECT 48.000 90.430 48.140 90.710 ;
        RECT 47.020 90.110 47.280 90.430 ;
        RECT 47.940 90.110 48.200 90.430 ;
        RECT 46.560 86.370 46.820 86.690 ;
        RECT 46.620 83.970 46.760 86.370 ;
        RECT 47.080 86.010 47.220 90.110 ;
        RECT 47.020 85.690 47.280 86.010 ;
        RECT 46.560 83.650 46.820 83.970 ;
        RECT 46.550 82.435 46.830 82.805 ;
        RECT 47.020 82.630 47.280 82.950 ;
        RECT 46.620 82.270 46.760 82.435 ;
        RECT 46.560 81.950 46.820 82.270 ;
        RECT 47.080 81.250 47.220 82.630 ;
        RECT 47.480 81.950 47.740 82.270 ;
        RECT 47.020 80.930 47.280 81.250 ;
        RECT 47.080 77.420 47.220 80.930 ;
        RECT 47.540 79.970 47.680 81.950 ;
        RECT 48.000 81.250 48.140 90.110 ;
        RECT 48.400 85.350 48.660 85.670 ;
        RECT 47.940 80.930 48.200 81.250 ;
        RECT 47.930 80.395 48.210 80.765 ;
        RECT 48.460 80.570 48.600 85.350 ;
        RECT 48.920 83.970 49.060 91.220 ;
        RECT 49.320 91.220 49.980 91.360 ;
        RECT 49.320 91.130 49.580 91.220 ;
        RECT 49.320 90.450 49.580 90.770 ;
        RECT 49.380 86.350 49.520 90.450 ;
        RECT 49.320 86.030 49.580 86.350 ;
        RECT 48.860 83.880 49.120 83.970 ;
        RECT 48.860 83.740 49.520 83.880 ;
        RECT 48.860 83.650 49.120 83.740 ;
        RECT 48.860 82.970 49.120 83.290 ;
        RECT 48.920 81.250 49.060 82.970 ;
        RECT 48.860 80.930 49.120 81.250 ;
        RECT 47.940 80.250 48.200 80.395 ;
        RECT 48.400 80.250 48.660 80.570 ;
        RECT 47.540 79.830 48.600 79.970 ;
        RECT 48.460 78.530 48.600 79.830 ;
        RECT 48.920 78.530 49.060 80.930 ;
        RECT 48.400 78.210 48.660 78.530 ;
        RECT 48.860 78.210 49.120 78.530 ;
        RECT 47.480 77.420 47.740 77.510 ;
        RECT 47.080 77.280 47.740 77.420 ;
        RECT 47.480 77.190 47.740 77.280 ;
        RECT 46.560 76.510 46.820 76.830 ;
        RECT 46.100 74.470 46.360 74.790 ;
        RECT 46.160 72.410 46.300 74.470 ;
        RECT 46.100 72.090 46.360 72.410 ;
        RECT 45.640 70.050 45.900 70.370 ;
        RECT 46.620 63.910 46.760 76.510 ;
        RECT 47.480 73.790 47.740 74.110 ;
        RECT 47.540 72.750 47.680 73.790 ;
        RECT 48.460 72.750 48.600 78.210 ;
        RECT 48.860 77.365 49.120 77.510 ;
        RECT 48.850 76.995 49.130 77.365 ;
        RECT 48.860 76.510 49.120 76.830 ;
        RECT 47.480 72.430 47.740 72.750 ;
        RECT 48.400 72.430 48.660 72.750 ;
        RECT 47.540 69.690 47.680 72.430 ;
        RECT 48.920 71.925 49.060 76.510 ;
        RECT 49.380 75.810 49.520 83.740 ;
        RECT 49.840 82.950 49.980 91.220 ;
        RECT 51.220 89.410 51.360 107.790 ;
        RECT 51.680 105.390 51.820 109.830 ;
        RECT 52.140 108.110 52.280 110.170 ;
        RECT 52.080 107.790 52.340 108.110 ;
        RECT 52.600 107.340 52.740 110.600 ;
        RECT 53.000 110.510 53.260 110.600 ;
        RECT 52.140 107.200 52.740 107.340 ;
        RECT 51.620 105.070 51.880 105.390 ;
        RECT 51.620 104.390 51.880 104.710 ;
        RECT 51.680 103.010 51.820 104.390 ;
        RECT 51.620 102.690 51.880 103.010 ;
        RECT 52.140 102.330 52.280 107.200 ;
        RECT 53.000 104.390 53.260 104.710 ;
        RECT 52.540 102.350 52.800 102.670 ;
        RECT 52.080 102.010 52.340 102.330 ;
        RECT 52.600 98.590 52.740 102.350 ;
        RECT 52.540 98.270 52.800 98.590 ;
        RECT 51.620 96.230 51.880 96.550 ;
        RECT 51.680 94.850 51.820 96.230 ;
        RECT 51.620 94.530 51.880 94.850 ;
        RECT 51.680 91.790 51.820 94.530 ;
        RECT 52.080 93.510 52.340 93.830 ;
        RECT 51.620 91.470 51.880 91.790 ;
        RECT 51.160 89.090 51.420 89.410 ;
        RECT 50.700 82.970 50.960 83.290 ;
        RECT 49.780 82.630 50.040 82.950 ;
        RECT 50.240 82.290 50.500 82.610 ;
        RECT 49.780 81.950 50.040 82.270 ;
        RECT 49.840 80.230 49.980 81.950 ;
        RECT 50.300 80.765 50.440 82.290 ;
        RECT 50.760 80.910 50.900 82.970 ;
        RECT 50.230 80.395 50.510 80.765 ;
        RECT 50.700 80.590 50.960 80.910 ;
        RECT 49.780 79.910 50.040 80.230 ;
        RECT 50.700 79.910 50.960 80.230 ;
        RECT 49.780 79.230 50.040 79.550 ;
        RECT 50.240 79.230 50.500 79.550 ;
        RECT 49.840 78.530 49.980 79.230 ;
        RECT 49.780 78.210 50.040 78.530 ;
        RECT 49.770 77.675 50.050 78.045 ;
        RECT 49.840 77.510 49.980 77.675 ;
        RECT 49.780 77.190 50.040 77.510 ;
        RECT 49.320 75.490 49.580 75.810 ;
        RECT 49.380 74.450 49.520 75.490 ;
        RECT 49.320 74.130 49.580 74.450 ;
        RECT 49.840 72.410 49.980 77.190 ;
        RECT 49.780 72.090 50.040 72.410 ;
        RECT 48.850 71.555 49.130 71.925 ;
        RECT 47.480 69.370 47.740 69.690 ;
        RECT 48.400 66.310 48.660 66.630 ;
        RECT 45.640 63.590 45.900 63.910 ;
        RECT 46.560 63.590 46.820 63.910 ;
        RECT 45.700 62.210 45.840 63.590 ;
        RECT 45.640 61.890 45.900 62.210 ;
        RECT 45.630 61.355 45.910 61.725 ;
        RECT 45.700 61.190 45.840 61.355 ;
        RECT 45.640 60.870 45.900 61.190 ;
        RECT 43.340 60.190 43.600 60.510 ;
        RECT 45.180 60.190 45.440 60.510 ;
        RECT 43.400 59.490 43.540 60.190 ;
        RECT 43.340 59.170 43.600 59.490 ;
        RECT 44.260 58.150 44.520 58.470 ;
        RECT 42.880 56.450 43.140 56.770 ;
        RECT 44.320 55.410 44.460 58.150 ;
        RECT 44.720 56.450 44.980 56.770 ;
        RECT 44.260 55.090 44.520 55.410 ;
        RECT 40.580 54.750 40.840 55.070 ;
        RECT 43.800 54.750 44.060 55.070 ;
        RECT 40.640 52.090 40.780 54.750 ;
        RECT 43.340 53.390 43.600 53.710 ;
        RECT 42.880 52.710 43.140 53.030 ;
        RECT 41.040 52.370 41.300 52.690 ;
        RECT 39.720 51.950 40.780 52.090 ;
        RECT 39.720 51.330 39.860 51.950 ;
        RECT 39.660 51.010 39.920 51.330 ;
        RECT 40.580 50.670 40.840 50.990 ;
        RECT 40.640 42.830 40.780 50.670 ;
        RECT 40.580 42.510 40.840 42.830 ;
        RECT 41.100 36.710 41.240 52.370 ;
        RECT 42.420 52.030 42.680 52.350 ;
        RECT 42.480 50.650 42.620 52.030 ;
        RECT 42.420 50.330 42.680 50.650 ;
        RECT 42.940 50.310 43.080 52.710 ;
        RECT 43.400 51.330 43.540 53.390 ;
        RECT 43.860 51.330 44.000 54.750 ;
        RECT 44.260 52.710 44.520 53.030 ;
        RECT 43.340 51.010 43.600 51.330 ;
        RECT 43.800 51.010 44.060 51.330 ;
        RECT 41.500 49.990 41.760 50.310 ;
        RECT 42.880 49.990 43.140 50.310 ;
        RECT 41.560 45.210 41.700 49.990 ;
        RECT 42.940 49.370 43.080 49.990 ;
        RECT 42.480 49.230 43.080 49.370 ;
        RECT 41.960 47.270 42.220 47.590 ;
        RECT 42.020 45.890 42.160 47.270 ;
        RECT 41.960 45.570 42.220 45.890 ;
        RECT 41.500 44.890 41.760 45.210 ;
        RECT 41.960 44.210 42.220 44.530 ;
        RECT 41.500 43.870 41.760 44.190 ;
        RECT 41.560 37.050 41.700 43.870 ;
        RECT 42.020 40.450 42.160 44.210 ;
        RECT 42.480 43.170 42.620 49.230 ;
        RECT 42.880 48.290 43.140 48.610 ;
        RECT 42.940 45.890 43.080 48.290 ;
        RECT 43.400 47.930 43.540 51.010 ;
        RECT 43.800 49.310 44.060 49.630 ;
        RECT 43.340 47.610 43.600 47.930 ;
        RECT 42.880 45.570 43.140 45.890 ;
        RECT 42.420 43.080 42.680 43.170 ;
        RECT 42.420 42.940 43.080 43.080 ;
        RECT 42.420 42.850 42.680 42.940 ;
        RECT 42.420 42.170 42.680 42.490 ;
        RECT 41.960 40.130 42.220 40.450 ;
        RECT 42.480 37.730 42.620 42.170 ;
        RECT 42.940 39.770 43.080 42.940 ;
        RECT 42.880 39.450 43.140 39.770 ;
        RECT 42.420 37.410 42.680 37.730 ;
        RECT 43.860 37.050 44.000 49.310 ;
        RECT 41.500 36.730 41.760 37.050 ;
        RECT 43.800 36.730 44.060 37.050 ;
        RECT 41.040 36.390 41.300 36.710 ;
        RECT 43.340 36.450 43.600 36.710 ;
        RECT 44.320 36.450 44.460 52.710 ;
        RECT 44.780 40.450 44.920 56.450 ;
        RECT 45.240 55.410 45.380 60.190 ;
        RECT 46.560 58.490 46.820 58.810 ;
        RECT 47.480 58.490 47.740 58.810 ;
        RECT 46.100 57.645 46.360 57.790 ;
        RECT 46.090 57.275 46.370 57.645 ;
        RECT 45.640 56.450 45.900 56.770 ;
        RECT 45.180 55.090 45.440 55.410 ;
        RECT 45.700 55.070 45.840 56.450 ;
        RECT 46.100 55.490 46.360 55.750 ;
        RECT 46.620 55.490 46.760 58.490 ;
        RECT 47.540 55.750 47.680 58.490 ;
        RECT 48.460 56.430 48.600 66.310 ;
        RECT 48.920 65.950 49.060 71.555 ;
        RECT 49.310 66.795 49.590 67.165 ;
        RECT 49.380 66.630 49.520 66.795 ;
        RECT 49.840 66.630 49.980 72.090 ;
        RECT 49.320 66.310 49.580 66.630 ;
        RECT 49.780 66.310 50.040 66.630 ;
        RECT 48.860 65.630 49.120 65.950 ;
        RECT 48.920 61.530 49.060 65.630 ;
        RECT 49.780 63.590 50.040 63.910 ;
        RECT 49.320 63.250 49.580 63.570 ;
        RECT 49.380 61.725 49.520 63.250 ;
        RECT 48.860 61.210 49.120 61.530 ;
        RECT 49.310 61.355 49.590 61.725 ;
        RECT 49.380 59.150 49.520 61.355 ;
        RECT 49.320 58.830 49.580 59.150 ;
        RECT 49.840 57.790 49.980 63.590 ;
        RECT 50.300 61.190 50.440 79.230 ;
        RECT 50.760 77.510 50.900 79.910 ;
        RECT 50.700 77.190 50.960 77.510 ;
        RECT 50.700 74.130 50.960 74.450 ;
        RECT 50.760 69.690 50.900 74.130 ;
        RECT 51.220 70.030 51.360 89.090 ;
        RECT 51.620 86.030 51.880 86.350 ;
        RECT 51.680 79.550 51.820 86.030 ;
        RECT 52.140 82.950 52.280 93.510 ;
        RECT 52.600 92.130 52.740 98.270 ;
        RECT 53.060 96.210 53.200 104.390 ;
        RECT 53.520 98.930 53.660 115.270 ;
        RECT 53.920 112.890 54.180 113.210 ;
        RECT 53.980 111.170 54.120 112.890 ;
        RECT 53.920 110.850 54.180 111.170 ;
        RECT 53.920 109.150 54.180 109.470 ;
        RECT 53.980 107.770 54.120 109.150 ;
        RECT 54.440 108.450 54.580 139.750 ;
        RECT 55.820 137.690 55.960 139.750 ;
        RECT 55.760 137.370 56.020 137.690 ;
        RECT 56.280 136.670 56.420 142.955 ;
        RECT 56.220 136.350 56.480 136.670 ;
        RECT 56.220 133.970 56.480 134.290 ;
        RECT 55.290 132.755 55.570 133.125 ;
        RECT 54.840 128.530 55.100 128.850 ;
        RECT 54.900 124.965 55.040 128.530 ;
        RECT 55.360 127.490 55.500 132.755 ;
        RECT 55.300 127.170 55.560 127.490 ;
        RECT 56.280 126.470 56.420 133.970 ;
        RECT 56.740 126.810 56.880 150.630 ;
        RECT 57.200 148.230 57.340 158.710 ;
        RECT 57.600 158.110 57.860 158.430 ;
        RECT 57.660 151.970 57.800 158.110 ;
        RECT 57.600 151.650 57.860 151.970 ;
        RECT 58.580 148.230 58.720 159.275 ;
        RECT 59.960 156.130 60.100 160.635 ;
        RECT 60.420 157.410 60.560 161.510 ;
        RECT 60.360 157.090 60.620 157.410 ;
        RECT 59.960 155.990 60.560 156.130 ;
        RECT 59.440 155.390 59.700 155.710 ;
        RECT 59.900 155.390 60.160 155.710 ;
        RECT 59.500 154.690 59.640 155.390 ;
        RECT 59.440 154.370 59.700 154.690 ;
        RECT 58.980 153.010 59.240 153.330 ;
        RECT 59.040 148.910 59.180 153.010 ;
        RECT 59.500 151.970 59.640 154.370 ;
        RECT 59.440 151.650 59.700 151.970 ;
        RECT 59.960 151.370 60.100 155.390 ;
        RECT 59.500 151.230 60.100 151.370 ;
        RECT 58.980 148.590 59.240 148.910 ;
        RECT 57.140 147.910 57.400 148.230 ;
        RECT 58.060 147.910 58.320 148.230 ;
        RECT 58.520 147.910 58.780 148.230 ;
        RECT 58.120 147.405 58.260 147.910 ;
        RECT 58.050 147.035 58.330 147.405 ;
        RECT 58.060 146.210 58.320 146.530 ;
        RECT 57.600 144.510 57.860 144.830 ;
        RECT 57.660 142.790 57.800 144.510 ;
        RECT 58.120 142.790 58.260 146.210 ;
        RECT 57.600 142.470 57.860 142.790 ;
        RECT 58.060 142.470 58.320 142.790 ;
        RECT 58.120 138.370 58.260 142.470 ;
        RECT 58.060 138.050 58.320 138.370 ;
        RECT 59.500 137.690 59.640 151.230 ;
        RECT 60.420 147.290 60.560 155.990 ;
        RECT 60.820 149.950 61.080 150.270 ;
        RECT 60.880 148.230 61.020 149.950 ;
        RECT 61.340 148.910 61.480 163.550 ;
        RECT 62.650 163.355 62.930 163.725 ;
        RECT 65.880 163.550 66.140 163.870 ;
        RECT 61.740 156.410 62.000 156.730 ;
        RECT 61.800 151.970 61.940 156.410 ;
        RECT 62.200 152.670 62.460 152.990 ;
        RECT 61.740 151.650 62.000 151.970 ;
        RECT 61.740 150.290 62.000 150.610 ;
        RECT 61.280 148.590 61.540 148.910 ;
        RECT 61.800 148.570 61.940 150.290 ;
        RECT 61.740 148.250 62.000 148.570 ;
        RECT 60.820 147.910 61.080 148.230 ;
        RECT 60.420 147.150 61.940 147.290 ;
        RECT 61.280 145.190 61.540 145.510 ;
        RECT 61.340 142.790 61.480 145.190 ;
        RECT 61.280 142.470 61.540 142.790 ;
        RECT 59.900 140.770 60.160 141.090 ;
        RECT 59.440 137.370 59.700 137.690 ;
        RECT 59.440 136.350 59.700 136.670 ;
        RECT 58.970 131.395 59.250 131.765 ;
        RECT 59.040 131.230 59.180 131.395 ;
        RECT 58.980 130.910 59.240 131.230 ;
        RECT 58.520 129.210 58.780 129.530 ;
        RECT 56.680 126.490 56.940 126.810 ;
        RECT 56.220 126.150 56.480 126.470 ;
        RECT 54.830 124.595 55.110 124.965 ;
        RECT 56.740 124.770 56.880 126.490 ;
        RECT 56.680 124.450 56.940 124.770 ;
        RECT 56.220 123.770 56.480 124.090 ;
        RECT 58.060 123.770 58.320 124.090 ;
        RECT 55.300 121.390 55.560 121.710 ;
        RECT 54.840 120.090 55.100 120.350 ;
        RECT 55.360 120.090 55.500 121.390 ;
        RECT 54.840 120.030 55.500 120.090 ;
        RECT 55.760 120.030 56.020 120.350 ;
        RECT 54.900 119.950 55.500 120.030 ;
        RECT 54.840 117.990 55.100 118.310 ;
        RECT 54.900 115.590 55.040 117.990 ;
        RECT 55.300 117.310 55.560 117.630 ;
        RECT 55.360 116.610 55.500 117.310 ;
        RECT 55.300 116.290 55.560 116.610 ;
        RECT 54.840 115.270 55.100 115.590 ;
        RECT 55.360 113.550 55.500 116.290 ;
        RECT 55.820 114.910 55.960 120.030 ;
        RECT 56.280 117.970 56.420 123.770 ;
        RECT 57.600 123.430 57.860 123.750 ;
        RECT 57.140 122.750 57.400 123.070 ;
        RECT 57.200 121.370 57.340 122.750 ;
        RECT 57.140 121.050 57.400 121.370 ;
        RECT 56.680 120.710 56.940 121.030 ;
        RECT 56.740 120.350 56.880 120.710 ;
        RECT 56.680 120.030 56.940 120.350 ;
        RECT 57.140 120.030 57.400 120.350 ;
        RECT 57.200 119.240 57.340 120.030 ;
        RECT 56.740 119.100 57.340 119.240 ;
        RECT 56.220 117.650 56.480 117.970 ;
        RECT 56.210 117.115 56.490 117.485 ;
        RECT 56.280 116.610 56.420 117.115 ;
        RECT 56.220 116.290 56.480 116.610 ;
        RECT 56.740 116.010 56.880 119.100 ;
        RECT 57.660 118.990 57.800 123.430 ;
        RECT 57.600 118.670 57.860 118.990 ;
        RECT 57.140 118.330 57.400 118.650 ;
        RECT 56.280 115.870 56.880 116.010 ;
        RECT 56.280 115.590 56.420 115.870 ;
        RECT 56.220 115.270 56.480 115.590 ;
        RECT 56.680 115.270 56.940 115.590 ;
        RECT 55.760 114.590 56.020 114.910 ;
        RECT 55.300 113.230 55.560 113.550 ;
        RECT 54.840 112.890 55.100 113.210 ;
        RECT 54.380 108.130 54.640 108.450 ;
        RECT 53.920 107.450 54.180 107.770 ;
        RECT 54.440 105.390 54.580 108.130 ;
        RECT 54.380 105.070 54.640 105.390 ;
        RECT 53.920 104.390 54.180 104.710 ;
        RECT 53.980 100.290 54.120 104.390 ;
        RECT 54.900 104.370 55.040 112.890 ;
        RECT 55.820 107.430 55.960 114.590 ;
        RECT 56.220 107.790 56.480 108.110 ;
        RECT 55.760 107.110 56.020 107.430 ;
        RECT 54.840 104.050 55.100 104.370 ;
        RECT 55.300 103.710 55.560 104.030 ;
        RECT 55.360 102.330 55.500 103.710 ;
        RECT 55.300 102.010 55.560 102.330 ;
        RECT 54.380 101.670 54.640 101.990 ;
        RECT 53.920 99.970 54.180 100.290 ;
        RECT 53.920 98.950 54.180 99.270 ;
        RECT 53.460 98.610 53.720 98.930 ;
        RECT 53.520 97.570 53.660 98.610 ;
        RECT 53.460 97.250 53.720 97.570 ;
        RECT 53.460 96.570 53.720 96.890 ;
        RECT 53.000 95.890 53.260 96.210 ;
        RECT 53.000 93.170 53.260 93.490 ;
        RECT 52.540 91.810 52.800 92.130 ;
        RECT 52.600 83.630 52.740 91.810 ;
        RECT 53.060 91.450 53.200 93.170 ;
        RECT 53.520 93.150 53.660 96.570 ;
        RECT 53.460 92.830 53.720 93.150 ;
        RECT 53.000 91.130 53.260 91.450 ;
        RECT 53.060 90.430 53.200 91.130 ;
        RECT 53.460 90.790 53.720 91.110 ;
        RECT 53.000 90.110 53.260 90.430 ;
        RECT 53.520 85.670 53.660 90.790 ;
        RECT 53.980 86.690 54.120 98.950 ;
        RECT 54.440 97.570 54.580 101.670 ;
        RECT 55.300 101.330 55.560 101.650 ;
        RECT 54.840 100.990 55.100 101.310 ;
        RECT 54.380 97.250 54.640 97.570 ;
        RECT 54.440 94.170 54.580 97.250 ;
        RECT 54.380 93.850 54.640 94.170 ;
        RECT 54.900 93.740 55.040 100.990 ;
        RECT 55.360 99.270 55.500 101.330 ;
        RECT 55.300 98.950 55.560 99.270 ;
        RECT 55.300 98.270 55.560 98.590 ;
        RECT 55.360 97.570 55.500 98.270 ;
        RECT 55.300 97.250 55.560 97.570 ;
        RECT 55.820 96.890 55.960 107.110 ;
        RECT 56.280 103.010 56.420 107.790 ;
        RECT 56.740 107.430 56.880 115.270 ;
        RECT 57.200 107.770 57.340 118.330 ;
        RECT 57.660 113.210 57.800 118.670 ;
        RECT 58.120 116.610 58.260 123.770 ;
        RECT 58.580 121.030 58.720 129.210 ;
        RECT 59.500 128.510 59.640 136.350 ;
        RECT 59.960 132.590 60.100 140.770 ;
        RECT 61.340 140.750 61.480 142.470 ;
        RECT 61.280 140.430 61.540 140.750 ;
        RECT 61.280 138.050 61.540 138.370 ;
        RECT 61.340 135.650 61.480 138.050 ;
        RECT 61.280 135.330 61.540 135.650 ;
        RECT 59.900 132.330 60.160 132.590 ;
        RECT 59.900 132.270 60.560 132.330 ;
        RECT 59.960 132.190 60.560 132.270 ;
        RECT 60.420 129.870 60.560 132.190 ;
        RECT 60.360 129.550 60.620 129.870 ;
        RECT 59.440 128.190 59.700 128.510 ;
        RECT 59.900 126.490 60.160 126.810 ;
        RECT 59.960 121.710 60.100 126.490 ;
        RECT 60.360 125.470 60.620 125.790 ;
        RECT 60.820 125.470 61.080 125.790 ;
        RECT 61.280 125.470 61.540 125.790 ;
        RECT 59.900 121.390 60.160 121.710 ;
        RECT 58.520 120.940 58.780 121.030 ;
        RECT 58.520 120.800 59.180 120.940 ;
        RECT 58.520 120.710 58.780 120.800 ;
        RECT 58.520 120.030 58.780 120.350 ;
        RECT 58.580 117.485 58.720 120.030 ;
        RECT 58.510 117.115 58.790 117.485 ;
        RECT 58.060 116.290 58.320 116.610 ;
        RECT 58.060 115.650 58.320 115.970 ;
        RECT 57.600 112.890 57.860 113.210 ;
        RECT 57.660 109.810 57.800 112.890 ;
        RECT 58.120 111.170 58.260 115.650 ;
        RECT 58.060 110.850 58.320 111.170 ;
        RECT 58.580 110.470 58.720 117.115 ;
        RECT 59.040 116.805 59.180 120.800 ;
        RECT 59.890 120.515 60.170 120.885 ;
        RECT 59.960 118.990 60.100 120.515 ;
        RECT 59.900 118.670 60.160 118.990 ;
        RECT 59.440 118.330 59.700 118.650 ;
        RECT 58.970 116.435 59.250 116.805 ;
        RECT 59.500 116.610 59.640 118.330 ;
        RECT 59.440 116.290 59.700 116.610 ;
        RECT 59.960 116.010 60.100 118.670 ;
        RECT 60.420 118.650 60.560 125.470 ;
        RECT 60.880 122.925 61.020 125.470 ;
        RECT 60.810 122.555 61.090 122.925 ;
        RECT 61.340 122.050 61.480 125.470 ;
        RECT 61.800 124.090 61.940 147.150 ;
        RECT 62.260 131.765 62.400 152.670 ;
        RECT 62.720 147.550 62.860 163.355 ;
        RECT 63.120 161.170 63.380 161.490 ;
        RECT 63.180 153.670 63.320 161.170 ;
        RECT 65.420 158.450 65.680 158.770 ;
        RECT 64.960 156.410 65.220 156.730 ;
        RECT 63.580 153.690 63.840 154.010 ;
        RECT 63.120 153.350 63.380 153.670 ;
        RECT 63.640 150.950 63.780 153.690 ;
        RECT 64.040 153.010 64.300 153.330 ;
        RECT 64.100 151.630 64.240 153.010 ;
        RECT 64.040 151.310 64.300 151.630 ;
        RECT 63.580 150.630 63.840 150.950 ;
        RECT 65.020 149.250 65.160 156.410 ;
        RECT 65.480 153.330 65.620 158.450 ;
        RECT 65.420 153.010 65.680 153.330 ;
        RECT 65.940 150.950 66.080 163.550 ;
        RECT 66.860 162.850 67.000 163.890 ;
        RECT 67.320 162.850 67.460 163.890 ;
        RECT 66.800 162.530 67.060 162.850 ;
        RECT 67.260 162.530 67.520 162.850 ;
        RECT 66.340 152.670 66.600 152.990 ;
        RECT 66.400 151.970 66.540 152.670 ;
        RECT 66.340 151.650 66.600 151.970 ;
        RECT 65.420 150.630 65.680 150.950 ;
        RECT 65.880 150.630 66.140 150.950 ;
        RECT 64.960 148.930 65.220 149.250 ;
        RECT 65.480 148.570 65.620 150.630 ;
        RECT 63.580 148.250 63.840 148.570 ;
        RECT 65.420 148.250 65.680 148.570 ;
        RECT 66.340 148.250 66.600 148.570 ;
        RECT 62.660 147.230 62.920 147.550 ;
        RECT 63.120 147.230 63.380 147.550 ;
        RECT 63.180 146.190 63.320 147.230 ;
        RECT 63.120 145.870 63.380 146.190 ;
        RECT 63.120 140.090 63.380 140.410 ;
        RECT 63.180 135.650 63.320 140.090 ;
        RECT 63.120 135.330 63.380 135.650 ;
        RECT 63.640 135.050 63.780 148.250 ;
        RECT 66.400 147.550 66.540 148.250 ;
        RECT 64.500 147.230 64.760 147.550 ;
        RECT 66.340 147.230 66.600 147.550 ;
        RECT 64.040 141.790 64.300 142.110 ;
        RECT 64.100 137.690 64.240 141.790 ;
        RECT 64.040 137.370 64.300 137.690 ;
        RECT 63.180 134.910 63.780 135.050 ;
        RECT 63.180 134.630 63.320 134.910 ;
        RECT 63.120 134.310 63.380 134.630 ;
        RECT 62.190 131.395 62.470 131.765 ;
        RECT 63.180 127.490 63.320 134.310 ;
        RECT 64.030 132.075 64.310 132.445 ;
        RECT 63.120 127.170 63.380 127.490 ;
        RECT 61.740 123.770 62.000 124.090 ;
        RECT 63.180 123.750 63.320 127.170 ;
        RECT 63.120 123.430 63.380 123.750 ;
        RECT 61.280 121.730 61.540 122.050 ;
        RECT 60.820 121.050 61.080 121.370 ;
        RECT 60.880 120.885 61.020 121.050 ;
        RECT 60.810 120.515 61.090 120.885 ;
        RECT 61.280 120.710 61.540 121.030 ;
        RECT 60.360 118.330 60.620 118.650 ;
        RECT 60.360 117.650 60.620 117.970 ;
        RECT 60.420 116.610 60.560 117.650 ;
        RECT 60.360 116.290 60.620 116.610 ;
        RECT 58.980 115.610 59.240 115.930 ;
        RECT 59.500 115.870 60.100 116.010 ;
        RECT 61.340 116.010 61.480 120.710 ;
        RECT 62.660 120.370 62.920 120.690 ;
        RECT 62.720 118.650 62.860 120.370 ;
        RECT 62.660 118.330 62.920 118.650 ;
        RECT 59.040 112.190 59.180 115.610 ;
        RECT 58.980 111.870 59.240 112.190 ;
        RECT 59.500 110.830 59.640 115.870 ;
        RECT 60.360 115.610 60.620 115.930 ;
        RECT 61.340 115.870 61.940 116.010 ;
        RECT 59.900 115.270 60.160 115.590 ;
        RECT 59.960 114.910 60.100 115.270 ;
        RECT 59.900 114.590 60.160 114.910 ;
        RECT 60.420 114.085 60.560 115.610 ;
        RECT 61.280 115.445 61.540 115.590 ;
        RECT 60.820 114.930 61.080 115.250 ;
        RECT 61.270 115.075 61.550 115.445 ;
        RECT 60.880 114.765 61.020 114.930 ;
        RECT 60.810 114.395 61.090 114.765 ;
        RECT 60.350 113.715 60.630 114.085 ;
        RECT 60.820 113.570 61.080 113.890 ;
        RECT 59.440 110.510 59.700 110.830 ;
        RECT 58.120 110.330 58.720 110.470 ;
        RECT 60.360 110.400 60.620 110.490 ;
        RECT 60.880 110.400 61.020 113.570 ;
        RECT 57.600 109.490 57.860 109.810 ;
        RECT 57.140 107.450 57.400 107.770 ;
        RECT 57.600 107.450 57.860 107.770 ;
        RECT 56.680 107.110 56.940 107.430 ;
        RECT 56.220 102.690 56.480 103.010 ;
        RECT 56.680 102.350 56.940 102.670 ;
        RECT 56.220 99.290 56.480 99.610 ;
        RECT 55.760 96.570 56.020 96.890 ;
        RECT 55.820 94.510 55.960 96.570 ;
        RECT 55.760 94.190 56.020 94.510 ;
        RECT 56.280 93.830 56.420 99.290 ;
        RECT 56.740 96.890 56.880 102.350 ;
        RECT 57.200 99.270 57.340 107.450 ;
        RECT 57.660 104.620 57.800 107.450 ;
        RECT 58.120 105.390 58.260 110.330 ;
        RECT 60.360 110.260 61.020 110.400 ;
        RECT 60.360 110.170 60.620 110.260 ;
        RECT 58.520 109.830 58.780 110.150 ;
        RECT 58.580 107.770 58.720 109.830 ;
        RECT 59.900 109.490 60.160 109.810 ;
        RECT 58.520 107.450 58.780 107.770 ;
        RECT 58.580 105.730 58.720 107.450 ;
        RECT 59.960 107.430 60.100 109.490 ;
        RECT 60.360 108.130 60.620 108.450 ;
        RECT 59.440 107.170 59.700 107.430 ;
        RECT 59.040 107.110 59.700 107.170 ;
        RECT 59.900 107.110 60.160 107.430 ;
        RECT 59.040 107.030 59.640 107.110 ;
        RECT 58.520 105.410 58.780 105.730 ;
        RECT 58.060 105.070 58.320 105.390 ;
        RECT 58.520 104.620 58.780 104.710 ;
        RECT 57.660 104.480 58.780 104.620 ;
        RECT 58.520 104.390 58.780 104.480 ;
        RECT 57.600 99.970 57.860 100.290 ;
        RECT 57.140 98.950 57.400 99.270 ;
        RECT 57.140 98.270 57.400 98.590 ;
        RECT 56.680 96.570 56.940 96.890 ;
        RECT 55.300 93.740 55.560 93.830 ;
        RECT 56.220 93.740 56.480 93.830 ;
        RECT 54.900 93.600 55.560 93.740 ;
        RECT 55.300 93.510 55.560 93.600 ;
        RECT 55.820 93.600 56.480 93.740 ;
        RECT 54.380 92.830 54.640 93.150 ;
        RECT 53.920 86.370 54.180 86.690 ;
        RECT 53.460 85.350 53.720 85.670 ;
        RECT 54.440 83.970 54.580 92.830 ;
        RECT 54.840 90.110 55.100 90.430 ;
        RECT 54.380 83.650 54.640 83.970 ;
        RECT 52.540 83.310 52.800 83.630 ;
        RECT 52.080 82.630 52.340 82.950 ;
        RECT 53.920 82.630 54.180 82.950 ;
        RECT 52.080 81.950 52.340 82.270 ;
        RECT 53.000 81.950 53.260 82.270 ;
        RECT 51.620 79.230 51.880 79.550 ;
        RECT 52.140 77.510 52.280 81.950 ;
        RECT 53.060 80.230 53.200 81.950 ;
        RECT 53.460 80.250 53.720 80.570 ;
        RECT 53.000 79.910 53.260 80.230 ;
        RECT 52.540 78.210 52.800 78.530 ;
        RECT 52.600 77.510 52.740 78.210 ;
        RECT 53.060 78.190 53.200 79.910 ;
        RECT 53.000 77.870 53.260 78.190 ;
        RECT 51.620 77.190 51.880 77.510 ;
        RECT 52.080 77.190 52.340 77.510 ;
        RECT 52.540 77.190 52.800 77.510 ;
        RECT 53.000 77.190 53.260 77.510 ;
        RECT 51.680 76.830 51.820 77.190 ;
        RECT 51.620 76.510 51.880 76.830 ;
        RECT 53.060 76.685 53.200 77.190 ;
        RECT 51.680 74.360 51.820 76.510 ;
        RECT 52.990 76.315 53.270 76.685 ;
        RECT 53.520 75.810 53.660 80.250 ;
        RECT 53.980 79.550 54.120 82.630 ;
        RECT 54.440 80.230 54.580 83.650 ;
        RECT 54.380 79.910 54.640 80.230 ;
        RECT 53.920 79.230 54.180 79.550 ;
        RECT 53.980 77.850 54.120 79.230 ;
        RECT 54.380 77.870 54.640 78.190 ;
        RECT 53.920 77.530 54.180 77.850 ;
        RECT 53.980 75.810 54.120 77.530 ;
        RECT 54.440 75.810 54.580 77.870 ;
        RECT 54.900 77.510 55.040 90.110 ;
        RECT 55.360 81.250 55.500 93.510 ;
        RECT 55.820 85.330 55.960 93.600 ;
        RECT 56.220 93.510 56.480 93.600 ;
        RECT 57.200 93.490 57.340 98.270 ;
        RECT 57.140 93.170 57.400 93.490 ;
        RECT 57.660 91.450 57.800 99.970 ;
        RECT 58.580 98.930 58.720 104.390 ;
        RECT 58.520 98.610 58.780 98.930 ;
        RECT 58.060 98.270 58.320 98.590 ;
        RECT 58.120 97.570 58.260 98.270 ;
        RECT 58.060 97.250 58.320 97.570 ;
        RECT 58.120 93.830 58.260 97.250 ;
        RECT 58.520 96.800 58.780 96.890 ;
        RECT 59.040 96.800 59.180 107.030 ;
        RECT 59.440 106.430 59.700 106.750 ;
        RECT 59.500 104.710 59.640 106.430 ;
        RECT 59.440 104.390 59.700 104.710 ;
        RECT 58.520 96.660 59.180 96.800 ;
        RECT 58.520 96.570 58.780 96.660 ;
        RECT 59.440 96.570 59.700 96.890 ;
        RECT 58.580 94.850 58.720 96.570 ;
        RECT 59.500 94.850 59.640 96.570 ;
        RECT 58.520 94.530 58.780 94.850 ;
        RECT 59.440 94.530 59.700 94.850 ;
        RECT 58.060 93.510 58.320 93.830 ;
        RECT 58.520 92.830 58.780 93.150 ;
        RECT 57.600 91.360 57.860 91.450 ;
        RECT 57.200 91.220 57.860 91.360 ;
        RECT 56.210 89.235 56.490 89.605 ;
        RECT 55.760 85.010 56.020 85.330 ;
        RECT 55.760 82.290 56.020 82.610 ;
        RECT 55.300 80.930 55.560 81.250 ;
        RECT 54.840 77.190 55.100 77.510 ;
        RECT 55.290 76.995 55.570 77.365 ;
        RECT 54.840 76.510 55.100 76.830 ;
        RECT 53.460 75.490 53.720 75.810 ;
        RECT 53.920 75.490 54.180 75.810 ;
        RECT 54.380 75.490 54.640 75.810 ;
        RECT 52.540 75.150 52.800 75.470 ;
        RECT 52.080 74.360 52.340 74.450 ;
        RECT 51.680 74.220 52.340 74.360 ;
        RECT 52.080 74.130 52.340 74.220 ;
        RECT 52.600 73.090 52.740 75.150 ;
        RECT 53.000 74.810 53.260 75.130 ;
        RECT 53.060 74.110 53.200 74.810 ;
        RECT 53.000 73.790 53.260 74.110 ;
        RECT 52.540 72.770 52.800 73.090 ;
        RECT 52.600 70.370 52.740 72.770 ;
        RECT 53.000 72.430 53.260 72.750 ;
        RECT 53.060 70.450 53.200 72.430 ;
        RECT 53.520 71.390 53.660 75.490 ;
        RECT 53.920 74.810 54.180 75.130 ;
        RECT 53.980 73.090 54.120 74.810 ;
        RECT 54.380 74.130 54.640 74.450 ;
        RECT 53.920 72.770 54.180 73.090 ;
        RECT 53.460 71.070 53.720 71.390 ;
        RECT 54.440 70.450 54.580 74.130 ;
        RECT 52.540 70.050 52.800 70.370 ;
        RECT 53.060 70.310 54.580 70.450 ;
        RECT 51.160 69.710 51.420 70.030 ;
        RECT 50.700 69.370 50.960 69.690 ;
        RECT 50.240 60.870 50.500 61.190 ;
        RECT 49.780 57.470 50.040 57.790 ;
        RECT 48.400 56.110 48.660 56.430 ;
        RECT 51.220 55.750 51.360 69.710 ;
        RECT 53.060 69.690 53.200 70.310 ;
        RECT 53.000 69.370 53.260 69.690 ;
        RECT 52.540 69.030 52.800 69.350 ;
        RECT 52.600 56.770 52.740 69.030 ;
        RECT 53.060 66.630 53.200 69.370 ;
        RECT 53.920 69.030 54.180 69.350 ;
        RECT 53.000 66.310 53.260 66.630 ;
        RECT 53.460 66.310 53.720 66.630 ;
        RECT 53.520 64.930 53.660 66.310 ;
        RECT 53.460 64.610 53.720 64.930 ;
        RECT 53.520 62.210 53.660 64.610 ;
        RECT 53.980 64.590 54.120 69.030 ;
        RECT 53.920 64.270 54.180 64.590 ;
        RECT 53.460 61.890 53.720 62.210 ;
        RECT 53.460 60.190 53.720 60.510 ;
        RECT 53.520 58.890 53.660 60.190 ;
        RECT 53.980 59.490 54.120 64.270 ;
        RECT 53.920 59.170 54.180 59.490 ;
        RECT 53.520 58.750 54.120 58.890 ;
        RECT 52.540 56.450 52.800 56.770 ;
        RECT 46.100 55.430 46.760 55.490 ;
        RECT 47.480 55.430 47.740 55.750 ;
        RECT 51.160 55.430 51.420 55.750 ;
        RECT 46.160 55.350 46.760 55.430 ;
        RECT 45.640 54.750 45.900 55.070 ;
        RECT 45.180 53.050 45.440 53.370 ;
        RECT 45.240 48.610 45.380 53.050 ;
        RECT 45.640 52.030 45.900 52.350 ;
        RECT 45.700 50.310 45.840 52.030 ;
        RECT 45.640 49.990 45.900 50.310 ;
        RECT 45.180 48.290 45.440 48.610 ;
        RECT 45.700 46.650 45.840 49.990 ;
        RECT 46.100 46.650 46.360 46.910 ;
        RECT 45.700 46.590 46.360 46.650 ;
        RECT 45.700 46.510 46.300 46.590 ;
        RECT 45.180 44.100 45.440 44.190 ;
        RECT 45.700 44.100 45.840 46.510 ;
        RECT 45.180 43.960 45.840 44.100 ;
        RECT 45.180 43.870 45.440 43.960 ;
        RECT 44.720 40.130 44.980 40.450 ;
        RECT 43.340 36.390 44.460 36.450 ;
        RECT 43.400 36.310 44.460 36.390 ;
        RECT 40.120 35.710 40.380 36.030 ;
        RECT 40.180 33.990 40.320 35.710 ;
        RECT 40.120 33.670 40.380 33.990 ;
        RECT 44.320 32.290 44.460 36.310 ;
        RECT 44.260 31.970 44.520 32.290 ;
        RECT 38.730 30.075 39.010 30.445 ;
        RECT 34.600 29.250 34.860 29.570 ;
        RECT 27.700 27.550 27.960 27.870 ;
        RECT 24.370 27.015 25.910 27.385 ;
        RECT 21.070 24.295 22.610 24.665 ;
        RECT 24.370 21.575 25.910 21.945 ;
        RECT 21.070 18.855 22.610 19.225 ;
        RECT 24.370 16.135 25.910 16.505 ;
        RECT 27.760 15.290 27.900 27.550 ;
        RECT 44.780 24.130 44.920 40.130 ;
        RECT 45.640 38.770 45.900 39.090 ;
        RECT 45.700 34.330 45.840 38.770 ;
        RECT 45.640 34.010 45.900 34.330 ;
        RECT 46.100 26.190 46.360 26.510 ;
        RECT 44.720 23.810 44.980 24.130 ;
        RECT 45.640 23.130 45.900 23.450 ;
        RECT 44.260 22.790 44.520 23.110 ;
        RECT 44.320 21.070 44.460 22.790 ;
        RECT 44.260 20.750 44.520 21.070 ;
        RECT 43.790 19.875 44.070 20.245 ;
        RECT 40.120 19.390 40.380 19.710 ;
        RECT 40.180 18.010 40.320 19.390 ;
        RECT 40.120 17.690 40.380 18.010 ;
        RECT 43.860 17.670 44.000 19.875 ;
        RECT 43.800 17.350 44.060 17.670 ;
        RECT 43.800 16.670 44.060 16.990 ;
        RECT 27.700 14.970 27.960 15.290 ;
        RECT 21.070 13.415 22.610 13.785 ;
        RECT 43.860 12.230 44.000 16.670 ;
        RECT 44.320 12.910 44.460 20.750 ;
        RECT 45.700 20.730 45.840 23.130 ;
        RECT 46.160 22.170 46.300 26.190 ;
        RECT 46.620 23.110 46.760 55.350 ;
        RECT 47.020 26.530 47.280 26.850 ;
        RECT 47.080 23.110 47.220 26.530 ;
        RECT 47.540 26.510 47.680 55.430 ;
        RECT 48.860 53.050 49.120 53.370 ;
        RECT 47.940 47.270 48.200 47.590 ;
        RECT 48.000 42.150 48.140 47.270 ;
        RECT 48.920 43.170 49.060 53.050 ;
        RECT 52.540 52.710 52.800 53.030 ;
        RECT 52.600 50.310 52.740 52.710 ;
        RECT 52.540 49.990 52.800 50.310 ;
        RECT 49.320 47.610 49.580 47.930 ;
        RECT 52.080 47.610 52.340 47.930 ;
        RECT 49.380 44.530 49.520 47.610 ;
        RECT 49.320 44.210 49.580 44.530 ;
        RECT 48.860 42.850 49.120 43.170 ;
        RECT 47.940 41.830 48.200 42.150 ;
        RECT 48.000 37.730 48.140 41.830 ;
        RECT 48.920 41.470 49.060 42.850 ;
        RECT 49.380 42.490 49.520 44.210 ;
        RECT 52.140 43.170 52.280 47.610 ;
        RECT 52.080 42.850 52.340 43.170 ;
        RECT 49.320 42.170 49.580 42.490 ;
        RECT 48.860 41.150 49.120 41.470 ;
        RECT 48.920 40.110 49.060 41.150 ;
        RECT 48.860 39.790 49.120 40.110 ;
        RECT 47.940 37.410 48.200 37.730 ;
        RECT 48.400 36.730 48.660 37.050 ;
        RECT 48.460 31.610 48.600 36.730 ;
        RECT 48.920 31.610 49.060 39.790 ;
        RECT 49.380 39.430 49.520 42.170 ;
        RECT 49.320 39.110 49.580 39.430 ;
        RECT 49.380 37.390 49.520 39.110 ;
        RECT 52.080 39.000 52.340 39.090 ;
        RECT 52.600 39.000 52.740 49.990 ;
        RECT 53.980 46.910 54.120 58.750 ;
        RECT 54.900 54.925 55.040 76.510 ;
        RECT 55.360 75.810 55.500 76.995 ;
        RECT 55.300 75.490 55.560 75.810 ;
        RECT 55.360 75.130 55.500 75.490 ;
        RECT 55.300 74.810 55.560 75.130 ;
        RECT 55.820 72.490 55.960 82.290 ;
        RECT 55.360 72.410 55.960 72.490 ;
        RECT 55.300 72.350 55.960 72.410 ;
        RECT 55.300 72.090 55.560 72.350 ;
        RECT 55.360 71.390 55.500 72.090 ;
        RECT 55.300 71.070 55.560 71.390 ;
        RECT 55.360 70.370 55.500 71.070 ;
        RECT 55.300 70.050 55.560 70.370 ;
        RECT 55.360 66.970 55.500 70.050 ;
        RECT 56.280 69.690 56.420 89.235 ;
        RECT 57.200 87.450 57.340 91.220 ;
        RECT 57.600 91.130 57.860 91.220 ;
        RECT 58.580 88.730 58.720 92.830 ;
        RECT 58.520 88.410 58.780 88.730 ;
        RECT 56.740 87.310 57.340 87.450 ;
        RECT 56.740 83.290 56.880 87.310 ;
        RECT 57.140 86.370 57.400 86.690 ;
        RECT 56.680 82.970 56.940 83.290 ;
        RECT 56.740 79.890 56.880 82.970 ;
        RECT 57.200 80.910 57.340 86.370 ;
        RECT 58.060 85.350 58.320 85.670 ;
        RECT 57.590 83.115 57.870 83.485 ;
        RECT 57.660 81.250 57.800 83.115 ;
        RECT 57.600 80.930 57.860 81.250 ;
        RECT 57.140 80.590 57.400 80.910 ;
        RECT 56.680 79.570 56.940 79.890 ;
        RECT 56.680 76.510 56.940 76.830 ;
        RECT 56.740 72.750 56.880 76.510 ;
        RECT 57.200 75.890 57.340 80.590 ;
        RECT 57.600 79.910 57.860 80.230 ;
        RECT 57.660 76.830 57.800 79.910 ;
        RECT 58.120 77.170 58.260 85.350 ;
        RECT 58.980 85.010 59.240 85.330 ;
        RECT 58.520 83.310 58.780 83.630 ;
        RECT 58.580 79.550 58.720 83.310 ;
        RECT 58.520 79.230 58.780 79.550 ;
        RECT 58.580 78.190 58.720 79.230 ;
        RECT 58.520 77.870 58.780 78.190 ;
        RECT 59.040 77.510 59.180 85.010 ;
        RECT 59.440 81.950 59.700 82.270 ;
        RECT 59.500 80.910 59.640 81.950 ;
        RECT 59.440 80.590 59.700 80.910 ;
        RECT 59.500 77.850 59.640 80.590 ;
        RECT 59.440 77.530 59.700 77.850 ;
        RECT 58.980 77.190 59.240 77.510 ;
        RECT 60.420 77.250 60.560 108.130 ;
        RECT 60.880 105.050 61.020 110.260 ;
        RECT 61.280 109.890 61.540 110.150 ;
        RECT 61.800 109.890 61.940 115.870 ;
        RECT 62.200 115.610 62.460 115.930 ;
        RECT 62.260 112.530 62.400 115.610 ;
        RECT 62.650 114.650 62.930 114.765 ;
        RECT 63.180 114.650 63.320 123.430 ;
        RECT 64.100 123.070 64.240 132.075 ;
        RECT 64.040 122.750 64.300 123.070 ;
        RECT 64.100 119.330 64.240 122.750 ;
        RECT 64.040 119.010 64.300 119.330 ;
        RECT 63.580 118.330 63.840 118.650 ;
        RECT 64.040 118.560 64.300 118.650 ;
        RECT 64.560 118.560 64.700 147.230 ;
        RECT 66.860 146.190 67.000 162.530 ;
        RECT 67.320 148.650 67.460 162.530 ;
        RECT 70.020 162.190 70.280 162.510 ;
        RECT 67.720 161.850 67.980 162.170 ;
        RECT 68.640 161.850 68.900 162.170 ;
        RECT 67.780 151.630 67.920 161.850 ;
        RECT 68.700 160.130 68.840 161.850 ;
        RECT 69.560 161.510 69.820 161.830 ;
        RECT 68.640 159.810 68.900 160.130 ;
        RECT 69.100 159.810 69.360 160.130 ;
        RECT 69.160 159.645 69.300 159.810 ;
        RECT 69.090 159.275 69.370 159.645 ;
        RECT 69.620 159.110 69.760 161.510 ;
        RECT 68.640 158.790 68.900 159.110 ;
        RECT 69.560 158.790 69.820 159.110 ;
        RECT 68.180 158.110 68.440 158.430 ;
        RECT 68.240 157.605 68.380 158.110 ;
        RECT 68.170 157.235 68.450 157.605 ;
        RECT 68.700 157.070 68.840 158.790 ;
        RECT 68.640 156.750 68.900 157.070 ;
        RECT 68.180 156.410 68.440 156.730 ;
        RECT 67.720 151.310 67.980 151.630 ;
        RECT 67.320 148.510 67.920 148.650 ;
        RECT 67.780 147.890 67.920 148.510 ;
        RECT 67.260 147.570 67.520 147.890 ;
        RECT 67.720 147.570 67.980 147.890 ;
        RECT 66.800 145.870 67.060 146.190 ;
        RECT 67.320 145.170 67.460 147.570 ;
        RECT 67.260 144.850 67.520 145.170 ;
        RECT 67.780 144.970 67.920 147.570 ;
        RECT 68.240 147.550 68.380 156.410 ;
        RECT 70.080 153.670 70.220 162.190 ;
        RECT 70.480 160.830 70.740 161.150 ;
        RECT 70.540 156.730 70.680 160.830 ;
        RECT 71.000 157.070 71.140 163.890 ;
        RECT 71.460 162.250 71.600 163.890 ;
        RECT 71.920 162.850 72.060 163.890 ;
        RECT 72.320 163.550 72.580 163.870 ;
        RECT 72.380 162.850 72.520 163.550 ;
        RECT 71.860 162.530 72.120 162.850 ;
        RECT 72.320 162.530 72.580 162.850 ;
        RECT 71.460 162.110 72.060 162.250 ;
        RECT 71.920 161.685 72.060 162.110 ;
        RECT 72.320 161.850 72.580 162.170 ;
        RECT 71.850 161.315 72.130 161.685 ;
        RECT 71.860 160.830 72.120 161.150 ;
        RECT 71.390 159.275 71.670 159.645 ;
        RECT 71.460 157.410 71.600 159.275 ;
        RECT 71.920 158.770 72.060 160.830 ;
        RECT 72.380 158.770 72.520 161.850 ;
        RECT 73.300 161.830 73.440 163.890 ;
        RECT 74.160 163.780 74.420 163.870 ;
        RECT 73.760 163.640 74.420 163.780 ;
        RECT 72.770 161.315 73.050 161.685 ;
        RECT 73.240 161.510 73.500 161.830 ;
        RECT 72.840 159.645 72.980 161.315 ;
        RECT 72.770 159.275 73.050 159.645 ;
        RECT 73.760 158.770 73.900 163.640 ;
        RECT 74.160 163.550 74.420 163.640 ;
        RECT 74.680 162.510 74.820 164.230 ;
        RECT 76.450 164.035 76.730 164.405 ;
        RECT 76.920 164.230 77.180 164.550 ;
        RECT 80.600 164.230 80.860 164.550 ;
        RECT 76.460 163.550 76.720 163.870 ;
        RECT 74.620 162.190 74.880 162.510 ;
        RECT 75.080 161.850 75.340 162.170 ;
        RECT 74.160 161.510 74.420 161.830 ;
        RECT 71.860 158.450 72.120 158.770 ;
        RECT 72.320 158.450 72.580 158.770 ;
        RECT 73.300 158.630 73.900 158.770 ;
        RECT 71.400 157.090 71.660 157.410 ;
        RECT 70.940 156.750 71.200 157.070 ;
        RECT 70.480 156.410 70.740 156.730 ;
        RECT 70.020 153.350 70.280 153.670 ;
        RECT 70.480 150.970 70.740 151.290 ;
        RECT 70.540 150.805 70.680 150.970 ;
        RECT 70.470 150.435 70.750 150.805 ;
        RECT 70.540 150.270 70.680 150.435 ;
        RECT 70.480 149.950 70.740 150.270 ;
        RECT 70.480 148.930 70.740 149.250 ;
        RECT 68.640 147.570 68.900 147.890 ;
        RECT 68.180 147.230 68.440 147.550 ;
        RECT 68.240 146.530 68.380 147.230 ;
        RECT 68.180 146.210 68.440 146.530 ;
        RECT 68.700 145.510 68.840 147.570 ;
        RECT 70.540 146.530 70.680 148.930 ;
        RECT 70.480 146.210 70.740 146.530 ;
        RECT 68.640 145.190 68.900 145.510 ;
        RECT 67.780 144.830 68.380 144.970 ;
        RECT 66.800 143.150 67.060 143.470 ;
        RECT 64.960 142.130 65.220 142.450 ;
        RECT 65.020 141.090 65.160 142.130 ;
        RECT 64.960 140.770 65.220 141.090 ;
        RECT 64.960 140.090 65.220 140.410 ;
        RECT 65.020 138.565 65.160 140.090 ;
        RECT 65.420 139.750 65.680 140.070 ;
        RECT 64.950 138.195 65.230 138.565 ;
        RECT 64.960 137.030 65.220 137.350 ;
        RECT 65.020 126.470 65.160 137.030 ;
        RECT 64.960 126.150 65.220 126.470 ;
        RECT 65.020 124.770 65.160 126.150 ;
        RECT 64.960 124.450 65.220 124.770 ;
        RECT 64.960 122.750 65.220 123.070 ;
        RECT 65.020 120.690 65.160 122.750 ;
        RECT 64.960 120.370 65.220 120.690 ;
        RECT 65.480 119.330 65.620 139.750 ;
        RECT 65.880 136.350 66.140 136.670 ;
        RECT 65.940 131.910 66.080 136.350 ;
        RECT 66.340 134.990 66.600 135.310 ;
        RECT 65.880 131.590 66.140 131.910 ;
        RECT 66.400 129.530 66.540 134.990 ;
        RECT 66.860 134.970 67.000 143.150 ;
        RECT 67.720 139.070 67.980 139.390 ;
        RECT 67.260 137.370 67.520 137.690 ;
        RECT 66.800 134.650 67.060 134.970 ;
        RECT 67.320 134.880 67.460 137.370 ;
        RECT 67.780 137.350 67.920 139.070 ;
        RECT 67.720 137.030 67.980 137.350 ;
        RECT 67.320 134.740 67.920 134.880 ;
        RECT 67.250 134.115 67.530 134.485 ;
        RECT 67.320 133.950 67.460 134.115 ;
        RECT 67.260 133.630 67.520 133.950 ;
        RECT 67.320 131.230 67.460 133.630 ;
        RECT 66.800 130.910 67.060 131.230 ;
        RECT 67.260 130.910 67.520 131.230 ;
        RECT 66.860 129.870 67.000 130.910 ;
        RECT 66.800 129.550 67.060 129.870 ;
        RECT 67.320 129.530 67.460 130.910 ;
        RECT 66.340 129.210 66.600 129.530 ;
        RECT 67.260 129.210 67.520 129.530 ;
        RECT 65.880 121.730 66.140 122.050 ;
        RECT 64.960 119.010 65.220 119.330 ;
        RECT 65.420 119.010 65.680 119.330 ;
        RECT 64.040 118.420 64.700 118.560 ;
        RECT 64.040 118.330 64.300 118.420 ;
        RECT 63.640 115.250 63.780 118.330 ;
        RECT 64.100 118.165 64.240 118.330 ;
        RECT 64.030 117.795 64.310 118.165 ;
        RECT 65.020 117.370 65.160 119.010 ;
        RECT 65.420 118.330 65.680 118.650 ;
        RECT 64.560 117.230 65.160 117.370 ;
        RECT 64.040 115.270 64.300 115.590 ;
        RECT 63.580 114.930 63.840 115.250 ;
        RECT 62.650 114.510 63.320 114.650 ;
        RECT 62.650 114.395 62.930 114.510 ;
        RECT 62.200 112.210 62.460 112.530 ;
        RECT 62.190 110.995 62.470 111.365 ;
        RECT 62.260 110.490 62.400 110.995 ;
        RECT 62.200 110.170 62.460 110.490 ;
        RECT 61.280 109.830 61.940 109.890 ;
        RECT 61.340 109.750 61.940 109.830 ;
        RECT 61.340 108.110 61.480 109.750 ;
        RECT 62.720 109.380 62.860 114.395 ;
        RECT 61.800 109.240 62.860 109.380 ;
        RECT 61.800 108.450 61.940 109.240 ;
        RECT 61.740 108.130 62.000 108.450 ;
        RECT 61.280 107.790 61.540 108.110 ;
        RECT 61.740 107.500 62.000 107.820 ;
        RECT 61.800 106.490 61.940 107.500 ;
        RECT 63.120 107.450 63.380 107.770 ;
        RECT 61.340 106.350 61.940 106.490 ;
        RECT 60.820 104.730 61.080 105.050 ;
        RECT 60.880 102.670 61.020 104.730 ;
        RECT 61.340 104.710 61.480 106.350 ;
        RECT 61.730 105.555 62.010 105.925 ;
        RECT 63.180 105.730 63.320 107.450 ;
        RECT 61.740 105.410 62.000 105.555 ;
        RECT 63.120 105.410 63.380 105.730 ;
        RECT 61.280 104.620 61.540 104.710 ;
        RECT 61.280 104.480 61.940 104.620 ;
        RECT 61.280 104.390 61.540 104.480 ;
        RECT 60.820 102.350 61.080 102.670 ;
        RECT 60.820 101.670 61.080 101.990 ;
        RECT 60.880 97.085 61.020 101.670 ;
        RECT 61.800 100.290 61.940 104.480 ;
        RECT 63.120 104.390 63.380 104.710 ;
        RECT 62.200 103.710 62.460 104.030 ;
        RECT 61.740 99.970 62.000 100.290 ;
        RECT 61.280 99.630 61.540 99.950 ;
        RECT 60.810 96.715 61.090 97.085 ;
        RECT 61.340 96.890 61.480 99.630 ;
        RECT 61.740 96.910 62.000 97.230 ;
        RECT 60.820 96.570 61.080 96.715 ;
        RECT 61.280 96.570 61.540 96.890 ;
        RECT 61.280 93.510 61.540 93.830 ;
        RECT 61.340 91.790 61.480 93.510 ;
        RECT 61.280 91.470 61.540 91.790 ;
        RECT 60.820 91.130 61.080 91.450 ;
        RECT 60.880 89.410 61.020 91.130 ;
        RECT 61.800 89.410 61.940 96.910 ;
        RECT 60.820 89.090 61.080 89.410 ;
        RECT 61.740 89.090 62.000 89.410 ;
        RECT 61.280 85.690 61.540 86.010 ;
        RECT 61.340 84.900 61.480 85.690 ;
        RECT 61.800 85.670 61.940 89.090 ;
        RECT 61.740 85.350 62.000 85.670 ;
        RECT 61.340 84.760 61.940 84.900 ;
        RECT 61.280 80.250 61.540 80.570 ;
        RECT 61.340 78.045 61.480 80.250 ;
        RECT 61.270 77.675 61.550 78.045 ;
        RECT 61.800 77.510 61.940 84.760 ;
        RECT 62.260 82.950 62.400 103.710 ;
        RECT 62.660 95.550 62.920 95.870 ;
        RECT 62.720 93.830 62.860 95.550 ;
        RECT 63.180 94.850 63.320 104.390 ;
        RECT 63.640 96.890 63.780 114.930 ;
        RECT 64.100 105.390 64.240 115.270 ;
        RECT 64.040 105.070 64.300 105.390 ;
        RECT 64.560 104.710 64.700 117.230 ;
        RECT 64.960 115.610 65.220 115.930 ;
        RECT 65.020 113.210 65.160 115.610 ;
        RECT 64.960 112.890 65.220 113.210 ;
        RECT 64.960 110.510 65.220 110.830 ;
        RECT 65.020 110.005 65.160 110.510 ;
        RECT 64.950 109.635 65.230 110.005 ;
        RECT 64.960 105.070 65.220 105.390 ;
        RECT 64.500 104.390 64.760 104.710 ;
        RECT 64.500 103.710 64.760 104.030 ;
        RECT 64.560 102.330 64.700 103.710 ;
        RECT 64.500 102.010 64.760 102.330 ;
        RECT 64.500 99.630 64.760 99.950 ;
        RECT 63.580 96.570 63.840 96.890 ;
        RECT 63.120 94.530 63.380 94.850 ;
        RECT 62.660 93.510 62.920 93.830 ;
        RECT 64.560 88.050 64.700 99.630 ;
        RECT 64.500 87.730 64.760 88.050 ;
        RECT 64.560 86.010 64.700 87.730 ;
        RECT 64.500 85.690 64.760 86.010 ;
        RECT 65.020 85.410 65.160 105.070 ;
        RECT 65.480 99.950 65.620 118.330 ;
        RECT 65.940 118.310 66.080 121.730 ;
        RECT 65.880 117.990 66.140 118.310 ;
        RECT 65.880 114.590 66.140 114.910 ;
        RECT 65.940 105.050 66.080 114.590 ;
        RECT 66.400 109.810 66.540 129.210 ;
        RECT 66.800 125.470 67.060 125.790 ;
        RECT 67.780 125.530 67.920 134.740 ;
        RECT 68.240 132.250 68.380 144.830 ;
        RECT 68.640 144.510 68.900 144.830 ;
        RECT 68.700 141.090 68.840 144.510 ;
        RECT 68.640 140.770 68.900 141.090 ;
        RECT 68.180 131.930 68.440 132.250 ;
        RECT 66.860 124.770 67.000 125.470 ;
        RECT 67.320 125.390 67.920 125.530 ;
        RECT 66.800 124.450 67.060 124.770 ;
        RECT 67.320 116.610 67.460 125.390 ;
        RECT 67.720 124.450 67.980 124.770 ;
        RECT 67.260 116.290 67.520 116.610 ;
        RECT 67.260 115.610 67.520 115.930 ;
        RECT 66.800 114.590 67.060 114.910 ;
        RECT 66.860 110.150 67.000 114.590 ;
        RECT 67.320 111.170 67.460 115.610 ;
        RECT 67.260 110.850 67.520 111.170 ;
        RECT 67.780 110.470 67.920 124.450 ;
        RECT 68.240 121.710 68.380 131.930 ;
        RECT 69.100 131.765 69.360 131.910 ;
        RECT 69.090 131.395 69.370 131.765 ;
        RECT 69.560 131.250 69.820 131.570 ;
        RECT 69.620 128.510 69.760 131.250 ;
        RECT 69.560 128.190 69.820 128.510 ;
        RECT 69.100 126.490 69.360 126.810 ;
        RECT 68.640 123.770 68.900 124.090 ;
        RECT 68.180 121.390 68.440 121.710 ;
        RECT 68.240 121.030 68.380 121.390 ;
        RECT 68.180 120.710 68.440 121.030 ;
        RECT 68.180 116.290 68.440 116.610 ;
        RECT 68.240 111.170 68.380 116.290 ;
        RECT 68.180 110.850 68.440 111.170 ;
        RECT 67.780 110.330 68.380 110.470 ;
        RECT 66.800 109.830 67.060 110.150 ;
        RECT 66.340 109.490 66.600 109.810 ;
        RECT 66.340 106.430 66.600 106.750 ;
        RECT 66.400 105.050 66.540 106.430 ;
        RECT 65.880 104.730 66.140 105.050 ;
        RECT 66.340 104.730 66.600 105.050 ;
        RECT 65.880 102.350 66.140 102.670 ;
        RECT 65.420 99.630 65.680 99.950 ;
        RECT 65.420 98.270 65.680 98.590 ;
        RECT 65.480 96.550 65.620 98.270 ;
        RECT 65.940 97.230 66.080 102.350 ;
        RECT 67.720 98.610 67.980 98.930 ;
        RECT 65.880 96.910 66.140 97.230 ;
        RECT 65.420 96.230 65.680 96.550 ;
        RECT 66.340 92.830 66.600 93.150 ;
        RECT 65.410 91.955 65.690 92.325 ;
        RECT 65.480 86.690 65.620 91.955 ;
        RECT 65.420 86.370 65.680 86.690 ;
        RECT 66.400 86.010 66.540 92.830 ;
        RECT 66.800 90.110 67.060 90.430 ;
        RECT 66.860 88.390 67.000 90.110 ;
        RECT 66.800 88.070 67.060 88.390 ;
        RECT 66.340 85.690 66.600 86.010 ;
        RECT 63.640 85.270 65.160 85.410 ;
        RECT 63.120 84.670 63.380 84.990 ;
        RECT 62.200 82.630 62.460 82.950 ;
        RECT 58.060 76.850 58.320 77.170 ;
        RECT 57.600 76.510 57.860 76.830 ;
        RECT 57.200 75.750 57.800 75.890 ;
        RECT 57.140 75.150 57.400 75.470 ;
        RECT 56.680 72.430 56.940 72.750 ;
        RECT 57.200 72.070 57.340 75.150 ;
        RECT 57.140 71.750 57.400 72.070 ;
        RECT 56.220 69.370 56.480 69.690 ;
        RECT 57.660 67.310 57.800 75.750 ;
        RECT 58.120 75.210 58.260 76.850 ;
        RECT 59.040 75.810 59.180 77.190 ;
        RECT 59.960 77.110 60.560 77.250 ;
        RECT 61.740 77.190 62.000 77.510 ;
        RECT 62.260 77.420 62.400 82.630 ;
        RECT 62.660 81.950 62.920 82.270 ;
        RECT 62.720 80.230 62.860 81.950 ;
        RECT 62.660 79.910 62.920 80.230 ;
        RECT 62.660 77.420 62.920 77.510 ;
        RECT 62.260 77.280 62.920 77.420 ;
        RECT 62.660 77.190 62.920 77.280 ;
        RECT 58.980 75.490 59.240 75.810 ;
        RECT 58.120 75.130 58.720 75.210 ;
        RECT 58.120 75.070 58.780 75.130 ;
        RECT 58.520 74.810 58.780 75.070 ;
        RECT 58.970 74.955 59.250 75.325 ;
        RECT 58.980 74.810 59.240 74.955 ;
        RECT 58.060 74.470 58.320 74.790 ;
        RECT 58.120 72.070 58.260 74.470 ;
        RECT 58.580 72.410 58.720 74.810 ;
        RECT 59.960 72.490 60.100 77.110 ;
        RECT 60.360 76.510 60.620 76.830 ;
        RECT 60.420 74.790 60.560 76.510 ;
        RECT 61.800 75.130 61.940 77.190 ;
        RECT 63.180 76.830 63.320 84.670 ;
        RECT 62.660 76.685 62.920 76.830 ;
        RECT 62.650 76.315 62.930 76.685 ;
        RECT 63.120 76.510 63.380 76.830 ;
        RECT 61.740 74.810 62.000 75.130 ;
        RECT 60.360 74.470 60.620 74.790 ;
        RECT 62.200 74.130 62.460 74.450 ;
        RECT 60.820 73.790 61.080 74.110 ;
        RECT 61.740 73.790 62.000 74.110 ;
        RECT 58.520 72.090 58.780 72.410 ;
        RECT 59.960 72.350 60.560 72.490 ;
        RECT 58.060 71.925 58.320 72.070 ;
        RECT 58.050 71.555 58.330 71.925 ;
        RECT 59.440 71.810 59.700 72.070 ;
        RECT 59.440 71.750 60.100 71.810 ;
        RECT 59.500 71.670 60.100 71.750 ;
        RECT 57.600 66.990 57.860 67.310 ;
        RECT 55.300 66.650 55.560 66.970 ;
        RECT 59.960 66.630 60.100 71.670 ;
        RECT 60.420 69.690 60.560 72.350 ;
        RECT 60.880 71.730 61.020 73.790 ;
        RECT 60.820 71.410 61.080 71.730 ;
        RECT 60.360 69.370 60.620 69.690 ;
        RECT 59.900 66.310 60.160 66.630 ;
        RECT 58.980 65.630 59.240 65.950 ;
        RECT 57.600 62.910 57.860 63.230 ;
        RECT 57.140 60.870 57.400 61.190 ;
        RECT 57.200 58.810 57.340 60.870 ;
        RECT 57.660 59.150 57.800 62.910 ;
        RECT 59.040 61.530 59.180 65.630 ;
        RECT 59.960 61.530 60.100 66.310 ;
        RECT 60.420 64.590 60.560 69.370 ;
        RECT 60.820 68.350 61.080 68.670 ;
        RECT 61.280 68.350 61.540 68.670 ;
        RECT 60.880 64.930 61.020 68.350 ;
        RECT 61.340 66.630 61.480 68.350 ;
        RECT 61.280 66.310 61.540 66.630 ;
        RECT 60.820 64.610 61.080 64.930 ;
        RECT 60.360 64.270 60.620 64.590 ;
        RECT 60.420 63.910 60.560 64.270 ;
        RECT 61.800 64.250 61.940 73.790 ;
        RECT 62.260 69.350 62.400 74.130 ;
        RECT 62.200 69.030 62.460 69.350 ;
        RECT 61.740 63.930 62.000 64.250 ;
        RECT 63.180 63.910 63.320 76.510 ;
        RECT 60.360 63.590 60.620 63.910 ;
        RECT 63.120 63.590 63.380 63.910 ;
        RECT 61.740 63.250 62.000 63.570 ;
        RECT 61.280 62.910 61.540 63.230 ;
        RECT 58.980 61.210 59.240 61.530 ;
        RECT 59.900 61.210 60.160 61.530 ;
        RECT 59.440 60.870 59.700 61.190 ;
        RECT 58.520 60.190 58.780 60.510 ;
        RECT 57.600 58.830 57.860 59.150 ;
        RECT 57.140 58.490 57.400 58.810 ;
        RECT 58.580 55.750 58.720 60.190 ;
        RECT 59.500 59.490 59.640 60.870 ;
        RECT 61.340 60.850 61.480 62.910 ;
        RECT 61.280 60.530 61.540 60.850 ;
        RECT 61.270 59.995 61.550 60.365 ;
        RECT 59.440 59.170 59.700 59.490 ;
        RECT 60.360 58.490 60.620 58.810 ;
        RECT 58.520 55.430 58.780 55.750 ;
        RECT 54.830 54.555 55.110 54.925 ;
        RECT 54.840 52.030 55.100 52.350 ;
        RECT 53.920 46.590 54.180 46.910 ;
        RECT 53.980 43.170 54.120 46.590 ;
        RECT 53.920 42.850 54.180 43.170 ;
        RECT 54.900 42.150 55.040 52.030 ;
        RECT 57.140 49.650 57.400 49.970 ;
        RECT 57.600 49.650 57.860 49.970 ;
        RECT 57.200 45.890 57.340 49.650 ;
        RECT 57.660 47.930 57.800 49.650 ;
        RECT 57.600 47.610 57.860 47.930 ;
        RECT 57.140 45.570 57.400 45.890 ;
        RECT 58.580 44.870 58.720 55.430 ;
        RECT 60.420 55.410 60.560 58.490 ;
        RECT 60.360 55.090 60.620 55.410 ;
        RECT 60.420 53.370 60.560 55.090 ;
        RECT 60.360 53.050 60.620 53.370 ;
        RECT 60.420 49.970 60.560 53.050 ;
        RECT 60.360 49.650 60.620 49.970 ;
        RECT 60.350 47.755 60.630 48.125 ;
        RECT 59.900 44.890 60.160 45.210 ;
        RECT 58.520 44.550 58.780 44.870 ;
        RECT 55.760 43.870 56.020 44.190 ;
        RECT 59.440 43.870 59.700 44.190 ;
        RECT 54.840 41.830 55.100 42.150 ;
        RECT 53.460 41.150 53.720 41.470 ;
        RECT 52.080 38.860 52.740 39.000 ;
        RECT 52.080 38.770 52.340 38.860 ;
        RECT 53.000 38.770 53.260 39.090 ;
        RECT 49.780 38.430 50.040 38.750 ;
        RECT 49.320 37.070 49.580 37.390 ;
        RECT 48.400 31.290 48.660 31.610 ;
        RECT 48.860 31.290 49.120 31.610 ;
        RECT 47.480 26.190 47.740 26.510 ;
        RECT 47.480 25.170 47.740 25.490 ;
        RECT 47.540 23.110 47.680 25.170 ;
        RECT 49.380 23.110 49.520 37.070 ;
        RECT 49.840 31.610 49.980 38.430 ;
        RECT 52.140 36.030 52.280 38.770 ;
        RECT 52.080 35.710 52.340 36.030 ;
        RECT 50.240 32.990 50.500 33.310 ;
        RECT 49.780 31.290 50.040 31.610 ;
        RECT 50.300 31.270 50.440 32.990 ;
        RECT 50.240 30.950 50.500 31.270 ;
        RECT 49.780 30.270 50.040 30.590 ;
        RECT 49.840 28.550 49.980 30.270 ;
        RECT 53.060 29.570 53.200 38.770 ;
        RECT 53.520 33.990 53.660 41.150 ;
        RECT 53.920 35.710 54.180 36.030 ;
        RECT 53.980 33.990 54.120 35.710 ;
        RECT 53.460 33.670 53.720 33.990 ;
        RECT 53.920 33.670 54.180 33.990 ;
        RECT 54.900 32.290 55.040 41.830 ;
        RECT 55.300 40.130 55.560 40.450 ;
        RECT 55.360 34.330 55.500 40.130 ;
        RECT 55.820 37.050 55.960 43.870 ;
        RECT 59.500 42.490 59.640 43.870 ;
        RECT 59.440 42.170 59.700 42.490 ;
        RECT 56.220 41.150 56.480 41.470 ;
        RECT 58.980 41.150 59.240 41.470 ;
        RECT 56.280 39.430 56.420 41.150 ;
        RECT 58.520 40.130 58.780 40.450 ;
        RECT 56.220 39.110 56.480 39.430 ;
        RECT 56.680 37.410 56.940 37.730 ;
        RECT 55.760 36.730 56.020 37.050 ;
        RECT 55.300 34.010 55.560 34.330 ;
        RECT 55.820 33.650 55.960 36.730 ;
        RECT 56.740 35.010 56.880 37.410 ;
        RECT 58.060 36.730 58.320 37.050 ;
        RECT 58.120 35.010 58.260 36.730 ;
        RECT 56.680 34.920 56.940 35.010 ;
        RECT 56.280 34.780 56.940 34.920 ;
        RECT 55.760 33.330 56.020 33.650 ;
        RECT 56.280 32.290 56.420 34.780 ;
        RECT 56.680 34.690 56.940 34.780 ;
        RECT 58.060 34.690 58.320 35.010 ;
        RECT 54.840 31.970 55.100 32.290 ;
        RECT 56.220 31.970 56.480 32.290 ;
        RECT 55.760 31.290 56.020 31.610 ;
        RECT 55.300 30.950 55.560 31.270 ;
        RECT 54.380 30.270 54.640 30.590 ;
        RECT 53.000 29.250 53.260 29.570 ;
        RECT 54.440 28.550 54.580 30.270 ;
        RECT 49.780 28.230 50.040 28.550 ;
        RECT 53.920 28.230 54.180 28.550 ;
        RECT 54.380 28.230 54.640 28.550 ;
        RECT 53.980 26.850 54.120 28.230 ;
        RECT 53.920 26.530 54.180 26.850 ;
        RECT 54.440 26.170 54.580 28.230 ;
        RECT 54.840 27.550 55.100 27.870 ;
        RECT 54.380 25.850 54.640 26.170 ;
        RECT 46.560 22.790 46.820 23.110 ;
        RECT 47.020 22.790 47.280 23.110 ;
        RECT 47.480 22.790 47.740 23.110 ;
        RECT 49.320 22.790 49.580 23.110 ;
        RECT 46.160 22.030 46.760 22.170 ;
        RECT 46.620 21.070 46.760 22.030 ;
        RECT 46.560 20.750 46.820 21.070 ;
        RECT 45.640 20.410 45.900 20.730 ;
        RECT 44.720 19.390 44.980 19.710 ;
        RECT 44.780 15.630 44.920 19.390 ;
        RECT 45.700 17.330 45.840 20.410 ;
        RECT 46.100 17.350 46.360 17.670 ;
        RECT 45.640 17.010 45.900 17.330 ;
        RECT 46.160 15.970 46.300 17.350 ;
        RECT 46.100 15.650 46.360 15.970 ;
        RECT 44.720 15.310 44.980 15.630 ;
        RECT 44.260 12.590 44.520 12.910 ;
        RECT 46.160 12.230 46.300 15.650 ;
        RECT 46.620 12.570 46.760 20.750 ;
        RECT 47.080 20.390 47.220 22.790 ;
        RECT 47.940 22.110 48.200 22.430 ;
        RECT 48.000 20.730 48.140 22.110 ;
        RECT 48.860 20.750 49.120 21.070 ;
        RECT 47.940 20.410 48.200 20.730 ;
        RECT 47.020 20.070 47.280 20.390 ;
        RECT 48.920 18.690 49.060 20.750 ;
        RECT 49.380 20.390 49.520 22.790 ;
        RECT 53.920 22.110 54.180 22.430 ;
        RECT 52.080 20.410 52.340 20.730 ;
        RECT 49.320 20.070 49.580 20.390 ;
        RECT 48.860 18.370 49.120 18.690 ;
        RECT 49.380 18.010 49.520 20.070 ;
        RECT 49.320 17.690 49.580 18.010 ;
        RECT 52.140 15.970 52.280 20.410 ;
        RECT 53.980 18.090 54.120 22.110 ;
        RECT 54.440 19.710 54.580 25.850 ;
        RECT 54.900 21.410 55.040 27.550 ;
        RECT 55.360 26.510 55.500 30.950 ;
        RECT 55.300 26.190 55.560 26.510 ;
        RECT 55.820 25.150 55.960 31.290 ;
        RECT 56.280 31.270 56.420 31.970 ;
        RECT 56.220 30.950 56.480 31.270 ;
        RECT 58.580 30.590 58.720 40.130 ;
        RECT 59.040 39.430 59.180 41.150 ;
        RECT 58.980 39.110 59.240 39.430 ;
        RECT 59.500 33.310 59.640 42.170 ;
        RECT 59.440 32.990 59.700 33.310 ;
        RECT 58.520 30.270 58.780 30.590 ;
        RECT 56.210 28.715 56.490 29.085 ;
        RECT 55.760 24.830 56.020 25.150 ;
        RECT 55.820 24.130 55.960 24.830 ;
        RECT 55.760 23.810 56.020 24.130 ;
        RECT 54.840 21.090 55.100 21.410 ;
        RECT 54.380 19.390 54.640 19.710 ;
        RECT 54.440 18.690 54.580 19.390 ;
        RECT 54.380 18.370 54.640 18.690 ;
        RECT 53.980 17.950 54.580 18.090 ;
        RECT 52.080 15.650 52.340 15.970 ;
        RECT 54.440 14.950 54.580 17.950 ;
        RECT 54.900 14.950 55.040 21.090 ;
        RECT 55.820 17.330 55.960 23.810 ;
        RECT 56.280 20.050 56.420 28.715 ;
        RECT 58.580 28.550 58.720 30.270 ;
        RECT 59.500 28.970 59.640 32.990 ;
        RECT 59.960 32.290 60.100 44.890 ;
        RECT 59.900 31.970 60.160 32.290 ;
        RECT 60.420 29.570 60.560 47.755 ;
        RECT 61.340 46.910 61.480 59.995 ;
        RECT 61.800 59.150 61.940 63.250 ;
        RECT 61.740 58.830 62.000 59.150 ;
        RECT 63.180 56.850 63.320 63.590 ;
        RECT 63.640 61.045 63.780 85.270 ;
        RECT 64.960 83.650 65.220 83.970 ;
        RECT 64.500 81.950 64.760 82.270 ;
        RECT 64.560 77.170 64.700 81.950 ;
        RECT 64.500 76.850 64.760 77.170 ;
        RECT 64.560 71.730 64.700 76.850 ;
        RECT 65.020 76.830 65.160 83.650 ;
        RECT 65.420 82.630 65.680 82.950 ;
        RECT 66.340 82.630 66.600 82.950 ;
        RECT 67.260 82.630 67.520 82.950 ;
        RECT 65.480 79.970 65.620 82.630 ;
        RECT 66.400 81.445 66.540 82.630 ;
        RECT 66.800 81.950 67.060 82.270 ;
        RECT 66.330 81.075 66.610 81.445 ;
        RECT 66.340 80.250 66.600 80.570 ;
        RECT 65.480 79.830 66.080 79.970 ;
        RECT 65.940 79.550 66.080 79.830 ;
        RECT 65.880 79.230 66.140 79.550 ;
        RECT 66.400 77.170 66.540 80.250 ;
        RECT 66.860 77.170 67.000 81.950 ;
        RECT 67.320 80.910 67.460 82.630 ;
        RECT 67.260 80.590 67.520 80.910 ;
        RECT 67.260 79.910 67.520 80.230 ;
        RECT 66.340 76.850 66.600 77.170 ;
        RECT 66.800 76.850 67.060 77.170 ;
        RECT 64.960 76.510 65.220 76.830 ;
        RECT 64.500 71.410 64.760 71.730 ;
        RECT 64.040 71.070 64.300 71.390 ;
        RECT 64.100 70.370 64.240 71.070 ;
        RECT 64.040 70.050 64.300 70.370 ;
        RECT 65.020 67.650 65.160 76.510 ;
        RECT 66.340 74.470 66.600 74.790 ;
        RECT 66.400 71.390 66.540 74.470 ;
        RECT 66.860 72.410 67.000 76.850 ;
        RECT 66.800 72.090 67.060 72.410 ;
        RECT 66.340 71.070 66.600 71.390 ;
        RECT 66.800 71.300 67.060 71.390 ;
        RECT 67.320 71.300 67.460 79.910 ;
        RECT 66.800 71.160 67.460 71.300 ;
        RECT 66.800 71.070 67.060 71.160 ;
        RECT 66.400 70.030 66.540 71.070 ;
        RECT 66.340 69.710 66.600 70.030 ;
        RECT 64.960 67.330 65.220 67.650 ;
        RECT 63.570 60.675 63.850 61.045 ;
        RECT 63.180 56.710 64.240 56.850 ;
        RECT 63.580 54.750 63.840 55.070 ;
        RECT 62.200 49.310 62.460 49.630 ;
        RECT 62.260 48.270 62.400 49.310 ;
        RECT 62.200 47.950 62.460 48.270 ;
        RECT 61.280 46.590 61.540 46.910 ;
        RECT 61.280 45.230 61.540 45.550 ;
        RECT 60.820 44.890 61.080 45.210 ;
        RECT 60.880 40.450 61.020 44.890 ;
        RECT 60.820 40.130 61.080 40.450 ;
        RECT 60.820 38.770 61.080 39.090 ;
        RECT 60.880 34.330 61.020 38.770 ;
        RECT 60.820 34.010 61.080 34.330 ;
        RECT 60.360 29.250 60.620 29.570 ;
        RECT 59.500 28.830 60.560 28.970 ;
        RECT 58.520 28.230 58.780 28.550 ;
        RECT 57.600 27.550 57.860 27.870 ;
        RECT 57.140 22.790 57.400 23.110 ;
        RECT 56.220 19.730 56.480 20.050 ;
        RECT 55.760 17.010 56.020 17.330 ;
        RECT 56.280 15.970 56.420 19.730 ;
        RECT 57.200 18.010 57.340 22.790 ;
        RECT 57.140 17.690 57.400 18.010 ;
        RECT 57.660 17.330 57.800 27.550 ;
        RECT 58.580 26.170 58.720 28.230 ;
        RECT 59.890 26.675 60.170 27.045 ;
        RECT 59.900 26.530 60.160 26.675 ;
        RECT 58.520 25.850 58.780 26.170 ;
        RECT 60.420 25.830 60.560 28.830 ;
        RECT 61.340 28.550 61.480 45.230 ;
        RECT 62.260 44.530 62.400 47.950 ;
        RECT 63.120 47.610 63.380 47.930 ;
        RECT 62.200 44.210 62.460 44.530 ;
        RECT 62.660 44.210 62.920 44.530 ;
        RECT 61.740 43.870 62.000 44.190 ;
        RECT 61.800 42.150 61.940 43.870 ;
        RECT 61.740 41.830 62.000 42.150 ;
        RECT 62.720 39.770 62.860 44.210 ;
        RECT 63.180 43.170 63.320 47.610 ;
        RECT 63.120 42.850 63.380 43.170 ;
        RECT 63.640 42.570 63.780 54.750 ;
        RECT 64.100 42.830 64.240 56.710 ;
        RECT 66.340 56.680 66.600 56.770 ;
        RECT 66.860 56.680 67.000 71.070 ;
        RECT 67.780 63.570 67.920 98.610 ;
        RECT 68.240 88.390 68.380 110.330 ;
        RECT 68.700 105.730 68.840 123.770 ;
        RECT 69.160 121.370 69.300 126.490 ;
        RECT 70.540 126.470 70.680 146.210 ;
        RECT 71.000 128.510 71.140 156.750 ;
        RECT 72.780 154.030 73.040 154.350 ;
        RECT 71.860 153.350 72.120 153.670 ;
        RECT 71.400 153.010 71.660 153.330 ;
        RECT 71.460 151.290 71.600 153.010 ;
        RECT 71.400 150.970 71.660 151.290 ;
        RECT 71.460 147.970 71.600 150.970 ;
        RECT 71.920 148.570 72.060 153.350 ;
        RECT 72.840 151.290 72.980 154.030 ;
        RECT 73.300 153.670 73.440 158.630 ;
        RECT 74.220 154.090 74.360 161.510 ;
        RECT 74.610 161.315 74.890 161.685 ;
        RECT 74.680 161.150 74.820 161.315 ;
        RECT 74.620 160.830 74.880 161.150 ;
        RECT 74.620 158.790 74.880 159.110 ;
        RECT 73.760 153.950 74.360 154.090 ;
        RECT 73.240 153.350 73.500 153.670 ;
        RECT 72.780 150.970 73.040 151.290 ;
        RECT 72.320 150.630 72.580 150.950 ;
        RECT 71.860 148.250 72.120 148.570 ;
        RECT 71.460 147.830 72.060 147.970 ;
        RECT 71.400 147.230 71.660 147.550 ;
        RECT 71.460 142.790 71.600 147.230 ;
        RECT 71.920 142.790 72.060 147.830 ;
        RECT 72.380 145.850 72.520 150.630 ;
        RECT 72.840 147.550 72.980 150.970 ;
        RECT 72.780 147.230 73.040 147.550 ;
        RECT 72.320 145.530 72.580 145.850 ;
        RECT 72.380 143.810 72.520 145.530 ;
        RECT 72.840 145.250 72.980 147.230 ;
        RECT 73.240 146.210 73.500 146.530 ;
        RECT 73.300 145.850 73.440 146.210 ;
        RECT 73.240 145.530 73.500 145.850 ;
        RECT 72.840 145.110 73.440 145.250 ;
        RECT 72.780 144.510 73.040 144.830 ;
        RECT 72.320 143.490 72.580 143.810 ;
        RECT 72.840 143.470 72.980 144.510 ;
        RECT 72.780 143.150 73.040 143.470 ;
        RECT 73.300 143.130 73.440 145.110 ;
        RECT 73.240 142.810 73.500 143.130 ;
        RECT 71.400 142.470 71.660 142.790 ;
        RECT 71.860 142.470 72.120 142.790 ;
        RECT 73.760 142.530 73.900 153.950 ;
        RECT 74.680 153.670 74.820 158.790 ;
        RECT 74.620 153.350 74.880 153.670 ;
        RECT 74.160 153.010 74.420 153.330 ;
        RECT 74.220 149.250 74.360 153.010 ;
        RECT 74.680 151.290 74.820 153.350 ;
        RECT 75.140 151.290 75.280 161.850 ;
        RECT 75.540 161.170 75.800 161.490 ;
        RECT 75.600 159.110 75.740 161.170 ;
        RECT 75.540 158.790 75.800 159.110 ;
        RECT 76.000 158.790 76.260 159.110 ;
        RECT 74.620 150.970 74.880 151.290 ;
        RECT 75.080 150.970 75.340 151.290 ;
        RECT 74.160 148.930 74.420 149.250 ;
        RECT 74.160 147.910 74.420 148.230 ;
        RECT 74.220 145.170 74.360 147.910 ;
        RECT 74.160 144.850 74.420 145.170 ;
        RECT 74.680 143.130 74.820 150.970 ;
        RECT 75.080 145.530 75.340 145.850 ;
        RECT 75.140 145.365 75.280 145.530 ;
        RECT 75.070 144.995 75.350 145.365 ;
        RECT 74.160 142.810 74.420 143.130 ;
        RECT 74.620 142.810 74.880 143.130 ;
        RECT 71.400 138.050 71.660 138.370 ;
        RECT 70.940 128.190 71.200 128.510 ;
        RECT 69.550 125.955 69.830 126.325 ;
        RECT 70.480 126.150 70.740 126.470 ;
        RECT 69.620 123.410 69.760 125.955 ;
        RECT 70.020 125.810 70.280 126.130 ;
        RECT 69.560 123.090 69.820 123.410 ;
        RECT 70.080 122.130 70.220 125.810 ;
        RECT 70.540 123.410 70.680 126.150 ;
        RECT 71.460 124.090 71.600 138.050 ;
        RECT 71.920 132.500 72.060 142.470 ;
        RECT 73.300 142.390 73.900 142.530 ;
        RECT 72.780 139.070 73.040 139.390 ;
        RECT 72.840 135.650 72.980 139.070 ;
        RECT 72.780 135.330 73.040 135.650 ;
        RECT 72.780 132.500 73.040 132.590 ;
        RECT 71.920 132.360 73.040 132.500 ;
        RECT 72.780 132.270 73.040 132.360 ;
        RECT 72.320 128.870 72.580 129.190 ;
        RECT 71.860 128.530 72.120 128.850 ;
        RECT 71.920 124.090 72.060 128.530 ;
        RECT 72.380 126.810 72.520 128.870 ;
        RECT 72.320 126.490 72.580 126.810 ;
        RECT 72.840 126.210 72.980 132.270 ;
        RECT 72.380 126.070 72.980 126.210 ;
        RECT 71.400 123.770 71.660 124.090 ;
        RECT 71.860 123.770 72.120 124.090 ;
        RECT 70.480 123.090 70.740 123.410 ;
        RECT 70.080 121.990 71.140 122.130 ;
        RECT 71.460 122.050 71.600 123.770 ;
        RECT 71.860 123.090 72.120 123.410 ;
        RECT 70.020 121.390 70.280 121.710 ;
        RECT 69.100 121.050 69.360 121.370 ;
        RECT 69.560 121.050 69.820 121.370 ;
        RECT 69.160 119.330 69.300 121.050 ;
        RECT 69.100 119.010 69.360 119.330 ;
        RECT 69.090 116.435 69.370 116.805 ;
        RECT 69.160 112.530 69.300 116.435 ;
        RECT 69.620 116.270 69.760 121.050 ;
        RECT 69.560 115.950 69.820 116.270 ;
        RECT 69.560 114.930 69.820 115.250 ;
        RECT 69.620 112.870 69.760 114.930 ;
        RECT 69.560 112.550 69.820 112.870 ;
        RECT 69.100 112.210 69.360 112.530 ;
        RECT 69.100 106.430 69.360 106.750 ;
        RECT 68.640 105.410 68.900 105.730 ;
        RECT 69.160 104.710 69.300 106.430 ;
        RECT 69.100 104.390 69.360 104.710 ;
        RECT 70.080 104.370 70.220 121.390 ;
        RECT 71.000 120.350 71.140 121.990 ;
        RECT 71.400 121.730 71.660 122.050 ;
        RECT 70.480 120.030 70.740 120.350 ;
        RECT 70.940 120.030 71.200 120.350 ;
        RECT 70.540 118.990 70.680 120.030 ;
        RECT 71.000 118.990 71.140 120.030 ;
        RECT 70.480 118.670 70.740 118.990 ;
        RECT 70.940 118.670 71.200 118.990 ;
        RECT 71.400 117.650 71.660 117.970 ;
        RECT 71.460 115.590 71.600 117.650 ;
        RECT 70.480 115.270 70.740 115.590 ;
        RECT 71.400 115.270 71.660 115.590 ;
        RECT 70.540 114.910 70.680 115.270 ;
        RECT 70.480 114.590 70.740 114.910 ;
        RECT 70.480 111.870 70.740 112.190 ;
        RECT 70.540 108.450 70.680 111.870 ;
        RECT 71.920 111.170 72.060 123.090 ;
        RECT 72.380 121.030 72.520 126.070 ;
        RECT 72.780 123.770 73.040 124.090 ;
        RECT 73.300 124.000 73.440 142.390 ;
        RECT 73.700 141.790 73.960 142.110 ;
        RECT 73.760 137.010 73.900 141.790 ;
        RECT 74.220 138.370 74.360 142.810 ;
        RECT 74.160 138.050 74.420 138.370 ;
        RECT 74.680 137.350 74.820 142.810 ;
        RECT 75.600 140.750 75.740 158.790 ;
        RECT 76.060 156.730 76.200 158.790 ;
        RECT 76.000 156.410 76.260 156.730 ;
        RECT 76.060 147.290 76.200 156.410 ;
        RECT 76.520 148.230 76.660 163.550 ;
        RECT 76.980 160.130 77.120 164.230 ;
        RECT 78.300 163.890 78.560 164.210 ;
        RECT 78.760 163.890 79.020 164.210 ;
        RECT 79.220 163.890 79.480 164.210 ;
        RECT 77.380 163.550 77.640 163.870 ;
        RECT 76.920 159.810 77.180 160.130 ;
        RECT 76.920 156.070 77.180 156.390 ;
        RECT 76.980 152.845 77.120 156.070 ;
        RECT 76.910 152.475 77.190 152.845 ;
        RECT 76.910 149.755 77.190 150.125 ;
        RECT 76.460 147.910 76.720 148.230 ;
        RECT 76.060 147.150 76.660 147.290 ;
        RECT 76.520 145.850 76.660 147.150 ;
        RECT 76.460 145.530 76.720 145.850 ;
        RECT 76.000 144.850 76.260 145.170 ;
        RECT 75.540 140.660 75.800 140.750 ;
        RECT 75.140 140.520 75.800 140.660 ;
        RECT 74.620 137.030 74.880 137.350 ;
        RECT 73.700 136.690 73.960 137.010 ;
        RECT 74.680 134.970 74.820 137.030 ;
        RECT 73.700 134.650 73.960 134.970 ;
        RECT 74.620 134.650 74.880 134.970 ;
        RECT 73.760 132.930 73.900 134.650 ;
        RECT 73.700 132.610 73.960 132.930 ;
        RECT 74.160 130.910 74.420 131.230 ;
        RECT 74.220 130.210 74.360 130.910 ;
        RECT 74.160 129.890 74.420 130.210 ;
        RECT 74.680 129.870 74.820 134.650 ;
        RECT 74.620 129.550 74.880 129.870 ;
        RECT 74.160 128.870 74.420 129.190 ;
        RECT 74.220 127.490 74.360 128.870 ;
        RECT 74.160 127.170 74.420 127.490 ;
        RECT 74.680 126.810 74.820 129.550 ;
        RECT 74.620 126.490 74.880 126.810 ;
        RECT 74.680 124.090 74.820 126.490 ;
        RECT 75.140 124.430 75.280 140.520 ;
        RECT 75.540 140.430 75.800 140.520 ;
        RECT 75.540 136.350 75.800 136.670 ;
        RECT 75.600 130.210 75.740 136.350 ;
        RECT 75.540 129.890 75.800 130.210 ;
        RECT 76.060 129.530 76.200 144.850 ;
        RECT 76.520 143.810 76.660 145.530 ;
        RECT 76.980 145.170 77.120 149.755 ;
        RECT 77.440 146.190 77.580 163.550 ;
        RECT 78.360 162.510 78.500 163.890 ;
        RECT 78.300 162.190 78.560 162.510 ;
        RECT 78.820 162.250 78.960 163.890 ;
        RECT 79.280 163.725 79.420 163.890 ;
        RECT 79.210 163.355 79.490 163.725 ;
        RECT 78.820 162.170 79.880 162.250 ;
        RECT 78.820 162.110 79.940 162.170 ;
        RECT 79.680 161.850 79.940 162.110 ;
        RECT 78.300 161.510 78.560 161.830 ;
        RECT 79.220 161.510 79.480 161.830 ;
        RECT 77.840 160.830 78.100 161.150 ;
        RECT 78.360 161.005 78.500 161.510 ;
        RECT 77.900 160.325 78.040 160.830 ;
        RECT 78.290 160.635 78.570 161.005 ;
        RECT 77.830 159.955 78.110 160.325 ;
        RECT 79.280 156.050 79.420 161.510 ;
        RECT 79.740 159.450 79.880 161.850 ;
        RECT 80.660 161.005 80.800 164.230 ;
        RECT 81.060 163.890 81.320 164.210 ;
        RECT 80.590 160.635 80.870 161.005 ;
        RECT 80.140 159.470 80.400 159.790 ;
        RECT 79.680 159.130 79.940 159.450 ;
        RECT 79.220 155.730 79.480 156.050 ;
        RECT 78.760 155.390 79.020 155.710 ;
        RECT 77.840 150.970 78.100 151.290 ;
        RECT 77.900 149.250 78.040 150.970 ;
        RECT 77.840 148.930 78.100 149.250 ;
        RECT 78.300 148.250 78.560 148.570 ;
        RECT 77.380 145.870 77.640 146.190 ;
        RECT 77.380 145.190 77.640 145.510 ;
        RECT 76.920 144.850 77.180 145.170 ;
        RECT 76.460 143.490 76.720 143.810 ;
        RECT 76.460 142.130 76.720 142.450 ;
        RECT 76.520 141.090 76.660 142.130 ;
        RECT 76.920 141.790 77.180 142.110 ;
        RECT 76.460 140.770 76.720 141.090 ;
        RECT 76.980 139.925 77.120 141.790 ;
        RECT 76.910 139.555 77.190 139.925 ;
        RECT 76.920 136.690 77.180 137.010 ;
        RECT 76.460 136.350 76.720 136.670 ;
        RECT 76.520 133.950 76.660 136.350 ;
        RECT 76.460 133.630 76.720 133.950 ;
        RECT 76.000 129.210 76.260 129.530 ;
        RECT 76.000 125.810 76.260 126.130 ;
        RECT 75.080 124.110 75.340 124.430 ;
        RECT 73.300 123.860 74.360 124.000 ;
        RECT 72.840 121.710 72.980 123.770 ;
        RECT 73.700 123.090 73.960 123.410 ;
        RECT 73.240 122.750 73.500 123.070 ;
        RECT 73.300 122.245 73.440 122.750 ;
        RECT 73.230 121.875 73.510 122.245 ;
        RECT 72.780 121.390 73.040 121.710 ;
        RECT 72.320 120.710 72.580 121.030 ;
        RECT 72.380 119.410 72.520 120.710 ;
        RECT 72.380 119.270 73.440 119.410 ;
        RECT 72.310 115.755 72.590 116.125 ;
        RECT 72.380 115.590 72.520 115.755 ;
        RECT 72.320 115.270 72.580 115.590 ;
        RECT 71.860 110.850 72.120 111.170 ;
        RECT 70.940 110.170 71.200 110.490 ;
        RECT 71.400 110.170 71.660 110.490 ;
        RECT 72.380 110.470 72.520 115.270 ;
        RECT 72.780 112.890 73.040 113.210 ;
        RECT 71.920 110.330 72.520 110.470 ;
        RECT 70.480 108.130 70.740 108.450 ;
        RECT 71.000 105.130 71.140 110.170 ;
        RECT 71.460 106.750 71.600 110.170 ;
        RECT 71.920 108.110 72.060 110.330 ;
        RECT 72.320 109.490 72.580 109.810 ;
        RECT 72.380 108.450 72.520 109.490 ;
        RECT 72.840 108.450 72.980 112.890 ;
        RECT 72.320 108.130 72.580 108.450 ;
        RECT 72.780 108.130 73.040 108.450 ;
        RECT 71.860 107.790 72.120 108.110 ;
        RECT 71.400 106.430 71.660 106.750 ;
        RECT 71.920 105.390 72.060 107.790 ;
        RECT 70.540 104.990 71.140 105.130 ;
        RECT 71.860 105.070 72.120 105.390 ;
        RECT 70.020 104.050 70.280 104.370 ;
        RECT 68.640 96.910 68.900 97.230 ;
        RECT 68.180 88.070 68.440 88.390 ;
        RECT 68.240 63.910 68.380 88.070 ;
        RECT 68.700 82.610 68.840 96.910 ;
        RECT 69.560 96.230 69.820 96.550 ;
        RECT 69.620 94.510 69.760 96.230 ;
        RECT 69.560 94.190 69.820 94.510 ;
        RECT 69.620 93.830 69.760 94.190 ;
        RECT 69.560 93.510 69.820 93.830 ;
        RECT 69.560 91.810 69.820 92.130 ;
        RECT 69.620 88.390 69.760 91.810 ;
        RECT 69.090 87.875 69.370 88.245 ;
        RECT 69.560 88.070 69.820 88.390 ;
        RECT 69.160 86.690 69.300 87.875 ;
        RECT 69.100 86.370 69.360 86.690 ;
        RECT 70.080 86.090 70.220 104.050 ;
        RECT 70.540 94.850 70.680 104.990 ;
        RECT 72.380 104.710 72.520 108.130 ;
        RECT 73.300 107.850 73.440 119.270 ;
        RECT 73.760 110.490 73.900 123.090 ;
        RECT 74.220 114.910 74.360 123.860 ;
        RECT 74.620 123.770 74.880 124.090 ;
        RECT 75.140 123.490 75.280 124.110 ;
        RECT 74.680 123.410 75.280 123.490 ;
        RECT 74.620 123.350 75.280 123.410 ;
        RECT 74.620 123.090 74.880 123.350 ;
        RECT 76.060 123.070 76.200 125.810 ;
        RECT 76.000 122.750 76.260 123.070 ;
        RECT 76.460 122.750 76.720 123.070 ;
        RECT 74.620 121.730 74.880 122.050 ;
        RECT 75.530 121.875 75.810 122.245 ;
        RECT 74.680 121.030 74.820 121.730 ;
        RECT 75.600 121.710 75.740 121.875 ;
        RECT 75.540 121.390 75.800 121.710 ;
        RECT 74.620 120.710 74.880 121.030 ;
        RECT 75.080 120.710 75.340 121.030 ;
        RECT 75.140 119.330 75.280 120.710 ;
        RECT 75.080 119.010 75.340 119.330 ;
        RECT 75.990 119.155 76.270 119.525 ;
        RECT 75.540 118.330 75.800 118.650 ;
        RECT 74.160 114.590 74.420 114.910 ;
        RECT 73.700 110.170 73.960 110.490 ;
        RECT 74.220 109.210 74.360 114.590 ;
        RECT 75.600 113.890 75.740 118.330 ;
        RECT 76.060 118.310 76.200 119.155 ;
        RECT 76.000 117.990 76.260 118.310 ;
        RECT 76.520 117.630 76.660 122.750 ;
        RECT 76.980 120.690 77.120 136.690 ;
        RECT 77.440 136.670 77.580 145.190 ;
        RECT 77.840 142.470 78.100 142.790 ;
        RECT 77.900 140.410 78.040 142.470 ;
        RECT 77.840 140.090 78.100 140.410 ;
        RECT 78.360 137.010 78.500 148.250 ;
        RECT 78.820 140.410 78.960 155.390 ;
        RECT 79.670 151.115 79.950 151.485 ;
        RECT 79.220 149.950 79.480 150.270 ;
        RECT 79.280 148.230 79.420 149.950 ;
        RECT 79.220 147.910 79.480 148.230 ;
        RECT 79.740 146.610 79.880 151.115 ;
        RECT 79.280 146.530 79.880 146.610 ;
        RECT 79.280 146.470 79.940 146.530 ;
        RECT 79.280 140.410 79.420 146.470 ;
        RECT 79.680 146.210 79.940 146.470 ;
        RECT 79.670 145.675 79.950 146.045 ;
        RECT 80.200 145.850 80.340 159.470 ;
        RECT 80.660 159.110 80.800 160.635 ;
        RECT 80.600 158.790 80.860 159.110 ;
        RECT 80.600 158.110 80.860 158.430 ;
        RECT 79.680 145.530 79.940 145.675 ;
        RECT 80.140 145.530 80.400 145.850 ;
        RECT 80.660 140.410 80.800 158.110 ;
        RECT 81.120 151.970 81.260 163.890 ;
        RECT 81.980 159.130 82.240 159.450 ;
        RECT 81.510 156.555 81.790 156.925 ;
        RECT 81.520 156.410 81.780 156.555 ;
        RECT 81.520 155.730 81.780 156.050 ;
        RECT 81.580 154.690 81.720 155.730 ;
        RECT 81.520 154.370 81.780 154.690 ;
        RECT 81.060 151.650 81.320 151.970 ;
        RECT 81.510 146.355 81.790 146.725 ;
        RECT 81.580 145.850 81.720 146.355 ;
        RECT 81.520 145.530 81.780 145.850 ;
        RECT 78.760 140.090 79.020 140.410 ;
        RECT 79.220 140.090 79.480 140.410 ;
        RECT 80.600 140.090 80.860 140.410 ;
        RECT 81.520 140.090 81.780 140.410 ;
        RECT 78.760 139.410 79.020 139.730 ;
        RECT 78.820 137.350 78.960 139.410 ;
        RECT 81.060 139.070 81.320 139.390 ;
        RECT 78.760 137.030 79.020 137.350 ;
        RECT 80.140 137.030 80.400 137.350 ;
        RECT 80.600 137.030 80.860 137.350 ;
        RECT 78.300 136.690 78.560 137.010 ;
        RECT 77.380 136.350 77.640 136.670 ;
        RECT 77.840 136.350 78.100 136.670 ;
        RECT 77.900 135.310 78.040 136.350 ;
        RECT 77.840 134.990 78.100 135.310 ;
        RECT 77.840 129.210 78.100 129.530 ;
        RECT 78.300 129.210 78.560 129.530 ;
        RECT 77.900 127.005 78.040 129.210 ;
        RECT 77.830 126.635 78.110 127.005 ;
        RECT 77.840 125.470 78.100 125.790 ;
        RECT 77.380 123.770 77.640 124.090 ;
        RECT 77.440 122.050 77.580 123.770 ;
        RECT 77.900 122.050 78.040 125.470 ;
        RECT 78.360 123.070 78.500 129.210 ;
        RECT 78.820 124.770 78.960 137.030 ;
        RECT 79.220 131.765 79.480 131.910 ;
        RECT 79.210 131.395 79.490 131.765 ;
        RECT 79.220 128.190 79.480 128.510 ;
        RECT 78.760 124.450 79.020 124.770 ;
        RECT 79.280 124.170 79.420 128.190 ;
        RECT 78.820 124.030 79.420 124.170 ;
        RECT 78.300 122.750 78.560 123.070 ;
        RECT 77.380 121.730 77.640 122.050 ;
        RECT 77.840 121.730 78.100 122.050 ;
        RECT 77.840 120.710 78.100 121.030 ;
        RECT 76.920 120.600 77.180 120.690 ;
        RECT 76.920 120.460 77.580 120.600 ;
        RECT 76.920 120.370 77.180 120.460 ;
        RECT 76.920 118.330 77.180 118.650 ;
        RECT 76.460 117.310 76.720 117.630 ;
        RECT 75.990 115.755 76.270 116.125 ;
        RECT 75.540 113.570 75.800 113.890 ;
        RECT 75.080 112.210 75.340 112.530 ;
        RECT 74.620 110.850 74.880 111.170 ;
        RECT 73.760 109.070 74.360 109.210 ;
        RECT 73.760 108.110 73.900 109.070 ;
        RECT 74.680 108.360 74.820 110.850 ;
        RECT 74.220 108.220 74.820 108.360 ;
        RECT 72.840 107.710 73.440 107.850 ;
        RECT 73.700 107.790 73.960 108.110 ;
        RECT 70.940 104.390 71.200 104.710 ;
        RECT 72.320 104.390 72.580 104.710 ;
        RECT 71.000 101.310 71.140 104.390 ;
        RECT 71.860 104.050 72.120 104.370 ;
        RECT 71.920 103.010 72.060 104.050 ;
        RECT 71.860 102.690 72.120 103.010 ;
        RECT 70.940 100.990 71.200 101.310 ;
        RECT 71.000 99.270 71.140 100.990 ;
        RECT 70.940 99.180 71.200 99.270 ;
        RECT 70.940 99.040 71.600 99.180 ;
        RECT 70.940 98.950 71.200 99.040 ;
        RECT 71.460 96.550 71.600 99.040 ;
        RECT 71.860 98.610 72.120 98.930 ;
        RECT 71.920 97.570 72.060 98.610 ;
        RECT 72.840 97.570 72.980 107.710 ;
        RECT 73.760 104.280 73.900 107.790 ;
        RECT 73.300 104.140 73.900 104.280 ;
        RECT 73.300 102.670 73.440 104.140 ;
        RECT 74.220 103.770 74.360 108.220 ;
        RECT 75.140 107.770 75.280 112.210 ;
        RECT 75.600 110.150 75.740 113.570 ;
        RECT 75.540 109.830 75.800 110.150 ;
        RECT 76.060 109.470 76.200 115.755 ;
        RECT 76.980 114.910 77.120 118.330 ;
        RECT 77.440 116.610 77.580 120.460 ;
        RECT 77.900 118.650 78.040 120.710 ;
        RECT 77.840 118.330 78.100 118.650 ;
        RECT 78.300 117.990 78.560 118.310 ;
        RECT 77.380 116.290 77.640 116.610 ;
        RECT 76.920 114.590 77.180 114.910 ;
        RECT 76.450 112.355 76.730 112.725 ;
        RECT 76.520 109.810 76.660 112.355 ;
        RECT 76.980 110.150 77.120 114.590 ;
        RECT 76.920 109.830 77.180 110.150 ;
        RECT 76.460 109.490 76.720 109.810 ;
        RECT 76.000 109.150 76.260 109.470 ;
        RECT 74.620 107.450 74.880 107.770 ;
        RECT 75.080 107.450 75.340 107.770 ;
        RECT 74.680 106.750 74.820 107.450 ;
        RECT 76.920 106.770 77.180 107.090 ;
        RECT 74.620 106.430 74.880 106.750 ;
        RECT 73.760 103.630 74.360 103.770 ;
        RECT 73.760 102.670 73.900 103.630 ;
        RECT 74.150 102.835 74.430 103.205 ;
        RECT 74.160 102.690 74.420 102.835 ;
        RECT 73.240 102.350 73.500 102.670 ;
        RECT 73.700 102.350 73.960 102.670 ;
        RECT 73.700 100.200 73.960 100.290 ;
        RECT 73.300 100.060 73.960 100.200 ;
        RECT 71.860 97.250 72.120 97.570 ;
        RECT 72.780 97.250 73.040 97.570 ;
        RECT 71.850 96.715 72.130 97.085 ;
        RECT 72.780 96.800 73.040 96.890 ;
        RECT 71.400 96.230 71.660 96.550 ;
        RECT 70.930 95.355 71.210 95.725 ;
        RECT 70.480 94.530 70.740 94.850 ;
        RECT 71.000 92.130 71.140 95.355 ;
        RECT 70.940 91.810 71.200 92.130 ;
        RECT 71.460 91.450 71.600 96.230 ;
        RECT 71.400 91.130 71.660 91.450 ;
        RECT 70.480 90.450 70.740 90.770 ;
        RECT 70.540 88.390 70.680 90.450 ;
        RECT 70.480 88.070 70.740 88.390 ;
        RECT 71.400 88.070 71.660 88.390 ;
        RECT 70.080 86.010 70.680 86.090 ;
        RECT 69.560 85.690 69.820 86.010 ;
        RECT 70.080 85.950 70.740 86.010 ;
        RECT 70.480 85.690 70.740 85.950 ;
        RECT 69.100 83.310 69.360 83.630 ;
        RECT 68.640 82.290 68.900 82.610 ;
        RECT 68.640 77.870 68.900 78.190 ;
        RECT 68.700 74.110 68.840 77.870 ;
        RECT 69.160 76.830 69.300 83.310 ;
        RECT 69.620 82.010 69.760 85.690 ;
        RECT 70.020 82.805 70.280 82.950 ;
        RECT 70.010 82.435 70.290 82.805 ;
        RECT 70.020 82.010 70.280 82.270 ;
        RECT 69.620 81.950 70.280 82.010 ;
        RECT 69.620 81.870 70.220 81.950 ;
        RECT 69.620 80.570 69.760 81.870 ;
        RECT 70.540 80.910 70.680 85.690 ;
        RECT 71.460 84.990 71.600 88.070 ;
        RECT 71.400 84.670 71.660 84.990 ;
        RECT 70.480 80.590 70.740 80.910 ;
        RECT 71.920 80.650 72.060 96.715 ;
        RECT 72.380 96.660 73.040 96.800 ;
        RECT 72.380 86.690 72.520 96.660 ;
        RECT 72.780 96.570 73.040 96.660 ;
        RECT 73.300 93.830 73.440 100.060 ;
        RECT 73.700 99.970 73.960 100.060 ;
        RECT 74.680 97.650 74.820 106.430 ;
        RECT 75.540 105.410 75.800 105.730 ;
        RECT 75.080 104.050 75.340 104.370 ;
        RECT 75.140 103.010 75.280 104.050 ;
        RECT 75.600 103.010 75.740 105.410 ;
        RECT 75.080 102.690 75.340 103.010 ;
        RECT 75.540 102.690 75.800 103.010 ;
        RECT 76.980 102.330 77.120 106.770 ;
        RECT 76.920 102.010 77.180 102.330 ;
        RECT 77.440 101.990 77.580 116.290 ;
        RECT 77.840 107.790 78.100 108.110 ;
        RECT 77.900 102.330 78.040 107.790 ;
        RECT 77.840 102.010 78.100 102.330 ;
        RECT 77.380 101.670 77.640 101.990 ;
        RECT 76.920 101.330 77.180 101.650 ;
        RECT 75.990 98.755 76.270 99.125 ;
        RECT 76.060 98.590 76.200 98.755 ;
        RECT 76.000 98.270 76.260 98.590 ;
        RECT 74.220 97.510 74.820 97.650 ;
        RECT 73.240 93.510 73.500 93.830 ;
        RECT 73.700 93.510 73.960 93.830 ;
        RECT 72.780 91.130 73.040 91.450 ;
        RECT 72.840 89.410 72.980 91.130 ;
        RECT 72.780 89.090 73.040 89.410 ;
        RECT 72.320 86.370 72.580 86.690 ;
        RECT 73.300 86.090 73.440 93.510 ;
        RECT 73.760 86.690 73.900 93.510 ;
        RECT 74.220 89.070 74.360 97.510 ;
        RECT 74.620 96.910 74.880 97.230 ;
        RECT 74.160 88.750 74.420 89.070 ;
        RECT 74.220 87.450 74.360 88.750 ;
        RECT 74.680 88.390 74.820 96.910 ;
        RECT 75.080 96.570 75.340 96.890 ;
        RECT 75.140 94.850 75.280 96.570 ;
        RECT 75.540 95.550 75.800 95.870 ;
        RECT 75.080 94.530 75.340 94.850 ;
        RECT 75.600 93.830 75.740 95.550 ;
        RECT 76.980 94.850 77.120 101.330 ;
        RECT 76.920 94.530 77.180 94.850 ;
        RECT 76.000 94.190 76.260 94.510 ;
        RECT 76.980 94.365 77.120 94.530 ;
        RECT 75.540 93.510 75.800 93.830 ;
        RECT 75.600 89.410 75.740 93.510 ;
        RECT 75.540 89.090 75.800 89.410 ;
        RECT 74.620 88.070 74.880 88.390 ;
        RECT 74.220 87.310 74.820 87.450 ;
        RECT 75.080 87.390 75.340 87.710 ;
        RECT 73.700 86.370 73.960 86.690 ;
        RECT 72.840 86.010 73.440 86.090 ;
        RECT 72.780 85.950 73.440 86.010 ;
        RECT 72.780 85.690 73.040 85.950 ;
        RECT 74.150 85.835 74.430 86.205 ;
        RECT 74.160 85.690 74.420 85.835 ;
        RECT 73.230 85.155 73.510 85.525 ;
        RECT 73.700 85.350 73.960 85.670 ;
        RECT 72.310 82.435 72.590 82.805 ;
        RECT 69.560 80.250 69.820 80.570 ;
        RECT 70.540 79.890 70.680 80.590 ;
        RECT 71.460 80.510 72.060 80.650 ;
        RECT 70.480 79.570 70.740 79.890 ;
        RECT 70.020 78.210 70.280 78.530 ;
        RECT 69.100 76.510 69.360 76.830 ;
        RECT 69.100 74.470 69.360 74.790 ;
        RECT 68.640 73.790 68.900 74.110 ;
        RECT 69.160 71.390 69.300 74.470 ;
        RECT 70.080 72.750 70.220 78.210 ;
        RECT 70.940 77.190 71.200 77.510 ;
        RECT 70.470 74.955 70.750 75.325 ;
        RECT 70.480 74.810 70.740 74.955 ;
        RECT 70.020 72.430 70.280 72.750 ;
        RECT 69.560 72.090 69.820 72.410 ;
        RECT 69.100 71.070 69.360 71.390 ;
        RECT 68.630 69.515 68.910 69.885 ;
        RECT 69.620 69.690 69.760 72.090 ;
        RECT 68.180 63.590 68.440 63.910 ;
        RECT 67.720 63.250 67.980 63.570 ;
        RECT 67.720 61.210 67.980 61.530 ;
        RECT 67.250 60.675 67.530 61.045 ;
        RECT 67.320 56.770 67.460 60.675 ;
        RECT 67.780 59.490 67.920 61.210 ;
        RECT 67.720 59.170 67.980 59.490 ;
        RECT 68.240 58.720 68.380 63.590 ;
        RECT 68.700 59.490 68.840 69.515 ;
        RECT 69.560 69.370 69.820 69.690 ;
        RECT 69.100 69.030 69.360 69.350 ;
        RECT 69.160 67.310 69.300 69.030 ;
        RECT 70.080 69.010 70.220 72.430 ;
        RECT 71.000 70.370 71.140 77.190 ;
        RECT 70.940 70.050 71.200 70.370 ;
        RECT 70.020 68.690 70.280 69.010 ;
        RECT 69.560 67.330 69.820 67.650 ;
        RECT 69.100 66.990 69.360 67.310 ;
        RECT 69.620 66.540 69.760 67.330 ;
        RECT 69.160 66.400 69.760 66.540 ;
        RECT 68.640 59.170 68.900 59.490 ;
        RECT 68.240 58.580 68.840 58.720 ;
        RECT 68.170 57.955 68.450 58.325 ;
        RECT 66.340 56.540 67.000 56.680 ;
        RECT 66.340 56.450 66.600 56.540 ;
        RECT 67.260 56.450 67.520 56.770 ;
        RECT 64.500 50.330 64.760 50.650 ;
        RECT 65.870 50.475 66.150 50.845 ;
        RECT 64.560 48.805 64.700 50.330 ;
        RECT 65.940 50.310 66.080 50.475 ;
        RECT 65.880 49.990 66.140 50.310 ;
        RECT 65.420 49.650 65.680 49.970 ;
        RECT 64.490 48.435 64.770 48.805 ;
        RECT 64.500 48.290 64.760 48.435 ;
        RECT 64.560 43.170 64.700 48.290 ;
        RECT 65.480 47.930 65.620 49.650 ;
        RECT 67.320 48.370 67.460 56.450 ;
        RECT 68.240 54.050 68.380 57.955 ;
        RECT 68.180 53.730 68.440 54.050 ;
        RECT 67.320 48.230 68.380 48.370 ;
        RECT 65.420 47.610 65.680 47.930 ;
        RECT 66.800 47.610 67.060 47.930 ;
        RECT 66.340 46.590 66.600 46.910 ;
        RECT 64.500 42.850 64.760 43.170 ;
        RECT 63.180 42.430 63.780 42.570 ;
        RECT 64.040 42.510 64.300 42.830 ;
        RECT 62.660 39.450 62.920 39.770 ;
        RECT 62.720 37.390 62.860 39.450 ;
        RECT 62.660 37.070 62.920 37.390 ;
        RECT 63.180 33.990 63.320 42.430 ;
        RECT 63.580 40.130 63.840 40.450 ;
        RECT 63.120 33.670 63.380 33.990 ;
        RECT 63.640 30.590 63.780 40.130 ;
        RECT 64.100 40.110 64.240 42.510 ;
        RECT 65.420 41.830 65.680 42.150 ;
        RECT 64.960 41.150 65.220 41.470 ;
        RECT 64.040 39.790 64.300 40.110 ;
        RECT 64.500 39.110 64.760 39.430 ;
        RECT 64.030 37.555 64.310 37.925 ;
        RECT 64.100 30.590 64.240 37.555 ;
        RECT 64.560 31.950 64.700 39.110 ;
        RECT 65.020 36.370 65.160 41.150 ;
        RECT 64.960 36.050 65.220 36.370 ;
        RECT 65.020 33.650 65.160 36.050 ;
        RECT 64.960 33.330 65.220 33.650 ;
        RECT 65.480 32.290 65.620 41.830 ;
        RECT 66.400 39.285 66.540 46.590 ;
        RECT 66.860 43.170 67.000 47.610 ;
        RECT 67.260 45.570 67.520 45.890 ;
        RECT 66.800 42.850 67.060 43.170 ;
        RECT 66.800 41.830 67.060 42.150 ;
        RECT 66.330 38.915 66.610 39.285 ;
        RECT 65.880 36.730 66.140 37.050 ;
        RECT 65.940 35.010 66.080 36.730 ;
        RECT 65.880 34.690 66.140 35.010 ;
        RECT 66.400 33.990 66.540 38.915 ;
        RECT 66.860 33.990 67.000 41.830 ;
        RECT 67.320 40.450 67.460 45.570 ;
        RECT 67.720 44.550 67.980 44.870 ;
        RECT 67.260 40.130 67.520 40.450 ;
        RECT 67.780 39.430 67.920 44.550 ;
        RECT 68.240 42.400 68.380 48.230 ;
        RECT 68.700 43.170 68.840 58.580 ;
        RECT 69.160 55.750 69.300 66.400 ;
        RECT 70.080 61.870 70.220 68.690 ;
        RECT 71.000 67.730 71.140 70.050 ;
        RECT 70.540 67.590 71.140 67.730 ;
        RECT 70.540 66.630 70.680 67.590 ;
        RECT 70.940 66.990 71.200 67.310 ;
        RECT 70.480 66.310 70.740 66.630 ;
        RECT 70.480 65.630 70.740 65.950 ;
        RECT 70.540 64.930 70.680 65.630 ;
        RECT 70.480 64.610 70.740 64.930 ;
        RECT 71.000 64.590 71.140 66.990 ;
        RECT 70.940 64.270 71.200 64.590 ;
        RECT 70.940 62.910 71.200 63.230 ;
        RECT 70.020 61.550 70.280 61.870 ;
        RECT 71.000 61.190 71.140 62.910 ;
        RECT 69.560 60.870 69.820 61.190 ;
        RECT 70.940 60.870 71.200 61.190 ;
        RECT 69.620 60.510 69.760 60.870 ;
        RECT 69.560 60.190 69.820 60.510 ;
        RECT 70.010 59.995 70.290 60.365 ;
        RECT 70.480 60.190 70.740 60.510 ;
        RECT 69.560 58.490 69.820 58.810 ;
        RECT 69.620 56.090 69.760 58.490 ;
        RECT 70.080 58.130 70.220 59.995 ;
        RECT 70.540 58.810 70.680 60.190 ;
        RECT 70.480 58.490 70.740 58.810 ;
        RECT 70.020 57.810 70.280 58.130 ;
        RECT 71.000 56.770 71.140 60.870 ;
        RECT 71.460 58.470 71.600 80.510 ;
        RECT 71.860 76.510 72.120 76.830 ;
        RECT 71.920 69.350 72.060 76.510 ;
        RECT 72.380 75.130 72.520 82.435 ;
        RECT 72.780 82.290 73.040 82.610 ;
        RECT 72.840 79.890 72.980 82.290 ;
        RECT 73.300 80.570 73.440 85.155 ;
        RECT 73.760 83.370 73.900 85.350 ;
        RECT 74.680 84.050 74.820 87.310 ;
        RECT 75.140 86.010 75.280 87.390 ;
        RECT 75.530 86.090 75.810 86.205 ;
        RECT 76.060 86.090 76.200 94.190 ;
        RECT 76.910 93.995 77.190 94.365 ;
        RECT 77.440 94.170 77.580 101.670 ;
        RECT 77.900 97.230 78.040 102.010 ;
        RECT 78.360 99.805 78.500 117.990 ;
        RECT 78.820 113.550 78.960 124.030 ;
        RECT 79.220 122.750 79.480 123.070 ;
        RECT 79.280 120.690 79.420 122.750 ;
        RECT 79.220 120.370 79.480 120.690 ;
        RECT 79.680 120.370 79.940 120.690 ;
        RECT 79.740 118.310 79.880 120.370 ;
        RECT 79.680 117.990 79.940 118.310 ;
        RECT 80.200 113.890 80.340 137.030 ;
        RECT 80.660 131.910 80.800 137.030 ;
        RECT 80.600 131.590 80.860 131.910 ;
        RECT 81.120 129.725 81.260 139.070 ;
        RECT 81.580 133.950 81.720 140.090 ;
        RECT 81.520 133.630 81.780 133.950 ;
        RECT 81.050 129.355 81.330 129.725 ;
        RECT 81.060 128.870 81.320 129.190 ;
        RECT 81.120 125.790 81.260 128.870 ;
        RECT 81.060 125.470 81.320 125.790 ;
        RECT 81.120 124.430 81.260 125.470 ;
        RECT 81.060 124.110 81.320 124.430 ;
        RECT 81.120 121.030 81.260 124.110 ;
        RECT 81.060 120.710 81.320 121.030 ;
        RECT 80.600 117.990 80.860 118.310 ;
        RECT 80.140 113.570 80.400 113.890 ;
        RECT 78.760 113.230 79.020 113.550 ;
        RECT 78.290 99.435 78.570 99.805 ;
        RECT 78.300 98.950 78.560 99.270 ;
        RECT 77.840 96.910 78.100 97.230 ;
        RECT 78.360 97.085 78.500 98.950 ;
        RECT 77.380 93.850 77.640 94.170 ;
        RECT 76.920 93.510 77.180 93.830 ;
        RECT 76.980 92.130 77.120 93.510 ;
        RECT 76.920 91.810 77.180 92.130 ;
        RECT 76.920 90.170 77.180 90.430 ;
        RECT 76.520 90.110 77.180 90.170 ;
        RECT 76.520 90.030 77.120 90.110 ;
        RECT 76.520 88.050 76.660 90.030 ;
        RECT 76.460 87.730 76.720 88.050 ;
        RECT 76.520 86.350 76.660 87.730 ;
        RECT 75.080 85.690 75.340 86.010 ;
        RECT 75.530 85.950 76.200 86.090 ;
        RECT 76.460 86.030 76.720 86.350 ;
        RECT 75.530 85.835 75.810 85.950 ;
        RECT 76.920 85.690 77.180 86.010 ;
        RECT 75.080 85.010 75.340 85.330 ;
        RECT 75.990 85.155 76.270 85.525 ;
        RECT 76.000 85.010 76.260 85.155 ;
        RECT 75.140 84.730 75.280 85.010 ;
        RECT 75.140 84.590 76.200 84.730 ;
        RECT 74.680 83.910 75.740 84.050 ;
        RECT 73.760 83.230 74.820 83.370 ;
        RECT 73.700 82.805 73.960 82.950 ;
        RECT 73.690 82.435 73.970 82.805 ;
        RECT 74.160 82.290 74.420 82.610 ;
        RECT 73.240 80.250 73.500 80.570 ;
        RECT 72.780 79.570 73.040 79.890 ;
        RECT 72.320 74.810 72.580 75.130 ;
        RECT 72.840 72.070 72.980 79.570 ;
        RECT 73.300 78.530 73.440 80.250 ;
        RECT 74.220 78.530 74.360 82.290 ;
        RECT 74.680 80.910 74.820 83.230 ;
        RECT 75.600 82.610 75.740 83.910 ;
        RECT 75.540 82.290 75.800 82.610 ;
        RECT 75.080 81.950 75.340 82.270 ;
        RECT 76.060 82.125 76.200 84.590 ;
        RECT 76.980 83.970 77.120 85.690 ;
        RECT 77.440 84.990 77.580 93.850 ;
        RECT 77.900 93.830 78.040 96.910 ;
        RECT 78.290 96.715 78.570 97.085 ;
        RECT 78.820 94.250 78.960 113.230 ;
        RECT 79.680 109.830 79.940 110.150 ;
        RECT 80.140 109.830 80.400 110.150 ;
        RECT 79.220 109.325 79.480 109.470 ;
        RECT 79.210 108.955 79.490 109.325 ;
        RECT 79.220 107.680 79.480 107.770 ;
        RECT 79.740 107.680 79.880 109.830 ;
        RECT 80.200 108.450 80.340 109.830 ;
        RECT 80.140 108.130 80.400 108.450 ;
        RECT 79.220 107.540 79.880 107.680 ;
        RECT 79.220 107.450 79.480 107.540 ;
        RECT 79.220 106.770 79.480 107.090 ;
        RECT 78.360 94.110 78.960 94.250 ;
        RECT 77.840 93.510 78.100 93.830 ;
        RECT 78.360 92.210 78.500 94.110 ;
        RECT 78.760 93.170 79.020 93.490 ;
        RECT 77.900 92.070 78.500 92.210 ;
        RECT 77.900 88.730 78.040 92.070 ;
        RECT 78.820 91.790 78.960 93.170 ;
        RECT 78.760 91.470 79.020 91.790 ;
        RECT 79.280 91.450 79.420 106.770 ;
        RECT 79.740 104.030 79.880 107.540 ;
        RECT 80.140 107.450 80.400 107.770 ;
        RECT 79.680 103.710 79.940 104.030 ;
        RECT 79.740 99.270 79.880 103.710 ;
        RECT 80.200 103.205 80.340 107.450 ;
        RECT 80.130 102.835 80.410 103.205 ;
        RECT 80.660 102.920 80.800 117.990 ;
        RECT 81.580 113.210 81.720 133.630 ;
        RECT 82.040 120.690 82.180 159.130 ;
        RECT 81.980 120.370 82.240 120.690 ;
        RECT 82.500 118.990 82.640 165.250 ;
        RECT 82.440 118.670 82.700 118.990 ;
        RECT 82.500 113.550 82.640 118.670 ;
        RECT 82.440 113.230 82.700 113.550 ;
        RECT 81.520 112.890 81.780 113.210 ;
        RECT 81.060 109.150 81.320 109.470 ;
        RECT 81.120 105.925 81.260 109.150 ;
        RECT 82.500 107.430 82.640 113.230 ;
        RECT 82.440 107.110 82.700 107.430 ;
        RECT 81.520 106.430 81.780 106.750 ;
        RECT 81.050 105.555 81.330 105.925 ;
        RECT 80.200 102.330 80.340 102.835 ;
        RECT 80.660 102.780 81.260 102.920 ;
        RECT 80.140 102.010 80.400 102.330 ;
        RECT 80.600 102.010 80.860 102.330 ;
        RECT 80.660 100.290 80.800 102.010 ;
        RECT 80.600 99.970 80.860 100.290 ;
        RECT 81.120 99.270 81.260 102.780 ;
        RECT 81.580 102.525 81.720 106.430 ;
        RECT 81.510 102.155 81.790 102.525 ;
        RECT 81.520 101.670 81.780 101.990 ;
        RECT 81.580 99.610 81.720 101.670 ;
        RECT 81.520 99.290 81.780 99.610 ;
        RECT 81.970 99.435 82.250 99.805 ;
        RECT 79.680 98.950 79.940 99.270 ;
        RECT 81.060 98.950 81.320 99.270 ;
        RECT 80.140 98.270 80.400 98.590 ;
        RECT 79.680 95.550 79.940 95.870 ;
        RECT 79.740 93.490 79.880 95.550 ;
        RECT 80.200 93.490 80.340 98.270 ;
        RECT 80.600 93.740 80.860 93.830 ;
        RECT 81.120 93.740 81.260 98.950 ;
        RECT 80.600 93.600 81.260 93.740 ;
        RECT 81.520 93.685 81.780 93.830 ;
        RECT 80.600 93.510 80.860 93.600 ;
        RECT 79.680 93.170 79.940 93.490 ;
        RECT 80.140 93.170 80.400 93.490 ;
        RECT 81.510 93.315 81.790 93.685 ;
        RECT 78.300 91.130 78.560 91.450 ;
        RECT 79.220 91.130 79.480 91.450 ;
        RECT 77.840 88.410 78.100 88.730 ;
        RECT 78.360 88.050 78.500 91.130 ;
        RECT 80.200 88.130 80.340 93.170 ;
        RECT 81.060 88.410 81.320 88.730 ;
        RECT 81.510 88.555 81.790 88.925 ;
        RECT 78.300 87.730 78.560 88.050 ;
        RECT 79.220 87.730 79.480 88.050 ;
        RECT 80.200 87.990 80.800 88.130 ;
        RECT 77.840 85.350 78.100 85.670 ;
        RECT 77.380 84.670 77.640 84.990 ;
        RECT 76.920 83.650 77.180 83.970 ;
        RECT 77.440 83.290 77.580 84.670 ;
        RECT 77.900 84.165 78.040 85.350 ;
        RECT 77.830 83.795 78.110 84.165 ;
        RECT 77.380 82.970 77.640 83.290 ;
        RECT 74.620 80.590 74.880 80.910 ;
        RECT 73.240 78.210 73.500 78.530 ;
        RECT 74.160 78.440 74.420 78.530 ;
        RECT 73.760 78.300 74.420 78.440 ;
        RECT 73.300 76.830 73.440 78.210 ;
        RECT 73.240 76.510 73.500 76.830 ;
        RECT 73.230 74.955 73.510 75.325 ;
        RECT 73.760 75.130 73.900 78.300 ;
        RECT 74.160 78.210 74.420 78.300 ;
        RECT 74.680 77.510 74.820 80.590 ;
        RECT 75.140 77.850 75.280 81.950 ;
        RECT 75.990 81.755 76.270 82.125 ;
        RECT 77.840 81.950 78.100 82.270 ;
        RECT 75.530 81.075 75.810 81.445 ;
        RECT 75.080 77.530 75.340 77.850 ;
        RECT 74.620 77.190 74.880 77.510 ;
        RECT 72.780 71.750 73.040 72.070 ;
        RECT 72.840 69.350 72.980 71.750 ;
        RECT 71.860 69.030 72.120 69.350 ;
        RECT 72.780 69.030 73.040 69.350 ;
        RECT 71.920 67.050 72.060 69.030 ;
        RECT 71.920 66.970 72.520 67.050 ;
        RECT 71.860 66.910 72.520 66.970 ;
        RECT 71.860 66.650 72.120 66.910 ;
        RECT 71.860 63.930 72.120 64.250 ;
        RECT 71.920 59.570 72.060 63.930 ;
        RECT 72.380 60.365 72.520 66.910 ;
        RECT 72.840 60.850 72.980 69.030 ;
        RECT 73.300 65.950 73.440 74.955 ;
        RECT 73.700 74.810 73.960 75.130 ;
        RECT 74.160 74.130 74.420 74.450 ;
        RECT 73.700 73.790 73.960 74.110 ;
        RECT 73.760 72.070 73.900 73.790 ;
        RECT 73.700 71.750 73.960 72.070 ;
        RECT 73.700 65.970 73.960 66.290 ;
        RECT 73.240 65.630 73.500 65.950 ;
        RECT 73.760 63.910 73.900 65.970 ;
        RECT 73.240 63.590 73.500 63.910 ;
        RECT 73.700 63.590 73.960 63.910 ;
        RECT 73.300 61.870 73.440 63.590 ;
        RECT 73.240 61.550 73.500 61.870 ;
        RECT 72.780 60.530 73.040 60.850 ;
        RECT 73.760 60.510 73.900 63.590 ;
        RECT 74.220 63.230 74.360 74.130 ;
        RECT 74.680 71.390 74.820 77.190 ;
        RECT 75.080 75.040 75.340 75.130 ;
        RECT 75.600 75.040 75.740 81.075 ;
        RECT 76.460 80.930 76.720 81.250 ;
        RECT 76.520 78.725 76.660 80.930 ;
        RECT 77.900 80.910 78.040 81.950 ;
        RECT 77.840 80.590 78.100 80.910 ;
        RECT 78.360 80.570 78.500 87.730 ;
        RECT 78.760 85.690 79.020 86.010 ;
        RECT 78.820 83.485 78.960 85.690 ;
        RECT 78.750 83.115 79.030 83.485 ;
        RECT 78.760 82.290 79.020 82.610 ;
        RECT 78.820 81.445 78.960 82.290 ;
        RECT 78.750 81.075 79.030 81.445 ;
        RECT 78.300 80.250 78.560 80.570 ;
        RECT 79.280 79.550 79.420 87.730 ;
        RECT 80.140 87.390 80.400 87.710 ;
        RECT 80.200 82.950 80.340 87.390 ;
        RECT 80.140 82.630 80.400 82.950 ;
        RECT 79.220 79.230 79.480 79.550 ;
        RECT 80.140 79.230 80.400 79.550 ;
        RECT 76.450 78.355 76.730 78.725 ;
        RECT 76.450 77.675 76.730 78.045 ;
        RECT 76.520 77.510 76.660 77.675 ;
        RECT 80.200 77.510 80.340 79.230 ;
        RECT 80.660 77.510 80.800 87.990 ;
        RECT 76.460 77.190 76.720 77.510 ;
        RECT 77.840 77.190 78.100 77.510 ;
        RECT 80.140 77.190 80.400 77.510 ;
        RECT 80.600 77.190 80.860 77.510 ;
        RECT 75.080 74.900 75.740 75.040 ;
        RECT 75.080 74.810 75.340 74.900 ;
        RECT 75.140 74.450 75.280 74.810 ;
        RECT 75.080 74.130 75.340 74.450 ;
        RECT 75.540 73.790 75.800 74.110 ;
        RECT 74.620 71.070 74.880 71.390 ;
        RECT 74.680 64.250 74.820 71.070 ;
        RECT 75.600 70.030 75.740 73.790 ;
        RECT 76.000 72.770 76.260 73.090 ;
        RECT 76.060 71.130 76.200 72.770 ;
        RECT 76.520 71.730 76.660 77.190 ;
        RECT 76.910 75.635 77.190 76.005 ;
        RECT 76.980 75.130 77.120 75.635 ;
        RECT 76.920 74.810 77.180 75.130 ;
        RECT 76.460 71.410 76.720 71.730 ;
        RECT 76.060 70.990 76.660 71.130 ;
        RECT 76.000 70.050 76.260 70.370 ;
        RECT 75.540 69.710 75.800 70.030 ;
        RECT 75.540 67.330 75.800 67.650 ;
        RECT 75.600 64.930 75.740 67.330 ;
        RECT 76.060 66.630 76.200 70.050 ;
        RECT 76.520 66.970 76.660 70.990 ;
        RECT 76.980 69.090 77.120 74.810 ;
        RECT 76.980 68.950 77.580 69.090 ;
        RECT 76.910 68.155 77.190 68.525 ;
        RECT 76.980 67.650 77.120 68.155 ;
        RECT 76.920 67.330 77.180 67.650 ;
        RECT 76.460 66.650 76.720 66.970 ;
        RECT 76.000 66.310 76.260 66.630 ;
        RECT 76.460 65.970 76.720 66.290 ;
        RECT 75.540 64.610 75.800 64.930 ;
        RECT 74.620 63.930 74.880 64.250 ;
        RECT 74.160 62.910 74.420 63.230 ;
        RECT 74.680 61.610 74.820 63.930 ;
        RECT 76.000 63.590 76.260 63.910 ;
        RECT 75.080 61.890 75.340 62.210 ;
        RECT 76.060 62.170 76.200 63.590 ;
        RECT 75.600 62.030 76.200 62.170 ;
        RECT 75.140 61.725 75.280 61.890 ;
        RECT 74.220 61.470 74.820 61.610 ;
        RECT 72.310 59.995 72.590 60.365 ;
        RECT 73.700 60.190 73.960 60.510 ;
        RECT 71.920 59.430 72.980 59.570 ;
        RECT 71.850 58.635 72.130 59.005 ;
        RECT 71.860 58.490 72.120 58.635 ;
        RECT 71.400 58.150 71.660 58.470 ;
        RECT 70.940 56.450 71.200 56.770 ;
        RECT 69.560 55.770 69.820 56.090 ;
        RECT 69.100 55.430 69.360 55.750 ;
        RECT 69.160 48.270 69.300 55.430 ;
        RECT 71.460 55.410 71.600 58.150 ;
        RECT 71.860 57.470 72.120 57.790 ;
        RECT 72.840 57.530 72.980 59.430 ;
        RECT 69.560 55.090 69.820 55.410 ;
        RECT 71.400 55.090 71.660 55.410 ;
        RECT 69.100 47.950 69.360 48.270 ;
        RECT 69.100 44.780 69.360 44.870 ;
        RECT 69.620 44.780 69.760 55.090 ;
        RECT 70.480 54.750 70.740 55.070 ;
        RECT 70.540 53.370 70.680 54.750 ;
        RECT 71.920 53.370 72.060 57.470 ;
        RECT 72.380 57.390 72.980 57.530 ;
        RECT 72.380 55.750 72.520 57.390 ;
        RECT 72.780 56.450 73.040 56.770 ;
        RECT 72.840 55.750 72.980 56.450 ;
        RECT 72.320 55.430 72.580 55.750 ;
        RECT 72.780 55.430 73.040 55.750 ;
        RECT 72.380 53.370 72.520 55.430 ;
        RECT 70.480 53.050 70.740 53.370 ;
        RECT 71.860 53.050 72.120 53.370 ;
        RECT 72.320 53.050 72.580 53.370 ;
        RECT 70.020 52.030 70.280 52.350 ;
        RECT 70.080 50.310 70.220 52.030 ;
        RECT 70.480 50.730 70.740 50.990 ;
        RECT 72.380 50.730 72.520 53.050 ;
        RECT 70.480 50.670 72.520 50.730 ;
        RECT 70.540 50.590 72.520 50.670 ;
        RECT 70.020 49.990 70.280 50.310 ;
        RECT 69.100 44.640 69.760 44.780 ;
        RECT 69.100 44.550 69.360 44.640 ;
        RECT 68.640 42.850 68.900 43.170 ;
        RECT 68.640 42.400 68.900 42.490 ;
        RECT 68.240 42.260 68.900 42.400 ;
        RECT 68.640 42.170 68.900 42.260 ;
        RECT 67.720 39.110 67.980 39.430 ;
        RECT 68.180 39.110 68.440 39.430 ;
        RECT 68.640 39.110 68.900 39.430 ;
        RECT 68.240 37.730 68.380 39.110 ;
        RECT 68.180 37.410 68.440 37.730 ;
        RECT 68.700 33.990 68.840 39.110 ;
        RECT 66.340 33.670 66.600 33.990 ;
        RECT 66.800 33.670 67.060 33.990 ;
        RECT 67.720 33.670 67.980 33.990 ;
        RECT 68.640 33.670 68.900 33.990 ;
        RECT 65.880 32.990 66.140 33.310 ;
        RECT 66.860 33.165 67.000 33.670 ;
        RECT 65.420 31.970 65.680 32.290 ;
        RECT 64.500 31.630 64.760 31.950 ;
        RECT 65.940 31.805 66.080 32.990 ;
        RECT 66.790 32.795 67.070 33.165 ;
        RECT 65.870 31.435 66.150 31.805 ;
        RECT 63.580 30.270 63.840 30.590 ;
        RECT 64.040 30.270 64.300 30.590 ;
        RECT 64.030 29.395 64.310 29.765 ;
        RECT 64.100 28.550 64.240 29.395 ;
        RECT 61.280 28.230 61.540 28.550 ;
        RECT 64.040 28.230 64.300 28.550 ;
        RECT 65.420 27.890 65.680 28.210 ;
        RECT 61.740 27.725 62.000 27.870 ;
        RECT 61.730 27.355 62.010 27.725 ;
        RECT 63.580 26.530 63.840 26.850 ;
        RECT 64.950 26.675 65.230 27.045 ;
        RECT 60.360 25.510 60.620 25.830 ;
        RECT 60.820 25.510 61.080 25.830 ;
        RECT 58.520 24.830 58.780 25.150 ;
        RECT 58.580 23.110 58.720 24.830 ;
        RECT 58.520 22.790 58.780 23.110 ;
        RECT 58.060 22.450 58.320 22.770 ;
        RECT 58.120 21.605 58.260 22.450 ;
        RECT 60.420 22.430 60.560 25.510 ;
        RECT 60.360 22.110 60.620 22.430 ;
        RECT 58.050 21.235 58.330 21.605 ;
        RECT 58.060 21.090 58.320 21.235 ;
        RECT 60.880 18.690 61.020 25.510 ;
        RECT 62.200 24.830 62.460 25.150 ;
        RECT 60.820 18.370 61.080 18.690 ;
        RECT 59.900 17.690 60.160 18.010 ;
        RECT 57.600 17.010 57.860 17.330 ;
        RECT 56.220 15.650 56.480 15.970 ;
        RECT 59.960 15.630 60.100 17.690 ;
        RECT 62.260 17.330 62.400 24.830 ;
        RECT 63.640 24.130 63.780 26.530 ;
        RECT 64.490 25.995 64.770 26.365 ;
        RECT 64.500 25.850 64.760 25.995 ;
        RECT 65.020 25.830 65.160 26.675 ;
        RECT 64.960 25.510 65.220 25.830 ;
        RECT 64.500 25.170 64.760 25.490 ;
        RECT 63.580 23.810 63.840 24.130 ;
        RECT 64.560 23.450 64.700 25.170 ;
        RECT 64.500 23.130 64.760 23.450 ;
        RECT 64.500 22.110 64.760 22.430 ;
        RECT 64.560 21.070 64.700 22.110 ;
        RECT 64.500 20.750 64.760 21.070 ;
        RECT 65.480 17.670 65.620 27.890 ;
        RECT 66.860 26.510 67.000 32.795 ;
        RECT 67.780 32.290 67.920 33.670 ;
        RECT 68.180 32.990 68.440 33.310 ;
        RECT 67.720 31.970 67.980 32.290 ;
        RECT 68.240 31.690 68.380 32.990 ;
        RECT 67.780 31.610 68.380 31.690 ;
        RECT 67.720 31.550 68.380 31.610 ;
        RECT 67.720 31.290 67.980 31.550 ;
        RECT 69.160 31.520 69.300 44.550 ;
        RECT 69.560 43.870 69.820 44.190 ;
        RECT 69.620 42.490 69.760 43.870 ;
        RECT 70.080 42.490 70.220 49.990 ;
        RECT 70.940 47.950 71.200 48.270 ;
        RECT 69.560 42.170 69.820 42.490 ;
        RECT 70.020 42.170 70.280 42.490 ;
        RECT 70.080 39.430 70.220 42.170 ;
        RECT 70.020 39.110 70.280 39.430 ;
        RECT 70.020 35.710 70.280 36.030 ;
        RECT 70.080 33.990 70.220 35.710 ;
        RECT 71.000 33.990 71.140 47.950 ;
        RECT 72.380 47.330 72.520 50.590 ;
        RECT 72.840 48.610 72.980 55.430 ;
        RECT 72.780 48.290 73.040 48.610 ;
        RECT 73.760 47.930 73.900 60.190 ;
        RECT 74.220 59.150 74.360 61.470 ;
        RECT 75.070 61.355 75.350 61.725 ;
        RECT 74.620 60.530 74.880 60.850 ;
        RECT 74.160 58.830 74.420 59.150 ;
        RECT 74.680 58.810 74.820 60.530 ;
        RECT 75.600 59.490 75.740 62.030 ;
        RECT 76.520 61.530 76.660 65.970 ;
        RECT 77.440 62.170 77.580 68.950 ;
        RECT 77.900 67.650 78.040 77.190 ;
        RECT 78.300 74.810 78.560 75.130 ;
        RECT 79.680 74.810 79.940 75.130 ;
        RECT 80.140 74.810 80.400 75.130 ;
        RECT 78.360 73.090 78.500 74.810 ;
        RECT 79.740 74.450 79.880 74.810 ;
        RECT 79.680 74.130 79.940 74.450 ;
        RECT 78.300 72.770 78.560 73.090 ;
        RECT 78.300 71.750 78.560 72.070 ;
        RECT 78.360 68.670 78.500 71.750 ;
        RECT 78.300 68.350 78.560 68.670 ;
        RECT 77.840 67.330 78.100 67.650 ;
        RECT 78.360 64.250 78.500 68.350 ;
        RECT 78.760 65.630 79.020 65.950 ;
        RECT 78.820 64.250 78.960 65.630 ;
        RECT 78.300 63.930 78.560 64.250 ;
        RECT 78.760 63.930 79.020 64.250 ;
        RECT 79.220 63.930 79.480 64.250 ;
        RECT 79.280 63.085 79.420 63.930 ;
        RECT 79.210 62.715 79.490 63.085 ;
        RECT 79.740 62.290 79.880 74.130 ;
        RECT 80.200 71.390 80.340 74.810 ;
        RECT 80.660 72.750 80.800 77.190 ;
        RECT 81.120 75.470 81.260 88.410 ;
        RECT 81.580 88.390 81.720 88.555 ;
        RECT 81.520 88.070 81.780 88.390 ;
        RECT 81.520 87.390 81.780 87.710 ;
        RECT 81.580 82.950 81.720 87.390 ;
        RECT 82.040 85.670 82.180 99.435 ;
        RECT 81.980 85.350 82.240 85.670 ;
        RECT 81.520 82.630 81.780 82.950 ;
        RECT 81.980 77.190 82.240 77.510 ;
        RECT 81.060 75.150 81.320 75.470 ;
        RECT 80.600 72.430 80.860 72.750 ;
        RECT 81.120 71.730 81.260 75.150 ;
        RECT 81.510 74.955 81.790 75.325 ;
        RECT 81.060 71.410 81.320 71.730 ;
        RECT 80.140 71.130 80.400 71.390 ;
        RECT 80.140 71.070 80.800 71.130 ;
        RECT 80.200 70.990 80.800 71.070 ;
        RECT 80.140 69.370 80.400 69.690 ;
        RECT 80.200 64.930 80.340 69.370 ;
        RECT 80.660 66.630 80.800 70.990 ;
        RECT 81.060 70.050 81.320 70.370 ;
        RECT 80.600 66.310 80.860 66.630 ;
        RECT 80.140 64.610 80.400 64.930 ;
        RECT 76.980 62.030 77.580 62.170 ;
        RECT 79.280 62.150 79.880 62.290 ;
        RECT 76.460 61.210 76.720 61.530 ;
        RECT 76.000 60.190 76.260 60.510 ;
        RECT 75.540 59.170 75.800 59.490 ;
        RECT 74.620 58.490 74.880 58.810 ;
        RECT 74.160 58.150 74.420 58.470 ;
        RECT 74.220 56.770 74.360 58.150 ;
        RECT 74.160 56.450 74.420 56.770 ;
        RECT 74.680 56.090 74.820 58.490 ;
        RECT 75.540 57.530 75.800 57.790 ;
        RECT 75.140 57.470 75.800 57.530 ;
        RECT 75.140 57.390 75.740 57.470 ;
        RECT 74.620 55.770 74.880 56.090 ;
        RECT 74.680 53.030 74.820 55.770 ;
        RECT 75.140 54.050 75.280 57.390 ;
        RECT 76.060 55.750 76.200 60.190 ;
        RECT 76.000 55.430 76.260 55.750 ;
        RECT 76.460 55.090 76.720 55.410 ;
        RECT 76.520 54.050 76.660 55.090 ;
        RECT 75.080 53.730 75.340 54.050 ;
        RECT 76.460 53.730 76.720 54.050 ;
        RECT 76.980 53.280 77.120 62.030 ;
        RECT 77.380 61.045 77.640 61.190 ;
        RECT 77.370 60.675 77.650 61.045 ;
        RECT 78.300 60.870 78.560 61.190 ;
        RECT 78.760 61.100 79.020 61.190 ;
        RECT 79.280 61.100 79.420 62.150 ;
        RECT 79.680 61.210 79.940 61.530 ;
        RECT 78.760 60.960 79.420 61.100 ;
        RECT 78.760 60.870 79.020 60.960 ;
        RECT 77.840 60.190 78.100 60.510 ;
        RECT 77.900 59.005 78.040 60.190 ;
        RECT 77.830 58.635 78.110 59.005 ;
        RECT 77.380 53.280 77.640 53.370 ;
        RECT 76.980 53.140 77.640 53.280 ;
        RECT 77.380 53.050 77.640 53.140 ;
        RECT 74.160 52.710 74.420 53.030 ;
        RECT 74.620 52.710 74.880 53.030 ;
        RECT 74.220 49.630 74.360 52.710 ;
        RECT 76.000 52.030 76.260 52.350 ;
        RECT 76.060 51.525 76.200 52.030 ;
        RECT 75.990 51.155 76.270 51.525 ;
        RECT 76.460 51.010 76.720 51.330 ;
        RECT 74.160 49.310 74.420 49.630 ;
        RECT 74.220 48.270 74.360 49.310 ;
        RECT 74.160 47.950 74.420 48.270 ;
        RECT 73.700 47.610 73.960 47.930 ;
        RECT 75.080 47.610 75.340 47.930 ;
        RECT 71.920 47.190 72.520 47.330 ;
        RECT 71.920 41.810 72.060 47.190 ;
        RECT 72.770 47.075 73.050 47.445 ;
        RECT 72.780 46.930 73.040 47.075 ;
        RECT 72.320 46.590 72.580 46.910 ;
        RECT 73.240 46.590 73.500 46.910 ;
        RECT 72.380 45.550 72.520 46.590 ;
        RECT 72.320 45.230 72.580 45.550 ;
        RECT 73.300 42.830 73.440 46.590 ;
        RECT 73.240 42.510 73.500 42.830 ;
        RECT 71.860 41.490 72.120 41.810 ;
        RECT 71.920 39.430 72.060 41.490 ;
        RECT 71.400 39.110 71.660 39.430 ;
        RECT 71.860 39.110 72.120 39.430 ;
        RECT 72.320 39.285 72.580 39.430 ;
        RECT 70.020 33.670 70.280 33.990 ;
        RECT 70.940 33.670 71.200 33.990 ;
        RECT 69.560 31.520 69.820 31.610 ;
        RECT 69.160 31.380 69.820 31.520 ;
        RECT 69.560 31.290 69.820 31.380 ;
        RECT 67.780 28.210 67.920 31.290 ;
        RECT 68.180 31.010 68.440 31.270 ;
        RECT 68.180 30.950 69.300 31.010 ;
        RECT 68.240 30.870 69.300 30.950 ;
        RECT 69.160 30.590 69.300 30.870 ;
        RECT 68.640 30.270 68.900 30.590 ;
        RECT 69.100 30.270 69.360 30.590 ;
        RECT 67.720 27.890 67.980 28.210 ;
        RECT 68.180 27.550 68.440 27.870 ;
        RECT 66.800 26.190 67.060 26.510 ;
        RECT 68.240 25.490 68.380 27.550 ;
        RECT 68.700 26.250 68.840 30.270 ;
        RECT 69.620 28.890 69.760 31.290 ;
        RECT 70.080 31.270 70.220 33.670 ;
        RECT 70.020 30.950 70.280 31.270 ;
        RECT 70.480 30.950 70.740 31.270 ;
        RECT 69.560 28.570 69.820 28.890 ;
        RECT 69.100 27.890 69.360 28.210 ;
        RECT 69.160 27.045 69.300 27.890 ;
        RECT 69.090 26.675 69.370 27.045 ;
        RECT 69.100 26.250 69.360 26.510 ;
        RECT 68.700 26.190 69.360 26.250 ;
        RECT 68.700 26.110 69.300 26.190 ;
        RECT 69.560 25.850 69.820 26.170 ;
        RECT 69.620 25.490 69.760 25.850 ;
        RECT 68.180 25.170 68.440 25.490 ;
        RECT 69.560 25.170 69.820 25.490 ;
        RECT 66.800 24.830 67.060 25.150 ;
        RECT 66.860 20.730 67.000 24.830 ;
        RECT 69.100 20.750 69.360 21.070 ;
        RECT 66.800 20.410 67.060 20.730 ;
        RECT 65.420 17.350 65.680 17.670 ;
        RECT 62.200 17.010 62.460 17.330 ;
        RECT 69.160 15.630 69.300 20.750 ;
        RECT 69.620 18.350 69.760 25.170 ;
        RECT 69.560 18.030 69.820 18.350 ;
        RECT 69.560 17.010 69.820 17.330 ;
        RECT 69.620 15.970 69.760 17.010 ;
        RECT 69.560 15.650 69.820 15.970 ;
        RECT 59.900 15.310 60.160 15.630 ;
        RECT 69.100 15.310 69.360 15.630 ;
        RECT 54.380 14.630 54.640 14.950 ;
        RECT 54.840 14.630 55.100 14.950 ;
        RECT 54.440 12.910 54.580 14.630 ;
        RECT 69.100 14.290 69.360 14.610 ;
        RECT 54.380 12.590 54.640 12.910 ;
        RECT 46.560 12.250 46.820 12.570 ;
        RECT 69.160 12.230 69.300 14.290 ;
        RECT 69.620 12.230 69.760 15.650 ;
        RECT 70.080 12.230 70.220 30.950 ;
        RECT 70.540 29.570 70.680 30.950 ;
        RECT 70.480 29.250 70.740 29.570 ;
        RECT 71.000 29.230 71.140 33.670 ;
        RECT 71.460 32.290 71.600 39.110 ;
        RECT 72.310 38.915 72.590 39.285 ;
        RECT 73.760 39.170 73.900 47.610 ;
        RECT 74.620 44.550 74.880 44.870 ;
        RECT 74.160 43.870 74.420 44.190 ;
        RECT 74.680 43.930 74.820 44.550 ;
        RECT 75.140 44.530 75.280 47.610 ;
        RECT 76.000 44.610 76.260 44.870 ;
        RECT 76.520 44.725 76.660 51.010 ;
        RECT 75.600 44.550 76.260 44.610 ;
        RECT 75.080 44.210 75.340 44.530 ;
        RECT 75.600 44.470 76.200 44.550 ;
        RECT 74.220 42.830 74.360 43.870 ;
        RECT 74.680 43.790 75.280 43.930 ;
        RECT 74.160 42.510 74.420 42.830 ;
        RECT 74.620 41.830 74.880 42.150 ;
        RECT 74.160 39.790 74.420 40.110 ;
        RECT 73.300 39.030 73.900 39.170 ;
        RECT 72.780 35.710 73.040 36.030 ;
        RECT 72.320 34.690 72.580 35.010 ;
        RECT 72.380 34.525 72.520 34.690 ;
        RECT 72.310 34.155 72.590 34.525 ;
        RECT 72.840 33.650 72.980 35.710 ;
        RECT 73.300 33.990 73.440 39.030 ;
        RECT 74.220 38.750 74.360 39.790 ;
        RECT 74.680 39.770 74.820 41.830 ;
        RECT 74.620 39.450 74.880 39.770 ;
        RECT 73.700 38.430 73.960 38.750 ;
        RECT 74.160 38.430 74.420 38.750 ;
        RECT 73.760 37.050 73.900 38.430 ;
        RECT 74.680 37.390 74.820 39.450 ;
        RECT 75.140 38.750 75.280 43.790 ;
        RECT 75.600 39.090 75.740 44.470 ;
        RECT 76.450 44.355 76.730 44.725 ;
        RECT 76.920 44.550 77.180 44.870 ;
        RECT 76.000 41.150 76.260 41.470 ;
        RECT 76.060 39.430 76.200 41.150 ;
        RECT 76.000 39.110 76.260 39.430 ;
        RECT 75.540 38.770 75.800 39.090 ;
        RECT 75.080 38.430 75.340 38.750 ;
        RECT 74.620 37.070 74.880 37.390 ;
        RECT 73.700 36.730 73.960 37.050 ;
        RECT 74.680 34.330 74.820 37.070 ;
        RECT 74.620 34.010 74.880 34.330 ;
        RECT 73.240 33.670 73.500 33.990 ;
        RECT 71.860 33.330 72.120 33.650 ;
        RECT 72.780 33.330 73.040 33.650 ;
        RECT 71.400 31.970 71.660 32.290 ;
        RECT 71.920 31.610 72.060 33.330 ;
        RECT 72.320 32.990 72.580 33.310 ;
        RECT 72.380 31.950 72.520 32.990 ;
        RECT 73.300 31.950 73.440 33.670 ;
        RECT 72.320 31.630 72.580 31.950 ;
        RECT 73.240 31.630 73.500 31.950 ;
        RECT 71.860 31.290 72.120 31.610 ;
        RECT 72.780 31.290 73.040 31.610 ;
        RECT 70.940 28.910 71.200 29.230 ;
        RECT 70.940 28.460 71.200 28.550 ;
        RECT 70.940 28.320 72.520 28.460 ;
        RECT 70.940 28.230 71.200 28.320 ;
        RECT 70.940 27.780 71.200 27.870 ;
        RECT 71.860 27.780 72.120 27.870 ;
        RECT 70.940 27.640 72.120 27.780 ;
        RECT 70.940 27.550 71.200 27.640 ;
        RECT 70.940 25.510 71.200 25.830 ;
        RECT 71.000 18.690 71.140 25.510 ;
        RECT 71.460 24.130 71.600 27.640 ;
        RECT 71.860 27.550 72.120 27.640 ;
        RECT 71.860 25.850 72.120 26.170 ;
        RECT 71.920 25.150 72.060 25.850 ;
        RECT 71.860 24.830 72.120 25.150 ;
        RECT 71.400 23.810 71.660 24.130 ;
        RECT 71.860 22.790 72.120 23.110 ;
        RECT 70.940 18.370 71.200 18.690 ;
        RECT 70.480 16.670 70.740 16.990 ;
        RECT 70.540 15.290 70.680 16.670 ;
        RECT 71.000 15.290 71.140 18.370 ;
        RECT 71.920 17.670 72.060 22.790 ;
        RECT 72.380 19.710 72.520 28.320 ;
        RECT 72.840 28.210 72.980 31.290 ;
        RECT 73.300 28.550 73.440 31.630 ;
        RECT 73.690 30.075 73.970 30.445 ;
        RECT 73.760 29.230 73.900 30.075 ;
        RECT 73.700 28.910 73.960 29.230 ;
        RECT 73.240 28.230 73.500 28.550 ;
        RECT 72.780 27.890 73.040 28.210 ;
        RECT 73.690 28.035 73.970 28.405 ;
        RECT 73.700 27.890 73.960 28.035 ;
        RECT 74.160 27.550 74.420 27.870 ;
        RECT 74.220 26.250 74.360 27.550 ;
        RECT 72.840 26.110 74.360 26.250 ;
        RECT 72.320 19.390 72.580 19.710 ;
        RECT 71.400 17.350 71.660 17.670 ;
        RECT 71.860 17.350 72.120 17.670 ;
        RECT 71.460 15.290 71.600 17.350 ;
        RECT 70.480 14.970 70.740 15.290 ;
        RECT 70.940 14.970 71.200 15.290 ;
        RECT 71.400 14.970 71.660 15.290 ;
        RECT 72.380 14.610 72.520 19.390 ;
        RECT 72.840 15.970 72.980 26.110 ;
        RECT 73.240 25.510 73.500 25.830 ;
        RECT 73.300 23.110 73.440 25.510 ;
        RECT 73.700 24.830 73.960 25.150 ;
        RECT 73.240 22.790 73.500 23.110 ;
        RECT 73.760 22.770 73.900 24.830 ;
        RECT 74.680 23.110 74.820 34.010 ;
        RECT 75.070 31.435 75.350 31.805 ;
        RECT 75.080 31.280 75.340 31.435 ;
        RECT 75.080 30.270 75.340 30.590 ;
        RECT 75.140 28.210 75.280 30.270 ;
        RECT 75.080 27.890 75.340 28.210 ;
        RECT 74.620 22.790 74.880 23.110 ;
        RECT 73.700 22.450 73.960 22.770 ;
        RECT 74.680 21.070 74.820 22.790 ;
        RECT 74.620 20.750 74.880 21.070 ;
        RECT 73.690 19.875 73.970 20.245 ;
        RECT 72.780 15.650 73.040 15.970 ;
        RECT 73.760 15.630 73.900 19.875 ;
        RECT 74.680 18.010 74.820 20.750 ;
        RECT 75.140 20.050 75.280 27.890 ;
        RECT 75.600 26.170 75.740 38.770 ;
        RECT 75.990 34.155 76.270 34.525 ;
        RECT 76.060 32.290 76.200 34.155 ;
        RECT 76.450 32.795 76.730 33.165 ;
        RECT 76.000 31.970 76.260 32.290 ;
        RECT 76.045 31.520 76.305 31.610 ;
        RECT 76.520 31.520 76.660 32.795 ;
        RECT 76.980 31.805 77.120 44.550 ;
        RECT 76.045 31.380 76.660 31.520 ;
        RECT 76.910 31.435 77.190 31.805 ;
        RECT 76.045 31.290 76.305 31.380 ;
        RECT 75.990 30.755 76.270 31.125 ;
        RECT 76.000 30.610 76.260 30.755 ;
        RECT 76.520 29.230 76.660 31.380 ;
        RECT 76.460 28.910 76.720 29.230 ;
        RECT 76.460 27.550 76.720 27.870 ;
        RECT 75.990 26.675 76.270 27.045 ;
        RECT 76.060 26.170 76.200 26.675 ;
        RECT 75.540 25.850 75.800 26.170 ;
        RECT 76.000 25.850 76.260 26.170 ;
        RECT 75.600 25.490 75.740 25.850 ;
        RECT 75.540 25.170 75.800 25.490 ;
        RECT 75.990 20.555 76.270 20.925 ;
        RECT 75.080 19.730 75.340 20.050 ;
        RECT 74.620 17.690 74.880 18.010 ;
        RECT 74.150 17.155 74.430 17.525 ;
        RECT 73.700 15.310 73.960 15.630 ;
        RECT 72.780 14.970 73.040 15.290 ;
        RECT 72.320 14.290 72.580 14.610 ;
        RECT 72.840 12.910 72.980 14.970 ;
        RECT 73.760 14.270 73.900 15.310 ;
        RECT 73.240 13.950 73.500 14.270 ;
        RECT 73.700 13.950 73.960 14.270 ;
        RECT 72.780 12.590 73.040 12.910 ;
        RECT 73.300 12.230 73.440 13.950 ;
        RECT 73.760 12.230 73.900 13.950 ;
        RECT 74.220 13.250 74.360 17.155 ;
        RECT 74.680 15.290 74.820 17.690 ;
        RECT 74.620 14.970 74.880 15.290 ;
        RECT 76.060 13.250 76.200 20.555 ;
        RECT 76.520 15.630 76.660 27.550 ;
        RECT 76.980 26.850 77.120 31.435 ;
        RECT 77.440 29.085 77.580 53.050 ;
        RECT 77.900 49.630 78.040 58.635 ;
        RECT 77.840 49.310 78.100 49.630 ;
        RECT 78.360 48.270 78.500 60.870 ;
        RECT 78.820 55.070 78.960 60.870 ;
        RECT 79.740 56.430 79.880 61.210 ;
        RECT 80.140 60.530 80.400 60.850 ;
        RECT 80.200 57.790 80.340 60.530 ;
        RECT 80.140 57.470 80.400 57.790 ;
        RECT 79.680 56.110 79.940 56.430 ;
        RECT 78.760 54.750 79.020 55.070 ;
        RECT 79.220 53.730 79.480 54.050 ;
        RECT 78.750 50.475 79.030 50.845 ;
        RECT 78.300 47.950 78.560 48.270 ;
        RECT 78.820 44.870 78.960 50.475 ;
        RECT 79.280 44.870 79.420 53.730 ;
        RECT 79.740 47.590 79.880 56.110 ;
        RECT 80.660 50.310 80.800 66.310 ;
        RECT 81.120 65.125 81.260 70.050 ;
        RECT 81.050 64.755 81.330 65.125 ;
        RECT 81.060 60.190 81.320 60.510 ;
        RECT 81.120 56.770 81.260 60.190 ;
        RECT 81.060 56.450 81.320 56.770 ;
        RECT 81.050 54.555 81.330 54.925 ;
        RECT 80.600 49.990 80.860 50.310 ;
        RECT 80.600 49.310 80.860 49.630 ;
        RECT 80.660 48.270 80.800 49.310 ;
        RECT 80.600 47.950 80.860 48.270 ;
        RECT 80.140 47.610 80.400 47.930 ;
        RECT 79.680 47.270 79.940 47.590 ;
        RECT 78.760 44.550 79.020 44.870 ;
        RECT 79.220 44.550 79.480 44.870 ;
        RECT 78.820 43.170 78.960 44.550 ;
        RECT 79.680 44.210 79.940 44.530 ;
        RECT 78.760 42.850 79.020 43.170 ;
        RECT 78.760 42.170 79.020 42.490 ;
        RECT 77.840 33.330 78.100 33.650 ;
        RECT 77.900 32.290 78.040 33.330 ;
        RECT 77.840 31.970 78.100 32.290 ;
        RECT 78.290 32.115 78.570 32.485 ;
        RECT 78.300 31.970 78.560 32.115 ;
        RECT 78.820 31.610 78.960 42.170 ;
        RECT 79.740 33.310 79.880 44.210 ;
        RECT 80.200 40.450 80.340 47.610 ;
        RECT 80.660 44.530 80.800 47.950 ;
        RECT 81.120 45.890 81.260 54.555 ;
        RECT 81.580 51.330 81.720 74.955 ;
        RECT 82.040 60.850 82.180 77.190 ;
        RECT 81.980 60.530 82.240 60.850 ;
        RECT 81.520 51.010 81.780 51.330 ;
        RECT 81.060 45.570 81.320 45.890 ;
        RECT 80.600 44.210 80.860 44.530 ;
        RECT 81.050 40.955 81.330 41.325 ;
        RECT 80.140 40.130 80.400 40.450 ;
        RECT 80.200 37.050 80.340 40.130 ;
        RECT 81.120 37.730 81.260 40.955 ;
        RECT 81.520 38.430 81.780 38.750 ;
        RECT 81.060 37.410 81.320 37.730 ;
        RECT 80.140 36.730 80.400 37.050 ;
        RECT 79.680 32.990 79.940 33.310 ;
        RECT 80.200 32.290 80.340 36.730 ;
        RECT 81.060 32.990 81.320 33.310 ;
        RECT 80.140 31.970 80.400 32.290 ;
        RECT 81.120 31.610 81.260 32.990 ;
        RECT 78.760 31.290 79.020 31.610 ;
        RECT 80.140 31.290 80.400 31.610 ;
        RECT 81.060 31.290 81.320 31.610 ;
        RECT 80.200 29.570 80.340 31.290 ;
        RECT 81.120 29.765 81.260 31.290 ;
        RECT 80.140 29.250 80.400 29.570 ;
        RECT 81.050 29.395 81.330 29.765 ;
        RECT 77.370 28.715 77.650 29.085 ;
        RECT 78.290 28.715 78.570 29.085 ;
        RECT 78.360 28.550 78.500 28.715 ;
        RECT 78.300 28.230 78.560 28.550 ;
        RECT 79.220 28.230 79.480 28.550 ;
        RECT 79.680 28.230 79.940 28.550 ;
        RECT 80.600 28.230 80.860 28.550 ;
        RECT 76.920 26.530 77.180 26.850 ;
        RECT 76.980 26.170 77.120 26.530 ;
        RECT 76.920 25.850 77.180 26.170 ;
        RECT 76.980 25.150 77.120 25.850 ;
        RECT 76.920 24.830 77.180 25.150 ;
        RECT 77.380 24.830 77.640 25.150 ;
        RECT 77.440 20.730 77.580 24.830 ;
        RECT 79.280 23.790 79.420 28.230 ;
        RECT 79.220 23.470 79.480 23.790 ;
        RECT 77.840 22.110 78.100 22.430 ;
        RECT 77.380 20.410 77.640 20.730 ;
        RECT 77.900 17.670 78.040 22.110 ;
        RECT 78.290 19.875 78.570 20.245 ;
        RECT 78.360 18.690 78.500 19.875 ;
        RECT 78.300 18.370 78.560 18.690 ;
        RECT 77.840 17.350 78.100 17.670 ;
        RECT 76.460 15.310 76.720 15.630 ;
        RECT 74.160 12.930 74.420 13.250 ;
        RECT 76.000 12.930 76.260 13.250 ;
        RECT 78.360 12.230 78.500 18.370 ;
        RECT 79.280 17.330 79.420 23.470 ;
        RECT 79.220 17.010 79.480 17.330 ;
        RECT 79.740 15.970 79.880 28.230 ;
        RECT 80.660 26.170 80.800 28.230 ;
        RECT 80.600 25.850 80.860 26.170 ;
        RECT 80.660 23.110 80.800 25.850 ;
        RECT 81.050 23.955 81.330 24.325 ;
        RECT 80.140 22.790 80.400 23.110 ;
        RECT 80.600 22.790 80.860 23.110 ;
        RECT 79.680 15.650 79.940 15.970 ;
        RECT 80.200 13.250 80.340 22.790 ;
        RECT 81.120 13.250 81.260 23.955 ;
        RECT 81.580 22.770 81.720 38.430 ;
        RECT 81.520 22.450 81.780 22.770 ;
        RECT 80.140 12.930 80.400 13.250 ;
        RECT 81.060 12.930 81.320 13.250 ;
        RECT 35.520 11.910 35.780 12.230 ;
        RECT 43.800 11.910 44.060 12.230 ;
        RECT 46.100 11.910 46.360 12.230 ;
        RECT 69.100 11.910 69.360 12.230 ;
        RECT 69.560 11.910 69.820 12.230 ;
        RECT 70.020 11.910 70.280 12.230 ;
        RECT 73.240 11.910 73.500 12.230 ;
        RECT 73.700 11.910 73.960 12.230 ;
        RECT 78.300 11.910 78.560 12.230 ;
        RECT 24.370 10.695 25.910 11.065 ;
        RECT 35.580 4.000 35.720 11.910 ;
        RECT 38.740 11.570 39.000 11.890 ;
        RECT 48.400 11.570 48.660 11.890 ;
        RECT 38.800 4.000 38.940 11.570 ;
        RECT 41.960 11.230 42.220 11.550 ;
        RECT 45.180 11.230 45.440 11.550 ;
        RECT 42.020 4.000 42.160 11.230 ;
        RECT 45.240 4.000 45.380 11.230 ;
        RECT 48.460 4.000 48.600 11.570 ;
        RECT 64.500 11.230 64.760 11.550 ;
        RECT 67.720 11.230 67.980 11.550 ;
        RECT 70.940 11.230 71.200 11.550 ;
        RECT 64.560 4.000 64.700 11.230 ;
        RECT 67.780 4.000 67.920 11.230 ;
        RECT 71.000 4.000 71.140 11.230 ;
      LAYER met3 ;
        RECT 21.050 165.755 22.630 166.085 ;
        RECT 64.005 164.370 64.335 164.385 ;
        RECT 76.425 164.370 76.755 164.385 ;
        RECT 64.005 164.070 76.755 164.370 ;
        RECT 64.005 164.055 64.335 164.070 ;
        RECT 76.425 164.055 76.755 164.070 ;
        RECT 62.625 163.690 62.955 163.705 ;
        RECT 79.185 163.690 79.515 163.705 ;
        RECT 62.625 163.390 79.515 163.690 ;
        RECT 62.625 163.375 62.955 163.390 ;
        RECT 79.185 163.375 79.515 163.390 ;
        RECT 24.350 163.035 25.930 163.365 ;
        RECT 71.825 161.650 72.155 161.665 ;
        RECT 72.745 161.650 73.075 161.665 ;
        RECT 74.585 161.650 74.915 161.665 ;
        RECT 71.825 161.350 74.915 161.650 ;
        RECT 71.825 161.335 72.155 161.350 ;
        RECT 72.745 161.335 73.075 161.350 ;
        RECT 74.585 161.335 74.915 161.350 ;
        RECT 59.865 160.970 60.195 160.985 ;
        RECT 78.265 160.970 78.595 160.985 ;
        RECT 80.565 160.970 80.895 160.985 ;
        RECT 59.865 160.670 80.895 160.970 ;
        RECT 59.865 160.655 60.195 160.670 ;
        RECT 78.265 160.655 78.595 160.670 ;
        RECT 80.565 160.655 80.895 160.670 ;
        RECT 21.050 160.315 22.630 160.645 ;
        RECT 77.805 160.290 78.135 160.305 ;
        RECT 61.950 159.990 78.135 160.290 ;
        RECT 35.025 159.610 35.355 159.625 ;
        RECT 40.750 159.610 41.130 159.620 ;
        RECT 35.025 159.310 41.130 159.610 ;
        RECT 35.025 159.295 35.355 159.310 ;
        RECT 40.750 159.300 41.130 159.310 ;
        RECT 58.485 159.610 58.815 159.625 ;
        RECT 61.950 159.610 62.250 159.990 ;
        RECT 77.805 159.975 78.135 159.990 ;
        RECT 58.485 159.310 62.250 159.610 ;
        RECT 69.065 159.620 69.395 159.625 ;
        RECT 69.065 159.610 69.650 159.620 ;
        RECT 71.365 159.610 71.695 159.625 ;
        RECT 72.745 159.610 73.075 159.625 ;
        RECT 69.065 159.310 69.850 159.610 ;
        RECT 71.365 159.310 73.075 159.610 ;
        RECT 58.485 159.295 58.815 159.310 ;
        RECT 69.065 159.300 69.650 159.310 ;
        RECT 69.065 159.295 69.395 159.300 ;
        RECT 71.365 159.295 71.695 159.310 ;
        RECT 72.745 159.295 73.075 159.310 ;
        RECT 35.945 158.930 36.275 158.945 ;
        RECT 38.910 158.930 39.290 158.940 ;
        RECT 35.945 158.630 39.290 158.930 ;
        RECT 35.945 158.615 36.275 158.630 ;
        RECT 38.910 158.620 39.290 158.630 ;
        RECT 24.350 157.595 25.930 157.925 ;
        RECT 67.430 157.570 67.810 157.580 ;
        RECT 68.145 157.570 68.475 157.585 ;
        RECT 67.430 157.270 68.475 157.570 ;
        RECT 67.430 157.260 67.810 157.270 ;
        RECT 68.145 157.255 68.475 157.270 ;
        RECT 4.000 156.580 4.330 156.900 ;
        RECT 81.485 156.890 81.815 156.905 ;
        RECT 81.485 156.590 84.945 156.890 ;
        RECT 81.485 156.575 81.815 156.590 ;
        RECT 21.050 154.875 22.630 155.205 ;
        RECT 52.505 153.490 52.835 153.505 ;
        RECT 52.505 153.190 84.945 153.490 ;
        RECT 52.505 153.175 52.835 153.190 ;
        RECT 71.110 152.810 71.490 152.820 ;
        RECT 76.885 152.810 77.215 152.825 ;
        RECT 71.110 152.510 77.215 152.810 ;
        RECT 71.110 152.500 71.490 152.510 ;
        RECT 76.885 152.495 77.215 152.510 ;
        RECT 24.350 152.155 25.930 152.485 ;
        RECT 53.885 152.140 54.215 152.145 ;
        RECT 53.630 152.130 54.215 152.140 ;
        RECT 53.430 151.830 76.050 152.130 ;
        RECT 53.630 151.820 54.215 151.830 ;
        RECT 53.885 151.815 54.215 151.820 ;
        RECT 75.750 151.450 76.050 151.830 ;
        RECT 79.645 151.450 79.975 151.465 ;
        RECT 75.750 151.150 79.975 151.450 ;
        RECT 79.645 151.135 79.975 151.150 ;
        RECT 0.525 150.770 0.855 150.785 ;
        RECT 70.445 150.780 70.775 150.785 ;
        RECT 3.950 150.770 4.330 150.780 ;
        RECT 0.525 150.470 4.330 150.770 ;
        RECT 0.525 150.455 0.855 150.470 ;
        RECT 3.950 150.460 4.330 150.470 ;
        RECT 70.190 150.770 70.775 150.780 ;
        RECT 70.190 150.470 71.000 150.770 ;
        RECT 70.190 150.460 70.775 150.470 ;
        RECT 70.445 150.455 70.775 150.460 ;
        RECT 76.885 150.090 77.215 150.105 ;
        RECT 76.885 149.790 84.945 150.090 ;
        RECT 76.885 149.775 77.215 149.790 ;
        RECT 21.050 149.435 22.630 149.765 ;
        RECT 34.565 148.730 34.895 148.745 ;
        RECT 36.405 148.730 36.735 148.745 ;
        RECT 40.545 148.730 40.875 148.745 ;
        RECT 34.565 148.430 40.875 148.730 ;
        RECT 34.565 148.415 34.895 148.430 ;
        RECT 36.405 148.415 36.735 148.430 ;
        RECT 40.545 148.415 40.875 148.430 ;
        RECT 58.025 147.370 58.355 147.385 ;
        RECT 60.070 147.370 60.450 147.380 ;
        RECT 58.025 147.070 60.450 147.370 ;
        RECT 58.025 147.055 58.355 147.070 ;
        RECT 60.070 147.060 60.450 147.070 ;
        RECT 24.350 146.715 25.930 147.045 ;
        RECT 81.485 146.690 81.815 146.705 ;
        RECT 81.485 146.390 84.945 146.690 ;
        RECT 81.485 146.375 81.815 146.390 ;
        RECT 47.190 146.010 47.570 146.020 ;
        RECT 79.645 146.010 79.975 146.025 ;
        RECT 47.190 145.710 79.975 146.010 ;
        RECT 47.190 145.700 47.570 145.710 ;
        RECT 79.645 145.695 79.975 145.710 ;
        RECT 59.150 145.330 59.530 145.340 ;
        RECT 75.045 145.330 75.375 145.345 ;
        RECT 59.150 145.030 75.375 145.330 ;
        RECT 59.150 145.020 59.530 145.030 ;
        RECT 75.045 145.015 75.375 145.030 ;
        RECT 21.050 143.995 22.630 144.325 ;
        RECT 56.185 143.290 56.515 143.305 ;
        RECT 56.185 142.990 84.945 143.290 ;
        RECT 56.185 142.975 56.515 142.990 ;
        RECT 24.350 141.275 25.930 141.605 ;
        RECT 76.885 139.890 77.215 139.905 ;
        RECT 76.885 139.590 84.945 139.890 ;
        RECT 76.885 139.575 77.215 139.590 ;
        RECT 21.050 138.555 22.630 138.885 ;
        RECT 62.830 138.530 63.210 138.540 ;
        RECT 64.925 138.530 65.255 138.545 ;
        RECT 62.830 138.230 65.255 138.530 ;
        RECT 62.830 138.220 63.210 138.230 ;
        RECT 64.925 138.215 65.255 138.230 ;
        RECT 69.270 136.490 69.650 136.500 ;
        RECT 69.270 136.190 84.945 136.490 ;
        RECT 69.270 136.180 69.650 136.190 ;
        RECT 24.350 135.835 25.930 136.165 ;
        RECT 13.865 135.130 14.195 135.145 ;
        RECT 23.985 135.130 24.315 135.145 ;
        RECT 29.505 135.130 29.835 135.145 ;
        RECT 13.865 134.830 29.835 135.130 ;
        RECT 13.865 134.815 14.195 134.830 ;
        RECT 23.985 134.815 24.315 134.830 ;
        RECT 29.505 134.815 29.835 134.830 ;
        RECT 14.325 134.450 14.655 134.465 ;
        RECT 25.365 134.450 25.695 134.465 ;
        RECT 67.225 134.460 67.555 134.465 ;
        RECT 67.225 134.450 67.810 134.460 ;
        RECT 14.325 134.150 25.695 134.450 ;
        RECT 67.000 134.150 67.810 134.450 ;
        RECT 14.325 134.135 14.655 134.150 ;
        RECT 25.365 134.135 25.695 134.150 ;
        RECT 67.225 134.140 67.810 134.150 ;
        RECT 67.225 134.135 67.555 134.140 ;
        RECT 15.245 133.770 15.575 133.785 ;
        RECT 17.545 133.770 17.875 133.785 ;
        RECT 15.245 133.470 17.875 133.770 ;
        RECT 15.245 133.455 15.575 133.470 ;
        RECT 17.545 133.455 17.875 133.470 ;
        RECT 21.050 133.115 22.630 133.445 ;
        RECT 55.265 133.090 55.595 133.105 ;
        RECT 55.265 132.790 84.945 133.090 ;
        RECT 55.265 132.775 55.595 132.790 ;
        RECT 12.945 132.410 13.275 132.425 ;
        RECT 13.865 132.410 14.195 132.425 ;
        RECT 12.945 132.110 14.195 132.410 ;
        RECT 12.945 132.095 13.275 132.110 ;
        RECT 13.865 132.095 14.195 132.110 ;
        RECT 64.005 132.410 64.335 132.425 ;
        RECT 71.110 132.410 71.490 132.420 ;
        RECT 64.005 132.110 71.490 132.410 ;
        RECT 64.005 132.095 64.335 132.110 ;
        RECT 71.110 132.100 71.490 132.110 ;
        RECT 58.945 131.730 59.275 131.745 ;
        RECT 62.165 131.730 62.495 131.745 ;
        RECT 69.065 131.730 69.395 131.745 ;
        RECT 58.945 131.430 69.395 131.730 ;
        RECT 58.945 131.415 59.275 131.430 ;
        RECT 62.165 131.415 62.495 131.430 ;
        RECT 69.065 131.415 69.395 131.430 ;
        RECT 73.870 131.730 74.250 131.740 ;
        RECT 79.185 131.730 79.515 131.745 ;
        RECT 73.870 131.430 79.515 131.730 ;
        RECT 73.870 131.420 74.250 131.430 ;
        RECT 79.185 131.415 79.515 131.430 ;
        RECT 24.350 130.395 25.930 130.725 ;
        RECT 81.025 129.690 81.355 129.705 ;
        RECT 81.025 129.390 84.945 129.690 ;
        RECT 81.025 129.375 81.355 129.390 ;
        RECT 21.050 127.675 22.630 128.005 ;
        RECT 38.245 127.650 38.575 127.665 ;
        RECT 40.545 127.660 40.875 127.665 ;
        RECT 38.910 127.650 39.290 127.660 ;
        RECT 40.545 127.650 41.130 127.660 ;
        RECT 38.245 127.350 39.290 127.650 ;
        RECT 40.320 127.350 41.130 127.650 ;
        RECT 38.245 127.335 38.575 127.350 ;
        RECT 38.910 127.340 39.290 127.350 ;
        RECT 40.545 127.340 41.130 127.350 ;
        RECT 40.545 127.335 40.875 127.340 ;
        RECT 4.205 126.970 4.535 126.985 ;
        RECT 3.990 126.655 4.535 126.970 ;
        RECT 72.950 126.970 73.330 126.980 ;
        RECT 77.805 126.970 78.135 126.985 ;
        RECT 72.950 126.670 78.135 126.970 ;
        RECT 72.950 126.660 73.330 126.670 ;
        RECT 77.805 126.655 78.135 126.670 ;
        RECT 3.990 126.440 4.290 126.655 ;
        RECT 4.000 125.990 4.290 126.440 ;
        RECT 69.525 126.290 69.855 126.305 ;
        RECT 69.525 125.990 84.945 126.290 ;
        RECT 69.525 125.975 69.855 125.990 ;
        RECT 24.350 124.955 25.930 125.285 ;
        RECT 54.805 124.940 55.135 124.945 ;
        RECT 54.550 124.930 55.135 124.940 ;
        RECT 54.350 124.630 55.135 124.930 ;
        RECT 54.550 124.620 55.135 124.630 ;
        RECT 60.990 124.930 61.370 124.940 ;
        RECT 70.190 124.930 70.570 124.940 ;
        RECT 60.990 124.630 70.570 124.930 ;
        RECT 60.990 124.620 61.370 124.630 ;
        RECT 70.190 124.620 70.570 124.630 ;
        RECT 54.805 124.615 55.135 124.620 ;
        RECT 60.785 122.890 61.115 122.905 ;
        RECT 60.785 122.590 84.945 122.890 ;
        RECT 60.785 122.575 61.115 122.590 ;
        RECT 21.050 122.235 22.630 122.565 ;
        RECT 73.205 122.210 73.535 122.225 ;
        RECT 75.505 122.210 75.835 122.225 ;
        RECT 73.205 121.910 75.835 122.210 ;
        RECT 73.205 121.895 73.535 121.910 ;
        RECT 75.505 121.895 75.835 121.910 ;
        RECT 19.845 121.540 20.175 121.545 ;
        RECT 19.590 121.530 20.175 121.540 ;
        RECT 19.390 121.230 20.175 121.530 ;
        RECT 19.590 121.220 20.175 121.230 ;
        RECT 19.845 121.215 20.175 121.220 ;
        RECT 15.910 120.850 16.290 120.860 ;
        RECT 17.085 120.850 17.415 120.865 ;
        RECT 15.910 120.550 17.415 120.850 ;
        RECT 15.910 120.540 16.290 120.550 ;
        RECT 17.085 120.535 17.415 120.550 ;
        RECT 59.865 120.850 60.195 120.865 ;
        RECT 60.785 120.850 61.115 120.865 ;
        RECT 59.865 120.550 61.115 120.850 ;
        RECT 59.865 120.535 60.195 120.550 ;
        RECT 60.785 120.535 61.115 120.550 ;
        RECT 24.350 119.515 25.930 119.845 ;
        RECT 75.965 119.490 76.295 119.505 ;
        RECT 75.965 119.190 84.945 119.490 ;
        RECT 75.965 119.175 76.295 119.190 ;
        RECT 64.005 118.130 64.335 118.145 ;
        RECT 64.670 118.130 65.050 118.140 ;
        RECT 64.005 117.830 65.050 118.130 ;
        RECT 64.005 117.815 64.335 117.830 ;
        RECT 64.670 117.820 65.050 117.830 ;
        RECT 56.185 117.450 56.515 117.465 ;
        RECT 58.485 117.450 58.815 117.465 ;
        RECT 56.185 117.150 58.815 117.450 ;
        RECT 56.185 117.135 56.515 117.150 ;
        RECT 58.485 117.135 58.815 117.150 ;
        RECT 21.050 116.795 22.630 117.125 ;
        RECT 51.585 116.770 51.915 116.785 ;
        RECT 58.945 116.770 59.275 116.785 ;
        RECT 69.065 116.770 69.395 116.785 ;
        RECT 51.585 116.470 69.395 116.770 ;
        RECT 51.585 116.455 51.915 116.470 ;
        RECT 58.945 116.455 59.275 116.470 ;
        RECT 69.065 116.455 69.395 116.470 ;
        RECT 72.285 116.090 72.615 116.105 ;
        RECT 73.870 116.090 74.250 116.100 ;
        RECT 72.285 115.790 74.250 116.090 ;
        RECT 72.285 115.775 72.615 115.790 ;
        RECT 73.870 115.780 74.250 115.790 ;
        RECT 75.965 116.090 76.295 116.105 ;
        RECT 75.965 115.790 84.945 116.090 ;
        RECT 75.965 115.775 76.295 115.790 ;
        RECT 45.350 115.410 45.730 115.420 ;
        RECT 47.445 115.410 47.775 115.425 ;
        RECT 45.350 115.110 47.775 115.410 ;
        RECT 45.350 115.100 45.730 115.110 ;
        RECT 47.445 115.095 47.775 115.110 ;
        RECT 58.230 115.410 58.610 115.420 ;
        RECT 61.245 115.410 61.575 115.425 ;
        RECT 58.230 115.110 61.575 115.410 ;
        RECT 58.230 115.100 58.610 115.110 ;
        RECT 61.245 115.095 61.575 115.110 ;
        RECT 60.785 114.730 61.115 114.745 ;
        RECT 62.625 114.730 62.955 114.745 ;
        RECT 60.785 114.430 62.955 114.730 ;
        RECT 60.785 114.415 61.115 114.430 ;
        RECT 62.625 114.415 62.955 114.430 ;
        RECT 24.350 114.075 25.930 114.405 ;
        RECT 57.310 114.050 57.690 114.060 ;
        RECT 60.325 114.050 60.655 114.065 ;
        RECT 57.310 113.750 60.655 114.050 ;
        RECT 57.310 113.740 57.690 113.750 ;
        RECT 60.325 113.735 60.655 113.750 ;
        RECT 76.425 112.690 76.755 112.705 ;
        RECT 76.425 112.390 84.945 112.690 ;
        RECT 76.425 112.375 76.755 112.390 ;
        RECT 21.050 111.355 22.630 111.685 ;
        RECT 48.365 111.330 48.695 111.345 ;
        RECT 62.165 111.330 62.495 111.345 ;
        RECT 48.365 111.030 62.495 111.330 ;
        RECT 48.365 111.015 48.695 111.030 ;
        RECT 62.165 111.015 62.495 111.030 ;
        RECT 59.150 110.650 59.530 110.660 ;
        RECT 73.870 110.650 74.250 110.660 ;
        RECT 59.150 110.350 74.250 110.650 ;
        RECT 59.150 110.340 59.530 110.350 ;
        RECT 73.870 110.340 74.250 110.350 ;
        RECT 64.925 109.970 65.255 109.985 ;
        RECT 65.590 109.970 65.970 109.980 ;
        RECT 64.925 109.670 65.970 109.970 ;
        RECT 64.925 109.655 65.255 109.670 ;
        RECT 65.590 109.660 65.970 109.670 ;
        RECT 79.185 109.290 79.515 109.305 ;
        RECT 79.185 108.990 84.945 109.290 ;
        RECT 79.185 108.975 79.515 108.990 ;
        RECT 24.350 108.635 25.930 108.965 ;
        RECT 60.070 107.250 60.450 107.260 ;
        RECT 67.430 107.250 67.810 107.260 ;
        RECT 60.070 106.950 67.810 107.250 ;
        RECT 60.070 106.940 60.450 106.950 ;
        RECT 67.430 106.940 67.810 106.950 ;
        RECT 4.205 106.570 4.535 106.585 ;
        RECT 3.990 106.255 4.535 106.570 ;
        RECT 3.990 106.040 4.290 106.255 ;
        RECT 4.000 105.590 4.290 106.040 ;
        RECT 21.050 105.915 22.630 106.245 ;
        RECT 61.705 105.890 62.035 105.905 ;
        RECT 62.830 105.890 63.210 105.900 ;
        RECT 61.705 105.590 63.210 105.890 ;
        RECT 61.705 105.575 62.035 105.590 ;
        RECT 62.830 105.580 63.210 105.590 ;
        RECT 81.025 105.890 81.355 105.905 ;
        RECT 81.025 105.590 84.945 105.890 ;
        RECT 81.025 105.575 81.355 105.590 ;
        RECT 11.105 104.530 11.435 104.545 ;
        RECT 14.325 104.530 14.655 104.545 ;
        RECT 11.105 104.230 14.655 104.530 ;
        RECT 11.105 104.215 11.435 104.230 ;
        RECT 14.325 104.215 14.655 104.230 ;
        RECT 46.270 103.850 46.650 103.860 ;
        RECT 46.985 103.850 47.315 103.865 ;
        RECT 46.270 103.550 47.315 103.850 ;
        RECT 46.270 103.540 46.650 103.550 ;
        RECT 46.985 103.535 47.315 103.550 ;
        RECT 24.350 103.195 25.930 103.525 ;
        RECT 19.590 103.170 19.970 103.180 ;
        RECT 20.765 103.170 21.095 103.185 ;
        RECT 19.590 102.870 21.095 103.170 ;
        RECT 19.590 102.860 19.970 102.870 ;
        RECT 20.765 102.855 21.095 102.870 ;
        RECT 74.125 103.170 74.455 103.185 ;
        RECT 80.105 103.170 80.435 103.185 ;
        RECT 74.125 102.870 80.435 103.170 ;
        RECT 74.125 102.855 74.455 102.870 ;
        RECT 80.105 102.855 80.435 102.870 ;
        RECT 81.485 102.490 81.815 102.505 ;
        RECT 81.485 102.190 84.945 102.490 ;
        RECT 81.485 102.175 81.815 102.190 ;
        RECT 21.050 100.475 22.630 100.805 ;
        RECT 78.265 99.770 78.595 99.785 ;
        RECT 81.945 99.770 82.275 99.785 ;
        RECT 78.265 99.470 82.275 99.770 ;
        RECT 78.265 99.455 78.595 99.470 ;
        RECT 81.945 99.455 82.275 99.470 ;
        RECT 25.825 99.090 26.155 99.105 ;
        RECT 26.745 99.090 27.075 99.105 ;
        RECT 25.825 98.790 27.075 99.090 ;
        RECT 25.825 98.775 26.155 98.790 ;
        RECT 26.745 98.775 27.075 98.790 ;
        RECT 75.965 99.090 76.295 99.105 ;
        RECT 75.965 98.790 84.945 99.090 ;
        RECT 75.965 98.775 76.295 98.790 ;
        RECT 24.350 97.755 25.930 98.085 ;
        RECT 25.825 97.050 26.155 97.065 ;
        RECT 29.965 97.050 30.295 97.065 ;
        RECT 60.785 97.060 61.115 97.065 ;
        RECT 60.785 97.050 61.370 97.060 ;
        RECT 25.825 96.750 30.295 97.050 ;
        RECT 60.560 96.750 61.370 97.050 ;
        RECT 25.825 96.735 26.155 96.750 ;
        RECT 29.965 96.735 30.295 96.750 ;
        RECT 60.785 96.740 61.370 96.750 ;
        RECT 71.825 97.050 72.155 97.065 ;
        RECT 78.265 97.050 78.595 97.065 ;
        RECT 71.825 96.750 78.595 97.050 ;
        RECT 60.785 96.735 61.115 96.740 ;
        RECT 71.825 96.735 72.155 96.750 ;
        RECT 78.265 96.735 78.595 96.750 ;
        RECT 19.590 96.370 19.970 96.380 ;
        RECT 21.225 96.370 21.555 96.385 ;
        RECT 19.590 96.070 21.555 96.370 ;
        RECT 19.590 96.060 19.970 96.070 ;
        RECT 21.225 96.055 21.555 96.070 ;
        RECT 70.905 95.690 71.235 95.705 ;
        RECT 70.905 95.390 84.945 95.690 ;
        RECT 70.905 95.375 71.235 95.390 ;
        RECT 21.050 95.035 22.630 95.365 ;
        RECT 76.885 94.340 77.215 94.345 ;
        RECT 76.630 94.330 77.215 94.340 ;
        RECT 76.430 94.030 77.215 94.330 ;
        RECT 76.630 94.020 77.215 94.030 ;
        RECT 76.885 94.015 77.215 94.020 ;
        RECT 68.350 93.650 68.730 93.660 ;
        RECT 81.485 93.650 81.815 93.665 ;
        RECT 68.350 93.350 81.815 93.650 ;
        RECT 68.350 93.340 68.730 93.350 ;
        RECT 81.485 93.335 81.815 93.350 ;
        RECT 24.350 92.315 25.930 92.645 ;
        RECT 65.385 92.290 65.715 92.305 ;
        RECT 65.385 91.990 84.945 92.290 ;
        RECT 65.385 91.975 65.715 91.990 ;
        RECT 21.050 89.595 22.630 89.925 ;
        RECT 56.185 89.570 56.515 89.585 ;
        RECT 65.590 89.570 65.970 89.580 ;
        RECT 56.185 89.270 65.970 89.570 ;
        RECT 56.185 89.255 56.515 89.270 ;
        RECT 65.590 89.260 65.970 89.270 ;
        RECT 53.630 88.890 54.010 88.900 ;
        RECT 81.485 88.890 81.815 88.905 ;
        RECT 53.630 88.590 81.815 88.890 ;
        RECT 53.630 88.580 54.010 88.590 ;
        RECT 81.485 88.575 81.815 88.590 ;
        RECT 82.190 88.590 84.945 88.890 ;
        RECT 12.025 88.210 12.355 88.225 ;
        RECT 19.385 88.210 19.715 88.225 ;
        RECT 12.025 87.910 19.715 88.210 ;
        RECT 12.025 87.895 12.355 87.910 ;
        RECT 19.385 87.895 19.715 87.910 ;
        RECT 69.065 88.210 69.395 88.225 ;
        RECT 82.190 88.210 82.490 88.590 ;
        RECT 69.065 87.910 82.490 88.210 ;
        RECT 69.065 87.895 69.395 87.910 ;
        RECT 24.350 86.875 25.930 87.205 ;
        RECT 15.705 86.180 16.035 86.185 ;
        RECT 15.705 86.170 16.290 86.180 ;
        RECT 74.125 86.170 74.455 86.185 ;
        RECT 75.505 86.170 75.835 86.185 ;
        RECT 15.480 85.870 16.290 86.170 ;
        RECT 15.705 85.860 16.290 85.870 ;
        RECT 73.910 85.870 75.835 86.170 ;
        RECT 15.705 85.855 16.035 85.860 ;
        RECT 73.910 85.855 74.455 85.870 ;
        RECT 75.505 85.855 75.835 85.870 ;
        RECT 73.205 85.490 73.535 85.505 ;
        RECT 73.910 85.490 74.210 85.855 ;
        RECT 73.205 85.190 74.210 85.490 ;
        RECT 75.965 85.490 76.295 85.505 ;
        RECT 75.965 85.190 84.945 85.490 ;
        RECT 73.205 85.175 73.535 85.190 ;
        RECT 75.965 85.175 76.295 85.190 ;
        RECT 21.050 84.155 22.630 84.485 ;
        RECT 71.110 84.130 71.490 84.140 ;
        RECT 77.805 84.130 78.135 84.145 ;
        RECT 71.110 83.830 78.135 84.130 ;
        RECT 71.110 83.820 71.490 83.830 ;
        RECT 77.805 83.815 78.135 83.830 ;
        RECT 54.550 83.450 54.930 83.460 ;
        RECT 57.565 83.450 57.895 83.465 ;
        RECT 54.550 83.150 57.895 83.450 ;
        RECT 54.550 83.140 54.930 83.150 ;
        RECT 57.565 83.135 57.895 83.150 ;
        RECT 74.790 83.450 75.170 83.460 ;
        RECT 78.725 83.450 79.055 83.465 ;
        RECT 74.790 83.150 79.055 83.450 ;
        RECT 74.790 83.140 75.170 83.150 ;
        RECT 78.725 83.135 79.055 83.150 ;
        RECT 46.525 82.780 46.855 82.785 ;
        RECT 46.270 82.770 46.855 82.780 ;
        RECT 46.070 82.470 46.855 82.770 ;
        RECT 46.270 82.460 46.855 82.470 ;
        RECT 46.525 82.455 46.855 82.460 ;
        RECT 69.985 82.770 70.315 82.785 ;
        RECT 72.285 82.770 72.615 82.785 ;
        RECT 73.665 82.770 73.995 82.785 ;
        RECT 69.985 82.470 73.995 82.770 ;
        RECT 69.985 82.455 70.315 82.470 ;
        RECT 72.285 82.455 72.615 82.470 ;
        RECT 73.665 82.455 73.995 82.470 ;
        RECT 75.965 82.090 76.295 82.105 ;
        RECT 75.965 81.790 84.945 82.090 ;
        RECT 75.965 81.775 76.295 81.790 ;
        RECT 24.350 81.435 25.930 81.765 ;
        RECT 66.305 81.410 66.635 81.425 ;
        RECT 75.505 81.410 75.835 81.425 ;
        RECT 78.725 81.410 79.055 81.425 ;
        RECT 66.305 81.110 79.055 81.410 ;
        RECT 66.305 81.095 66.635 81.110 ;
        RECT 75.505 81.095 75.835 81.110 ;
        RECT 78.725 81.095 79.055 81.110 ;
        RECT 47.905 80.730 48.235 80.745 ;
        RECT 50.205 80.730 50.535 80.745 ;
        RECT 47.905 80.430 50.535 80.730 ;
        RECT 47.905 80.415 48.235 80.430 ;
        RECT 49.990 80.415 50.535 80.430 ;
        RECT 21.050 78.715 22.630 79.045 ;
        RECT 14.325 78.690 14.655 78.705 ;
        RECT 15.910 78.690 16.290 78.700 ;
        RECT 14.325 78.390 16.290 78.690 ;
        RECT 14.325 78.375 14.655 78.390 ;
        RECT 15.910 78.380 16.290 78.390 ;
        RECT 49.990 78.025 50.290 80.415 ;
        RECT 76.425 78.690 76.755 78.705 ;
        RECT 76.425 78.390 84.945 78.690 ;
        RECT 76.425 78.375 76.755 78.390 ;
        RECT 13.405 78.010 13.735 78.025 ;
        RECT 16.165 78.010 16.495 78.025 ;
        RECT 25.825 78.010 26.155 78.025 ;
        RECT 13.405 77.710 26.155 78.010 ;
        RECT 13.405 77.695 13.735 77.710 ;
        RECT 16.165 77.695 16.495 77.710 ;
        RECT 25.825 77.695 26.155 77.710 ;
        RECT 44.225 78.010 44.555 78.025 ;
        RECT 49.745 78.010 50.290 78.025 ;
        RECT 44.225 77.710 50.290 78.010 ;
        RECT 61.245 78.010 61.575 78.025 ;
        RECT 76.425 78.020 76.755 78.025 ;
        RECT 76.425 78.010 77.010 78.020 ;
        RECT 61.245 77.710 77.010 78.010 ;
        RECT 44.225 77.695 44.555 77.710 ;
        RECT 49.745 77.695 50.075 77.710 ;
        RECT 61.245 77.695 61.575 77.710 ;
        RECT 76.425 77.700 77.010 77.710 ;
        RECT 76.425 77.695 76.755 77.700 ;
        RECT 15.705 77.330 16.035 77.345 ;
        RECT 20.305 77.330 20.635 77.345 ;
        RECT 15.705 77.030 20.635 77.330 ;
        RECT 15.705 77.015 16.035 77.030 ;
        RECT 20.305 77.015 20.635 77.030 ;
        RECT 23.270 77.330 23.650 77.340 ;
        RECT 24.445 77.330 24.775 77.345 ;
        RECT 23.270 77.030 24.775 77.330 ;
        RECT 23.270 77.020 23.650 77.030 ;
        RECT 24.445 77.015 24.775 77.030 ;
        RECT 25.365 77.330 25.695 77.345 ;
        RECT 48.825 77.330 49.155 77.345 ;
        RECT 55.265 77.330 55.595 77.345 ;
        RECT 25.365 77.030 29.130 77.330 ;
        RECT 25.365 77.015 25.695 77.030 ;
        RECT 28.830 76.665 29.130 77.030 ;
        RECT 48.825 77.030 55.595 77.330 ;
        RECT 48.825 77.015 49.155 77.030 ;
        RECT 55.265 77.015 55.595 77.030 ;
        RECT 28.830 76.660 29.375 76.665 ;
        RECT 28.790 76.650 29.375 76.660 ;
        RECT 43.765 76.650 44.095 76.665 ;
        RECT 52.965 76.650 53.295 76.665 ;
        RECT 28.790 76.350 29.600 76.650 ;
        RECT 43.765 76.350 53.295 76.650 ;
        RECT 28.790 76.340 29.375 76.350 ;
        RECT 29.045 76.335 29.375 76.340 ;
        RECT 43.765 76.335 44.095 76.350 ;
        RECT 52.965 76.335 53.295 76.350 ;
        RECT 62.625 76.650 62.955 76.665 ;
        RECT 63.750 76.650 64.130 76.660 ;
        RECT 62.625 76.350 64.130 76.650 ;
        RECT 62.625 76.335 62.955 76.350 ;
        RECT 63.750 76.340 64.130 76.350 ;
        RECT 24.350 75.995 25.930 76.325 ;
        RECT 60.990 75.970 61.370 75.980 ;
        RECT 76.885 75.970 77.215 75.985 ;
        RECT 60.990 75.670 77.215 75.970 ;
        RECT 60.990 75.660 61.370 75.670 ;
        RECT 76.885 75.655 77.215 75.670 ;
        RECT 58.945 75.290 59.275 75.305 ;
        RECT 60.070 75.290 60.450 75.300 ;
        RECT 58.945 74.990 60.450 75.290 ;
        RECT 58.945 74.975 59.275 74.990 ;
        RECT 60.070 74.980 60.450 74.990 ;
        RECT 70.445 75.290 70.775 75.305 ;
        RECT 71.110 75.290 71.490 75.300 ;
        RECT 73.205 75.290 73.535 75.305 ;
        RECT 70.445 74.990 73.535 75.290 ;
        RECT 70.445 74.975 70.775 74.990 ;
        RECT 71.110 74.980 71.490 74.990 ;
        RECT 73.205 74.975 73.535 74.990 ;
        RECT 81.485 75.290 81.815 75.305 ;
        RECT 81.485 74.990 84.945 75.290 ;
        RECT 81.485 74.975 81.815 74.990 ;
        RECT 21.050 73.275 22.630 73.605 ;
        RECT 16.830 71.890 17.210 71.900 ;
        RECT 31.805 71.890 32.135 71.905 ;
        RECT 33.645 71.890 33.975 71.905 ;
        RECT 16.830 71.590 33.975 71.890 ;
        RECT 16.830 71.580 17.210 71.590 ;
        RECT 31.805 71.575 32.135 71.590 ;
        RECT 33.645 71.575 33.975 71.590 ;
        RECT 48.825 71.890 49.155 71.905 ;
        RECT 58.025 71.890 58.355 71.905 ;
        RECT 48.825 71.590 58.355 71.890 ;
        RECT 48.825 71.575 49.155 71.590 ;
        RECT 58.025 71.575 58.355 71.590 ;
        RECT 69.540 71.590 84.945 71.890 ;
        RECT 24.350 70.555 25.930 70.885 ;
        RECT 18.005 69.850 18.335 69.865 ;
        RECT 18.670 69.850 19.050 69.860 ;
        RECT 23.985 69.850 24.315 69.865 ;
        RECT 18.005 69.550 24.315 69.850 ;
        RECT 18.005 69.535 18.335 69.550 ;
        RECT 18.670 69.540 19.050 69.550 ;
        RECT 23.985 69.535 24.315 69.550 ;
        RECT 68.605 69.850 68.935 69.865 ;
        RECT 69.540 69.850 69.840 71.590 ;
        RECT 68.605 69.550 69.840 69.850 ;
        RECT 68.605 69.535 68.935 69.550 ;
        RECT 18.005 68.490 18.335 68.505 ;
        RECT 19.590 68.490 19.970 68.500 ;
        RECT 18.005 68.190 19.970 68.490 ;
        RECT 18.005 68.175 18.335 68.190 ;
        RECT 19.590 68.180 19.970 68.190 ;
        RECT 76.885 68.490 77.215 68.505 ;
        RECT 76.885 68.190 84.945 68.490 ;
        RECT 76.885 68.175 77.215 68.190 ;
        RECT 21.050 67.835 22.630 68.165 ;
        RECT 17.085 66.815 17.415 67.145 ;
        RECT 19.385 67.130 19.715 67.145 ;
        RECT 21.225 67.130 21.555 67.145 ;
        RECT 19.385 66.830 21.555 67.130 ;
        RECT 19.385 66.815 19.715 66.830 ;
        RECT 21.225 66.815 21.555 66.830 ;
        RECT 49.285 67.130 49.615 67.145 ;
        RECT 58.230 67.130 58.610 67.140 ;
        RECT 49.285 66.830 58.610 67.130 ;
        RECT 49.285 66.815 49.615 66.830 ;
        RECT 58.230 66.820 58.610 66.830 ;
        RECT 17.100 66.450 17.400 66.815 ;
        RECT 21.225 66.450 21.555 66.465 ;
        RECT 17.100 66.150 21.555 66.450 ;
        RECT 21.225 66.135 21.555 66.150 ;
        RECT 24.350 65.115 25.930 65.445 ;
        RECT 81.025 65.090 81.355 65.105 ;
        RECT 81.025 64.790 84.945 65.090 ;
        RECT 81.025 64.775 81.355 64.790 ;
        RECT 24.445 64.410 24.775 64.425 ;
        RECT 28.790 64.410 29.170 64.420 ;
        RECT 24.445 64.110 29.170 64.410 ;
        RECT 24.445 64.095 24.775 64.110 ;
        RECT 28.790 64.100 29.170 64.110 ;
        RECT 72.030 63.050 72.410 63.060 ;
        RECT 79.185 63.050 79.515 63.065 ;
        RECT 72.030 62.750 79.515 63.050 ;
        RECT 72.030 62.740 72.410 62.750 ;
        RECT 79.185 62.735 79.515 62.750 ;
        RECT 21.050 62.395 22.630 62.725 ;
        RECT 24.905 62.370 25.235 62.385 ;
        RECT 32.265 62.370 32.595 62.385 ;
        RECT 24.905 62.070 32.595 62.370 ;
        RECT 24.905 62.055 25.235 62.070 ;
        RECT 32.265 62.055 32.595 62.070 ;
        RECT 17.085 61.700 17.415 61.705 ;
        RECT 45.605 61.700 45.935 61.705 ;
        RECT 16.830 61.690 17.415 61.700 ;
        RECT 45.350 61.690 45.935 61.700 ;
        RECT 49.285 61.690 49.615 61.705 ;
        RECT 16.830 61.390 17.640 61.690 ;
        RECT 45.150 61.390 49.615 61.690 ;
        RECT 16.830 61.380 17.415 61.390 ;
        RECT 45.350 61.380 45.935 61.390 ;
        RECT 17.085 61.375 17.415 61.380 ;
        RECT 45.605 61.375 45.935 61.380 ;
        RECT 49.285 61.375 49.615 61.390 ;
        RECT 75.045 61.690 75.375 61.705 ;
        RECT 75.045 61.390 84.945 61.690 ;
        RECT 75.045 61.375 75.375 61.390 ;
        RECT 63.545 61.010 63.875 61.025 ;
        RECT 61.950 60.710 63.875 61.010 ;
        RECT 14.325 60.330 14.655 60.345 ;
        RECT 20.765 60.330 21.095 60.345 ;
        RECT 14.325 60.030 21.095 60.330 ;
        RECT 14.325 60.015 14.655 60.030 ;
        RECT 20.765 60.015 21.095 60.030 ;
        RECT 61.245 60.330 61.575 60.345 ;
        RECT 61.950 60.330 62.250 60.710 ;
        RECT 63.545 60.695 63.875 60.710 ;
        RECT 67.225 61.010 67.555 61.025 ;
        RECT 77.345 61.010 77.675 61.025 ;
        RECT 67.225 60.710 77.675 61.010 ;
        RECT 67.225 60.695 67.555 60.710 ;
        RECT 77.345 60.695 77.675 60.710 ;
        RECT 61.245 60.030 62.250 60.330 ;
        RECT 69.985 60.330 70.315 60.345 ;
        RECT 72.285 60.330 72.615 60.345 ;
        RECT 69.985 60.030 72.615 60.330 ;
        RECT 61.245 60.015 61.575 60.030 ;
        RECT 69.985 60.015 70.315 60.030 ;
        RECT 72.285 60.015 72.615 60.030 ;
        RECT 24.350 59.675 25.930 60.005 ;
        RECT 71.825 58.970 72.155 58.985 ;
        RECT 77.805 58.970 78.135 58.985 ;
        RECT 71.825 58.670 78.135 58.970 ;
        RECT 71.825 58.655 72.155 58.670 ;
        RECT 77.805 58.655 78.135 58.670 ;
        RECT 68.145 58.290 68.475 58.305 ;
        RECT 68.145 57.990 84.945 58.290 ;
        RECT 68.145 57.975 68.475 57.990 ;
        RECT 45.350 57.610 45.730 57.620 ;
        RECT 46.065 57.610 46.395 57.625 ;
        RECT 45.350 57.310 46.395 57.610 ;
        RECT 45.350 57.300 45.730 57.310 ;
        RECT 46.065 57.295 46.395 57.310 ;
        RECT 21.050 56.955 22.630 57.285 ;
        RECT 18.670 56.250 19.050 56.260 ;
        RECT 22.605 56.250 22.935 56.265 ;
        RECT 18.670 55.950 22.935 56.250 ;
        RECT 18.670 55.940 19.050 55.950 ;
        RECT 22.605 55.935 22.935 55.950 ;
        RECT 54.805 54.890 55.135 54.905 ;
        RECT 62.830 54.890 63.210 54.900 ;
        RECT 54.805 54.590 63.210 54.890 ;
        RECT 54.805 54.575 55.135 54.590 ;
        RECT 62.830 54.580 63.210 54.590 ;
        RECT 81.025 54.890 81.355 54.905 ;
        RECT 81.025 54.590 84.945 54.890 ;
        RECT 81.025 54.575 81.355 54.590 ;
        RECT 24.350 54.235 25.930 54.565 ;
        RECT 23.270 53.530 23.650 53.540 ;
        RECT 24.905 53.530 25.235 53.545 ;
        RECT 23.270 53.230 25.235 53.530 ;
        RECT 23.270 53.220 23.650 53.230 ;
        RECT 24.905 53.215 25.235 53.230 ;
        RECT 21.050 51.515 22.630 51.845 ;
        RECT 75.965 51.490 76.295 51.505 ;
        RECT 75.965 51.190 84.945 51.490 ;
        RECT 75.965 51.175 76.295 51.190 ;
        RECT 65.845 50.810 66.175 50.825 ;
        RECT 68.350 50.810 68.730 50.820 ;
        RECT 78.725 50.810 79.055 50.825 ;
        RECT 65.845 50.510 79.055 50.810 ;
        RECT 65.845 50.495 66.175 50.510 ;
        RECT 68.350 50.500 68.730 50.510 ;
        RECT 78.725 50.495 79.055 50.510 ;
        RECT 24.350 48.795 25.930 49.125 ;
        RECT 64.465 48.780 64.795 48.785 ;
        RECT 64.465 48.770 65.050 48.780 ;
        RECT 64.240 48.470 65.050 48.770 ;
        RECT 64.465 48.460 65.050 48.470 ;
        RECT 64.465 48.455 64.795 48.460 ;
        RECT 60.325 48.090 60.655 48.105 ;
        RECT 60.325 47.790 84.945 48.090 ;
        RECT 60.325 47.775 60.655 47.790 ;
        RECT 67.430 47.410 67.810 47.420 ;
        RECT 72.745 47.410 73.075 47.425 ;
        RECT 67.430 47.110 73.075 47.410 ;
        RECT 67.430 47.100 67.810 47.110 ;
        RECT 72.745 47.095 73.075 47.110 ;
        RECT 21.050 46.075 22.630 46.405 ;
        RECT 76.425 44.690 76.755 44.705 ;
        RECT 76.425 44.390 84.945 44.690 ;
        RECT 76.425 44.375 76.755 44.390 ;
        RECT 24.350 43.355 25.930 43.685 ;
        RECT 81.025 41.290 81.355 41.305 ;
        RECT 81.025 40.990 84.945 41.290 ;
        RECT 81.025 40.975 81.355 40.990 ;
        RECT 21.050 40.635 22.630 40.965 ;
        RECT 26.285 39.250 26.615 39.265 ;
        RECT 66.305 39.250 66.635 39.265 ;
        RECT 72.285 39.250 72.615 39.265 ;
        RECT 26.285 38.950 27.290 39.250 ;
        RECT 26.285 38.935 26.615 38.950 ;
        RECT 24.350 37.915 25.930 38.245 ;
        RECT 20.305 37.210 20.635 37.225 ;
        RECT 25.825 37.210 26.155 37.225 ;
        RECT 26.990 37.210 27.290 38.950 ;
        RECT 66.305 38.950 72.615 39.250 ;
        RECT 66.305 38.935 66.635 38.950 ;
        RECT 72.285 38.935 72.615 38.950 ;
        RECT 64.005 37.890 64.335 37.905 ;
        RECT 64.005 37.590 84.945 37.890 ;
        RECT 64.005 37.575 64.335 37.590 ;
        RECT 20.305 36.910 27.290 37.210 ;
        RECT 20.305 36.895 20.635 36.910 ;
        RECT 25.825 36.895 26.155 36.910 ;
        RECT 21.050 35.195 22.630 35.525 ;
        RECT 72.285 34.490 72.615 34.505 ;
        RECT 72.950 34.490 73.330 34.500 ;
        RECT 72.285 34.190 73.330 34.490 ;
        RECT 72.285 34.175 72.615 34.190 ;
        RECT 72.950 34.180 73.330 34.190 ;
        RECT 75.965 34.490 76.295 34.505 ;
        RECT 75.965 34.190 84.945 34.490 ;
        RECT 75.965 34.175 76.295 34.190 ;
        RECT 14.785 33.810 15.115 33.825 ;
        RECT 26.745 33.810 27.075 33.825 ;
        RECT 14.785 33.510 27.075 33.810 ;
        RECT 14.785 33.495 15.115 33.510 ;
        RECT 26.745 33.495 27.075 33.510 ;
        RECT 66.765 33.130 67.095 33.145 ;
        RECT 76.425 33.130 76.755 33.145 ;
        RECT 66.765 32.830 76.755 33.130 ;
        RECT 66.765 32.815 67.095 32.830 ;
        RECT 76.425 32.815 76.755 32.830 ;
        RECT 24.350 32.475 25.930 32.805 ;
        RECT 47.190 32.450 47.570 32.460 ;
        RECT 78.265 32.450 78.595 32.465 ;
        RECT 47.190 32.150 78.595 32.450 ;
        RECT 47.190 32.140 47.570 32.150 ;
        RECT 78.265 32.135 78.595 32.150 ;
        RECT 65.845 31.770 66.175 31.785 ;
        RECT 75.045 31.770 75.375 31.785 ;
        RECT 76.885 31.770 77.215 31.785 ;
        RECT 65.845 31.470 77.215 31.770 ;
        RECT 65.845 31.455 66.175 31.470 ;
        RECT 75.045 31.455 75.375 31.470 ;
        RECT 76.885 31.455 77.215 31.470 ;
        RECT 75.965 31.090 76.295 31.105 ;
        RECT 75.965 30.790 84.945 31.090 ;
        RECT 75.965 30.775 76.295 30.790 ;
        RECT 38.705 30.410 39.035 30.425 ;
        RECT 73.665 30.410 73.995 30.425 ;
        RECT 38.705 30.110 73.995 30.410 ;
        RECT 38.705 30.095 39.035 30.110 ;
        RECT 73.665 30.095 73.995 30.110 ;
        RECT 21.050 29.755 22.630 30.085 ;
        RECT 64.005 29.730 64.335 29.745 ;
        RECT 81.025 29.730 81.355 29.745 ;
        RECT 64.005 29.430 81.355 29.730 ;
        RECT 64.005 29.415 64.335 29.430 ;
        RECT 81.025 29.415 81.355 29.430 ;
        RECT 56.185 29.050 56.515 29.065 ;
        RECT 77.345 29.050 77.675 29.065 ;
        RECT 78.265 29.050 78.595 29.065 ;
        RECT 56.185 28.750 78.595 29.050 ;
        RECT 56.185 28.735 56.515 28.750 ;
        RECT 77.345 28.735 77.675 28.750 ;
        RECT 78.265 28.735 78.595 28.750 ;
        RECT 73.665 28.380 73.995 28.385 ;
        RECT 73.665 28.370 74.250 28.380 ;
        RECT 73.440 28.070 74.250 28.370 ;
        RECT 73.665 28.060 74.250 28.070 ;
        RECT 73.665 28.055 73.995 28.060 ;
        RECT 61.705 27.690 62.035 27.705 ;
        RECT 61.705 27.390 84.945 27.690 ;
        RECT 61.705 27.375 62.035 27.390 ;
        RECT 24.350 27.035 25.930 27.365 ;
        RECT 59.865 27.020 60.195 27.025 ;
        RECT 59.865 27.010 60.450 27.020 ;
        RECT 59.640 26.710 60.450 27.010 ;
        RECT 59.865 26.700 60.450 26.710 ;
        RECT 62.830 27.010 63.210 27.020 ;
        RECT 64.925 27.010 65.255 27.025 ;
        RECT 62.830 26.710 65.255 27.010 ;
        RECT 62.830 26.700 63.210 26.710 ;
        RECT 59.865 26.695 60.195 26.700 ;
        RECT 64.925 26.695 65.255 26.710 ;
        RECT 69.065 27.010 69.395 27.025 ;
        RECT 75.965 27.010 76.295 27.025 ;
        RECT 69.065 26.710 76.295 27.010 ;
        RECT 69.065 26.695 69.395 26.710 ;
        RECT 75.965 26.695 76.295 26.710 ;
        RECT 63.750 26.330 64.130 26.340 ;
        RECT 64.465 26.330 64.795 26.345 ;
        RECT 63.750 26.030 64.795 26.330 ;
        RECT 63.750 26.020 64.130 26.030 ;
        RECT 64.465 26.015 64.795 26.030 ;
        RECT 21.050 24.315 22.630 24.645 ;
        RECT 81.025 24.290 81.355 24.305 ;
        RECT 81.025 23.990 84.945 24.290 ;
        RECT 81.025 23.975 81.355 23.990 ;
        RECT 24.350 21.595 25.930 21.925 ;
        RECT 57.310 21.570 57.690 21.580 ;
        RECT 58.025 21.570 58.355 21.585 ;
        RECT 57.310 21.270 58.355 21.570 ;
        RECT 57.310 21.260 57.690 21.270 ;
        RECT 58.025 21.255 58.355 21.270 ;
        RECT 75.965 20.890 76.295 20.905 ;
        RECT 75.965 20.590 84.945 20.890 ;
        RECT 75.965 20.575 76.295 20.590 ;
        RECT 43.765 20.210 44.095 20.225 ;
        RECT 45.350 20.210 45.730 20.220 ;
        RECT 43.765 19.910 45.730 20.210 ;
        RECT 43.765 19.895 44.095 19.910 ;
        RECT 45.350 19.900 45.730 19.910 ;
        RECT 72.030 20.210 72.410 20.220 ;
        RECT 73.665 20.210 73.995 20.225 ;
        RECT 72.030 19.910 73.995 20.210 ;
        RECT 72.030 19.900 72.410 19.910 ;
        RECT 73.665 19.895 73.995 19.910 ;
        RECT 74.790 20.210 75.170 20.220 ;
        RECT 78.265 20.210 78.595 20.225 ;
        RECT 74.790 19.910 78.595 20.210 ;
        RECT 74.790 19.900 75.170 19.910 ;
        RECT 78.265 19.895 78.595 19.910 ;
        RECT 21.050 18.875 22.630 19.205 ;
        RECT 74.125 17.490 74.455 17.505 ;
        RECT 74.125 17.190 84.945 17.490 ;
        RECT 74.125 17.175 74.455 17.190 ;
        RECT 24.350 16.155 25.930 16.485 ;
        RECT 21.050 13.435 22.630 13.765 ;
        RECT 24.350 10.715 25.930 11.045 ;
      LAYER met4 ;
        RECT 40.775 159.295 41.105 159.625 ;
        RECT 69.295 159.295 69.625 159.625 ;
        RECT 38.935 158.615 39.265 158.945 ;
        RECT 3.975 156.575 4.305 156.905 ;
        RECT 3.990 150.785 4.290 156.575 ;
        RECT 3.975 150.455 4.305 150.785 ;
        RECT 38.950 127.665 39.250 158.615 ;
        RECT 40.790 127.665 41.090 159.295 ;
        RECT 67.455 157.255 67.785 157.585 ;
        RECT 53.655 151.815 53.985 152.145 ;
        RECT 47.215 145.695 47.545 146.025 ;
        RECT 38.935 127.335 39.265 127.665 ;
        RECT 40.775 127.335 41.105 127.665 ;
        RECT 19.615 121.215 19.945 121.545 ;
        RECT 15.935 120.535 16.265 120.865 ;
        RECT 15.950 86.185 16.250 120.535 ;
        RECT 19.630 103.185 19.930 121.215 ;
        RECT 45.375 115.095 45.705 115.425 ;
        RECT 19.615 102.855 19.945 103.185 ;
        RECT 19.615 96.055 19.945 96.385 ;
        RECT 15.935 85.855 16.265 86.185 ;
        RECT 15.950 78.705 16.250 85.855 ;
        RECT 15.935 78.375 16.265 78.705 ;
        RECT 15.950 76.650 16.250 78.375 ;
        RECT 15.950 76.350 17.170 76.650 ;
        RECT 16.870 71.905 17.170 76.350 ;
        RECT 16.855 71.575 17.185 71.905 ;
        RECT 16.870 61.705 17.170 71.575 ;
        RECT 18.695 69.535 19.025 69.865 ;
        RECT 16.855 61.375 17.185 61.705 ;
        RECT 18.710 56.265 19.010 69.535 ;
        RECT 19.630 68.505 19.930 96.055 ;
        RECT 23.295 77.015 23.625 77.345 ;
        RECT 19.615 68.175 19.945 68.505 ;
        RECT 18.695 55.935 19.025 56.265 ;
        RECT 23.310 53.545 23.610 77.015 ;
        RECT 28.815 76.335 29.145 76.665 ;
        RECT 28.830 64.425 29.130 76.335 ;
        RECT 28.815 64.095 29.145 64.425 ;
        RECT 45.390 61.705 45.690 115.095 ;
        RECT 46.295 103.535 46.625 103.865 ;
        RECT 46.310 82.785 46.610 103.535 ;
        RECT 46.295 82.455 46.625 82.785 ;
        RECT 45.375 61.375 45.705 61.705 ;
        RECT 45.375 57.295 45.705 57.625 ;
        RECT 23.295 53.215 23.625 53.545 ;
        RECT 45.390 20.225 45.690 57.295 ;
        RECT 47.230 32.465 47.530 145.695 ;
        RECT 53.670 88.905 53.970 151.815 ;
        RECT 60.095 147.055 60.425 147.385 ;
        RECT 59.175 145.015 59.505 145.345 ;
        RECT 54.575 124.615 54.905 124.945 ;
        RECT 53.655 88.575 53.985 88.905 ;
        RECT 54.590 83.465 54.890 124.615 ;
        RECT 58.255 115.095 58.585 115.425 ;
        RECT 57.335 113.735 57.665 114.065 ;
        RECT 54.575 83.135 54.905 83.465 ;
        RECT 47.215 32.135 47.545 32.465 ;
        RECT 57.350 21.585 57.650 113.735 ;
        RECT 58.270 67.145 58.570 115.095 ;
        RECT 59.190 110.665 59.490 145.015 ;
        RECT 59.175 110.335 59.505 110.665 ;
        RECT 60.110 107.265 60.410 147.055 ;
        RECT 62.855 138.215 63.185 138.545 ;
        RECT 61.015 124.615 61.345 124.945 ;
        RECT 60.095 106.935 60.425 107.265 ;
        RECT 61.030 100.450 61.330 124.615 ;
        RECT 62.870 105.905 63.170 138.215 ;
        RECT 67.470 134.465 67.770 157.255 ;
        RECT 69.310 136.505 69.610 159.295 ;
        RECT 71.135 152.495 71.465 152.825 ;
        RECT 70.215 150.455 70.545 150.785 ;
        RECT 69.295 136.175 69.625 136.505 ;
        RECT 67.455 134.135 67.785 134.465 ;
        RECT 70.230 124.945 70.530 150.455 ;
        RECT 71.150 132.425 71.450 152.495 ;
        RECT 71.135 132.095 71.465 132.425 ;
        RECT 73.895 131.415 74.225 131.745 ;
        RECT 72.975 126.655 73.305 126.985 ;
        RECT 70.215 124.615 70.545 124.945 ;
        RECT 64.695 117.815 65.025 118.145 ;
        RECT 62.855 105.575 63.185 105.905 ;
        RECT 60.110 100.150 61.330 100.450 ;
        RECT 60.110 75.305 60.410 100.150 ;
        RECT 61.015 96.735 61.345 97.065 ;
        RECT 61.030 75.985 61.330 96.735 ;
        RECT 63.775 76.335 64.105 76.665 ;
        RECT 61.015 75.655 61.345 75.985 ;
        RECT 60.095 74.975 60.425 75.305 ;
        RECT 58.255 66.815 58.585 67.145 ;
        RECT 60.110 27.025 60.410 74.975 ;
        RECT 62.855 54.575 63.185 54.905 ;
        RECT 62.870 27.025 63.170 54.575 ;
        RECT 60.095 26.695 60.425 27.025 ;
        RECT 62.855 26.695 63.185 27.025 ;
        RECT 63.790 26.345 64.090 76.335 ;
        RECT 64.710 48.785 65.010 117.815 ;
        RECT 65.615 109.655 65.945 109.985 ;
        RECT 65.630 89.585 65.930 109.655 ;
        RECT 67.455 106.935 67.785 107.265 ;
        RECT 65.615 89.255 65.945 89.585 ;
        RECT 64.695 48.455 65.025 48.785 ;
        RECT 67.470 47.425 67.770 106.935 ;
        RECT 68.375 93.335 68.705 93.665 ;
        RECT 68.390 50.825 68.690 93.335 ;
        RECT 71.135 83.815 71.465 84.145 ;
        RECT 71.150 75.305 71.450 83.815 ;
        RECT 71.135 74.975 71.465 75.305 ;
        RECT 72.055 62.735 72.385 63.065 ;
        RECT 68.375 50.495 68.705 50.825 ;
        RECT 67.455 47.095 67.785 47.425 ;
        RECT 63.775 26.015 64.105 26.345 ;
        RECT 57.335 21.255 57.665 21.585 ;
        RECT 72.070 20.225 72.370 62.735 ;
        RECT 72.990 34.505 73.290 126.655 ;
        RECT 73.910 116.105 74.210 131.415 ;
        RECT 73.895 115.775 74.225 116.105 ;
        RECT 73.895 110.335 74.225 110.665 ;
        RECT 72.975 34.175 73.305 34.505 ;
        RECT 73.910 28.385 74.210 110.335 ;
        RECT 76.655 94.015 76.985 94.345 ;
        RECT 74.815 83.135 75.145 83.465 ;
        RECT 73.895 28.055 74.225 28.385 ;
        RECT 74.830 20.225 75.130 83.135 ;
        RECT 76.670 78.025 76.970 94.015 ;
        RECT 76.655 77.695 76.985 78.025 ;
        RECT 45.375 19.895 45.705 20.225 ;
        RECT 72.055 19.895 72.385 20.225 ;
        RECT 74.815 19.895 75.145 20.225 ;
  END
END main
END LIBRARY

