VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 12.560 47.315 48.820 48.920 ;
      LAYER pwell ;
        RECT 12.755 46.115 14.125 46.925 ;
        RECT 14.135 46.115 19.645 46.925 ;
        RECT 21.060 46.795 22.405 47.025 ;
        RECT 20.575 46.115 22.405 46.795 ;
        RECT 22.545 46.115 25.545 47.025 ;
        RECT 25.645 46.200 26.075 46.985 ;
        RECT 29.670 46.795 30.590 47.025 ;
        RECT 27.125 46.115 30.590 46.795 ;
        RECT 31.615 46.795 32.960 47.025 ;
        RECT 36.110 46.795 37.030 47.025 ;
        RECT 31.615 46.115 33.445 46.795 ;
        RECT 33.565 46.115 37.030 46.795 ;
        RECT 37.135 46.115 38.505 46.895 ;
        RECT 38.525 46.200 38.955 46.985 ;
        RECT 39.895 46.795 41.240 47.025 ;
        RECT 39.895 46.115 41.725 46.795 ;
        RECT 41.735 46.115 43.105 46.925 ;
        RECT 43.115 46.115 44.485 46.895 ;
        RECT 44.495 46.115 45.865 46.895 ;
        RECT 45.875 46.115 47.245 46.895 ;
        RECT 47.255 46.115 48.625 46.925 ;
        RECT 12.895 45.905 13.065 46.115 ;
        RECT 14.275 45.905 14.445 46.115 ;
        RECT 17.950 45.955 18.070 46.065 ;
        RECT 19.805 45.960 19.965 46.070 ;
        RECT 20.715 45.925 20.885 46.115 ;
        RECT 25.315 45.905 25.485 46.115 ;
        RECT 25.775 45.905 25.945 46.095 ;
        RECT 26.245 45.960 26.405 46.070 ;
        RECT 27.155 45.925 27.325 46.115 ;
        RECT 30.845 45.960 31.005 46.070 ;
        RECT 33.135 45.925 33.305 46.115 ;
        RECT 33.595 45.925 33.765 46.115 ;
        RECT 37.285 46.095 37.455 46.115 ;
        RECT 34.975 45.925 35.145 46.095 ;
        RECT 34.975 45.905 35.140 45.925 ;
        RECT 35.435 45.905 35.605 46.095 ;
        RECT 37.275 45.925 37.455 46.095 ;
        RECT 37.275 45.905 37.445 45.925 ;
        RECT 39.115 45.905 39.285 46.095 ;
        RECT 41.415 45.925 41.585 46.115 ;
        RECT 41.875 45.925 42.045 46.115 ;
        RECT 42.335 45.905 42.505 46.095 ;
        RECT 44.175 45.925 44.345 46.115 ;
        RECT 45.555 45.925 45.725 46.115 ;
        RECT 46.925 45.905 47.095 46.115 ;
        RECT 48.315 45.905 48.485 46.115 ;
        RECT 12.755 45.095 14.125 45.905 ;
        RECT 14.135 45.095 17.805 45.905 ;
        RECT 18.315 45.225 25.625 45.905 ;
        RECT 25.635 45.225 32.945 45.905 ;
        RECT 18.315 44.995 19.665 45.225 ;
        RECT 21.200 45.005 22.110 45.225 ;
        RECT 29.150 45.005 30.060 45.225 ;
        RECT 31.595 44.995 32.945 45.225 ;
        RECT 33.305 45.225 35.140 45.905 ;
        RECT 35.295 45.225 37.125 45.905 ;
        RECT 33.305 44.995 34.235 45.225 ;
        RECT 35.780 44.995 37.125 45.225 ;
        RECT 37.145 44.995 38.495 45.905 ;
        RECT 38.525 45.035 38.955 45.820 ;
        RECT 39.055 44.995 42.055 45.905 ;
        RECT 42.305 45.225 45.770 45.905 ;
        RECT 44.850 44.995 45.770 45.225 ;
        RECT 45.875 45.125 47.245 45.905 ;
        RECT 47.255 45.095 48.625 45.905 ;
      LAYER nwell ;
        RECT 12.560 41.875 48.820 44.705 ;
      LAYER pwell ;
        RECT 12.755 40.675 14.125 41.485 ;
        RECT 17.650 41.355 18.560 41.575 ;
        RECT 20.095 41.355 21.445 41.585 ;
        RECT 14.135 40.675 21.445 41.355 ;
        RECT 21.590 41.355 22.510 41.585 ;
        RECT 21.590 40.675 25.055 41.355 ;
        RECT 25.645 40.760 26.075 41.545 ;
        RECT 26.095 41.355 27.025 41.585 ;
        RECT 31.745 41.355 32.675 41.585 ;
        RECT 26.095 40.675 29.995 41.355 ;
        RECT 30.840 40.675 32.675 41.355 ;
        RECT 33.005 40.675 34.355 41.585 ;
        RECT 37.890 41.355 38.800 41.575 ;
        RECT 40.335 41.355 41.685 41.585 ;
        RECT 43.245 41.355 44.175 41.585 ;
        RECT 34.375 40.675 41.685 41.355 ;
        RECT 42.340 40.675 44.175 41.355 ;
        RECT 44.495 40.675 45.865 41.455 ;
        RECT 45.875 40.675 47.245 41.455 ;
        RECT 47.255 40.675 48.625 41.485 ;
        RECT 12.895 40.465 13.065 40.675 ;
        RECT 14.275 40.485 14.445 40.675 ;
        RECT 15.655 40.465 15.825 40.655 ;
        RECT 16.390 40.465 16.560 40.655 ;
        RECT 20.255 40.465 20.425 40.655 ;
        RECT 24.855 40.485 25.025 40.675 ;
        RECT 25.310 40.515 25.430 40.625 ;
        RECT 26.510 40.485 26.680 40.675 ;
        RECT 30.840 40.655 31.005 40.675 ;
        RECT 30.375 40.625 30.545 40.655 ;
        RECT 30.370 40.515 30.545 40.625 ;
        RECT 30.375 40.465 30.545 40.515 ;
        RECT 30.835 40.485 31.005 40.655 ;
        RECT 34.055 40.465 34.225 40.675 ;
        RECT 34.515 40.465 34.685 40.675 ;
        RECT 42.340 40.655 42.505 40.675 ;
        RECT 12.755 39.655 14.125 40.465 ;
        RECT 14.135 39.785 15.965 40.465 ;
        RECT 15.975 39.785 19.875 40.465 ;
        RECT 14.135 39.555 15.480 39.785 ;
        RECT 15.975 39.555 16.905 39.785 ;
        RECT 20.115 39.655 21.485 40.465 ;
        RECT 21.580 39.785 30.685 40.465 ;
        RECT 30.790 39.785 34.255 40.465 ;
        RECT 30.790 39.555 31.710 39.785 ;
        RECT 34.375 39.655 35.745 40.465 ;
        RECT 35.900 40.435 36.070 40.655 ;
        RECT 39.115 40.465 39.285 40.655 ;
        RECT 41.870 40.515 41.990 40.625 ;
        RECT 42.335 40.485 42.505 40.655 ;
        RECT 42.795 40.465 42.965 40.655 ;
        RECT 44.635 40.485 44.805 40.675 ;
        RECT 46.485 40.510 46.645 40.620 ;
        RECT 46.925 40.485 47.095 40.675 ;
        RECT 48.315 40.465 48.485 40.675 ;
        RECT 37.560 40.435 38.505 40.465 ;
        RECT 35.755 39.755 38.505 40.435 ;
        RECT 37.560 39.555 38.505 39.755 ;
        RECT 38.525 39.595 38.955 40.380 ;
        RECT 39.055 39.555 42.505 40.465 ;
        RECT 42.735 39.555 46.185 40.465 ;
        RECT 47.255 39.655 48.625 40.465 ;
      LAYER nwell ;
        RECT 12.560 36.435 48.820 39.265 ;
      LAYER pwell ;
        RECT 12.755 35.235 14.125 36.045 ;
        RECT 14.135 35.915 15.065 36.145 ;
        RECT 21.790 35.915 22.700 36.135 ;
        RECT 24.235 35.915 25.585 36.145 ;
        RECT 14.135 35.235 18.035 35.915 ;
        RECT 18.275 35.235 25.585 35.915 ;
        RECT 25.645 35.320 26.075 36.105 ;
        RECT 29.610 35.915 30.520 36.135 ;
        RECT 32.055 35.915 33.405 36.145 ;
        RECT 26.095 35.235 33.405 35.915 ;
        RECT 33.915 35.915 35.280 36.145 ;
        RECT 33.915 35.235 37.125 35.915 ;
        RECT 38.135 35.235 41.135 36.145 ;
        RECT 41.275 35.235 42.625 36.145 ;
        RECT 43.195 35.235 46.645 36.145 ;
        RECT 47.255 35.235 48.625 36.045 ;
        RECT 12.895 35.025 13.065 35.235 ;
        RECT 14.550 35.045 14.720 35.235 ;
        RECT 18.415 35.045 18.585 35.235 ;
        RECT 21.175 35.025 21.345 35.215 ;
        RECT 21.635 35.025 21.805 35.215 ;
        RECT 24.390 35.075 24.510 35.185 ;
        RECT 24.855 35.025 25.025 35.215 ;
        RECT 26.235 35.045 26.405 35.235 ;
        RECT 33.590 35.075 33.710 35.185 ;
        RECT 36.810 35.045 36.980 35.235 ;
        RECT 37.275 35.025 37.445 35.215 ;
        RECT 37.745 35.070 37.905 35.180 ;
        RECT 38.195 35.045 38.365 35.235 ;
        RECT 41.420 35.215 41.590 35.235 ;
        RECT 12.755 34.215 14.125 35.025 ;
        RECT 14.175 34.345 21.485 35.025 ;
        RECT 14.175 34.115 15.525 34.345 ;
        RECT 17.060 34.125 17.970 34.345 ;
        RECT 21.495 34.215 24.245 35.025 ;
        RECT 24.715 34.345 33.820 35.025 ;
        RECT 34.010 34.345 37.475 35.025 ;
        RECT 39.110 34.995 39.280 35.215 ;
        RECT 41.415 35.045 41.590 35.215 ;
        RECT 42.790 35.075 42.910 35.185 ;
        RECT 43.255 35.045 43.425 35.235 ;
        RECT 44.170 35.075 44.290 35.185 ;
        RECT 41.415 35.025 41.585 35.045 ;
        RECT 45.550 35.025 45.720 35.215 ;
        RECT 46.935 35.185 47.105 35.215 ;
        RECT 46.930 35.075 47.105 35.185 ;
        RECT 46.935 35.025 47.105 35.075 ;
        RECT 48.315 35.025 48.485 35.235 ;
        RECT 40.310 34.995 41.265 35.025 ;
        RECT 34.010 34.115 34.930 34.345 ;
        RECT 38.525 34.155 38.955 34.940 ;
        RECT 38.985 34.315 41.265 34.995 ;
        RECT 40.310 34.115 41.265 34.315 ;
        RECT 41.275 34.215 44.025 35.025 ;
        RECT 44.515 34.115 45.865 35.025 ;
        RECT 45.875 34.245 47.245 35.025 ;
        RECT 47.255 34.215 48.625 35.025 ;
      LAYER nwell ;
        RECT 12.560 30.995 48.820 33.825 ;
      LAYER pwell ;
        RECT 12.755 29.795 14.125 30.605 ;
        RECT 14.135 29.795 15.505 30.605 ;
        RECT 18.170 30.475 19.090 30.705 ;
        RECT 15.625 29.795 19.090 30.475 ;
        RECT 19.290 30.475 20.210 30.705 ;
        RECT 19.290 29.795 22.755 30.475 ;
        RECT 22.875 29.795 25.625 30.605 ;
        RECT 25.645 29.880 26.075 30.665 ;
        RECT 26.115 29.795 27.465 30.705 ;
        RECT 27.545 29.795 31.605 30.705 ;
        RECT 31.710 30.475 32.630 30.705 ;
        RECT 31.710 29.795 35.175 30.475 ;
        RECT 35.295 29.795 36.665 30.605 ;
        RECT 36.675 30.505 37.625 30.705 ;
        RECT 36.675 29.825 40.345 30.505 ;
        RECT 36.675 29.795 37.625 29.825 ;
        RECT 12.895 29.585 13.065 29.795 ;
        RECT 14.275 29.605 14.445 29.795 ;
        RECT 15.655 29.585 15.825 29.795 ;
        RECT 16.110 29.635 16.230 29.745 ;
        RECT 16.850 29.585 17.020 29.775 ;
        RECT 20.715 29.585 20.885 29.775 ;
        RECT 22.555 29.605 22.725 29.795 ;
        RECT 23.015 29.605 23.185 29.795 ;
        RECT 27.150 29.605 27.320 29.795 ;
        RECT 28.350 29.585 28.520 29.775 ;
        RECT 31.295 29.605 31.465 29.795 ;
        RECT 34.975 29.605 35.145 29.795 ;
        RECT 35.435 29.585 35.605 29.795 ;
        RECT 35.895 29.585 36.065 29.775 ;
        RECT 40.030 29.605 40.200 29.825 ;
        RECT 40.355 29.795 41.705 30.705 ;
        RECT 41.735 29.795 43.105 30.575 ;
        RECT 43.255 29.795 46.705 30.705 ;
        RECT 47.255 29.795 48.625 30.605 ;
        RECT 40.500 29.605 40.670 29.795 ;
        RECT 41.885 29.775 42.055 29.795 ;
        RECT 41.870 29.605 42.055 29.775 ;
        RECT 42.345 29.630 42.505 29.740 ;
        RECT 41.870 29.585 42.040 29.605 ;
        RECT 46.475 29.585 46.645 29.795 ;
        RECT 46.930 29.635 47.050 29.745 ;
        RECT 48.315 29.585 48.485 29.795 ;
        RECT 12.755 28.775 14.125 29.585 ;
        RECT 14.135 28.905 15.965 29.585 ;
        RECT 16.435 28.905 20.335 29.585 ;
        RECT 20.575 28.905 27.885 29.585 ;
        RECT 14.135 28.675 15.480 28.905 ;
        RECT 16.435 28.675 17.365 28.905 ;
        RECT 24.090 28.685 25.000 28.905 ;
        RECT 26.535 28.675 27.885 28.905 ;
        RECT 27.935 28.905 31.835 29.585 ;
        RECT 32.170 28.905 35.635 29.585 ;
        RECT 27.935 28.675 28.865 28.905 ;
        RECT 32.170 28.675 33.090 28.905 ;
        RECT 35.755 28.775 38.505 29.585 ;
        RECT 38.525 28.715 38.955 29.500 ;
        RECT 39.265 28.675 42.185 29.585 ;
        RECT 43.255 28.675 46.705 29.585 ;
        RECT 47.255 28.775 48.625 29.585 ;
      LAYER nwell ;
        RECT 12.560 25.555 48.820 28.385 ;
      LAYER pwell ;
        RECT 12.755 24.355 14.125 25.165 ;
        RECT 17.650 25.035 18.560 25.255 ;
        RECT 20.095 25.035 21.445 25.265 ;
        RECT 14.135 24.355 21.445 25.035 ;
        RECT 21.495 24.355 25.165 25.165 ;
        RECT 25.645 24.440 26.075 25.225 ;
        RECT 29.610 25.035 30.520 25.255 ;
        RECT 32.055 25.035 33.405 25.265 ;
        RECT 35.300 25.035 36.665 25.265 ;
        RECT 26.095 24.355 33.405 25.035 ;
        RECT 33.455 24.355 36.665 25.035 ;
        RECT 36.675 24.355 39.425 25.165 ;
        RECT 42.550 25.035 43.470 25.265 ;
        RECT 40.005 24.355 43.470 25.035 ;
        RECT 43.655 24.355 46.655 25.265 ;
        RECT 47.255 24.355 48.625 25.165 ;
        RECT 12.895 24.145 13.065 24.355 ;
        RECT 14.275 24.165 14.445 24.355 ;
        RECT 15.655 24.145 15.825 24.335 ;
        RECT 16.125 24.190 16.285 24.300 ;
        RECT 17.035 24.145 17.205 24.335 ;
        RECT 20.725 24.190 20.885 24.300 ;
        RECT 21.635 24.145 21.805 24.355 ;
        RECT 25.310 24.195 25.430 24.305 ;
        RECT 26.235 24.165 26.405 24.355 ;
        RECT 28.720 24.145 28.890 24.335 ;
        RECT 29.455 24.145 29.625 24.335 ;
        RECT 31.295 24.145 31.465 24.335 ;
        RECT 33.600 24.165 33.770 24.355 ;
        RECT 36.815 24.165 36.985 24.355 ;
        RECT 39.390 24.145 39.560 24.335 ;
        RECT 39.570 24.195 39.690 24.305 ;
        RECT 40.035 24.165 40.205 24.355 ;
        RECT 43.255 24.145 43.425 24.335 ;
        RECT 43.715 24.165 43.885 24.355 ;
        RECT 12.755 23.335 14.125 24.145 ;
        RECT 14.135 23.465 15.965 24.145 ;
        RECT 17.005 23.465 20.470 24.145 ;
        RECT 21.605 23.465 25.070 24.145 ;
        RECT 25.405 23.465 29.305 24.145 ;
        RECT 14.135 23.235 15.480 23.465 ;
        RECT 19.550 23.235 20.470 23.465 ;
        RECT 24.150 23.235 25.070 23.465 ;
        RECT 28.375 23.235 29.305 23.465 ;
        RECT 29.315 23.335 31.145 24.145 ;
        RECT 31.155 23.465 38.465 24.145 ;
        RECT 34.670 23.245 35.580 23.465 ;
        RECT 37.115 23.235 38.465 23.465 ;
        RECT 38.525 23.275 38.955 24.060 ;
        RECT 38.975 23.465 42.875 24.145 ;
        RECT 38.975 23.235 39.905 23.465 ;
        RECT 43.115 23.365 44.485 24.145 ;
        RECT 44.495 24.115 45.440 24.145 ;
        RECT 46.930 24.115 47.100 24.335 ;
        RECT 48.315 24.145 48.485 24.355 ;
        RECT 44.495 23.435 47.245 24.115 ;
        RECT 44.495 23.235 45.440 23.435 ;
        RECT 47.255 23.335 48.625 24.145 ;
      LAYER nwell ;
        RECT 12.560 20.115 48.820 22.945 ;
      LAYER pwell ;
        RECT 12.755 18.915 14.125 19.725 ;
        RECT 14.175 19.595 15.525 19.825 ;
        RECT 17.060 19.595 17.970 19.815 ;
        RECT 14.175 18.915 21.485 19.595 ;
        RECT 21.495 18.915 25.165 19.725 ;
        RECT 25.645 19.000 26.075 19.785 ;
        RECT 26.095 18.915 35.200 19.595 ;
        RECT 35.295 18.915 36.665 19.725 ;
        RECT 36.675 18.915 38.045 19.695 ;
        RECT 38.055 18.915 39.425 19.695 ;
        RECT 39.435 18.915 40.805 19.695 ;
        RECT 40.815 18.915 42.185 19.695 ;
        RECT 42.215 18.915 43.565 19.825 ;
        RECT 43.655 18.915 47.105 19.825 ;
        RECT 47.255 18.915 48.625 19.725 ;
        RECT 12.895 18.705 13.065 18.915 ;
        RECT 15.655 18.705 15.825 18.895 ;
        RECT 16.125 18.750 16.285 18.860 ;
        RECT 17.310 18.705 17.480 18.895 ;
        RECT 21.175 18.705 21.345 18.915 ;
        RECT 21.635 18.725 21.805 18.915 ;
        RECT 24.855 18.705 25.025 18.895 ;
        RECT 25.310 18.755 25.430 18.865 ;
        RECT 26.235 18.725 26.405 18.915 ;
        RECT 33.135 18.705 33.305 18.895 ;
        RECT 33.870 18.705 34.040 18.895 ;
        RECT 35.435 18.725 35.605 18.915 ;
        RECT 36.815 18.725 36.985 18.915 ;
        RECT 37.745 18.750 37.905 18.860 ;
        RECT 38.195 18.725 38.365 18.915 ;
        RECT 39.575 18.725 39.745 18.915 ;
        RECT 40.955 18.725 41.125 18.915 ;
        RECT 42.335 18.705 42.505 18.895 ;
        RECT 42.805 18.750 42.965 18.860 ;
        RECT 43.250 18.725 43.420 18.915 ;
        RECT 43.715 18.725 43.885 18.915 ;
        RECT 46.015 18.705 46.185 18.895 ;
        RECT 46.485 18.750 46.645 18.860 ;
        RECT 48.315 18.705 48.485 18.915 ;
        RECT 12.755 17.895 14.125 18.705 ;
        RECT 14.135 18.025 15.965 18.705 ;
        RECT 16.895 18.025 20.795 18.705 ;
        RECT 14.135 17.795 15.480 18.025 ;
        RECT 16.895 17.795 17.825 18.025 ;
        RECT 21.035 17.895 24.705 18.705 ;
        RECT 24.715 17.895 26.085 18.705 ;
        RECT 26.135 18.025 33.445 18.705 ;
        RECT 33.455 18.025 37.355 18.705 ;
        RECT 26.135 17.795 27.485 18.025 ;
        RECT 29.020 17.805 29.930 18.025 ;
        RECT 33.455 17.795 34.385 18.025 ;
        RECT 38.525 17.835 38.955 18.620 ;
        RECT 39.070 18.025 42.535 18.705 ;
        RECT 39.070 17.795 39.990 18.025 ;
        RECT 43.575 17.795 46.325 18.705 ;
        RECT 47.255 17.895 48.625 18.705 ;
      LAYER nwell ;
        RECT 12.560 14.675 48.820 17.505 ;
      LAYER pwell ;
        RECT 12.755 13.475 14.125 14.285 ;
        RECT 14.135 13.475 19.645 14.285 ;
        RECT 19.655 13.475 23.325 14.285 ;
        RECT 24.280 14.155 25.625 14.385 ;
        RECT 23.795 13.475 25.625 14.155 ;
        RECT 25.645 13.560 26.075 14.345 ;
        RECT 26.555 14.155 27.900 14.385 ;
        RECT 31.910 14.155 32.820 14.375 ;
        RECT 34.355 14.155 35.705 14.385 ;
        RECT 26.555 13.475 28.385 14.155 ;
        RECT 28.395 13.475 35.705 14.155 ;
        RECT 35.755 14.155 37.100 14.385 ;
        RECT 35.755 13.475 37.585 14.155 ;
        RECT 38.525 13.560 38.955 14.345 ;
        RECT 40.380 14.155 41.725 14.385 ;
        RECT 39.895 13.475 41.725 14.155 ;
        RECT 41.735 13.475 43.105 14.255 ;
        RECT 45.855 14.155 46.785 14.385 ;
        RECT 44.035 13.475 46.785 14.155 ;
        RECT 47.255 13.475 48.625 14.285 ;
        RECT 12.895 13.285 13.065 13.475 ;
        RECT 14.275 13.285 14.445 13.475 ;
        RECT 19.795 13.285 19.965 13.475 ;
        RECT 23.470 13.315 23.590 13.425 ;
        RECT 23.935 13.285 24.105 13.475 ;
        RECT 26.230 13.315 26.350 13.425 ;
        RECT 28.075 13.285 28.245 13.475 ;
        RECT 28.535 13.285 28.705 13.475 ;
        RECT 37.275 13.285 37.445 13.475 ;
        RECT 37.745 13.320 37.905 13.430 ;
        RECT 39.125 13.320 39.285 13.430 ;
        RECT 40.035 13.285 40.205 13.475 ;
        RECT 42.785 13.285 42.955 13.475 ;
        RECT 43.265 13.320 43.425 13.430 ;
        RECT 44.175 13.285 44.345 13.475 ;
        RECT 46.930 13.315 47.050 13.425 ;
        RECT 48.315 13.285 48.485 13.475 ;
      LAYER li1 ;
        RECT 12.750 48.645 48.630 48.815 ;
        RECT 12.835 47.555 14.045 48.645 ;
        RECT 14.215 48.210 19.560 48.645 ;
        RECT 12.835 46.845 13.355 47.385 ;
        RECT 13.525 47.015 14.045 47.555 ;
        RECT 12.835 46.095 14.045 46.845 ;
        RECT 15.800 46.640 16.140 47.470 ;
        RECT 17.620 46.960 17.970 48.210 ;
        RECT 20.745 47.715 20.915 48.475 ;
        RECT 21.130 47.885 21.460 48.645 ;
        RECT 20.745 47.545 21.460 47.715 ;
        RECT 21.630 47.570 21.885 48.475 ;
        RECT 20.655 46.995 21.010 47.365 ;
        RECT 21.290 47.335 21.460 47.545 ;
        RECT 21.290 47.005 21.545 47.335 ;
        RECT 21.290 46.815 21.460 47.005 ;
        RECT 21.715 46.840 21.885 47.570 ;
        RECT 22.060 47.495 22.320 48.645 ;
        RECT 22.505 47.845 22.835 48.645 ;
        RECT 23.015 48.305 24.445 48.475 ;
        RECT 23.015 47.675 23.265 48.305 ;
        RECT 22.495 47.505 23.265 47.675 ;
        RECT 20.745 46.645 21.460 46.815 ;
        RECT 14.215 46.095 19.560 46.640 ;
        RECT 20.745 46.265 20.915 46.645 ;
        RECT 21.130 46.095 21.460 46.475 ;
        RECT 21.630 46.265 21.885 46.840 ;
        RECT 22.060 46.095 22.320 46.935 ;
        RECT 22.495 46.835 22.665 47.505 ;
        RECT 22.835 47.005 23.240 47.335 ;
        RECT 23.455 47.005 23.705 48.135 ;
        RECT 23.905 47.335 24.105 48.135 ;
        RECT 24.275 47.625 24.445 48.305 ;
        RECT 24.615 47.795 24.930 48.645 ;
        RECT 25.105 47.845 25.545 48.475 ;
        RECT 24.275 47.455 25.065 47.625 ;
        RECT 23.905 47.005 24.150 47.335 ;
        RECT 24.335 47.005 24.725 47.285 ;
        RECT 24.895 47.005 25.065 47.455 ;
        RECT 25.235 46.835 25.545 47.845 ;
        RECT 25.715 47.480 26.005 48.645 ;
        RECT 27.210 48.015 27.495 48.475 ;
        RECT 27.665 48.185 27.935 48.645 ;
        RECT 27.210 47.795 28.165 48.015 ;
        RECT 27.095 47.065 27.785 47.625 ;
        RECT 27.955 46.895 28.165 47.795 ;
        RECT 22.495 46.265 22.985 46.835 ;
        RECT 23.155 46.665 24.315 46.835 ;
        RECT 23.155 46.265 23.385 46.665 ;
        RECT 23.555 46.095 23.975 46.495 ;
        RECT 24.145 46.265 24.315 46.665 ;
        RECT 24.485 46.095 24.935 46.835 ;
        RECT 25.105 46.275 25.545 46.835 ;
        RECT 25.715 46.095 26.005 46.820 ;
        RECT 27.210 46.725 28.165 46.895 ;
        RECT 28.335 47.625 28.735 48.475 ;
        RECT 28.925 48.015 29.205 48.475 ;
        RECT 29.725 48.185 30.050 48.645 ;
        RECT 28.925 47.795 30.050 48.015 ;
        RECT 28.335 47.065 29.430 47.625 ;
        RECT 29.600 47.335 30.050 47.795 ;
        RECT 30.220 47.505 30.605 48.475 ;
        RECT 27.210 46.265 27.495 46.725 ;
        RECT 27.665 46.095 27.935 46.555 ;
        RECT 28.335 46.265 28.735 47.065 ;
        RECT 29.600 47.005 30.155 47.335 ;
        RECT 29.600 46.895 30.050 47.005 ;
        RECT 28.925 46.725 30.050 46.895 ;
        RECT 30.325 46.835 30.605 47.505 ;
        RECT 31.700 47.495 31.960 48.645 ;
        RECT 32.135 47.570 32.390 48.475 ;
        RECT 32.560 47.885 32.890 48.645 ;
        RECT 33.105 47.715 33.275 48.475 ;
        RECT 33.650 48.015 33.935 48.475 ;
        RECT 34.105 48.185 34.375 48.645 ;
        RECT 33.650 47.795 34.605 48.015 ;
        RECT 28.925 46.265 29.205 46.725 ;
        RECT 29.725 46.095 30.050 46.555 ;
        RECT 30.220 46.265 30.605 46.835 ;
        RECT 31.700 46.095 31.960 46.935 ;
        RECT 32.135 46.840 32.305 47.570 ;
        RECT 32.560 47.545 33.275 47.715 ;
        RECT 32.560 47.335 32.730 47.545 ;
        RECT 32.475 47.005 32.730 47.335 ;
        RECT 32.135 46.265 32.390 46.840 ;
        RECT 32.560 46.815 32.730 47.005 ;
        RECT 33.010 46.995 33.365 47.365 ;
        RECT 33.535 47.065 34.225 47.625 ;
        RECT 34.395 46.895 34.605 47.795 ;
        RECT 32.560 46.645 33.275 46.815 ;
        RECT 32.560 46.095 32.890 46.475 ;
        RECT 33.105 46.265 33.275 46.645 ;
        RECT 33.650 46.725 34.605 46.895 ;
        RECT 34.775 47.625 35.175 48.475 ;
        RECT 35.365 48.015 35.645 48.475 ;
        RECT 36.165 48.185 36.490 48.645 ;
        RECT 35.365 47.795 36.490 48.015 ;
        RECT 34.775 47.065 35.870 47.625 ;
        RECT 36.040 47.335 36.490 47.795 ;
        RECT 36.660 47.505 37.045 48.475 ;
        RECT 37.295 47.715 37.475 48.475 ;
        RECT 37.655 47.885 37.985 48.645 ;
        RECT 37.295 47.545 37.970 47.715 ;
        RECT 38.155 47.570 38.425 48.475 ;
        RECT 33.650 46.265 33.935 46.725 ;
        RECT 34.105 46.095 34.375 46.555 ;
        RECT 34.775 46.265 35.175 47.065 ;
        RECT 36.040 47.005 36.595 47.335 ;
        RECT 36.040 46.895 36.490 47.005 ;
        RECT 35.365 46.725 36.490 46.895 ;
        RECT 36.765 46.835 37.045 47.505 ;
        RECT 37.800 47.400 37.970 47.545 ;
        RECT 37.235 46.995 37.575 47.365 ;
        RECT 37.800 47.070 38.075 47.400 ;
        RECT 35.365 46.265 35.645 46.725 ;
        RECT 36.165 46.095 36.490 46.555 ;
        RECT 36.660 46.265 37.045 46.835 ;
        RECT 37.800 46.815 37.970 47.070 ;
        RECT 37.305 46.645 37.970 46.815 ;
        RECT 38.245 46.770 38.425 47.570 ;
        RECT 38.595 47.480 38.885 48.645 ;
        RECT 39.980 47.495 40.240 48.645 ;
        RECT 40.415 47.570 40.670 48.475 ;
        RECT 40.840 47.885 41.170 48.645 ;
        RECT 41.385 47.715 41.555 48.475 ;
        RECT 37.305 46.265 37.475 46.645 ;
        RECT 37.655 46.095 37.985 46.475 ;
        RECT 38.165 46.265 38.425 46.770 ;
        RECT 38.595 46.095 38.885 46.820 ;
        RECT 39.980 46.095 40.240 46.935 ;
        RECT 40.415 46.840 40.585 47.570 ;
        RECT 40.840 47.545 41.555 47.715 ;
        RECT 41.815 47.555 43.025 48.645 ;
        RECT 40.840 47.335 41.010 47.545 ;
        RECT 40.755 47.005 41.010 47.335 ;
        RECT 40.415 46.265 40.670 46.840 ;
        RECT 40.840 46.815 41.010 47.005 ;
        RECT 41.290 46.995 41.645 47.365 ;
        RECT 41.815 46.845 42.335 47.385 ;
        RECT 42.505 47.015 43.025 47.555 ;
        RECT 43.195 47.570 43.465 48.475 ;
        RECT 43.635 47.885 43.965 48.645 ;
        RECT 44.145 47.715 44.315 48.475 ;
        RECT 40.840 46.645 41.555 46.815 ;
        RECT 40.840 46.095 41.170 46.475 ;
        RECT 41.385 46.265 41.555 46.645 ;
        RECT 41.815 46.095 43.025 46.845 ;
        RECT 43.195 46.770 43.365 47.570 ;
        RECT 43.650 47.545 44.315 47.715 ;
        RECT 44.575 47.570 44.845 48.475 ;
        RECT 45.015 47.885 45.345 48.645 ;
        RECT 45.525 47.715 45.695 48.475 ;
        RECT 43.650 47.400 43.820 47.545 ;
        RECT 43.535 47.070 43.820 47.400 ;
        RECT 43.650 46.815 43.820 47.070 ;
        RECT 44.055 46.995 44.385 47.365 ;
        RECT 43.195 46.265 43.455 46.770 ;
        RECT 43.650 46.645 44.315 46.815 ;
        RECT 43.635 46.095 43.965 46.475 ;
        RECT 44.145 46.265 44.315 46.645 ;
        RECT 44.575 46.770 44.745 47.570 ;
        RECT 45.030 47.545 45.695 47.715 ;
        RECT 45.955 47.570 46.225 48.475 ;
        RECT 46.395 47.885 46.725 48.645 ;
        RECT 46.905 47.715 47.085 48.475 ;
        RECT 45.030 47.400 45.200 47.545 ;
        RECT 44.915 47.070 45.200 47.400 ;
        RECT 45.030 46.815 45.200 47.070 ;
        RECT 45.435 46.995 45.765 47.365 ;
        RECT 44.575 46.265 44.835 46.770 ;
        RECT 45.030 46.645 45.695 46.815 ;
        RECT 45.015 46.095 45.345 46.475 ;
        RECT 45.525 46.265 45.695 46.645 ;
        RECT 45.955 46.770 46.135 47.570 ;
        RECT 46.410 47.545 47.085 47.715 ;
        RECT 47.335 47.555 48.545 48.645 ;
        RECT 46.410 47.400 46.580 47.545 ;
        RECT 46.305 47.070 46.580 47.400 ;
        RECT 46.410 46.815 46.580 47.070 ;
        RECT 46.805 46.995 47.145 47.365 ;
        RECT 47.335 47.015 47.855 47.555 ;
        RECT 48.025 46.845 48.545 47.385 ;
        RECT 45.955 46.265 46.215 46.770 ;
        RECT 46.410 46.645 47.075 46.815 ;
        RECT 46.395 46.095 46.725 46.475 ;
        RECT 46.905 46.265 47.075 46.645 ;
        RECT 47.335 46.095 48.545 46.845 ;
        RECT 12.750 45.925 48.630 46.095 ;
        RECT 12.835 45.175 14.045 45.925 ;
        RECT 12.835 44.635 13.355 45.175 ;
        RECT 14.215 45.155 17.725 45.925 ;
        RECT 18.405 45.270 18.735 45.705 ;
        RECT 18.905 45.315 19.075 45.925 ;
        RECT 18.355 45.185 18.735 45.270 ;
        RECT 19.245 45.185 19.575 45.710 ;
        RECT 19.835 45.395 20.045 45.925 ;
        RECT 20.320 45.475 21.105 45.645 ;
        RECT 21.275 45.475 21.680 45.645 ;
        RECT 13.525 44.465 14.045 45.005 ;
        RECT 14.215 44.635 15.865 45.155 ;
        RECT 18.355 45.145 18.580 45.185 ;
        RECT 16.035 44.465 17.725 44.985 ;
        RECT 12.835 43.375 14.045 44.465 ;
        RECT 14.215 43.375 17.725 44.465 ;
        RECT 18.355 44.565 18.525 45.145 ;
        RECT 19.245 45.015 19.445 45.185 ;
        RECT 20.320 45.015 20.490 45.475 ;
        RECT 18.695 44.685 19.445 45.015 ;
        RECT 19.615 44.685 20.490 45.015 ;
        RECT 18.355 44.515 18.570 44.565 ;
        RECT 18.355 44.435 18.745 44.515 ;
        RECT 18.415 43.590 18.745 44.435 ;
        RECT 19.255 44.480 19.445 44.685 ;
        RECT 18.915 43.375 19.085 44.385 ;
        RECT 19.255 44.105 20.150 44.480 ;
        RECT 19.255 43.545 19.595 44.105 ;
        RECT 19.825 43.375 20.140 43.875 ;
        RECT 20.320 43.845 20.490 44.685 ;
        RECT 20.660 44.975 21.125 45.305 ;
        RECT 21.510 45.245 21.680 45.475 ;
        RECT 21.860 45.425 22.230 45.925 ;
        RECT 22.550 45.475 23.225 45.645 ;
        RECT 23.420 45.475 23.755 45.645 ;
        RECT 20.660 44.015 20.980 44.975 ;
        RECT 21.510 44.945 22.340 45.245 ;
        RECT 21.150 44.045 21.340 44.765 ;
        RECT 21.510 43.875 21.680 44.945 ;
        RECT 22.140 44.915 22.340 44.945 ;
        RECT 21.850 44.695 22.020 44.765 ;
        RECT 22.550 44.695 22.720 45.475 ;
        RECT 23.585 45.335 23.755 45.475 ;
        RECT 23.925 45.465 24.175 45.925 ;
        RECT 21.850 44.525 22.720 44.695 ;
        RECT 22.890 45.055 23.415 45.275 ;
        RECT 23.585 45.205 23.810 45.335 ;
        RECT 21.850 44.435 22.360 44.525 ;
        RECT 20.320 43.675 21.205 43.845 ;
        RECT 21.430 43.545 21.680 43.875 ;
        RECT 21.850 43.375 22.020 44.175 ;
        RECT 22.190 43.820 22.360 44.435 ;
        RECT 22.890 44.355 23.060 45.055 ;
        RECT 22.530 43.990 23.060 44.355 ;
        RECT 23.230 44.290 23.470 44.885 ;
        RECT 23.640 44.100 23.810 45.205 ;
        RECT 23.980 44.345 24.260 45.295 ;
        RECT 23.505 43.970 23.810 44.100 ;
        RECT 22.190 43.650 23.295 43.820 ;
        RECT 23.505 43.545 23.755 43.970 ;
        RECT 23.925 43.375 24.190 43.835 ;
        RECT 24.430 43.545 24.615 45.665 ;
        RECT 24.785 45.545 25.115 45.925 ;
        RECT 25.285 45.375 25.455 45.665 ;
        RECT 24.790 45.205 25.455 45.375 ;
        RECT 25.805 45.375 25.975 45.665 ;
        RECT 26.145 45.545 26.475 45.925 ;
        RECT 25.805 45.205 26.470 45.375 ;
        RECT 24.790 44.215 25.020 45.205 ;
        RECT 25.190 44.385 25.540 45.035 ;
        RECT 25.720 44.385 26.070 45.035 ;
        RECT 26.240 44.215 26.470 45.205 ;
        RECT 24.790 44.045 25.455 44.215 ;
        RECT 24.785 43.375 25.115 43.875 ;
        RECT 25.285 43.545 25.455 44.045 ;
        RECT 25.805 44.045 26.470 44.215 ;
        RECT 25.805 43.545 25.975 44.045 ;
        RECT 26.145 43.375 26.475 43.875 ;
        RECT 26.645 43.545 26.830 45.665 ;
        RECT 27.085 45.465 27.335 45.925 ;
        RECT 27.505 45.475 27.840 45.645 ;
        RECT 28.035 45.475 28.710 45.645 ;
        RECT 27.505 45.335 27.675 45.475 ;
        RECT 27.000 44.345 27.280 45.295 ;
        RECT 27.450 45.205 27.675 45.335 ;
        RECT 27.450 44.100 27.620 45.205 ;
        RECT 27.845 45.055 28.370 45.275 ;
        RECT 27.790 44.290 28.030 44.885 ;
        RECT 28.200 44.355 28.370 45.055 ;
        RECT 28.540 44.695 28.710 45.475 ;
        RECT 29.030 45.425 29.400 45.925 ;
        RECT 29.580 45.475 29.985 45.645 ;
        RECT 30.155 45.475 30.940 45.645 ;
        RECT 29.580 45.245 29.750 45.475 ;
        RECT 28.920 44.945 29.750 45.245 ;
        RECT 30.135 44.975 30.600 45.305 ;
        RECT 28.920 44.915 29.120 44.945 ;
        RECT 29.240 44.695 29.410 44.765 ;
        RECT 28.540 44.525 29.410 44.695 ;
        RECT 28.900 44.435 29.410 44.525 ;
        RECT 27.450 43.970 27.755 44.100 ;
        RECT 28.200 43.990 28.730 44.355 ;
        RECT 27.070 43.375 27.335 43.835 ;
        RECT 27.505 43.545 27.755 43.970 ;
        RECT 28.900 43.820 29.070 44.435 ;
        RECT 27.965 43.650 29.070 43.820 ;
        RECT 29.240 43.375 29.410 44.175 ;
        RECT 29.580 43.875 29.750 44.945 ;
        RECT 29.920 44.045 30.110 44.765 ;
        RECT 30.280 44.015 30.600 44.975 ;
        RECT 30.770 45.015 30.940 45.475 ;
        RECT 31.215 45.395 31.425 45.925 ;
        RECT 31.685 45.185 32.015 45.710 ;
        RECT 32.185 45.315 32.355 45.925 ;
        RECT 32.525 45.270 32.855 45.705 ;
        RECT 32.525 45.185 32.905 45.270 ;
        RECT 31.815 45.015 32.015 45.185 ;
        RECT 32.680 45.145 32.905 45.185 ;
        RECT 30.770 44.685 31.645 45.015 ;
        RECT 31.815 44.685 32.565 45.015 ;
        RECT 29.580 43.545 29.830 43.875 ;
        RECT 30.770 43.845 30.940 44.685 ;
        RECT 31.815 44.480 32.005 44.685 ;
        RECT 32.735 44.565 32.905 45.145 ;
        RECT 32.690 44.515 32.905 44.565 ;
        RECT 31.110 44.105 32.005 44.480 ;
        RECT 32.515 44.435 32.905 44.515 ;
        RECT 33.110 45.185 33.725 45.755 ;
        RECT 33.895 45.415 34.110 45.925 ;
        RECT 34.340 45.415 34.620 45.745 ;
        RECT 34.800 45.415 35.040 45.925 ;
        RECT 30.055 43.675 30.940 43.845 ;
        RECT 31.120 43.375 31.435 43.875 ;
        RECT 31.665 43.545 32.005 44.105 ;
        RECT 32.175 43.375 32.345 44.385 ;
        RECT 32.515 43.590 32.845 44.435 ;
        RECT 33.110 44.165 33.425 45.185 ;
        RECT 33.595 44.515 33.765 45.015 ;
        RECT 34.015 44.685 34.280 45.245 ;
        RECT 34.450 44.515 34.620 45.415 ;
        RECT 35.465 45.375 35.635 45.755 ;
        RECT 35.850 45.545 36.180 45.925 ;
        RECT 34.790 44.685 35.145 45.245 ;
        RECT 35.465 45.205 36.180 45.375 ;
        RECT 35.375 44.655 35.730 45.025 ;
        RECT 36.010 45.015 36.180 45.205 ;
        RECT 36.350 45.180 36.605 45.755 ;
        RECT 36.010 44.685 36.265 45.015 ;
        RECT 33.595 44.345 35.020 44.515 ;
        RECT 36.010 44.475 36.180 44.685 ;
        RECT 33.110 43.545 33.645 44.165 ;
        RECT 33.815 43.375 34.145 44.175 ;
        RECT 34.630 44.170 35.020 44.345 ;
        RECT 35.465 44.305 36.180 44.475 ;
        RECT 36.435 44.450 36.605 45.180 ;
        RECT 36.780 45.085 37.040 45.925 ;
        RECT 37.255 45.105 37.485 45.925 ;
        RECT 37.655 45.125 37.985 45.755 ;
        RECT 37.235 44.685 37.565 44.935 ;
        RECT 37.735 44.525 37.985 45.125 ;
        RECT 38.155 45.105 38.365 45.925 ;
        RECT 38.595 45.200 38.885 45.925 ;
        RECT 39.055 45.185 39.495 45.745 ;
        RECT 39.665 45.185 40.115 45.925 ;
        RECT 40.285 45.355 40.455 45.755 ;
        RECT 40.625 45.525 41.045 45.925 ;
        RECT 41.215 45.355 41.445 45.755 ;
        RECT 40.285 45.185 41.445 45.355 ;
        RECT 41.615 45.185 42.105 45.755 ;
        RECT 35.465 43.545 35.635 44.305 ;
        RECT 35.850 43.375 36.180 44.135 ;
        RECT 36.350 43.545 36.605 44.450 ;
        RECT 36.780 43.375 37.040 44.525 ;
        RECT 37.255 43.375 37.485 44.515 ;
        RECT 37.655 43.545 37.985 44.525 ;
        RECT 38.155 43.375 38.365 44.515 ;
        RECT 38.595 43.375 38.885 44.540 ;
        RECT 39.055 44.175 39.365 45.185 ;
        RECT 39.535 44.565 39.705 45.015 ;
        RECT 39.875 44.735 40.265 45.015 ;
        RECT 40.450 44.685 40.695 45.015 ;
        RECT 39.535 44.395 40.325 44.565 ;
        RECT 39.055 43.545 39.495 44.175 ;
        RECT 39.670 43.375 39.985 44.225 ;
        RECT 40.155 43.715 40.325 44.395 ;
        RECT 40.495 43.885 40.695 44.685 ;
        RECT 40.895 43.885 41.145 45.015 ;
        RECT 41.360 44.685 41.765 45.015 ;
        RECT 41.935 44.515 42.105 45.185 ;
        RECT 42.390 45.295 42.675 45.755 ;
        RECT 42.845 45.465 43.115 45.925 ;
        RECT 42.390 45.125 43.345 45.295 ;
        RECT 41.335 44.345 42.105 44.515 ;
        RECT 42.275 44.395 42.965 44.955 ;
        RECT 41.335 43.715 41.585 44.345 ;
        RECT 43.135 44.225 43.345 45.125 ;
        RECT 40.155 43.545 41.585 43.715 ;
        RECT 41.765 43.375 42.095 44.175 ;
        RECT 42.390 44.005 43.345 44.225 ;
        RECT 43.515 44.955 43.915 45.755 ;
        RECT 44.105 45.295 44.385 45.755 ;
        RECT 44.905 45.465 45.230 45.925 ;
        RECT 44.105 45.125 45.230 45.295 ;
        RECT 45.400 45.185 45.785 45.755 ;
        RECT 44.780 45.015 45.230 45.125 ;
        RECT 43.515 44.395 44.610 44.955 ;
        RECT 44.780 44.685 45.335 45.015 ;
        RECT 42.390 43.545 42.675 44.005 ;
        RECT 42.845 43.375 43.115 43.835 ;
        RECT 43.515 43.545 43.915 44.395 ;
        RECT 44.780 44.225 45.230 44.685 ;
        RECT 45.505 44.515 45.785 45.185 ;
        RECT 44.105 44.005 45.230 44.225 ;
        RECT 44.105 43.545 44.385 44.005 ;
        RECT 44.905 43.375 45.230 43.835 ;
        RECT 45.400 43.545 45.785 44.515 ;
        RECT 45.955 45.250 46.215 45.755 ;
        RECT 46.395 45.545 46.725 45.925 ;
        RECT 46.905 45.375 47.075 45.755 ;
        RECT 45.955 44.450 46.135 45.250 ;
        RECT 46.410 45.205 47.075 45.375 ;
        RECT 46.410 44.950 46.580 45.205 ;
        RECT 47.335 45.175 48.545 45.925 ;
        RECT 46.305 44.620 46.580 44.950 ;
        RECT 46.805 44.655 47.145 45.025 ;
        RECT 46.410 44.475 46.580 44.620 ;
        RECT 45.955 43.545 46.225 44.450 ;
        RECT 46.410 44.305 47.085 44.475 ;
        RECT 46.395 43.375 46.725 44.135 ;
        RECT 46.905 43.545 47.085 44.305 ;
        RECT 47.335 44.465 47.855 45.005 ;
        RECT 48.025 44.635 48.545 45.175 ;
        RECT 47.335 43.375 48.545 44.465 ;
        RECT 12.750 43.205 48.630 43.375 ;
        RECT 12.835 42.115 14.045 43.205 ;
        RECT 14.305 42.535 14.475 43.035 ;
        RECT 14.645 42.705 14.975 43.205 ;
        RECT 14.305 42.365 14.970 42.535 ;
        RECT 12.835 41.405 13.355 41.945 ;
        RECT 13.525 41.575 14.045 42.115 ;
        RECT 14.220 41.545 14.570 42.195 ;
        RECT 12.835 40.655 14.045 41.405 ;
        RECT 14.740 41.375 14.970 42.365 ;
        RECT 14.305 41.205 14.970 41.375 ;
        RECT 14.305 40.915 14.475 41.205 ;
        RECT 14.645 40.655 14.975 41.035 ;
        RECT 15.145 40.915 15.330 43.035 ;
        RECT 15.570 42.745 15.835 43.205 ;
        RECT 16.005 42.610 16.255 43.035 ;
        RECT 16.465 42.760 17.570 42.930 ;
        RECT 15.950 42.480 16.255 42.610 ;
        RECT 15.500 41.285 15.780 42.235 ;
        RECT 15.950 41.375 16.120 42.480 ;
        RECT 16.290 41.695 16.530 42.290 ;
        RECT 16.700 42.225 17.230 42.590 ;
        RECT 16.700 41.525 16.870 42.225 ;
        RECT 17.400 42.145 17.570 42.760 ;
        RECT 17.740 42.405 17.910 43.205 ;
        RECT 18.080 42.705 18.330 43.035 ;
        RECT 18.555 42.735 19.440 42.905 ;
        RECT 17.400 42.055 17.910 42.145 ;
        RECT 15.950 41.245 16.175 41.375 ;
        RECT 16.345 41.305 16.870 41.525 ;
        RECT 17.040 41.885 17.910 42.055 ;
        RECT 15.585 40.655 15.835 41.115 ;
        RECT 16.005 41.105 16.175 41.245 ;
        RECT 17.040 41.105 17.210 41.885 ;
        RECT 17.740 41.815 17.910 41.885 ;
        RECT 17.420 41.635 17.620 41.665 ;
        RECT 18.080 41.635 18.250 42.705 ;
        RECT 18.420 41.815 18.610 42.535 ;
        RECT 17.420 41.335 18.250 41.635 ;
        RECT 18.780 41.605 19.100 42.565 ;
        RECT 16.005 40.935 16.340 41.105 ;
        RECT 16.535 40.935 17.210 41.105 ;
        RECT 17.530 40.655 17.900 41.155 ;
        RECT 18.080 41.105 18.250 41.335 ;
        RECT 18.635 41.275 19.100 41.605 ;
        RECT 19.270 41.895 19.440 42.735 ;
        RECT 19.620 42.705 19.935 43.205 ;
        RECT 20.165 42.475 20.505 43.035 ;
        RECT 19.610 42.100 20.505 42.475 ;
        RECT 20.675 42.195 20.845 43.205 ;
        RECT 20.315 41.895 20.505 42.100 ;
        RECT 21.015 42.145 21.345 42.990 ;
        RECT 21.015 42.065 21.405 42.145 ;
        RECT 21.190 42.015 21.405 42.065 ;
        RECT 19.270 41.565 20.145 41.895 ;
        RECT 20.315 41.565 21.065 41.895 ;
        RECT 19.270 41.105 19.440 41.565 ;
        RECT 20.315 41.395 20.515 41.565 ;
        RECT 21.235 41.435 21.405 42.015 ;
        RECT 21.180 41.395 21.405 41.435 ;
        RECT 18.080 40.935 18.485 41.105 ;
        RECT 18.655 40.935 19.440 41.105 ;
        RECT 19.715 40.655 19.925 41.185 ;
        RECT 20.185 40.870 20.515 41.395 ;
        RECT 21.025 41.310 21.405 41.395 ;
        RECT 21.575 42.065 21.960 43.035 ;
        RECT 22.130 42.745 22.455 43.205 ;
        RECT 22.975 42.575 23.255 43.035 ;
        RECT 22.130 42.355 23.255 42.575 ;
        RECT 21.575 41.395 21.855 42.065 ;
        RECT 22.130 41.895 22.580 42.355 ;
        RECT 23.445 42.185 23.845 43.035 ;
        RECT 24.245 42.745 24.515 43.205 ;
        RECT 24.685 42.575 24.970 43.035 ;
        RECT 22.025 41.565 22.580 41.895 ;
        RECT 22.750 41.625 23.845 42.185 ;
        RECT 22.130 41.455 22.580 41.565 ;
        RECT 20.685 40.655 20.855 41.265 ;
        RECT 21.025 40.875 21.355 41.310 ;
        RECT 21.575 40.825 21.960 41.395 ;
        RECT 22.130 41.285 23.255 41.455 ;
        RECT 22.130 40.655 22.455 41.115 ;
        RECT 22.975 40.825 23.255 41.285 ;
        RECT 23.445 40.825 23.845 41.625 ;
        RECT 24.015 42.355 24.970 42.575 ;
        RECT 24.015 41.455 24.225 42.355 ;
        RECT 24.395 41.625 25.085 42.185 ;
        RECT 25.715 42.040 26.005 43.205 ;
        RECT 26.180 42.065 26.515 43.035 ;
        RECT 26.685 42.065 26.855 43.205 ;
        RECT 27.025 42.865 29.055 43.035 ;
        RECT 24.015 41.285 24.970 41.455 ;
        RECT 26.180 41.395 26.350 42.065 ;
        RECT 27.025 41.895 27.195 42.865 ;
        RECT 26.520 41.565 26.775 41.895 ;
        RECT 27.000 41.565 27.195 41.895 ;
        RECT 27.365 42.525 28.490 42.695 ;
        RECT 26.605 41.395 26.775 41.565 ;
        RECT 27.365 41.395 27.535 42.525 ;
        RECT 24.245 40.655 24.515 41.115 ;
        RECT 24.685 40.825 24.970 41.285 ;
        RECT 25.715 40.655 26.005 41.380 ;
        RECT 26.180 40.825 26.435 41.395 ;
        RECT 26.605 41.225 27.535 41.395 ;
        RECT 27.705 42.185 28.715 42.355 ;
        RECT 27.705 41.385 27.875 42.185 ;
        RECT 28.080 41.845 28.355 41.985 ;
        RECT 28.075 41.675 28.355 41.845 ;
        RECT 27.360 41.190 27.535 41.225 ;
        RECT 26.605 40.655 26.935 41.055 ;
        RECT 27.360 40.825 27.890 41.190 ;
        RECT 28.080 40.825 28.355 41.675 ;
        RECT 28.525 40.825 28.715 42.185 ;
        RECT 28.885 42.200 29.055 42.865 ;
        RECT 29.225 42.445 29.395 43.205 ;
        RECT 29.630 42.445 30.145 42.855 ;
        RECT 28.885 42.010 29.635 42.200 ;
        RECT 29.805 41.635 30.145 42.445 ;
        RECT 30.960 42.235 31.350 42.410 ;
        RECT 31.835 42.405 32.165 43.205 ;
        RECT 32.335 42.415 32.870 43.035 ;
        RECT 30.960 42.065 32.385 42.235 ;
        RECT 28.915 41.465 30.145 41.635 ;
        RECT 28.895 40.655 29.405 41.190 ;
        RECT 29.625 40.860 29.870 41.465 ;
        RECT 30.835 41.335 31.190 41.895 ;
        RECT 31.360 41.165 31.530 42.065 ;
        RECT 31.700 41.335 31.965 41.895 ;
        RECT 32.215 41.565 32.385 42.065 ;
        RECT 32.555 41.395 32.870 42.415 ;
        RECT 33.135 42.065 33.345 43.205 ;
        RECT 33.515 42.055 33.845 43.035 ;
        RECT 34.015 42.065 34.245 43.205 ;
        RECT 34.545 42.535 34.715 43.035 ;
        RECT 34.885 42.705 35.215 43.205 ;
        RECT 34.545 42.365 35.210 42.535 ;
        RECT 30.940 40.655 31.180 41.165 ;
        RECT 31.360 40.835 31.640 41.165 ;
        RECT 31.870 40.655 32.085 41.165 ;
        RECT 32.255 40.825 32.870 41.395 ;
        RECT 33.135 40.655 33.345 41.475 ;
        RECT 33.515 41.455 33.765 42.055 ;
        RECT 33.935 41.645 34.265 41.895 ;
        RECT 34.460 41.545 34.810 42.195 ;
        RECT 33.515 40.825 33.845 41.455 ;
        RECT 34.015 40.655 34.245 41.475 ;
        RECT 34.980 41.375 35.210 42.365 ;
        RECT 34.545 41.205 35.210 41.375 ;
        RECT 34.545 40.915 34.715 41.205 ;
        RECT 34.885 40.655 35.215 41.035 ;
        RECT 35.385 40.915 35.570 43.035 ;
        RECT 35.810 42.745 36.075 43.205 ;
        RECT 36.245 42.610 36.495 43.035 ;
        RECT 36.705 42.760 37.810 42.930 ;
        RECT 36.190 42.480 36.495 42.610 ;
        RECT 35.740 41.285 36.020 42.235 ;
        RECT 36.190 41.375 36.360 42.480 ;
        RECT 36.530 41.695 36.770 42.290 ;
        RECT 36.940 42.225 37.470 42.590 ;
        RECT 36.940 41.525 37.110 42.225 ;
        RECT 37.640 42.145 37.810 42.760 ;
        RECT 37.980 42.405 38.150 43.205 ;
        RECT 38.320 42.705 38.570 43.035 ;
        RECT 38.795 42.735 39.680 42.905 ;
        RECT 37.640 42.055 38.150 42.145 ;
        RECT 36.190 41.245 36.415 41.375 ;
        RECT 36.585 41.305 37.110 41.525 ;
        RECT 37.280 41.885 38.150 42.055 ;
        RECT 35.825 40.655 36.075 41.115 ;
        RECT 36.245 41.105 36.415 41.245 ;
        RECT 37.280 41.105 37.450 41.885 ;
        RECT 37.980 41.815 38.150 41.885 ;
        RECT 37.660 41.635 37.860 41.665 ;
        RECT 38.320 41.635 38.490 42.705 ;
        RECT 38.660 41.815 38.850 42.535 ;
        RECT 37.660 41.335 38.490 41.635 ;
        RECT 39.020 41.605 39.340 42.565 ;
        RECT 36.245 40.935 36.580 41.105 ;
        RECT 36.775 40.935 37.450 41.105 ;
        RECT 37.770 40.655 38.140 41.155 ;
        RECT 38.320 41.105 38.490 41.335 ;
        RECT 38.875 41.275 39.340 41.605 ;
        RECT 39.510 41.895 39.680 42.735 ;
        RECT 39.860 42.705 40.175 43.205 ;
        RECT 40.405 42.475 40.745 43.035 ;
        RECT 39.850 42.100 40.745 42.475 ;
        RECT 40.915 42.195 41.085 43.205 ;
        RECT 40.555 41.895 40.745 42.100 ;
        RECT 41.255 42.145 41.585 42.990 ;
        RECT 42.460 42.235 42.850 42.410 ;
        RECT 43.335 42.405 43.665 43.205 ;
        RECT 43.835 42.415 44.370 43.035 ;
        RECT 41.255 42.065 41.645 42.145 ;
        RECT 42.460 42.065 43.885 42.235 ;
        RECT 41.430 42.015 41.645 42.065 ;
        RECT 39.510 41.565 40.385 41.895 ;
        RECT 40.555 41.565 41.305 41.895 ;
        RECT 39.510 41.105 39.680 41.565 ;
        RECT 40.555 41.395 40.755 41.565 ;
        RECT 41.475 41.435 41.645 42.015 ;
        RECT 41.420 41.395 41.645 41.435 ;
        RECT 38.320 40.935 38.725 41.105 ;
        RECT 38.895 40.935 39.680 41.105 ;
        RECT 39.955 40.655 40.165 41.185 ;
        RECT 40.425 40.870 40.755 41.395 ;
        RECT 41.265 41.310 41.645 41.395 ;
        RECT 42.335 41.335 42.690 41.895 ;
        RECT 40.925 40.655 41.095 41.265 ;
        RECT 41.265 40.875 41.595 41.310 ;
        RECT 42.860 41.165 43.030 42.065 ;
        RECT 43.200 41.335 43.465 41.895 ;
        RECT 43.715 41.565 43.885 42.065 ;
        RECT 44.055 41.395 44.370 42.415 ;
        RECT 44.665 42.275 44.835 43.035 ;
        RECT 45.015 42.445 45.345 43.205 ;
        RECT 44.665 42.105 45.330 42.275 ;
        RECT 45.515 42.130 45.785 43.035 ;
        RECT 45.160 41.960 45.330 42.105 ;
        RECT 44.595 41.555 44.925 41.925 ;
        RECT 45.160 41.630 45.445 41.960 ;
        RECT 42.440 40.655 42.680 41.165 ;
        RECT 42.860 40.835 43.140 41.165 ;
        RECT 43.370 40.655 43.585 41.165 ;
        RECT 43.755 40.825 44.370 41.395 ;
        RECT 45.160 41.375 45.330 41.630 ;
        RECT 44.665 41.205 45.330 41.375 ;
        RECT 45.615 41.330 45.785 42.130 ;
        RECT 44.665 40.825 44.835 41.205 ;
        RECT 45.015 40.655 45.345 41.035 ;
        RECT 45.525 40.825 45.785 41.330 ;
        RECT 45.955 42.130 46.225 43.035 ;
        RECT 46.395 42.445 46.725 43.205 ;
        RECT 46.905 42.275 47.085 43.035 ;
        RECT 45.955 41.330 46.135 42.130 ;
        RECT 46.410 42.105 47.085 42.275 ;
        RECT 47.335 42.115 48.545 43.205 ;
        RECT 46.410 41.960 46.580 42.105 ;
        RECT 46.305 41.630 46.580 41.960 ;
        RECT 46.410 41.375 46.580 41.630 ;
        RECT 46.805 41.555 47.145 41.925 ;
        RECT 47.335 41.575 47.855 42.115 ;
        RECT 48.025 41.405 48.545 41.945 ;
        RECT 45.955 40.825 46.215 41.330 ;
        RECT 46.410 41.205 47.075 41.375 ;
        RECT 46.395 40.655 46.725 41.035 ;
        RECT 46.905 40.825 47.075 41.205 ;
        RECT 47.335 40.655 48.545 41.405 ;
        RECT 12.750 40.485 48.630 40.655 ;
        RECT 12.835 39.735 14.045 40.485 ;
        RECT 12.835 39.195 13.355 39.735 ;
        RECT 14.220 39.645 14.480 40.485 ;
        RECT 14.655 39.740 14.910 40.315 ;
        RECT 15.080 40.105 15.410 40.485 ;
        RECT 15.625 39.935 15.795 40.315 ;
        RECT 15.080 39.765 15.795 39.935 ;
        RECT 13.525 39.025 14.045 39.565 ;
        RECT 12.835 37.935 14.045 39.025 ;
        RECT 14.220 37.935 14.480 39.085 ;
        RECT 14.655 39.010 14.825 39.740 ;
        RECT 15.080 39.575 15.250 39.765 ;
        RECT 16.060 39.745 16.315 40.315 ;
        RECT 16.485 40.085 16.815 40.485 ;
        RECT 17.240 39.950 17.770 40.315 ;
        RECT 17.960 40.145 18.235 40.315 ;
        RECT 17.955 39.975 18.235 40.145 ;
        RECT 17.240 39.915 17.415 39.950 ;
        RECT 16.485 39.745 17.415 39.915 ;
        RECT 14.995 39.245 15.250 39.575 ;
        RECT 15.080 39.035 15.250 39.245 ;
        RECT 15.530 39.215 15.885 39.585 ;
        RECT 16.060 39.075 16.230 39.745 ;
        RECT 16.485 39.575 16.655 39.745 ;
        RECT 16.400 39.245 16.655 39.575 ;
        RECT 16.880 39.245 17.075 39.575 ;
        RECT 14.655 38.105 14.910 39.010 ;
        RECT 15.080 38.865 15.795 39.035 ;
        RECT 15.080 37.935 15.410 38.695 ;
        RECT 15.625 38.105 15.795 38.865 ;
        RECT 16.060 38.105 16.395 39.075 ;
        RECT 16.565 37.935 16.735 39.075 ;
        RECT 16.905 38.275 17.075 39.245 ;
        RECT 17.245 38.615 17.415 39.745 ;
        RECT 17.585 38.955 17.755 39.755 ;
        RECT 17.960 39.155 18.235 39.975 ;
        RECT 18.405 38.955 18.595 40.315 ;
        RECT 18.775 39.950 19.285 40.485 ;
        RECT 19.505 39.675 19.750 40.280 ;
        RECT 20.195 39.735 21.405 40.485 ;
        RECT 21.665 40.005 21.965 40.485 ;
        RECT 22.135 39.835 22.395 40.290 ;
        RECT 22.565 40.005 22.825 40.485 ;
        RECT 23.005 39.835 23.265 40.290 ;
        RECT 23.435 40.005 23.685 40.485 ;
        RECT 23.865 39.835 24.125 40.290 ;
        RECT 24.295 40.005 24.545 40.485 ;
        RECT 24.725 39.835 24.985 40.290 ;
        RECT 25.155 40.005 25.400 40.485 ;
        RECT 25.570 39.835 25.845 40.290 ;
        RECT 26.015 40.005 26.260 40.485 ;
        RECT 26.430 39.835 26.690 40.290 ;
        RECT 26.860 40.005 27.120 40.485 ;
        RECT 27.290 39.835 27.550 40.290 ;
        RECT 27.720 40.005 27.980 40.485 ;
        RECT 28.150 39.835 28.410 40.290 ;
        RECT 28.580 39.925 28.840 40.485 ;
        RECT 18.795 39.505 20.025 39.675 ;
        RECT 17.585 38.785 18.595 38.955 ;
        RECT 18.765 38.940 19.515 39.130 ;
        RECT 17.245 38.445 18.370 38.615 ;
        RECT 18.765 38.275 18.935 38.940 ;
        RECT 19.685 38.695 20.025 39.505 ;
        RECT 20.195 39.195 20.715 39.735 ;
        RECT 21.665 39.665 28.410 39.835 ;
        RECT 20.885 39.025 21.405 39.565 ;
        RECT 16.905 38.105 18.935 38.275 ;
        RECT 19.105 37.935 19.275 38.695 ;
        RECT 19.510 38.285 20.025 38.695 ;
        RECT 20.195 37.935 21.405 39.025 ;
        RECT 21.665 39.075 22.830 39.665 ;
        RECT 29.010 39.495 29.260 40.305 ;
        RECT 29.440 39.960 29.700 40.485 ;
        RECT 29.870 39.495 30.120 40.305 ;
        RECT 30.300 39.975 30.605 40.485 ;
        RECT 23.000 39.245 30.120 39.495 ;
        RECT 30.290 39.245 30.605 39.805 ;
        RECT 30.775 39.745 31.160 40.315 ;
        RECT 31.330 40.025 31.655 40.485 ;
        RECT 32.175 39.855 32.455 40.315 ;
        RECT 21.665 38.850 28.410 39.075 ;
        RECT 21.665 37.935 21.935 38.680 ;
        RECT 22.105 38.110 22.395 38.850 ;
        RECT 23.005 38.835 28.410 38.850 ;
        RECT 22.565 37.940 22.820 38.665 ;
        RECT 23.005 38.110 23.265 38.835 ;
        RECT 23.435 37.940 23.680 38.665 ;
        RECT 23.865 38.110 24.125 38.835 ;
        RECT 24.295 37.940 24.540 38.665 ;
        RECT 24.725 38.110 24.985 38.835 ;
        RECT 25.155 37.940 25.400 38.665 ;
        RECT 25.570 38.110 25.830 38.835 ;
        RECT 26.000 37.940 26.260 38.665 ;
        RECT 26.430 38.110 26.690 38.835 ;
        RECT 26.860 37.940 27.120 38.665 ;
        RECT 27.290 38.110 27.550 38.835 ;
        RECT 27.720 37.940 27.980 38.665 ;
        RECT 28.150 38.110 28.410 38.835 ;
        RECT 28.580 37.940 28.840 38.735 ;
        RECT 29.010 38.110 29.260 39.245 ;
        RECT 22.565 37.935 28.840 37.940 ;
        RECT 29.440 37.935 29.700 38.745 ;
        RECT 29.875 38.105 30.120 39.245 ;
        RECT 30.775 39.075 31.055 39.745 ;
        RECT 31.330 39.685 32.455 39.855 ;
        RECT 31.330 39.575 31.780 39.685 ;
        RECT 31.225 39.245 31.780 39.575 ;
        RECT 32.645 39.515 33.045 40.315 ;
        RECT 33.445 40.025 33.715 40.485 ;
        RECT 33.885 39.855 34.170 40.315 ;
        RECT 30.300 37.935 30.595 38.745 ;
        RECT 30.775 38.105 31.160 39.075 ;
        RECT 31.330 38.785 31.780 39.245 ;
        RECT 31.950 38.955 33.045 39.515 ;
        RECT 31.330 38.565 32.455 38.785 ;
        RECT 31.330 37.935 31.655 38.395 ;
        RECT 32.175 38.105 32.455 38.565 ;
        RECT 32.645 38.105 33.045 38.955 ;
        RECT 33.215 39.685 34.170 39.855 ;
        RECT 34.455 39.735 35.665 40.485 ;
        RECT 35.845 39.985 36.175 40.485 ;
        RECT 36.375 39.915 36.545 40.265 ;
        RECT 36.745 40.085 37.075 40.485 ;
        RECT 37.245 39.915 37.415 40.265 ;
        RECT 37.585 40.085 37.965 40.485 ;
        RECT 33.215 38.785 33.425 39.685 ;
        RECT 33.595 38.955 34.285 39.515 ;
        RECT 34.455 39.195 34.975 39.735 ;
        RECT 35.145 39.025 35.665 39.565 ;
        RECT 35.840 39.245 36.190 39.815 ;
        RECT 36.375 39.745 37.985 39.915 ;
        RECT 38.155 39.810 38.425 40.155 ;
        RECT 37.815 39.575 37.985 39.745 ;
        RECT 33.215 38.565 34.170 38.785 ;
        RECT 33.445 37.935 33.715 38.395 ;
        RECT 33.885 38.105 34.170 38.565 ;
        RECT 34.455 37.935 35.665 39.025 ;
        RECT 35.840 38.785 36.160 39.075 ;
        RECT 36.360 38.955 37.070 39.575 ;
        RECT 37.240 39.245 37.645 39.575 ;
        RECT 37.815 39.245 38.085 39.575 ;
        RECT 37.815 39.075 37.985 39.245 ;
        RECT 38.255 39.075 38.425 39.810 ;
        RECT 38.595 39.760 38.885 40.485 ;
        RECT 39.055 39.745 39.415 40.120 ;
        RECT 39.680 39.745 39.850 40.485 ;
        RECT 40.130 39.915 40.300 40.120 ;
        RECT 40.130 39.745 40.670 39.915 ;
        RECT 37.260 38.905 37.985 39.075 ;
        RECT 37.260 38.785 37.430 38.905 ;
        RECT 35.840 38.615 37.430 38.785 ;
        RECT 35.840 38.155 37.495 38.445 ;
        RECT 37.665 37.935 37.945 38.735 ;
        RECT 38.155 38.105 38.425 39.075 ;
        RECT 38.595 37.935 38.885 39.100 ;
        RECT 39.055 39.090 39.310 39.745 ;
        RECT 39.480 39.245 39.830 39.575 ;
        RECT 40.000 39.245 40.330 39.575 ;
        RECT 39.055 38.105 39.395 39.090 ;
        RECT 39.565 38.705 39.830 39.245 ;
        RECT 40.500 39.045 40.670 39.745 ;
        RECT 40.045 38.875 40.670 39.045 ;
        RECT 40.840 39.115 41.010 40.315 ;
        RECT 41.240 39.835 41.570 40.315 ;
        RECT 41.740 40.015 41.910 40.485 ;
        RECT 42.080 39.835 42.410 40.300 ;
        RECT 41.240 39.665 42.410 39.835 ;
        RECT 42.735 39.745 43.095 40.120 ;
        RECT 43.360 39.745 43.530 40.485 ;
        RECT 43.810 39.915 43.980 40.120 ;
        RECT 43.810 39.745 44.350 39.915 ;
        RECT 41.180 39.285 41.750 39.495 ;
        RECT 41.920 39.285 42.565 39.495 ;
        RECT 40.840 38.705 41.545 39.115 ;
        RECT 42.735 39.090 42.990 39.745 ;
        RECT 43.160 39.245 43.510 39.575 ;
        RECT 43.680 39.245 44.010 39.575 ;
        RECT 39.565 38.535 41.545 38.705 ;
        RECT 39.565 37.935 39.975 38.365 ;
        RECT 40.720 37.935 41.050 38.355 ;
        RECT 41.220 38.105 41.545 38.535 ;
        RECT 42.020 37.935 42.350 39.035 ;
        RECT 42.735 38.105 43.075 39.090 ;
        RECT 43.245 38.705 43.510 39.245 ;
        RECT 44.180 39.045 44.350 39.745 ;
        RECT 43.725 38.875 44.350 39.045 ;
        RECT 44.520 39.115 44.690 40.315 ;
        RECT 44.920 39.835 45.250 40.315 ;
        RECT 45.420 40.015 45.590 40.485 ;
        RECT 45.760 39.835 46.090 40.300 ;
        RECT 44.920 39.665 46.090 39.835 ;
        RECT 47.335 39.735 48.545 40.485 ;
        RECT 44.860 39.285 45.430 39.495 ;
        RECT 45.600 39.285 46.245 39.495 ;
        RECT 44.520 38.705 45.225 39.115 ;
        RECT 43.245 38.535 45.225 38.705 ;
        RECT 43.245 37.935 43.655 38.365 ;
        RECT 44.400 37.935 44.730 38.355 ;
        RECT 44.900 38.105 45.225 38.535 ;
        RECT 45.700 37.935 46.030 39.035 ;
        RECT 47.335 39.025 47.855 39.565 ;
        RECT 48.025 39.195 48.545 39.735 ;
        RECT 47.335 37.935 48.545 39.025 ;
        RECT 12.750 37.765 48.630 37.935 ;
        RECT 12.835 36.675 14.045 37.765 ;
        RECT 12.835 35.965 13.355 36.505 ;
        RECT 13.525 36.135 14.045 36.675 ;
        RECT 14.220 36.625 14.555 37.595 ;
        RECT 14.725 36.625 14.895 37.765 ;
        RECT 15.065 37.425 17.095 37.595 ;
        RECT 12.835 35.215 14.045 35.965 ;
        RECT 14.220 35.955 14.390 36.625 ;
        RECT 15.065 36.455 15.235 37.425 ;
        RECT 14.560 36.125 14.815 36.455 ;
        RECT 15.040 36.125 15.235 36.455 ;
        RECT 15.405 37.085 16.530 37.255 ;
        RECT 14.645 35.955 14.815 36.125 ;
        RECT 15.405 35.955 15.575 37.085 ;
        RECT 14.220 35.385 14.475 35.955 ;
        RECT 14.645 35.785 15.575 35.955 ;
        RECT 15.745 36.745 16.755 36.915 ;
        RECT 15.745 35.945 15.915 36.745 ;
        RECT 15.400 35.750 15.575 35.785 ;
        RECT 14.645 35.215 14.975 35.615 ;
        RECT 15.400 35.385 15.930 35.750 ;
        RECT 16.120 35.725 16.395 36.545 ;
        RECT 16.115 35.555 16.395 35.725 ;
        RECT 16.120 35.385 16.395 35.555 ;
        RECT 16.565 35.385 16.755 36.745 ;
        RECT 16.925 36.760 17.095 37.425 ;
        RECT 17.265 37.005 17.435 37.765 ;
        RECT 17.670 37.005 18.185 37.415 ;
        RECT 16.925 36.570 17.675 36.760 ;
        RECT 17.845 36.195 18.185 37.005 ;
        RECT 18.445 37.095 18.615 37.595 ;
        RECT 18.785 37.265 19.115 37.765 ;
        RECT 18.445 36.925 19.110 37.095 ;
        RECT 16.955 36.025 18.185 36.195 ;
        RECT 18.360 36.105 18.710 36.755 ;
        RECT 16.935 35.215 17.445 35.750 ;
        RECT 17.665 35.420 17.910 36.025 ;
        RECT 18.880 35.935 19.110 36.925 ;
        RECT 18.445 35.765 19.110 35.935 ;
        RECT 18.445 35.475 18.615 35.765 ;
        RECT 18.785 35.215 19.115 35.595 ;
        RECT 19.285 35.475 19.470 37.595 ;
        RECT 19.710 37.305 19.975 37.765 ;
        RECT 20.145 37.170 20.395 37.595 ;
        RECT 20.605 37.320 21.710 37.490 ;
        RECT 20.090 37.040 20.395 37.170 ;
        RECT 19.640 35.845 19.920 36.795 ;
        RECT 20.090 35.935 20.260 37.040 ;
        RECT 20.430 36.255 20.670 36.850 ;
        RECT 20.840 36.785 21.370 37.150 ;
        RECT 20.840 36.085 21.010 36.785 ;
        RECT 21.540 36.705 21.710 37.320 ;
        RECT 21.880 36.965 22.050 37.765 ;
        RECT 22.220 37.265 22.470 37.595 ;
        RECT 22.695 37.295 23.580 37.465 ;
        RECT 21.540 36.615 22.050 36.705 ;
        RECT 20.090 35.805 20.315 35.935 ;
        RECT 20.485 35.865 21.010 36.085 ;
        RECT 21.180 36.445 22.050 36.615 ;
        RECT 19.725 35.215 19.975 35.675 ;
        RECT 20.145 35.665 20.315 35.805 ;
        RECT 21.180 35.665 21.350 36.445 ;
        RECT 21.880 36.375 22.050 36.445 ;
        RECT 21.560 36.195 21.760 36.225 ;
        RECT 22.220 36.195 22.390 37.265 ;
        RECT 22.560 36.375 22.750 37.095 ;
        RECT 21.560 35.895 22.390 36.195 ;
        RECT 22.920 36.165 23.240 37.125 ;
        RECT 20.145 35.495 20.480 35.665 ;
        RECT 20.675 35.495 21.350 35.665 ;
        RECT 21.670 35.215 22.040 35.715 ;
        RECT 22.220 35.665 22.390 35.895 ;
        RECT 22.775 35.835 23.240 36.165 ;
        RECT 23.410 36.455 23.580 37.295 ;
        RECT 23.760 37.265 24.075 37.765 ;
        RECT 24.305 37.035 24.645 37.595 ;
        RECT 23.750 36.660 24.645 37.035 ;
        RECT 24.815 36.755 24.985 37.765 ;
        RECT 24.455 36.455 24.645 36.660 ;
        RECT 25.155 36.705 25.485 37.550 ;
        RECT 25.155 36.625 25.545 36.705 ;
        RECT 25.330 36.575 25.545 36.625 ;
        RECT 25.715 36.600 26.005 37.765 ;
        RECT 26.265 37.095 26.435 37.595 ;
        RECT 26.605 37.265 26.935 37.765 ;
        RECT 26.265 36.925 26.930 37.095 ;
        RECT 23.410 36.125 24.285 36.455 ;
        RECT 24.455 36.125 25.205 36.455 ;
        RECT 23.410 35.665 23.580 36.125 ;
        RECT 24.455 35.955 24.655 36.125 ;
        RECT 25.375 35.995 25.545 36.575 ;
        RECT 26.180 36.105 26.530 36.755 ;
        RECT 25.320 35.955 25.545 35.995 ;
        RECT 22.220 35.495 22.625 35.665 ;
        RECT 22.795 35.495 23.580 35.665 ;
        RECT 23.855 35.215 24.065 35.745 ;
        RECT 24.325 35.430 24.655 35.955 ;
        RECT 25.165 35.870 25.545 35.955 ;
        RECT 24.825 35.215 24.995 35.825 ;
        RECT 25.165 35.435 25.495 35.870 ;
        RECT 25.715 35.215 26.005 35.940 ;
        RECT 26.700 35.935 26.930 36.925 ;
        RECT 26.265 35.765 26.930 35.935 ;
        RECT 26.265 35.475 26.435 35.765 ;
        RECT 26.605 35.215 26.935 35.595 ;
        RECT 27.105 35.475 27.290 37.595 ;
        RECT 27.530 37.305 27.795 37.765 ;
        RECT 27.965 37.170 28.215 37.595 ;
        RECT 28.425 37.320 29.530 37.490 ;
        RECT 27.910 37.040 28.215 37.170 ;
        RECT 27.460 35.845 27.740 36.795 ;
        RECT 27.910 35.935 28.080 37.040 ;
        RECT 28.250 36.255 28.490 36.850 ;
        RECT 28.660 36.785 29.190 37.150 ;
        RECT 28.660 36.085 28.830 36.785 ;
        RECT 29.360 36.705 29.530 37.320 ;
        RECT 29.700 36.965 29.870 37.765 ;
        RECT 30.040 37.265 30.290 37.595 ;
        RECT 30.515 37.295 31.400 37.465 ;
        RECT 29.360 36.615 29.870 36.705 ;
        RECT 27.910 35.805 28.135 35.935 ;
        RECT 28.305 35.865 28.830 36.085 ;
        RECT 29.000 36.445 29.870 36.615 ;
        RECT 27.545 35.215 27.795 35.675 ;
        RECT 27.965 35.665 28.135 35.805 ;
        RECT 29.000 35.665 29.170 36.445 ;
        RECT 29.700 36.375 29.870 36.445 ;
        RECT 29.380 36.195 29.580 36.225 ;
        RECT 30.040 36.195 30.210 37.265 ;
        RECT 30.380 36.375 30.570 37.095 ;
        RECT 29.380 35.895 30.210 36.195 ;
        RECT 30.740 36.165 31.060 37.125 ;
        RECT 27.965 35.495 28.300 35.665 ;
        RECT 28.495 35.495 29.170 35.665 ;
        RECT 29.490 35.215 29.860 35.715 ;
        RECT 30.040 35.665 30.210 35.895 ;
        RECT 30.595 35.835 31.060 36.165 ;
        RECT 31.230 36.455 31.400 37.295 ;
        RECT 31.580 37.265 31.895 37.765 ;
        RECT 32.125 37.035 32.465 37.595 ;
        RECT 31.570 36.660 32.465 37.035 ;
        RECT 32.635 36.755 32.805 37.765 ;
        RECT 32.275 36.455 32.465 36.660 ;
        RECT 32.975 36.705 33.305 37.550 ;
        RECT 33.995 36.810 34.265 37.765 ;
        RECT 34.450 36.710 34.755 37.495 ;
        RECT 34.935 37.295 35.620 37.765 ;
        RECT 34.930 36.775 35.625 37.085 ;
        RECT 32.975 36.625 33.365 36.705 ;
        RECT 33.150 36.575 33.365 36.625 ;
        RECT 31.230 36.125 32.105 36.455 ;
        RECT 32.275 36.125 33.025 36.455 ;
        RECT 31.230 35.665 31.400 36.125 ;
        RECT 32.275 35.955 32.475 36.125 ;
        RECT 33.195 35.995 33.365 36.575 ;
        RECT 33.140 35.955 33.365 35.995 ;
        RECT 30.040 35.495 30.445 35.665 ;
        RECT 30.615 35.495 31.400 35.665 ;
        RECT 31.675 35.215 31.885 35.745 ;
        RECT 32.145 35.430 32.475 35.955 ;
        RECT 32.985 35.870 33.365 35.955 ;
        RECT 34.450 35.905 34.625 36.710 ;
        RECT 35.800 36.605 36.085 37.550 ;
        RECT 36.285 37.315 36.615 37.765 ;
        RECT 36.785 37.145 36.955 37.575 ;
        RECT 35.225 36.455 36.085 36.605 ;
        RECT 34.795 36.435 36.085 36.455 ;
        RECT 36.275 36.915 36.955 37.145 ;
        RECT 38.135 36.965 38.575 37.595 ;
        RECT 34.795 36.075 35.785 36.435 ;
        RECT 36.275 36.265 36.510 36.915 ;
        RECT 32.645 35.215 32.815 35.825 ;
        RECT 32.985 35.435 33.315 35.870 ;
        RECT 33.995 35.215 34.265 35.850 ;
        RECT 34.450 35.385 34.685 35.905 ;
        RECT 35.615 35.740 35.785 36.075 ;
        RECT 35.955 35.935 36.510 36.265 ;
        RECT 36.295 35.785 36.510 35.935 ;
        RECT 36.680 36.065 36.980 36.745 ;
        RECT 36.680 35.895 36.985 36.065 ;
        RECT 38.135 35.955 38.445 36.965 ;
        RECT 38.750 36.915 39.065 37.765 ;
        RECT 39.235 37.425 40.665 37.595 ;
        RECT 39.235 36.745 39.405 37.425 ;
        RECT 38.615 36.575 39.405 36.745 ;
        RECT 38.615 36.125 38.785 36.575 ;
        RECT 39.575 36.455 39.775 37.255 ;
        RECT 38.955 36.125 39.345 36.405 ;
        RECT 39.530 36.125 39.775 36.455 ;
        RECT 39.975 36.125 40.225 37.255 ;
        RECT 40.415 36.795 40.665 37.425 ;
        RECT 40.845 36.965 41.175 37.765 ;
        RECT 41.365 36.795 41.695 37.580 ;
        RECT 40.415 36.625 41.185 36.795 ;
        RECT 41.365 36.625 42.045 36.795 ;
        RECT 42.225 36.625 42.555 37.765 ;
        RECT 40.440 36.125 40.845 36.455 ;
        RECT 41.015 35.955 41.185 36.625 ;
        RECT 41.355 36.205 41.705 36.455 ;
        RECT 41.875 36.025 42.045 36.625 ;
        RECT 43.195 36.610 43.535 37.595 ;
        RECT 43.705 37.335 44.115 37.765 ;
        RECT 44.860 37.345 45.190 37.765 ;
        RECT 45.360 37.165 45.685 37.595 ;
        RECT 43.705 36.995 45.685 37.165 ;
        RECT 42.215 36.205 42.565 36.455 ;
        RECT 34.855 35.215 35.255 35.710 ;
        RECT 35.615 35.545 36.015 35.740 ;
        RECT 35.845 35.400 36.015 35.545 ;
        RECT 36.295 35.410 36.535 35.785 ;
        RECT 36.705 35.215 37.035 35.720 ;
        RECT 38.135 35.395 38.575 35.955 ;
        RECT 38.745 35.215 39.195 35.955 ;
        RECT 39.365 35.785 40.525 35.955 ;
        RECT 39.365 35.385 39.535 35.785 ;
        RECT 39.705 35.215 40.125 35.615 ;
        RECT 40.295 35.385 40.525 35.785 ;
        RECT 40.695 35.385 41.185 35.955 ;
        RECT 41.375 35.215 41.615 36.025 ;
        RECT 41.785 35.385 42.115 36.025 ;
        RECT 42.285 35.215 42.555 36.025 ;
        RECT 43.195 35.955 43.450 36.610 ;
        RECT 43.705 36.455 43.970 36.995 ;
        RECT 44.185 36.655 44.810 36.825 ;
        RECT 43.620 36.125 43.970 36.455 ;
        RECT 44.140 36.125 44.470 36.455 ;
        RECT 44.640 35.955 44.810 36.655 ;
        RECT 43.195 35.580 43.555 35.955 ;
        RECT 43.820 35.215 43.990 35.955 ;
        RECT 44.270 35.785 44.810 35.955 ;
        RECT 44.980 36.585 45.685 36.995 ;
        RECT 46.160 36.665 46.490 37.765 ;
        RECT 47.335 36.675 48.545 37.765 ;
        RECT 44.270 35.580 44.440 35.785 ;
        RECT 44.980 35.385 45.150 36.585 ;
        RECT 45.320 36.205 45.890 36.415 ;
        RECT 46.060 36.205 46.705 36.415 ;
        RECT 47.335 36.135 47.855 36.675 ;
        RECT 45.380 35.865 46.550 36.035 ;
        RECT 48.025 35.965 48.545 36.505 ;
        RECT 45.380 35.385 45.710 35.865 ;
        RECT 45.880 35.215 46.050 35.685 ;
        RECT 46.220 35.400 46.550 35.865 ;
        RECT 47.335 35.215 48.545 35.965 ;
        RECT 12.750 35.045 48.630 35.215 ;
        RECT 12.835 34.295 14.045 35.045 ;
        RECT 14.265 34.390 14.595 34.825 ;
        RECT 14.765 34.435 14.935 35.045 ;
        RECT 14.215 34.305 14.595 34.390 ;
        RECT 15.105 34.305 15.435 34.830 ;
        RECT 15.695 34.515 15.905 35.045 ;
        RECT 16.180 34.595 16.965 34.765 ;
        RECT 17.135 34.595 17.540 34.765 ;
        RECT 12.835 33.755 13.355 34.295 ;
        RECT 14.215 34.265 14.440 34.305 ;
        RECT 13.525 33.585 14.045 34.125 ;
        RECT 12.835 32.495 14.045 33.585 ;
        RECT 14.215 33.685 14.385 34.265 ;
        RECT 15.105 34.135 15.305 34.305 ;
        RECT 16.180 34.135 16.350 34.595 ;
        RECT 14.555 33.805 15.305 34.135 ;
        RECT 15.475 33.805 16.350 34.135 ;
        RECT 14.215 33.635 14.430 33.685 ;
        RECT 14.215 33.555 14.605 33.635 ;
        RECT 14.275 32.710 14.605 33.555 ;
        RECT 15.115 33.600 15.305 33.805 ;
        RECT 14.775 32.495 14.945 33.505 ;
        RECT 15.115 33.225 16.010 33.600 ;
        RECT 15.115 32.665 15.455 33.225 ;
        RECT 15.685 32.495 16.000 32.995 ;
        RECT 16.180 32.965 16.350 33.805 ;
        RECT 16.520 34.095 16.985 34.425 ;
        RECT 17.370 34.365 17.540 34.595 ;
        RECT 17.720 34.545 18.090 35.045 ;
        RECT 18.410 34.595 19.085 34.765 ;
        RECT 19.280 34.595 19.615 34.765 ;
        RECT 16.520 33.135 16.840 34.095 ;
        RECT 17.370 34.065 18.200 34.365 ;
        RECT 17.010 33.165 17.200 33.885 ;
        RECT 17.370 32.995 17.540 34.065 ;
        RECT 18.000 34.035 18.200 34.065 ;
        RECT 17.710 33.815 17.880 33.885 ;
        RECT 18.410 33.815 18.580 34.595 ;
        RECT 19.445 34.455 19.615 34.595 ;
        RECT 19.785 34.585 20.035 35.045 ;
        RECT 17.710 33.645 18.580 33.815 ;
        RECT 18.750 34.175 19.275 34.395 ;
        RECT 19.445 34.325 19.670 34.455 ;
        RECT 17.710 33.555 18.220 33.645 ;
        RECT 16.180 32.795 17.065 32.965 ;
        RECT 17.290 32.665 17.540 32.995 ;
        RECT 17.710 32.495 17.880 33.295 ;
        RECT 18.050 32.940 18.220 33.555 ;
        RECT 18.750 33.475 18.920 34.175 ;
        RECT 18.390 33.110 18.920 33.475 ;
        RECT 19.090 33.410 19.330 34.005 ;
        RECT 19.500 33.220 19.670 34.325 ;
        RECT 19.840 33.465 20.120 34.415 ;
        RECT 19.365 33.090 19.670 33.220 ;
        RECT 18.050 32.770 19.155 32.940 ;
        RECT 19.365 32.665 19.615 33.090 ;
        RECT 19.785 32.495 20.050 32.955 ;
        RECT 20.290 32.665 20.475 34.785 ;
        RECT 20.645 34.665 20.975 35.045 ;
        RECT 21.145 34.495 21.315 34.785 ;
        RECT 20.650 34.325 21.315 34.495 ;
        RECT 20.650 33.335 20.880 34.325 ;
        RECT 21.575 34.275 24.165 35.045 ;
        RECT 24.795 34.535 25.100 35.045 ;
        RECT 21.050 33.505 21.400 34.155 ;
        RECT 21.575 33.755 22.785 34.275 ;
        RECT 22.955 33.585 24.165 34.105 ;
        RECT 24.795 33.805 25.110 34.365 ;
        RECT 25.280 34.055 25.530 34.865 ;
        RECT 25.700 34.520 25.960 35.045 ;
        RECT 26.140 34.055 26.390 34.865 ;
        RECT 26.560 34.485 26.820 35.045 ;
        RECT 26.990 34.395 27.250 34.850 ;
        RECT 27.420 34.565 27.680 35.045 ;
        RECT 27.850 34.395 28.110 34.850 ;
        RECT 28.280 34.565 28.540 35.045 ;
        RECT 28.710 34.395 28.970 34.850 ;
        RECT 29.140 34.565 29.385 35.045 ;
        RECT 29.555 34.395 29.830 34.850 ;
        RECT 30.000 34.565 30.245 35.045 ;
        RECT 30.415 34.395 30.675 34.850 ;
        RECT 30.855 34.565 31.105 35.045 ;
        RECT 31.275 34.395 31.535 34.850 ;
        RECT 31.715 34.565 31.965 35.045 ;
        RECT 32.135 34.395 32.395 34.850 ;
        RECT 32.575 34.565 32.835 35.045 ;
        RECT 33.005 34.395 33.265 34.850 ;
        RECT 33.435 34.565 33.735 35.045 ;
        RECT 26.990 34.225 33.735 34.395 ;
        RECT 25.280 33.805 32.400 34.055 ;
        RECT 20.650 33.165 21.315 33.335 ;
        RECT 20.645 32.495 20.975 32.995 ;
        RECT 21.145 32.665 21.315 33.165 ;
        RECT 21.575 32.495 24.165 33.585 ;
        RECT 24.805 32.495 25.100 33.305 ;
        RECT 25.280 32.665 25.525 33.805 ;
        RECT 25.700 32.495 25.960 33.305 ;
        RECT 26.140 32.670 26.390 33.805 ;
        RECT 32.570 33.635 33.735 34.225 ;
        RECT 26.990 33.410 33.735 33.635 ;
        RECT 33.995 34.305 34.380 34.875 ;
        RECT 34.550 34.585 34.875 35.045 ;
        RECT 35.395 34.415 35.675 34.875 ;
        RECT 33.995 33.635 34.275 34.305 ;
        RECT 34.550 34.245 35.675 34.415 ;
        RECT 34.550 34.135 35.000 34.245 ;
        RECT 34.445 33.805 35.000 34.135 ;
        RECT 35.865 34.075 36.265 34.875 ;
        RECT 36.665 34.585 36.935 35.045 ;
        RECT 37.105 34.415 37.390 34.875 ;
        RECT 26.990 33.395 32.395 33.410 ;
        RECT 26.560 32.500 26.820 33.295 ;
        RECT 26.990 32.670 27.250 33.395 ;
        RECT 27.420 32.500 27.680 33.225 ;
        RECT 27.850 32.670 28.110 33.395 ;
        RECT 28.280 32.500 28.540 33.225 ;
        RECT 28.710 32.670 28.970 33.395 ;
        RECT 29.140 32.500 29.400 33.225 ;
        RECT 29.570 32.670 29.830 33.395 ;
        RECT 30.000 32.500 30.245 33.225 ;
        RECT 30.415 32.670 30.675 33.395 ;
        RECT 30.860 32.500 31.105 33.225 ;
        RECT 31.275 32.670 31.535 33.395 ;
        RECT 31.720 32.500 31.965 33.225 ;
        RECT 32.135 32.670 32.395 33.395 ;
        RECT 32.580 32.500 32.835 33.225 ;
        RECT 33.005 32.670 33.295 33.410 ;
        RECT 26.560 32.495 32.835 32.500 ;
        RECT 33.465 32.495 33.735 33.240 ;
        RECT 33.995 32.665 34.380 33.635 ;
        RECT 34.550 33.345 35.000 33.805 ;
        RECT 35.170 33.515 36.265 34.075 ;
        RECT 34.550 33.125 35.675 33.345 ;
        RECT 34.550 32.495 34.875 32.955 ;
        RECT 35.395 32.665 35.675 33.125 ;
        RECT 35.865 32.665 36.265 33.515 ;
        RECT 36.435 34.245 37.390 34.415 ;
        RECT 38.595 34.320 38.885 35.045 ;
        RECT 39.070 34.475 39.325 34.825 ;
        RECT 39.495 34.645 39.825 35.045 ;
        RECT 39.995 34.475 40.165 34.825 ;
        RECT 40.335 34.645 40.715 35.045 ;
        RECT 39.070 34.305 40.735 34.475 ;
        RECT 40.905 34.370 41.180 34.715 ;
        RECT 36.435 33.345 36.645 34.245 ;
        RECT 40.565 34.135 40.735 34.305 ;
        RECT 36.815 33.515 37.505 34.075 ;
        RECT 39.055 33.805 39.400 34.135 ;
        RECT 39.570 33.805 40.395 34.135 ;
        RECT 40.565 33.805 40.840 34.135 ;
        RECT 36.435 33.125 37.390 33.345 ;
        RECT 36.665 32.495 36.935 32.955 ;
        RECT 37.105 32.665 37.390 33.125 ;
        RECT 38.595 32.495 38.885 33.660 ;
        RECT 39.075 33.345 39.400 33.635 ;
        RECT 39.570 33.515 39.765 33.805 ;
        RECT 40.565 33.635 40.735 33.805 ;
        RECT 41.010 33.635 41.180 34.370 ;
        RECT 41.355 34.275 43.945 35.045 ;
        RECT 41.355 33.755 42.565 34.275 ;
        RECT 44.585 34.235 44.855 35.045 ;
        RECT 45.025 34.235 45.355 34.875 ;
        RECT 45.525 34.235 45.765 35.045 ;
        RECT 45.955 34.370 46.215 34.875 ;
        RECT 46.395 34.665 46.725 35.045 ;
        RECT 46.905 34.495 47.075 34.875 ;
        RECT 40.075 33.465 40.735 33.635 ;
        RECT 40.075 33.345 40.245 33.465 ;
        RECT 39.075 33.175 40.245 33.345 ;
        RECT 39.055 32.715 40.245 33.005 ;
        RECT 40.415 32.495 40.695 33.295 ;
        RECT 40.905 32.665 41.180 33.635 ;
        RECT 42.735 33.585 43.945 34.105 ;
        RECT 44.575 33.805 44.925 34.055 ;
        RECT 45.095 33.635 45.265 34.235 ;
        RECT 45.435 33.805 45.785 34.055 ;
        RECT 41.355 32.495 43.945 33.585 ;
        RECT 44.585 32.495 44.915 33.635 ;
        RECT 45.095 33.465 45.775 33.635 ;
        RECT 45.445 32.680 45.775 33.465 ;
        RECT 45.955 33.570 46.125 34.370 ;
        RECT 46.410 34.325 47.075 34.495 ;
        RECT 46.410 34.070 46.580 34.325 ;
        RECT 47.335 34.295 48.545 35.045 ;
        RECT 46.295 33.740 46.580 34.070 ;
        RECT 46.815 33.775 47.145 34.145 ;
        RECT 46.410 33.595 46.580 33.740 ;
        RECT 45.955 32.665 46.225 33.570 ;
        RECT 46.410 33.425 47.075 33.595 ;
        RECT 46.395 32.495 46.725 33.255 ;
        RECT 46.905 32.665 47.075 33.425 ;
        RECT 47.335 33.585 47.855 34.125 ;
        RECT 48.025 33.755 48.545 34.295 ;
        RECT 47.335 32.495 48.545 33.585 ;
        RECT 12.750 32.325 48.630 32.495 ;
        RECT 12.835 31.235 14.045 32.325 ;
        RECT 14.215 31.235 15.425 32.325 ;
        RECT 15.710 31.695 15.995 32.155 ;
        RECT 16.165 31.865 16.435 32.325 ;
        RECT 15.710 31.475 16.665 31.695 ;
        RECT 12.835 30.525 13.355 31.065 ;
        RECT 13.525 30.695 14.045 31.235 ;
        RECT 14.215 30.525 14.735 31.065 ;
        RECT 14.905 30.695 15.425 31.235 ;
        RECT 15.595 30.745 16.285 31.305 ;
        RECT 16.455 30.575 16.665 31.475 ;
        RECT 12.835 29.775 14.045 30.525 ;
        RECT 14.215 29.775 15.425 30.525 ;
        RECT 15.710 30.405 16.665 30.575 ;
        RECT 16.835 31.305 17.235 32.155 ;
        RECT 17.425 31.695 17.705 32.155 ;
        RECT 18.225 31.865 18.550 32.325 ;
        RECT 17.425 31.475 18.550 31.695 ;
        RECT 16.835 30.745 17.930 31.305 ;
        RECT 18.100 31.015 18.550 31.475 ;
        RECT 18.720 31.185 19.105 32.155 ;
        RECT 15.710 29.945 15.995 30.405 ;
        RECT 16.165 29.775 16.435 30.235 ;
        RECT 16.835 29.945 17.235 30.745 ;
        RECT 18.100 30.685 18.655 31.015 ;
        RECT 18.100 30.575 18.550 30.685 ;
        RECT 17.425 30.405 18.550 30.575 ;
        RECT 18.825 30.515 19.105 31.185 ;
        RECT 17.425 29.945 17.705 30.405 ;
        RECT 18.225 29.775 18.550 30.235 ;
        RECT 18.720 29.945 19.105 30.515 ;
        RECT 19.275 31.185 19.660 32.155 ;
        RECT 19.830 31.865 20.155 32.325 ;
        RECT 20.675 31.695 20.955 32.155 ;
        RECT 19.830 31.475 20.955 31.695 ;
        RECT 19.275 30.515 19.555 31.185 ;
        RECT 19.830 31.015 20.280 31.475 ;
        RECT 21.145 31.305 21.545 32.155 ;
        RECT 21.945 31.865 22.215 32.325 ;
        RECT 22.385 31.695 22.670 32.155 ;
        RECT 19.725 30.685 20.280 31.015 ;
        RECT 20.450 30.745 21.545 31.305 ;
        RECT 19.830 30.575 20.280 30.685 ;
        RECT 19.275 29.945 19.660 30.515 ;
        RECT 19.830 30.405 20.955 30.575 ;
        RECT 19.830 29.775 20.155 30.235 ;
        RECT 20.675 29.945 20.955 30.405 ;
        RECT 21.145 29.945 21.545 30.745 ;
        RECT 21.715 31.475 22.670 31.695 ;
        RECT 21.715 30.575 21.925 31.475 ;
        RECT 22.095 30.745 22.785 31.305 ;
        RECT 22.955 31.235 25.545 32.325 ;
        RECT 21.715 30.405 22.670 30.575 ;
        RECT 21.945 29.775 22.215 30.235 ;
        RECT 22.385 29.945 22.670 30.405 ;
        RECT 22.955 30.545 24.165 31.065 ;
        RECT 24.335 30.715 25.545 31.235 ;
        RECT 25.715 31.160 26.005 32.325 ;
        RECT 26.185 31.185 26.515 32.325 ;
        RECT 27.045 31.355 27.375 32.140 ;
        RECT 26.695 31.185 27.375 31.355 ;
        RECT 27.675 31.205 28.005 32.325 ;
        RECT 26.175 30.765 26.525 31.015 ;
        RECT 26.695 30.585 26.865 31.185 ;
        RECT 27.035 30.765 27.385 31.015 ;
        RECT 27.615 30.765 28.125 31.015 ;
        RECT 28.335 30.765 28.705 32.080 ;
        RECT 28.875 30.765 29.205 32.080 ;
        RECT 29.415 30.765 29.745 32.080 ;
        RECT 30.015 31.435 30.265 32.155 ;
        RECT 30.435 31.605 30.765 32.325 ;
        RECT 30.015 31.145 30.765 31.435 ;
        RECT 31.000 31.145 31.525 32.155 ;
        RECT 30.505 30.975 30.765 31.145 ;
        RECT 29.915 30.765 30.335 30.975 ;
        RECT 30.505 30.765 31.085 30.975 ;
        RECT 30.505 30.595 30.875 30.765 ;
        RECT 22.955 29.775 25.545 30.545 ;
        RECT 25.715 29.775 26.005 30.500 ;
        RECT 26.185 29.775 26.455 30.585 ;
        RECT 26.625 29.945 26.955 30.585 ;
        RECT 27.125 29.775 27.365 30.585 ;
        RECT 27.655 30.425 29.955 30.595 ;
        RECT 27.655 29.945 27.985 30.425 ;
        RECT 28.155 29.775 28.485 30.235 ;
        RECT 28.700 29.945 29.030 30.425 ;
        RECT 29.230 29.775 29.560 30.235 ;
        RECT 29.785 30.105 29.955 30.425 ;
        RECT 30.125 30.405 30.875 30.595 ;
        RECT 31.255 30.575 31.525 31.145 ;
        RECT 30.125 29.960 30.455 30.405 ;
        RECT 30.725 29.775 30.895 30.235 ;
        RECT 31.185 29.945 31.525 30.575 ;
        RECT 31.695 31.185 32.080 32.155 ;
        RECT 32.250 31.865 32.575 32.325 ;
        RECT 33.095 31.695 33.375 32.155 ;
        RECT 32.250 31.475 33.375 31.695 ;
        RECT 31.695 30.515 31.975 31.185 ;
        RECT 32.250 31.015 32.700 31.475 ;
        RECT 33.565 31.305 33.965 32.155 ;
        RECT 34.365 31.865 34.635 32.325 ;
        RECT 34.805 31.695 35.090 32.155 ;
        RECT 32.145 30.685 32.700 31.015 ;
        RECT 32.870 30.745 33.965 31.305 ;
        RECT 32.250 30.575 32.700 30.685 ;
        RECT 31.695 29.945 32.080 30.515 ;
        RECT 32.250 30.405 33.375 30.575 ;
        RECT 32.250 29.775 32.575 30.235 ;
        RECT 33.095 29.945 33.375 30.405 ;
        RECT 33.565 29.945 33.965 30.745 ;
        RECT 34.135 31.475 35.090 31.695 ;
        RECT 34.135 30.575 34.345 31.475 ;
        RECT 34.515 30.745 35.205 31.305 ;
        RECT 35.375 31.235 36.585 32.325 ;
        RECT 34.135 30.405 35.090 30.575 ;
        RECT 34.365 29.775 34.635 30.235 ;
        RECT 34.805 29.945 35.090 30.405 ;
        RECT 35.375 30.525 35.895 31.065 ;
        RECT 36.065 30.695 36.585 31.235 ;
        RECT 36.755 31.185 37.030 32.155 ;
        RECT 37.240 31.525 37.520 32.325 ;
        RECT 37.690 31.815 39.740 32.105 ;
        RECT 37.690 31.475 39.320 31.645 ;
        RECT 37.690 31.355 37.860 31.475 ;
        RECT 37.200 31.185 37.860 31.355 ;
        RECT 35.375 29.775 36.585 30.525 ;
        RECT 36.755 30.450 36.925 31.185 ;
        RECT 37.200 31.015 37.370 31.185 ;
        RECT 37.095 30.685 37.370 31.015 ;
        RECT 37.540 30.685 37.920 31.015 ;
        RECT 38.090 30.685 38.830 31.305 ;
        RECT 39.000 31.185 39.320 31.475 ;
        RECT 39.515 31.015 39.755 31.610 ;
        RECT 39.925 31.250 40.265 32.325 ;
        RECT 40.445 31.355 40.775 32.140 ;
        RECT 40.445 31.185 41.125 31.355 ;
        RECT 41.305 31.185 41.635 32.325 ;
        RECT 41.895 31.395 42.075 32.155 ;
        RECT 42.255 31.565 42.585 32.325 ;
        RECT 41.895 31.225 42.570 31.395 ;
        RECT 42.755 31.250 43.025 32.155 ;
        RECT 39.100 30.685 39.755 31.015 ;
        RECT 37.200 30.515 37.370 30.685 ;
        RECT 36.755 30.105 37.030 30.450 ;
        RECT 37.200 30.345 38.785 30.515 ;
        RECT 37.220 29.775 37.600 30.175 ;
        RECT 37.770 29.995 37.940 30.345 ;
        RECT 38.110 29.775 38.440 30.175 ;
        RECT 38.615 29.995 38.785 30.345 ;
        RECT 38.985 29.775 39.315 30.275 ;
        RECT 39.510 29.995 39.755 30.685 ;
        RECT 39.925 30.445 40.265 31.015 ;
        RECT 40.435 30.765 40.785 31.015 ;
        RECT 40.955 30.585 41.125 31.185 ;
        RECT 42.400 31.080 42.570 31.225 ;
        RECT 41.295 30.765 41.645 31.015 ;
        RECT 41.835 30.675 42.175 31.045 ;
        RECT 42.400 30.750 42.675 31.080 ;
        RECT 39.925 29.775 40.265 30.275 ;
        RECT 40.455 29.775 40.695 30.585 ;
        RECT 40.865 29.945 41.195 30.585 ;
        RECT 41.365 29.775 41.635 30.585 ;
        RECT 42.400 30.495 42.570 30.750 ;
        RECT 41.905 30.325 42.570 30.495 ;
        RECT 42.845 30.450 43.025 31.250 ;
        RECT 43.410 31.225 43.740 32.325 ;
        RECT 44.215 31.725 44.540 32.155 ;
        RECT 44.710 31.905 45.040 32.325 ;
        RECT 45.785 31.895 46.195 32.325 ;
        RECT 44.215 31.555 46.195 31.725 ;
        RECT 44.215 31.145 44.920 31.555 ;
        RECT 43.195 30.765 43.840 30.975 ;
        RECT 44.010 30.765 44.580 30.975 ;
        RECT 41.905 29.945 42.075 30.325 ;
        RECT 42.255 29.775 42.585 30.155 ;
        RECT 42.765 29.945 43.025 30.450 ;
        RECT 43.350 30.425 44.520 30.595 ;
        RECT 43.350 29.960 43.680 30.425 ;
        RECT 43.850 29.775 44.020 30.245 ;
        RECT 44.190 29.945 44.520 30.425 ;
        RECT 44.750 29.945 44.920 31.145 ;
        RECT 45.090 31.215 45.715 31.385 ;
        RECT 45.090 30.515 45.260 31.215 ;
        RECT 45.930 31.015 46.195 31.555 ;
        RECT 46.365 31.170 46.705 32.155 ;
        RECT 45.430 30.685 45.760 31.015 ;
        RECT 45.930 30.685 46.280 31.015 ;
        RECT 46.450 30.515 46.705 31.170 ;
        RECT 47.335 31.235 48.545 32.325 ;
        RECT 47.335 30.695 47.855 31.235 ;
        RECT 48.025 30.525 48.545 31.065 ;
        RECT 45.090 30.345 45.630 30.515 ;
        RECT 45.460 30.140 45.630 30.345 ;
        RECT 45.910 29.775 46.080 30.515 ;
        RECT 46.345 30.140 46.705 30.515 ;
        RECT 47.335 29.775 48.545 30.525 ;
        RECT 12.750 29.605 48.630 29.775 ;
        RECT 12.835 28.855 14.045 29.605 ;
        RECT 12.835 28.315 13.355 28.855 ;
        RECT 14.220 28.765 14.480 29.605 ;
        RECT 14.655 28.860 14.910 29.435 ;
        RECT 15.080 29.225 15.410 29.605 ;
        RECT 15.625 29.055 15.795 29.435 ;
        RECT 15.080 28.885 15.795 29.055 ;
        RECT 13.525 28.145 14.045 28.685 ;
        RECT 12.835 27.055 14.045 28.145 ;
        RECT 14.220 27.055 14.480 28.205 ;
        RECT 14.655 28.130 14.825 28.860 ;
        RECT 15.080 28.695 15.250 28.885 ;
        RECT 16.520 28.865 16.775 29.435 ;
        RECT 16.945 29.205 17.275 29.605 ;
        RECT 17.700 29.070 18.230 29.435 ;
        RECT 18.420 29.265 18.695 29.435 ;
        RECT 18.415 29.095 18.695 29.265 ;
        RECT 17.700 29.035 17.875 29.070 ;
        RECT 16.945 28.865 17.875 29.035 ;
        RECT 14.995 28.365 15.250 28.695 ;
        RECT 15.080 28.155 15.250 28.365 ;
        RECT 15.530 28.335 15.885 28.705 ;
        RECT 16.520 28.195 16.690 28.865 ;
        RECT 16.945 28.695 17.115 28.865 ;
        RECT 16.860 28.365 17.115 28.695 ;
        RECT 17.340 28.365 17.535 28.695 ;
        RECT 14.655 27.225 14.910 28.130 ;
        RECT 15.080 27.985 15.795 28.155 ;
        RECT 15.080 27.055 15.410 27.815 ;
        RECT 15.625 27.225 15.795 27.985 ;
        RECT 16.520 27.225 16.855 28.195 ;
        RECT 17.025 27.055 17.195 28.195 ;
        RECT 17.365 27.395 17.535 28.365 ;
        RECT 17.705 27.735 17.875 28.865 ;
        RECT 18.045 28.075 18.215 28.875 ;
        RECT 18.420 28.275 18.695 29.095 ;
        RECT 18.865 28.075 19.055 29.435 ;
        RECT 19.235 29.070 19.745 29.605 ;
        RECT 19.965 28.795 20.210 29.400 ;
        RECT 20.745 29.055 20.915 29.345 ;
        RECT 21.085 29.225 21.415 29.605 ;
        RECT 20.745 28.885 21.410 29.055 ;
        RECT 19.255 28.625 20.485 28.795 ;
        RECT 18.045 27.905 19.055 28.075 ;
        RECT 19.225 28.060 19.975 28.250 ;
        RECT 17.705 27.565 18.830 27.735 ;
        RECT 19.225 27.395 19.395 28.060 ;
        RECT 20.145 27.815 20.485 28.625 ;
        RECT 20.660 28.065 21.010 28.715 ;
        RECT 21.180 27.895 21.410 28.885 ;
        RECT 17.365 27.225 19.395 27.395 ;
        RECT 19.565 27.055 19.735 27.815 ;
        RECT 19.970 27.405 20.485 27.815 ;
        RECT 20.745 27.725 21.410 27.895 ;
        RECT 20.745 27.225 20.915 27.725 ;
        RECT 21.085 27.055 21.415 27.555 ;
        RECT 21.585 27.225 21.770 29.345 ;
        RECT 22.025 29.145 22.275 29.605 ;
        RECT 22.445 29.155 22.780 29.325 ;
        RECT 22.975 29.155 23.650 29.325 ;
        RECT 22.445 29.015 22.615 29.155 ;
        RECT 21.940 28.025 22.220 28.975 ;
        RECT 22.390 28.885 22.615 29.015 ;
        RECT 22.390 27.780 22.560 28.885 ;
        RECT 22.785 28.735 23.310 28.955 ;
        RECT 22.730 27.970 22.970 28.565 ;
        RECT 23.140 28.035 23.310 28.735 ;
        RECT 23.480 28.375 23.650 29.155 ;
        RECT 23.970 29.105 24.340 29.605 ;
        RECT 24.520 29.155 24.925 29.325 ;
        RECT 25.095 29.155 25.880 29.325 ;
        RECT 24.520 28.925 24.690 29.155 ;
        RECT 23.860 28.625 24.690 28.925 ;
        RECT 25.075 28.655 25.540 28.985 ;
        RECT 23.860 28.595 24.060 28.625 ;
        RECT 24.180 28.375 24.350 28.445 ;
        RECT 23.480 28.205 24.350 28.375 ;
        RECT 23.840 28.115 24.350 28.205 ;
        RECT 22.390 27.650 22.695 27.780 ;
        RECT 23.140 27.670 23.670 28.035 ;
        RECT 22.010 27.055 22.275 27.515 ;
        RECT 22.445 27.225 22.695 27.650 ;
        RECT 23.840 27.500 24.010 28.115 ;
        RECT 22.905 27.330 24.010 27.500 ;
        RECT 24.180 27.055 24.350 27.855 ;
        RECT 24.520 27.555 24.690 28.625 ;
        RECT 24.860 27.725 25.050 28.445 ;
        RECT 25.220 27.695 25.540 28.655 ;
        RECT 25.710 28.695 25.880 29.155 ;
        RECT 26.155 29.075 26.365 29.605 ;
        RECT 26.625 28.865 26.955 29.390 ;
        RECT 27.125 28.995 27.295 29.605 ;
        RECT 27.465 28.950 27.795 29.385 ;
        RECT 27.465 28.865 27.845 28.950 ;
        RECT 26.755 28.695 26.955 28.865 ;
        RECT 27.620 28.825 27.845 28.865 ;
        RECT 25.710 28.365 26.585 28.695 ;
        RECT 26.755 28.365 27.505 28.695 ;
        RECT 24.520 27.225 24.770 27.555 ;
        RECT 25.710 27.525 25.880 28.365 ;
        RECT 26.755 28.160 26.945 28.365 ;
        RECT 27.675 28.245 27.845 28.825 ;
        RECT 27.630 28.195 27.845 28.245 ;
        RECT 26.050 27.785 26.945 28.160 ;
        RECT 27.455 28.115 27.845 28.195 ;
        RECT 28.020 28.865 28.275 29.435 ;
        RECT 28.445 29.205 28.775 29.605 ;
        RECT 29.200 29.070 29.730 29.435 ;
        RECT 29.200 29.035 29.375 29.070 ;
        RECT 28.445 28.865 29.375 29.035 ;
        RECT 28.020 28.195 28.190 28.865 ;
        RECT 28.445 28.695 28.615 28.865 ;
        RECT 28.360 28.365 28.615 28.695 ;
        RECT 28.840 28.365 29.035 28.695 ;
        RECT 24.995 27.355 25.880 27.525 ;
        RECT 26.060 27.055 26.375 27.555 ;
        RECT 26.605 27.225 26.945 27.785 ;
        RECT 27.115 27.055 27.285 28.065 ;
        RECT 27.455 27.270 27.785 28.115 ;
        RECT 28.020 27.225 28.355 28.195 ;
        RECT 28.525 27.055 28.695 28.195 ;
        RECT 28.865 27.395 29.035 28.365 ;
        RECT 29.205 27.735 29.375 28.865 ;
        RECT 29.545 28.075 29.715 28.875 ;
        RECT 29.920 28.585 30.195 29.435 ;
        RECT 29.915 28.415 30.195 28.585 ;
        RECT 29.920 28.275 30.195 28.415 ;
        RECT 30.365 28.075 30.555 29.435 ;
        RECT 30.735 29.070 31.245 29.605 ;
        RECT 31.465 28.795 31.710 29.400 ;
        RECT 32.155 28.865 32.540 29.435 ;
        RECT 32.710 29.145 33.035 29.605 ;
        RECT 33.555 28.975 33.835 29.435 ;
        RECT 30.755 28.625 31.985 28.795 ;
        RECT 29.545 27.905 30.555 28.075 ;
        RECT 30.725 28.060 31.475 28.250 ;
        RECT 29.205 27.565 30.330 27.735 ;
        RECT 30.725 27.395 30.895 28.060 ;
        RECT 31.645 27.815 31.985 28.625 ;
        RECT 28.865 27.225 30.895 27.395 ;
        RECT 31.065 27.055 31.235 27.815 ;
        RECT 31.470 27.405 31.985 27.815 ;
        RECT 32.155 28.195 32.435 28.865 ;
        RECT 32.710 28.805 33.835 28.975 ;
        RECT 32.710 28.695 33.160 28.805 ;
        RECT 32.605 28.365 33.160 28.695 ;
        RECT 34.025 28.635 34.425 29.435 ;
        RECT 34.825 29.145 35.095 29.605 ;
        RECT 35.265 28.975 35.550 29.435 ;
        RECT 32.155 27.225 32.540 28.195 ;
        RECT 32.710 27.905 33.160 28.365 ;
        RECT 33.330 28.075 34.425 28.635 ;
        RECT 32.710 27.685 33.835 27.905 ;
        RECT 32.710 27.055 33.035 27.515 ;
        RECT 33.555 27.225 33.835 27.685 ;
        RECT 34.025 27.225 34.425 28.075 ;
        RECT 34.595 28.805 35.550 28.975 ;
        RECT 35.835 28.835 38.425 29.605 ;
        RECT 38.595 28.880 38.885 29.605 ;
        RECT 39.385 29.205 39.715 29.605 ;
        RECT 39.885 29.035 40.215 29.375 ;
        RECT 41.265 29.205 41.595 29.605 ;
        RECT 39.230 28.865 41.595 29.035 ;
        RECT 41.765 28.880 42.095 29.390 ;
        RECT 34.595 27.905 34.805 28.805 ;
        RECT 34.975 28.075 35.665 28.635 ;
        RECT 35.835 28.315 37.045 28.835 ;
        RECT 37.215 28.145 38.425 28.665 ;
        RECT 34.595 27.685 35.550 27.905 ;
        RECT 34.825 27.055 35.095 27.515 ;
        RECT 35.265 27.225 35.550 27.685 ;
        RECT 35.835 27.055 38.425 28.145 ;
        RECT 38.595 27.055 38.885 28.220 ;
        RECT 39.230 27.865 39.400 28.865 ;
        RECT 41.425 28.695 41.595 28.865 ;
        RECT 39.570 28.035 39.815 28.695 ;
        RECT 40.030 28.035 40.295 28.695 ;
        RECT 40.490 28.035 40.775 28.695 ;
        RECT 40.950 28.365 41.255 28.695 ;
        RECT 41.425 28.365 41.735 28.695 ;
        RECT 40.950 28.035 41.165 28.365 ;
        RECT 39.230 27.695 39.685 27.865 ;
        RECT 39.355 27.265 39.685 27.695 ;
        RECT 39.865 27.695 41.155 27.865 ;
        RECT 39.865 27.275 40.115 27.695 ;
        RECT 40.345 27.055 40.675 27.525 ;
        RECT 40.905 27.275 41.155 27.695 ;
        RECT 41.345 27.055 41.595 28.195 ;
        RECT 41.905 28.115 42.095 28.880 ;
        RECT 43.350 28.955 43.680 29.420 ;
        RECT 43.850 29.135 44.020 29.605 ;
        RECT 44.190 28.955 44.520 29.435 ;
        RECT 43.350 28.785 44.520 28.955 ;
        RECT 43.195 28.405 43.840 28.615 ;
        RECT 44.010 28.405 44.580 28.615 ;
        RECT 44.750 28.235 44.920 29.435 ;
        RECT 45.460 29.035 45.630 29.240 ;
        RECT 41.765 27.265 42.095 28.115 ;
        RECT 43.410 27.055 43.740 28.155 ;
        RECT 44.215 27.825 44.920 28.235 ;
        RECT 45.090 28.865 45.630 29.035 ;
        RECT 45.910 28.865 46.080 29.605 ;
        RECT 46.475 29.240 46.645 29.265 ;
        RECT 46.345 28.865 46.705 29.240 ;
        RECT 45.090 28.165 45.260 28.865 ;
        RECT 45.430 28.365 45.760 28.695 ;
        RECT 45.930 28.365 46.280 28.695 ;
        RECT 45.090 27.995 45.715 28.165 ;
        RECT 45.930 27.825 46.195 28.365 ;
        RECT 46.450 28.210 46.705 28.865 ;
        RECT 47.335 28.855 48.545 29.605 ;
        RECT 44.215 27.655 46.195 27.825 ;
        RECT 44.215 27.225 44.540 27.655 ;
        RECT 44.710 27.055 45.040 27.475 ;
        RECT 45.785 27.055 46.195 27.485 ;
        RECT 46.365 27.225 46.705 28.210 ;
        RECT 47.335 28.145 47.855 28.685 ;
        RECT 48.025 28.315 48.545 28.855 ;
        RECT 47.335 27.055 48.545 28.145 ;
        RECT 12.750 26.885 48.630 27.055 ;
        RECT 12.835 25.795 14.045 26.885 ;
        RECT 14.305 26.215 14.475 26.715 ;
        RECT 14.645 26.385 14.975 26.885 ;
        RECT 14.305 26.045 14.970 26.215 ;
        RECT 12.835 25.085 13.355 25.625 ;
        RECT 13.525 25.255 14.045 25.795 ;
        RECT 14.220 25.225 14.570 25.875 ;
        RECT 12.835 24.335 14.045 25.085 ;
        RECT 14.740 25.055 14.970 26.045 ;
        RECT 14.305 24.885 14.970 25.055 ;
        RECT 14.305 24.595 14.475 24.885 ;
        RECT 14.645 24.335 14.975 24.715 ;
        RECT 15.145 24.595 15.330 26.715 ;
        RECT 15.570 26.425 15.835 26.885 ;
        RECT 16.005 26.290 16.255 26.715 ;
        RECT 16.465 26.440 17.570 26.610 ;
        RECT 15.950 26.160 16.255 26.290 ;
        RECT 15.500 24.965 15.780 25.915 ;
        RECT 15.950 25.055 16.120 26.160 ;
        RECT 16.290 25.375 16.530 25.970 ;
        RECT 16.700 25.905 17.230 26.270 ;
        RECT 16.700 25.205 16.870 25.905 ;
        RECT 17.400 25.825 17.570 26.440 ;
        RECT 17.740 26.085 17.910 26.885 ;
        RECT 18.080 26.385 18.330 26.715 ;
        RECT 18.555 26.415 19.440 26.585 ;
        RECT 17.400 25.735 17.910 25.825 ;
        RECT 15.950 24.925 16.175 25.055 ;
        RECT 16.345 24.985 16.870 25.205 ;
        RECT 17.040 25.565 17.910 25.735 ;
        RECT 15.585 24.335 15.835 24.795 ;
        RECT 16.005 24.785 16.175 24.925 ;
        RECT 17.040 24.785 17.210 25.565 ;
        RECT 17.740 25.495 17.910 25.565 ;
        RECT 17.420 25.315 17.620 25.345 ;
        RECT 18.080 25.315 18.250 26.385 ;
        RECT 18.420 25.495 18.610 26.215 ;
        RECT 17.420 25.015 18.250 25.315 ;
        RECT 18.780 25.285 19.100 26.245 ;
        RECT 16.005 24.615 16.340 24.785 ;
        RECT 16.535 24.615 17.210 24.785 ;
        RECT 17.530 24.335 17.900 24.835 ;
        RECT 18.080 24.785 18.250 25.015 ;
        RECT 18.635 24.955 19.100 25.285 ;
        RECT 19.270 25.575 19.440 26.415 ;
        RECT 19.620 26.385 19.935 26.885 ;
        RECT 20.165 26.155 20.505 26.715 ;
        RECT 19.610 25.780 20.505 26.155 ;
        RECT 20.675 25.875 20.845 26.885 ;
        RECT 20.315 25.575 20.505 25.780 ;
        RECT 21.015 25.825 21.345 26.670 ;
        RECT 21.015 25.745 21.405 25.825 ;
        RECT 21.575 25.795 25.085 26.885 ;
        RECT 21.190 25.695 21.405 25.745 ;
        RECT 19.270 25.245 20.145 25.575 ;
        RECT 20.315 25.245 21.065 25.575 ;
        RECT 19.270 24.785 19.440 25.245 ;
        RECT 20.315 25.075 20.515 25.245 ;
        RECT 21.235 25.115 21.405 25.695 ;
        RECT 21.180 25.075 21.405 25.115 ;
        RECT 18.080 24.615 18.485 24.785 ;
        RECT 18.655 24.615 19.440 24.785 ;
        RECT 19.715 24.335 19.925 24.865 ;
        RECT 20.185 24.550 20.515 25.075 ;
        RECT 21.025 24.990 21.405 25.075 ;
        RECT 21.575 25.105 23.225 25.625 ;
        RECT 23.395 25.275 25.085 25.795 ;
        RECT 25.715 25.720 26.005 26.885 ;
        RECT 26.265 26.215 26.435 26.715 ;
        RECT 26.605 26.385 26.935 26.885 ;
        RECT 26.265 26.045 26.930 26.215 ;
        RECT 26.180 25.225 26.530 25.875 ;
        RECT 20.685 24.335 20.855 24.945 ;
        RECT 21.025 24.555 21.355 24.990 ;
        RECT 21.575 24.335 25.085 25.105 ;
        RECT 25.715 24.335 26.005 25.060 ;
        RECT 26.700 25.055 26.930 26.045 ;
        RECT 26.265 24.885 26.930 25.055 ;
        RECT 26.265 24.595 26.435 24.885 ;
        RECT 26.605 24.335 26.935 24.715 ;
        RECT 27.105 24.595 27.290 26.715 ;
        RECT 27.530 26.425 27.795 26.885 ;
        RECT 27.965 26.290 28.215 26.715 ;
        RECT 28.425 26.440 29.530 26.610 ;
        RECT 27.910 26.160 28.215 26.290 ;
        RECT 27.460 24.965 27.740 25.915 ;
        RECT 27.910 25.055 28.080 26.160 ;
        RECT 28.250 25.375 28.490 25.970 ;
        RECT 28.660 25.905 29.190 26.270 ;
        RECT 28.660 25.205 28.830 25.905 ;
        RECT 29.360 25.825 29.530 26.440 ;
        RECT 29.700 26.085 29.870 26.885 ;
        RECT 30.040 26.385 30.290 26.715 ;
        RECT 30.515 26.415 31.400 26.585 ;
        RECT 29.360 25.735 29.870 25.825 ;
        RECT 27.910 24.925 28.135 25.055 ;
        RECT 28.305 24.985 28.830 25.205 ;
        RECT 29.000 25.565 29.870 25.735 ;
        RECT 27.545 24.335 27.795 24.795 ;
        RECT 27.965 24.785 28.135 24.925 ;
        RECT 29.000 24.785 29.170 25.565 ;
        RECT 29.700 25.495 29.870 25.565 ;
        RECT 29.380 25.315 29.580 25.345 ;
        RECT 30.040 25.315 30.210 26.385 ;
        RECT 30.380 25.495 30.570 26.215 ;
        RECT 29.380 25.015 30.210 25.315 ;
        RECT 30.740 25.285 31.060 26.245 ;
        RECT 27.965 24.615 28.300 24.785 ;
        RECT 28.495 24.615 29.170 24.785 ;
        RECT 29.490 24.335 29.860 24.835 ;
        RECT 30.040 24.785 30.210 25.015 ;
        RECT 30.595 24.955 31.060 25.285 ;
        RECT 31.230 25.575 31.400 26.415 ;
        RECT 31.580 26.385 31.895 26.885 ;
        RECT 32.125 26.155 32.465 26.715 ;
        RECT 31.570 25.780 32.465 26.155 ;
        RECT 32.635 25.875 32.805 26.885 ;
        RECT 32.275 25.575 32.465 25.780 ;
        RECT 32.975 25.825 33.305 26.670 ;
        RECT 33.625 26.265 33.795 26.695 ;
        RECT 33.965 26.435 34.295 26.885 ;
        RECT 33.625 26.035 34.305 26.265 ;
        RECT 32.975 25.745 33.365 25.825 ;
        RECT 33.150 25.695 33.365 25.745 ;
        RECT 33.595 25.695 33.900 25.865 ;
        RECT 31.230 25.245 32.105 25.575 ;
        RECT 32.275 25.245 33.025 25.575 ;
        RECT 31.230 24.785 31.400 25.245 ;
        RECT 32.275 25.075 32.475 25.245 ;
        RECT 33.195 25.115 33.365 25.695 ;
        RECT 33.140 25.075 33.365 25.115 ;
        RECT 30.040 24.615 30.445 24.785 ;
        RECT 30.615 24.615 31.400 24.785 ;
        RECT 31.675 24.335 31.885 24.865 ;
        RECT 32.145 24.550 32.475 25.075 ;
        RECT 32.985 24.990 33.365 25.075 ;
        RECT 33.600 25.015 33.900 25.695 ;
        RECT 34.070 25.385 34.305 26.035 ;
        RECT 34.495 25.725 34.780 26.670 ;
        RECT 34.960 26.415 35.645 26.885 ;
        RECT 34.955 25.895 35.650 26.205 ;
        RECT 35.825 25.830 36.130 26.615 ;
        RECT 36.315 25.930 36.585 26.885 ;
        RECT 34.495 25.575 35.355 25.725 ;
        RECT 34.495 25.555 35.785 25.575 ;
        RECT 34.070 25.055 34.625 25.385 ;
        RECT 34.795 25.195 35.785 25.555 ;
        RECT 32.645 24.335 32.815 24.945 ;
        RECT 32.985 24.555 33.315 24.990 ;
        RECT 34.070 24.905 34.285 25.055 ;
        RECT 33.545 24.335 33.875 24.840 ;
        RECT 34.045 24.530 34.285 24.905 ;
        RECT 34.795 24.860 34.965 25.195 ;
        RECT 35.955 25.025 36.130 25.830 ;
        RECT 36.755 25.795 39.345 26.885 ;
        RECT 40.090 26.255 40.375 26.715 ;
        RECT 40.545 26.425 40.815 26.885 ;
        RECT 40.090 26.035 41.045 26.255 ;
        RECT 34.565 24.665 34.965 24.860 ;
        RECT 34.565 24.520 34.735 24.665 ;
        RECT 35.325 24.335 35.725 24.830 ;
        RECT 35.895 24.505 36.130 25.025 ;
        RECT 36.755 25.105 37.965 25.625 ;
        RECT 38.135 25.275 39.345 25.795 ;
        RECT 39.975 25.305 40.665 25.865 ;
        RECT 40.835 25.135 41.045 26.035 ;
        RECT 36.315 24.335 36.585 24.970 ;
        RECT 36.755 24.335 39.345 25.105 ;
        RECT 40.090 24.965 41.045 25.135 ;
        RECT 41.215 25.865 41.615 26.715 ;
        RECT 41.805 26.255 42.085 26.715 ;
        RECT 42.605 26.425 42.930 26.885 ;
        RECT 41.805 26.035 42.930 26.255 ;
        RECT 41.215 25.305 42.310 25.865 ;
        RECT 42.480 25.575 42.930 26.035 ;
        RECT 43.100 25.745 43.485 26.715 ;
        RECT 40.090 24.505 40.375 24.965 ;
        RECT 40.545 24.335 40.815 24.795 ;
        RECT 41.215 24.505 41.615 25.305 ;
        RECT 42.480 25.245 43.035 25.575 ;
        RECT 42.480 25.135 42.930 25.245 ;
        RECT 41.805 24.965 42.930 25.135 ;
        RECT 43.205 25.075 43.485 25.745 ;
        RECT 41.805 24.505 42.085 24.965 ;
        RECT 42.605 24.335 42.930 24.795 ;
        RECT 43.100 24.505 43.485 25.075 ;
        RECT 43.655 26.085 44.095 26.715 ;
        RECT 43.655 25.075 43.965 26.085 ;
        RECT 44.270 26.035 44.585 26.885 ;
        RECT 44.755 26.545 46.185 26.715 ;
        RECT 44.755 25.865 44.925 26.545 ;
        RECT 44.135 25.695 44.925 25.865 ;
        RECT 44.135 25.245 44.305 25.695 ;
        RECT 45.095 25.575 45.295 26.375 ;
        RECT 44.475 25.245 44.865 25.525 ;
        RECT 45.050 25.245 45.295 25.575 ;
        RECT 45.495 25.245 45.745 26.375 ;
        RECT 45.935 25.915 46.185 26.545 ;
        RECT 46.365 26.085 46.695 26.885 ;
        RECT 45.935 25.745 46.705 25.915 ;
        RECT 45.960 25.245 46.365 25.575 ;
        RECT 46.535 25.075 46.705 25.745 ;
        RECT 47.335 25.795 48.545 26.885 ;
        RECT 47.335 25.255 47.855 25.795 ;
        RECT 48.025 25.085 48.545 25.625 ;
        RECT 43.655 24.515 44.095 25.075 ;
        RECT 44.265 24.335 44.715 25.075 ;
        RECT 44.885 24.905 46.045 25.075 ;
        RECT 44.885 24.505 45.055 24.905 ;
        RECT 45.225 24.335 45.645 24.735 ;
        RECT 45.815 24.505 46.045 24.905 ;
        RECT 46.215 24.505 46.705 25.075 ;
        RECT 47.335 24.335 48.545 25.085 ;
        RECT 12.750 24.165 48.630 24.335 ;
        RECT 12.835 23.415 14.045 24.165 ;
        RECT 12.835 22.875 13.355 23.415 ;
        RECT 14.220 23.325 14.480 24.165 ;
        RECT 14.655 23.420 14.910 23.995 ;
        RECT 15.080 23.785 15.410 24.165 ;
        RECT 15.625 23.615 15.795 23.995 ;
        RECT 15.080 23.445 15.795 23.615 ;
        RECT 17.090 23.535 17.375 23.995 ;
        RECT 17.545 23.705 17.815 24.165 ;
        RECT 13.525 22.705 14.045 23.245 ;
        RECT 12.835 21.615 14.045 22.705 ;
        RECT 14.220 21.615 14.480 22.765 ;
        RECT 14.655 22.690 14.825 23.420 ;
        RECT 15.080 23.255 15.250 23.445 ;
        RECT 17.090 23.365 18.045 23.535 ;
        RECT 14.995 22.925 15.250 23.255 ;
        RECT 15.080 22.715 15.250 22.925 ;
        RECT 15.530 22.895 15.885 23.265 ;
        RECT 14.655 21.785 14.910 22.690 ;
        RECT 15.080 22.545 15.795 22.715 ;
        RECT 16.975 22.635 17.665 23.195 ;
        RECT 15.080 21.615 15.410 22.375 ;
        RECT 15.625 21.785 15.795 22.545 ;
        RECT 17.835 22.465 18.045 23.365 ;
        RECT 17.090 22.245 18.045 22.465 ;
        RECT 18.215 23.195 18.615 23.995 ;
        RECT 18.805 23.535 19.085 23.995 ;
        RECT 19.605 23.705 19.930 24.165 ;
        RECT 18.805 23.365 19.930 23.535 ;
        RECT 20.100 23.425 20.485 23.995 ;
        RECT 19.480 23.255 19.930 23.365 ;
        RECT 18.215 22.635 19.310 23.195 ;
        RECT 19.480 22.925 20.035 23.255 ;
        RECT 17.090 21.785 17.375 22.245 ;
        RECT 17.545 21.615 17.815 22.075 ;
        RECT 18.215 21.785 18.615 22.635 ;
        RECT 19.480 22.465 19.930 22.925 ;
        RECT 20.205 22.755 20.485 23.425 ;
        RECT 21.690 23.535 21.975 23.995 ;
        RECT 22.145 23.705 22.415 24.165 ;
        RECT 21.690 23.365 22.645 23.535 ;
        RECT 18.805 22.245 19.930 22.465 ;
        RECT 18.805 21.785 19.085 22.245 ;
        RECT 19.605 21.615 19.930 22.075 ;
        RECT 20.100 21.785 20.485 22.755 ;
        RECT 21.575 22.635 22.265 23.195 ;
        RECT 22.435 22.465 22.645 23.365 ;
        RECT 21.690 22.245 22.645 22.465 ;
        RECT 22.815 23.195 23.215 23.995 ;
        RECT 23.405 23.535 23.685 23.995 ;
        RECT 24.205 23.705 24.530 24.165 ;
        RECT 23.405 23.365 24.530 23.535 ;
        RECT 24.700 23.425 25.085 23.995 ;
        RECT 24.080 23.255 24.530 23.365 ;
        RECT 22.815 22.635 23.910 23.195 ;
        RECT 24.080 22.925 24.635 23.255 ;
        RECT 21.690 21.785 21.975 22.245 ;
        RECT 22.145 21.615 22.415 22.075 ;
        RECT 22.815 21.785 23.215 22.635 ;
        RECT 24.080 22.465 24.530 22.925 ;
        RECT 24.805 22.755 25.085 23.425 ;
        RECT 25.530 23.355 25.775 23.960 ;
        RECT 25.995 23.630 26.505 24.165 ;
        RECT 23.405 22.245 24.530 22.465 ;
        RECT 23.405 21.785 23.685 22.245 ;
        RECT 24.205 21.615 24.530 22.075 ;
        RECT 24.700 21.785 25.085 22.755 ;
        RECT 25.255 23.185 26.485 23.355 ;
        RECT 25.255 22.375 25.595 23.185 ;
        RECT 25.765 22.620 26.515 22.810 ;
        RECT 25.255 21.965 25.770 22.375 ;
        RECT 26.005 21.615 26.175 22.375 ;
        RECT 26.345 21.955 26.515 22.620 ;
        RECT 26.685 22.635 26.875 23.995 ;
        RECT 27.045 23.145 27.320 23.995 ;
        RECT 27.510 23.630 28.040 23.995 ;
        RECT 28.465 23.765 28.795 24.165 ;
        RECT 27.865 23.595 28.040 23.630 ;
        RECT 27.045 22.975 27.325 23.145 ;
        RECT 27.045 22.835 27.320 22.975 ;
        RECT 27.525 22.635 27.695 23.435 ;
        RECT 26.685 22.465 27.695 22.635 ;
        RECT 27.865 23.425 28.795 23.595 ;
        RECT 28.965 23.425 29.220 23.995 ;
        RECT 27.865 22.295 28.035 23.425 ;
        RECT 28.625 23.255 28.795 23.425 ;
        RECT 26.910 22.125 28.035 22.295 ;
        RECT 28.205 22.925 28.400 23.255 ;
        RECT 28.625 22.925 28.880 23.255 ;
        RECT 28.205 21.955 28.375 22.925 ;
        RECT 29.050 22.755 29.220 23.425 ;
        RECT 29.395 23.395 31.065 24.165 ;
        RECT 31.325 23.615 31.495 23.905 ;
        RECT 31.665 23.785 31.995 24.165 ;
        RECT 31.325 23.445 31.990 23.615 ;
        RECT 29.395 22.875 30.145 23.395 ;
        RECT 26.345 21.785 28.375 21.955 ;
        RECT 28.545 21.615 28.715 22.755 ;
        RECT 28.885 21.785 29.220 22.755 ;
        RECT 30.315 22.705 31.065 23.225 ;
        RECT 29.395 21.615 31.065 22.705 ;
        RECT 31.240 22.625 31.590 23.275 ;
        RECT 31.760 22.455 31.990 23.445 ;
        RECT 31.325 22.285 31.990 22.455 ;
        RECT 31.325 21.785 31.495 22.285 ;
        RECT 31.665 21.615 31.995 22.115 ;
        RECT 32.165 21.785 32.350 23.905 ;
        RECT 32.605 23.705 32.855 24.165 ;
        RECT 33.025 23.715 33.360 23.885 ;
        RECT 33.555 23.715 34.230 23.885 ;
        RECT 33.025 23.575 33.195 23.715 ;
        RECT 32.520 22.585 32.800 23.535 ;
        RECT 32.970 23.445 33.195 23.575 ;
        RECT 32.970 22.340 33.140 23.445 ;
        RECT 33.365 23.295 33.890 23.515 ;
        RECT 33.310 22.530 33.550 23.125 ;
        RECT 33.720 22.595 33.890 23.295 ;
        RECT 34.060 22.935 34.230 23.715 ;
        RECT 34.550 23.665 34.920 24.165 ;
        RECT 35.100 23.715 35.505 23.885 ;
        RECT 35.675 23.715 36.460 23.885 ;
        RECT 35.100 23.485 35.270 23.715 ;
        RECT 34.440 23.185 35.270 23.485 ;
        RECT 35.655 23.215 36.120 23.545 ;
        RECT 34.440 23.155 34.640 23.185 ;
        RECT 34.760 22.935 34.930 23.005 ;
        RECT 34.060 22.765 34.930 22.935 ;
        RECT 34.420 22.675 34.930 22.765 ;
        RECT 32.970 22.210 33.275 22.340 ;
        RECT 33.720 22.230 34.250 22.595 ;
        RECT 32.590 21.615 32.855 22.075 ;
        RECT 33.025 21.785 33.275 22.210 ;
        RECT 34.420 22.060 34.590 22.675 ;
        RECT 33.485 21.890 34.590 22.060 ;
        RECT 34.760 21.615 34.930 22.415 ;
        RECT 35.100 22.115 35.270 23.185 ;
        RECT 35.440 22.285 35.630 23.005 ;
        RECT 35.800 22.255 36.120 23.215 ;
        RECT 36.290 23.255 36.460 23.715 ;
        RECT 36.735 23.635 36.945 24.165 ;
        RECT 37.205 23.425 37.535 23.950 ;
        RECT 37.705 23.555 37.875 24.165 ;
        RECT 38.045 23.510 38.375 23.945 ;
        RECT 38.045 23.425 38.425 23.510 ;
        RECT 38.595 23.440 38.885 24.165 ;
        RECT 37.335 23.255 37.535 23.425 ;
        RECT 38.200 23.385 38.425 23.425 ;
        RECT 36.290 22.925 37.165 23.255 ;
        RECT 37.335 22.925 38.085 23.255 ;
        RECT 35.100 21.785 35.350 22.115 ;
        RECT 36.290 22.085 36.460 22.925 ;
        RECT 37.335 22.720 37.525 22.925 ;
        RECT 38.255 22.805 38.425 23.385 ;
        RECT 38.210 22.755 38.425 22.805 ;
        RECT 39.060 23.425 39.315 23.995 ;
        RECT 39.485 23.765 39.815 24.165 ;
        RECT 40.240 23.630 40.770 23.995 ;
        RECT 40.960 23.825 41.235 23.995 ;
        RECT 40.955 23.655 41.235 23.825 ;
        RECT 40.240 23.595 40.415 23.630 ;
        RECT 39.485 23.425 40.415 23.595 ;
        RECT 36.630 22.345 37.525 22.720 ;
        RECT 38.035 22.675 38.425 22.755 ;
        RECT 35.575 21.915 36.460 22.085 ;
        RECT 36.640 21.615 36.955 22.115 ;
        RECT 37.185 21.785 37.525 22.345 ;
        RECT 37.695 21.615 37.865 22.625 ;
        RECT 38.035 21.830 38.365 22.675 ;
        RECT 38.595 21.615 38.885 22.780 ;
        RECT 39.060 22.755 39.230 23.425 ;
        RECT 39.485 23.255 39.655 23.425 ;
        RECT 39.400 22.925 39.655 23.255 ;
        RECT 39.880 22.925 40.075 23.255 ;
        RECT 39.060 21.785 39.395 22.755 ;
        RECT 39.565 21.615 39.735 22.755 ;
        RECT 39.905 21.955 40.075 22.925 ;
        RECT 40.245 22.295 40.415 23.425 ;
        RECT 40.585 22.635 40.755 23.435 ;
        RECT 40.960 22.835 41.235 23.655 ;
        RECT 41.405 22.635 41.595 23.995 ;
        RECT 41.775 23.630 42.285 24.165 ;
        RECT 42.505 23.355 42.750 23.960 ;
        RECT 43.285 23.615 43.455 23.995 ;
        RECT 43.635 23.785 43.965 24.165 ;
        RECT 43.285 23.445 43.950 23.615 ;
        RECT 44.145 23.490 44.405 23.995 ;
        RECT 41.795 23.185 43.025 23.355 ;
        RECT 40.585 22.465 41.595 22.635 ;
        RECT 41.765 22.620 42.515 22.810 ;
        RECT 40.245 22.125 41.370 22.295 ;
        RECT 41.765 21.955 41.935 22.620 ;
        RECT 42.685 22.375 43.025 23.185 ;
        RECT 43.215 22.895 43.545 23.265 ;
        RECT 43.780 23.190 43.950 23.445 ;
        RECT 43.780 22.860 44.065 23.190 ;
        RECT 43.780 22.715 43.950 22.860 ;
        RECT 39.905 21.785 41.935 21.955 ;
        RECT 42.105 21.615 42.275 22.375 ;
        RECT 42.510 21.965 43.025 22.375 ;
        RECT 43.285 22.545 43.950 22.715 ;
        RECT 44.235 22.690 44.405 23.490 ;
        RECT 43.285 21.785 43.455 22.545 ;
        RECT 43.635 21.615 43.965 22.375 ;
        RECT 44.135 21.785 44.405 22.690 ;
        RECT 44.575 23.490 44.845 23.835 ;
        RECT 45.035 23.765 45.415 24.165 ;
        RECT 45.585 23.595 45.755 23.945 ;
        RECT 45.925 23.765 46.255 24.165 ;
        RECT 46.455 23.595 46.625 23.945 ;
        RECT 46.825 23.665 47.155 24.165 ;
        RECT 44.575 22.755 44.745 23.490 ;
        RECT 45.015 23.425 46.625 23.595 ;
        RECT 45.015 23.255 45.185 23.425 ;
        RECT 44.915 22.925 45.185 23.255 ;
        RECT 45.355 22.925 45.760 23.255 ;
        RECT 45.015 22.755 45.185 22.925 ;
        RECT 44.575 21.785 44.845 22.755 ;
        RECT 45.015 22.585 45.740 22.755 ;
        RECT 45.930 22.635 46.640 23.255 ;
        RECT 46.810 22.925 47.160 23.495 ;
        RECT 47.335 23.415 48.545 24.165 ;
        RECT 45.570 22.465 45.740 22.585 ;
        RECT 46.840 22.465 47.160 22.755 ;
        RECT 45.055 21.615 45.335 22.415 ;
        RECT 45.570 22.295 47.160 22.465 ;
        RECT 47.335 22.705 47.855 23.245 ;
        RECT 48.025 22.875 48.545 23.415 ;
        RECT 45.505 21.835 47.160 22.125 ;
        RECT 47.335 21.615 48.545 22.705 ;
        RECT 12.750 21.445 48.630 21.615 ;
        RECT 12.835 20.355 14.045 21.445 ;
        RECT 14.275 20.385 14.605 21.230 ;
        RECT 14.775 20.435 14.945 21.445 ;
        RECT 15.115 20.715 15.455 21.275 ;
        RECT 15.685 20.945 16.000 21.445 ;
        RECT 16.180 20.975 17.065 21.145 ;
        RECT 12.835 19.645 13.355 20.185 ;
        RECT 13.525 19.815 14.045 20.355 ;
        RECT 14.215 20.305 14.605 20.385 ;
        RECT 15.115 20.340 16.010 20.715 ;
        RECT 14.215 20.255 14.430 20.305 ;
        RECT 14.215 19.675 14.385 20.255 ;
        RECT 15.115 20.135 15.305 20.340 ;
        RECT 16.180 20.135 16.350 20.975 ;
        RECT 17.290 20.945 17.540 21.275 ;
        RECT 14.555 19.805 15.305 20.135 ;
        RECT 15.475 19.805 16.350 20.135 ;
        RECT 12.835 18.895 14.045 19.645 ;
        RECT 14.215 19.635 14.440 19.675 ;
        RECT 15.105 19.635 15.305 19.805 ;
        RECT 14.215 19.550 14.595 19.635 ;
        RECT 14.265 19.115 14.595 19.550 ;
        RECT 14.765 18.895 14.935 19.505 ;
        RECT 15.105 19.110 15.435 19.635 ;
        RECT 15.695 18.895 15.905 19.425 ;
        RECT 16.180 19.345 16.350 19.805 ;
        RECT 16.520 19.845 16.840 20.805 ;
        RECT 17.010 20.055 17.200 20.775 ;
        RECT 17.370 19.875 17.540 20.945 ;
        RECT 17.710 20.645 17.880 21.445 ;
        RECT 18.050 21.000 19.155 21.170 ;
        RECT 18.050 20.385 18.220 21.000 ;
        RECT 19.365 20.850 19.615 21.275 ;
        RECT 19.785 20.985 20.050 21.445 ;
        RECT 18.390 20.465 18.920 20.830 ;
        RECT 19.365 20.720 19.670 20.850 ;
        RECT 17.710 20.295 18.220 20.385 ;
        RECT 17.710 20.125 18.580 20.295 ;
        RECT 17.710 20.055 17.880 20.125 ;
        RECT 18.000 19.875 18.200 19.905 ;
        RECT 16.520 19.515 16.985 19.845 ;
        RECT 17.370 19.575 18.200 19.875 ;
        RECT 17.370 19.345 17.540 19.575 ;
        RECT 16.180 19.175 16.965 19.345 ;
        RECT 17.135 19.175 17.540 19.345 ;
        RECT 17.720 18.895 18.090 19.395 ;
        RECT 18.410 19.345 18.580 20.125 ;
        RECT 18.750 19.765 18.920 20.465 ;
        RECT 19.090 19.935 19.330 20.530 ;
        RECT 18.750 19.545 19.275 19.765 ;
        RECT 19.500 19.615 19.670 20.720 ;
        RECT 19.445 19.485 19.670 19.615 ;
        RECT 19.840 19.525 20.120 20.475 ;
        RECT 19.445 19.345 19.615 19.485 ;
        RECT 18.410 19.175 19.085 19.345 ;
        RECT 19.280 19.175 19.615 19.345 ;
        RECT 19.785 18.895 20.035 19.355 ;
        RECT 20.290 19.155 20.475 21.275 ;
        RECT 20.645 20.945 20.975 21.445 ;
        RECT 21.145 20.775 21.315 21.275 ;
        RECT 20.650 20.605 21.315 20.775 ;
        RECT 20.650 19.615 20.880 20.605 ;
        RECT 21.050 19.785 21.400 20.435 ;
        RECT 21.575 20.355 25.085 21.445 ;
        RECT 21.575 19.665 23.225 20.185 ;
        RECT 23.395 19.835 25.085 20.355 ;
        RECT 25.715 20.280 26.005 21.445 ;
        RECT 26.185 20.635 26.480 21.445 ;
        RECT 26.660 20.135 26.905 21.275 ;
        RECT 27.080 20.635 27.340 21.445 ;
        RECT 27.940 21.440 34.215 21.445 ;
        RECT 27.520 20.135 27.770 21.270 ;
        RECT 27.940 20.645 28.200 21.440 ;
        RECT 28.370 20.545 28.630 21.270 ;
        RECT 28.800 20.715 29.060 21.440 ;
        RECT 29.230 20.545 29.490 21.270 ;
        RECT 29.660 20.715 29.920 21.440 ;
        RECT 30.090 20.545 30.350 21.270 ;
        RECT 30.520 20.715 30.780 21.440 ;
        RECT 30.950 20.545 31.210 21.270 ;
        RECT 31.380 20.715 31.625 21.440 ;
        RECT 31.795 20.545 32.055 21.270 ;
        RECT 32.240 20.715 32.485 21.440 ;
        RECT 32.655 20.545 32.915 21.270 ;
        RECT 33.100 20.715 33.345 21.440 ;
        RECT 33.515 20.545 33.775 21.270 ;
        RECT 33.960 20.715 34.215 21.440 ;
        RECT 28.370 20.530 33.775 20.545 ;
        RECT 34.385 20.530 34.675 21.270 ;
        RECT 34.845 20.700 35.115 21.445 ;
        RECT 28.370 20.305 35.115 20.530 ;
        RECT 35.375 20.355 36.585 21.445 ;
        RECT 20.650 19.445 21.315 19.615 ;
        RECT 20.645 18.895 20.975 19.275 ;
        RECT 21.145 19.155 21.315 19.445 ;
        RECT 21.575 18.895 25.085 19.665 ;
        RECT 25.715 18.895 26.005 19.620 ;
        RECT 26.175 19.575 26.490 20.135 ;
        RECT 26.660 19.885 33.780 20.135 ;
        RECT 26.175 18.895 26.480 19.405 ;
        RECT 26.660 19.075 26.910 19.885 ;
        RECT 27.080 18.895 27.340 19.420 ;
        RECT 27.520 19.075 27.770 19.885 ;
        RECT 33.950 19.715 35.115 20.305 ;
        RECT 28.370 19.545 35.115 19.715 ;
        RECT 35.375 19.645 35.895 20.185 ;
        RECT 36.065 19.815 36.585 20.355 ;
        RECT 36.845 20.515 37.015 21.275 ;
        RECT 37.195 20.685 37.525 21.445 ;
        RECT 36.845 20.345 37.510 20.515 ;
        RECT 37.695 20.370 37.965 21.275 ;
        RECT 37.340 20.200 37.510 20.345 ;
        RECT 36.775 19.795 37.105 20.165 ;
        RECT 37.340 19.870 37.625 20.200 ;
        RECT 27.940 18.895 28.200 19.455 ;
        RECT 28.370 19.090 28.630 19.545 ;
        RECT 28.800 18.895 29.060 19.375 ;
        RECT 29.230 19.090 29.490 19.545 ;
        RECT 29.660 18.895 29.920 19.375 ;
        RECT 30.090 19.090 30.350 19.545 ;
        RECT 30.520 18.895 30.765 19.375 ;
        RECT 30.935 19.090 31.210 19.545 ;
        RECT 31.380 18.895 31.625 19.375 ;
        RECT 31.795 19.090 32.055 19.545 ;
        RECT 32.235 18.895 32.485 19.375 ;
        RECT 32.655 19.090 32.915 19.545 ;
        RECT 33.095 18.895 33.345 19.375 ;
        RECT 33.515 19.090 33.775 19.545 ;
        RECT 33.955 18.895 34.215 19.375 ;
        RECT 34.385 19.090 34.645 19.545 ;
        RECT 34.815 18.895 35.115 19.375 ;
        RECT 35.375 18.895 36.585 19.645 ;
        RECT 37.340 19.615 37.510 19.870 ;
        RECT 36.845 19.445 37.510 19.615 ;
        RECT 37.795 19.570 37.965 20.370 ;
        RECT 38.225 20.515 38.395 21.275 ;
        RECT 38.575 20.685 38.905 21.445 ;
        RECT 38.225 20.345 38.890 20.515 ;
        RECT 39.075 20.370 39.345 21.275 ;
        RECT 38.720 20.200 38.890 20.345 ;
        RECT 38.155 19.795 38.485 20.165 ;
        RECT 38.720 19.870 39.005 20.200 ;
        RECT 38.720 19.615 38.890 19.870 ;
        RECT 36.845 19.065 37.015 19.445 ;
        RECT 37.195 18.895 37.525 19.275 ;
        RECT 37.705 19.065 37.965 19.570 ;
        RECT 38.225 19.445 38.890 19.615 ;
        RECT 39.175 19.570 39.345 20.370 ;
        RECT 39.605 20.515 39.775 21.275 ;
        RECT 39.955 20.685 40.285 21.445 ;
        RECT 39.605 20.345 40.270 20.515 ;
        RECT 40.455 20.370 40.725 21.275 ;
        RECT 40.100 20.200 40.270 20.345 ;
        RECT 39.535 19.795 39.865 20.165 ;
        RECT 40.100 19.870 40.385 20.200 ;
        RECT 40.100 19.615 40.270 19.870 ;
        RECT 38.225 19.065 38.395 19.445 ;
        RECT 38.575 18.895 38.905 19.275 ;
        RECT 39.085 19.065 39.345 19.570 ;
        RECT 39.605 19.445 40.270 19.615 ;
        RECT 40.555 19.570 40.725 20.370 ;
        RECT 40.985 20.515 41.155 21.275 ;
        RECT 41.335 20.685 41.665 21.445 ;
        RECT 40.985 20.345 41.650 20.515 ;
        RECT 41.835 20.370 42.105 21.275 ;
        RECT 41.480 20.200 41.650 20.345 ;
        RECT 40.915 19.795 41.245 20.165 ;
        RECT 41.480 19.870 41.765 20.200 ;
        RECT 41.480 19.615 41.650 19.870 ;
        RECT 39.605 19.065 39.775 19.445 ;
        RECT 39.955 18.895 40.285 19.275 ;
        RECT 40.465 19.065 40.725 19.570 ;
        RECT 40.985 19.445 41.650 19.615 ;
        RECT 41.935 19.570 42.105 20.370 ;
        RECT 42.285 20.305 42.615 21.445 ;
        RECT 43.145 20.475 43.475 21.260 ;
        RECT 42.795 20.305 43.475 20.475 ;
        RECT 42.275 19.885 42.625 20.135 ;
        RECT 42.795 19.705 42.965 20.305 ;
        RECT 43.655 20.290 43.995 21.275 ;
        RECT 44.165 21.015 44.575 21.445 ;
        RECT 45.320 21.025 45.650 21.445 ;
        RECT 45.820 20.845 46.145 21.275 ;
        RECT 44.165 20.675 46.145 20.845 ;
        RECT 43.135 19.885 43.485 20.135 ;
        RECT 40.985 19.065 41.155 19.445 ;
        RECT 41.335 18.895 41.665 19.275 ;
        RECT 41.845 19.065 42.105 19.570 ;
        RECT 42.285 18.895 42.555 19.705 ;
        RECT 42.725 19.065 43.055 19.705 ;
        RECT 43.225 18.895 43.465 19.705 ;
        RECT 43.655 19.635 43.910 20.290 ;
        RECT 44.165 20.135 44.430 20.675 ;
        RECT 44.645 20.335 45.270 20.505 ;
        RECT 44.080 19.805 44.430 20.135 ;
        RECT 44.600 19.805 44.930 20.135 ;
        RECT 45.100 19.635 45.270 20.335 ;
        RECT 43.655 19.260 44.015 19.635 ;
        RECT 44.280 18.895 44.450 19.635 ;
        RECT 44.730 19.465 45.270 19.635 ;
        RECT 45.440 20.265 46.145 20.675 ;
        RECT 46.620 20.345 46.950 21.445 ;
        RECT 47.335 20.355 48.545 21.445 ;
        RECT 44.730 19.260 44.900 19.465 ;
        RECT 45.440 19.065 45.610 20.265 ;
        RECT 45.780 19.885 46.350 20.095 ;
        RECT 46.520 19.885 47.165 20.095 ;
        RECT 47.335 19.815 47.855 20.355 ;
        RECT 45.840 19.545 47.010 19.715 ;
        RECT 48.025 19.645 48.545 20.185 ;
        RECT 45.840 19.065 46.170 19.545 ;
        RECT 46.340 18.895 46.510 19.365 ;
        RECT 46.680 19.080 47.010 19.545 ;
        RECT 47.335 18.895 48.545 19.645 ;
        RECT 12.750 18.725 48.630 18.895 ;
        RECT 12.835 17.975 14.045 18.725 ;
        RECT 12.835 17.435 13.355 17.975 ;
        RECT 14.220 17.885 14.480 18.725 ;
        RECT 14.655 17.980 14.910 18.555 ;
        RECT 15.080 18.345 15.410 18.725 ;
        RECT 15.625 18.175 15.795 18.555 ;
        RECT 15.080 18.005 15.795 18.175 ;
        RECT 13.525 17.265 14.045 17.805 ;
        RECT 12.835 16.175 14.045 17.265 ;
        RECT 14.220 16.175 14.480 17.325 ;
        RECT 14.655 17.250 14.825 17.980 ;
        RECT 15.080 17.815 15.250 18.005 ;
        RECT 16.980 17.985 17.235 18.555 ;
        RECT 17.405 18.325 17.735 18.725 ;
        RECT 18.160 18.190 18.690 18.555 ;
        RECT 18.880 18.385 19.155 18.555 ;
        RECT 18.875 18.215 19.155 18.385 ;
        RECT 18.160 18.155 18.335 18.190 ;
        RECT 17.405 17.985 18.335 18.155 ;
        RECT 14.995 17.485 15.250 17.815 ;
        RECT 15.080 17.275 15.250 17.485 ;
        RECT 15.530 17.455 15.885 17.825 ;
        RECT 16.980 17.315 17.150 17.985 ;
        RECT 17.405 17.815 17.575 17.985 ;
        RECT 17.320 17.485 17.575 17.815 ;
        RECT 17.800 17.485 17.995 17.815 ;
        RECT 14.655 16.345 14.910 17.250 ;
        RECT 15.080 17.105 15.795 17.275 ;
        RECT 15.080 16.175 15.410 16.935 ;
        RECT 15.625 16.345 15.795 17.105 ;
        RECT 16.980 16.345 17.315 17.315 ;
        RECT 17.485 16.175 17.655 17.315 ;
        RECT 17.825 16.515 17.995 17.485 ;
        RECT 18.165 16.855 18.335 17.985 ;
        RECT 18.505 17.195 18.675 17.995 ;
        RECT 18.880 17.395 19.155 18.215 ;
        RECT 19.325 17.195 19.515 18.555 ;
        RECT 19.695 18.190 20.205 18.725 ;
        RECT 20.425 17.915 20.670 18.520 ;
        RECT 21.115 17.955 24.625 18.725 ;
        RECT 24.795 17.975 26.005 18.725 ;
        RECT 26.225 18.070 26.555 18.505 ;
        RECT 26.725 18.115 26.895 18.725 ;
        RECT 26.175 17.985 26.555 18.070 ;
        RECT 27.065 17.985 27.395 18.510 ;
        RECT 27.655 18.195 27.865 18.725 ;
        RECT 28.140 18.275 28.925 18.445 ;
        RECT 29.095 18.275 29.500 18.445 ;
        RECT 19.715 17.745 20.945 17.915 ;
        RECT 18.505 17.025 19.515 17.195 ;
        RECT 19.685 17.180 20.435 17.370 ;
        RECT 18.165 16.685 19.290 16.855 ;
        RECT 19.685 16.515 19.855 17.180 ;
        RECT 20.605 16.935 20.945 17.745 ;
        RECT 21.115 17.435 22.765 17.955 ;
        RECT 22.935 17.265 24.625 17.785 ;
        RECT 24.795 17.435 25.315 17.975 ;
        RECT 26.175 17.945 26.400 17.985 ;
        RECT 25.485 17.265 26.005 17.805 ;
        RECT 17.825 16.345 19.855 16.515 ;
        RECT 20.025 16.175 20.195 16.935 ;
        RECT 20.430 16.525 20.945 16.935 ;
        RECT 21.115 16.175 24.625 17.265 ;
        RECT 24.795 16.175 26.005 17.265 ;
        RECT 26.175 17.365 26.345 17.945 ;
        RECT 27.065 17.815 27.265 17.985 ;
        RECT 28.140 17.815 28.310 18.275 ;
        RECT 26.515 17.485 27.265 17.815 ;
        RECT 27.435 17.485 28.310 17.815 ;
        RECT 26.175 17.315 26.390 17.365 ;
        RECT 26.175 17.235 26.565 17.315 ;
        RECT 26.235 16.390 26.565 17.235 ;
        RECT 27.075 17.280 27.265 17.485 ;
        RECT 26.735 16.175 26.905 17.185 ;
        RECT 27.075 16.905 27.970 17.280 ;
        RECT 27.075 16.345 27.415 16.905 ;
        RECT 27.645 16.175 27.960 16.675 ;
        RECT 28.140 16.645 28.310 17.485 ;
        RECT 28.480 17.775 28.945 18.105 ;
        RECT 29.330 18.045 29.500 18.275 ;
        RECT 29.680 18.225 30.050 18.725 ;
        RECT 30.370 18.275 31.045 18.445 ;
        RECT 31.240 18.275 31.575 18.445 ;
        RECT 28.480 16.815 28.800 17.775 ;
        RECT 29.330 17.745 30.160 18.045 ;
        RECT 28.970 16.845 29.160 17.565 ;
        RECT 29.330 16.675 29.500 17.745 ;
        RECT 29.960 17.715 30.160 17.745 ;
        RECT 29.670 17.495 29.840 17.565 ;
        RECT 30.370 17.495 30.540 18.275 ;
        RECT 31.405 18.135 31.575 18.275 ;
        RECT 31.745 18.265 31.995 18.725 ;
        RECT 29.670 17.325 30.540 17.495 ;
        RECT 30.710 17.855 31.235 18.075 ;
        RECT 31.405 18.005 31.630 18.135 ;
        RECT 29.670 17.235 30.180 17.325 ;
        RECT 28.140 16.475 29.025 16.645 ;
        RECT 29.250 16.345 29.500 16.675 ;
        RECT 29.670 16.175 29.840 16.975 ;
        RECT 30.010 16.620 30.180 17.235 ;
        RECT 30.710 17.155 30.880 17.855 ;
        RECT 30.350 16.790 30.880 17.155 ;
        RECT 31.050 17.090 31.290 17.685 ;
        RECT 31.460 16.900 31.630 18.005 ;
        RECT 31.800 17.145 32.080 18.095 ;
        RECT 31.325 16.770 31.630 16.900 ;
        RECT 30.010 16.450 31.115 16.620 ;
        RECT 31.325 16.345 31.575 16.770 ;
        RECT 31.745 16.175 32.010 16.635 ;
        RECT 32.250 16.345 32.435 18.465 ;
        RECT 32.605 18.345 32.935 18.725 ;
        RECT 33.105 18.175 33.275 18.465 ;
        RECT 32.610 18.005 33.275 18.175 ;
        RECT 32.610 17.015 32.840 18.005 ;
        RECT 33.540 17.985 33.795 18.555 ;
        RECT 33.965 18.325 34.295 18.725 ;
        RECT 34.720 18.190 35.250 18.555 ;
        RECT 34.720 18.155 34.895 18.190 ;
        RECT 33.965 17.985 34.895 18.155 ;
        RECT 33.010 17.185 33.360 17.835 ;
        RECT 33.540 17.315 33.710 17.985 ;
        RECT 33.965 17.815 34.135 17.985 ;
        RECT 33.880 17.485 34.135 17.815 ;
        RECT 34.360 17.485 34.555 17.815 ;
        RECT 32.610 16.845 33.275 17.015 ;
        RECT 32.605 16.175 32.935 16.675 ;
        RECT 33.105 16.345 33.275 16.845 ;
        RECT 33.540 16.345 33.875 17.315 ;
        RECT 34.045 16.175 34.215 17.315 ;
        RECT 34.385 16.515 34.555 17.485 ;
        RECT 34.725 16.855 34.895 17.985 ;
        RECT 35.065 17.195 35.235 17.995 ;
        RECT 35.440 17.705 35.715 18.555 ;
        RECT 35.435 17.535 35.715 17.705 ;
        RECT 35.440 17.395 35.715 17.535 ;
        RECT 35.885 17.195 36.075 18.555 ;
        RECT 36.255 18.190 36.765 18.725 ;
        RECT 36.985 17.915 37.230 18.520 ;
        RECT 38.595 18.000 38.885 18.725 ;
        RECT 39.055 17.985 39.440 18.555 ;
        RECT 39.610 18.265 39.935 18.725 ;
        RECT 40.455 18.095 40.735 18.555 ;
        RECT 36.275 17.745 37.505 17.915 ;
        RECT 35.065 17.025 36.075 17.195 ;
        RECT 36.245 17.180 36.995 17.370 ;
        RECT 34.725 16.685 35.850 16.855 ;
        RECT 36.245 16.515 36.415 17.180 ;
        RECT 37.165 16.935 37.505 17.745 ;
        RECT 34.385 16.345 36.415 16.515 ;
        RECT 36.585 16.175 36.755 16.935 ;
        RECT 36.990 16.525 37.505 16.935 ;
        RECT 38.595 16.175 38.885 17.340 ;
        RECT 39.055 17.315 39.335 17.985 ;
        RECT 39.610 17.925 40.735 18.095 ;
        RECT 39.610 17.815 40.060 17.925 ;
        RECT 39.505 17.485 40.060 17.815 ;
        RECT 40.925 17.755 41.325 18.555 ;
        RECT 41.725 18.265 41.995 18.725 ;
        RECT 42.165 18.095 42.450 18.555 ;
        RECT 39.055 16.345 39.440 17.315 ;
        RECT 39.610 17.025 40.060 17.485 ;
        RECT 40.230 17.195 41.325 17.755 ;
        RECT 39.610 16.805 40.735 17.025 ;
        RECT 39.610 16.175 39.935 16.635 ;
        RECT 40.455 16.345 40.735 16.805 ;
        RECT 40.925 16.345 41.325 17.195 ;
        RECT 41.495 17.925 42.450 18.095 ;
        RECT 43.655 18.095 43.995 18.555 ;
        RECT 44.165 18.265 44.335 18.725 ;
        RECT 44.965 18.290 45.325 18.555 ;
        RECT 44.970 18.285 45.325 18.290 ;
        RECT 44.975 18.275 45.325 18.285 ;
        RECT 44.980 18.270 45.325 18.275 ;
        RECT 44.985 18.260 45.325 18.270 ;
        RECT 45.565 18.265 45.735 18.725 ;
        RECT 44.990 18.255 45.325 18.260 ;
        RECT 45.000 18.245 45.325 18.255 ;
        RECT 45.010 18.235 45.325 18.245 ;
        RECT 44.505 18.095 44.835 18.175 ;
        RECT 41.495 17.025 41.705 17.925 ;
        RECT 43.655 17.905 44.835 18.095 ;
        RECT 45.025 18.095 45.325 18.235 ;
        RECT 45.025 17.905 45.735 18.095 ;
        RECT 41.875 17.195 42.565 17.755 ;
        RECT 43.655 17.535 43.985 17.735 ;
        RECT 44.295 17.715 44.625 17.735 ;
        RECT 44.175 17.535 44.625 17.715 ;
        RECT 43.655 17.195 43.885 17.535 ;
        RECT 41.495 16.805 42.450 17.025 ;
        RECT 41.725 16.175 41.995 16.635 ;
        RECT 42.165 16.345 42.450 16.805 ;
        RECT 43.665 16.175 43.995 16.895 ;
        RECT 44.175 16.420 44.390 17.535 ;
        RECT 44.795 17.505 45.265 17.735 ;
        RECT 45.450 17.335 45.735 17.905 ;
        RECT 45.905 17.780 46.245 18.555 ;
        RECT 47.335 17.975 48.545 18.725 ;
        RECT 44.585 17.120 45.735 17.335 ;
        RECT 44.585 16.345 44.915 17.120 ;
        RECT 45.085 16.175 45.795 16.950 ;
        RECT 45.965 16.345 46.245 17.780 ;
        RECT 47.335 17.265 47.855 17.805 ;
        RECT 48.025 17.435 48.545 17.975 ;
        RECT 47.335 16.175 48.545 17.265 ;
        RECT 12.750 16.005 48.630 16.175 ;
        RECT 12.835 14.915 14.045 16.005 ;
        RECT 14.215 15.570 19.560 16.005 ;
        RECT 12.835 14.205 13.355 14.745 ;
        RECT 13.525 14.375 14.045 14.915 ;
        RECT 12.835 13.455 14.045 14.205 ;
        RECT 15.800 14.000 16.140 14.830 ;
        RECT 17.620 14.320 17.970 15.570 ;
        RECT 19.735 14.915 23.245 16.005 ;
        RECT 19.735 14.225 21.385 14.745 ;
        RECT 21.555 14.395 23.245 14.915 ;
        RECT 23.965 15.075 24.135 15.835 ;
        RECT 24.350 15.245 24.680 16.005 ;
        RECT 23.965 14.905 24.680 15.075 ;
        RECT 24.850 14.930 25.105 15.835 ;
        RECT 23.875 14.355 24.230 14.725 ;
        RECT 24.510 14.695 24.680 14.905 ;
        RECT 24.510 14.365 24.765 14.695 ;
        RECT 14.215 13.455 19.560 14.000 ;
        RECT 19.735 13.455 23.245 14.225 ;
        RECT 24.510 14.175 24.680 14.365 ;
        RECT 24.935 14.200 25.105 14.930 ;
        RECT 25.280 14.855 25.540 16.005 ;
        RECT 25.715 14.840 26.005 16.005 ;
        RECT 26.640 14.855 26.900 16.005 ;
        RECT 27.075 14.930 27.330 15.835 ;
        RECT 27.500 15.245 27.830 16.005 ;
        RECT 28.045 15.075 28.215 15.835 ;
        RECT 28.565 15.335 28.735 15.835 ;
        RECT 28.905 15.505 29.235 16.005 ;
        RECT 28.565 15.165 29.230 15.335 ;
        RECT 23.965 14.005 24.680 14.175 ;
        RECT 23.965 13.625 24.135 14.005 ;
        RECT 24.350 13.455 24.680 13.835 ;
        RECT 24.850 13.625 25.105 14.200 ;
        RECT 25.280 13.455 25.540 14.295 ;
        RECT 25.715 13.455 26.005 14.180 ;
        RECT 26.640 13.455 26.900 14.295 ;
        RECT 27.075 14.200 27.245 14.930 ;
        RECT 27.500 14.905 28.215 15.075 ;
        RECT 27.500 14.695 27.670 14.905 ;
        RECT 27.415 14.365 27.670 14.695 ;
        RECT 27.075 13.625 27.330 14.200 ;
        RECT 27.500 14.175 27.670 14.365 ;
        RECT 27.950 14.355 28.305 14.725 ;
        RECT 28.480 14.345 28.830 14.995 ;
        RECT 29.000 14.175 29.230 15.165 ;
        RECT 27.500 14.005 28.215 14.175 ;
        RECT 27.500 13.455 27.830 13.835 ;
        RECT 28.045 13.625 28.215 14.005 ;
        RECT 28.565 14.005 29.230 14.175 ;
        RECT 28.565 13.715 28.735 14.005 ;
        RECT 28.905 13.455 29.235 13.835 ;
        RECT 29.405 13.715 29.590 15.835 ;
        RECT 29.830 15.545 30.095 16.005 ;
        RECT 30.265 15.410 30.515 15.835 ;
        RECT 30.725 15.560 31.830 15.730 ;
        RECT 30.210 15.280 30.515 15.410 ;
        RECT 29.760 14.085 30.040 15.035 ;
        RECT 30.210 14.175 30.380 15.280 ;
        RECT 30.550 14.495 30.790 15.090 ;
        RECT 30.960 15.025 31.490 15.390 ;
        RECT 30.960 14.325 31.130 15.025 ;
        RECT 31.660 14.945 31.830 15.560 ;
        RECT 32.000 15.205 32.170 16.005 ;
        RECT 32.340 15.505 32.590 15.835 ;
        RECT 32.815 15.535 33.700 15.705 ;
        RECT 31.660 14.855 32.170 14.945 ;
        RECT 30.210 14.045 30.435 14.175 ;
        RECT 30.605 14.105 31.130 14.325 ;
        RECT 31.300 14.685 32.170 14.855 ;
        RECT 29.845 13.455 30.095 13.915 ;
        RECT 30.265 13.905 30.435 14.045 ;
        RECT 31.300 13.905 31.470 14.685 ;
        RECT 32.000 14.615 32.170 14.685 ;
        RECT 31.680 14.435 31.880 14.465 ;
        RECT 32.340 14.435 32.510 15.505 ;
        RECT 32.680 14.615 32.870 15.335 ;
        RECT 31.680 14.135 32.510 14.435 ;
        RECT 33.040 14.405 33.360 15.365 ;
        RECT 30.265 13.735 30.600 13.905 ;
        RECT 30.795 13.735 31.470 13.905 ;
        RECT 31.790 13.455 32.160 13.955 ;
        RECT 32.340 13.905 32.510 14.135 ;
        RECT 32.895 14.075 33.360 14.405 ;
        RECT 33.530 14.695 33.700 15.535 ;
        RECT 33.880 15.505 34.195 16.005 ;
        RECT 34.425 15.275 34.765 15.835 ;
        RECT 33.870 14.900 34.765 15.275 ;
        RECT 34.935 14.995 35.105 16.005 ;
        RECT 34.575 14.695 34.765 14.900 ;
        RECT 35.275 14.945 35.605 15.790 ;
        RECT 35.275 14.865 35.665 14.945 ;
        RECT 35.450 14.815 35.665 14.865 ;
        RECT 35.840 14.855 36.100 16.005 ;
        RECT 36.275 14.930 36.530 15.835 ;
        RECT 36.700 15.245 37.030 16.005 ;
        RECT 37.245 15.075 37.415 15.835 ;
        RECT 33.530 14.365 34.405 14.695 ;
        RECT 34.575 14.365 35.325 14.695 ;
        RECT 33.530 13.905 33.700 14.365 ;
        RECT 34.575 14.195 34.775 14.365 ;
        RECT 35.495 14.235 35.665 14.815 ;
        RECT 35.440 14.195 35.665 14.235 ;
        RECT 32.340 13.735 32.745 13.905 ;
        RECT 32.915 13.735 33.700 13.905 ;
        RECT 33.975 13.455 34.185 13.985 ;
        RECT 34.445 13.670 34.775 14.195 ;
        RECT 35.285 14.110 35.665 14.195 ;
        RECT 34.945 13.455 35.115 14.065 ;
        RECT 35.285 13.675 35.615 14.110 ;
        RECT 35.840 13.455 36.100 14.295 ;
        RECT 36.275 14.200 36.445 14.930 ;
        RECT 36.700 14.905 37.415 15.075 ;
        RECT 36.700 14.695 36.870 14.905 ;
        RECT 38.595 14.840 38.885 16.005 ;
        RECT 40.065 15.075 40.235 15.835 ;
        RECT 40.450 15.245 40.780 16.005 ;
        RECT 40.065 14.905 40.780 15.075 ;
        RECT 40.950 14.930 41.205 15.835 ;
        RECT 36.615 14.365 36.870 14.695 ;
        RECT 36.275 13.625 36.530 14.200 ;
        RECT 36.700 14.175 36.870 14.365 ;
        RECT 37.150 14.355 37.505 14.725 ;
        RECT 39.975 14.355 40.330 14.725 ;
        RECT 40.610 14.695 40.780 14.905 ;
        RECT 40.610 14.365 40.865 14.695 ;
        RECT 36.700 14.005 37.415 14.175 ;
        RECT 36.700 13.455 37.030 13.835 ;
        RECT 37.245 13.625 37.415 14.005 ;
        RECT 38.595 13.455 38.885 14.180 ;
        RECT 40.610 14.175 40.780 14.365 ;
        RECT 41.035 14.200 41.205 14.930 ;
        RECT 41.380 14.855 41.640 16.005 ;
        RECT 41.815 14.930 42.085 15.835 ;
        RECT 42.255 15.245 42.585 16.005 ;
        RECT 42.765 15.075 42.945 15.835 ;
        RECT 44.205 15.385 44.375 15.815 ;
        RECT 44.545 15.555 44.875 16.005 ;
        RECT 44.205 15.155 44.880 15.385 ;
        RECT 40.065 14.005 40.780 14.175 ;
        RECT 40.065 13.625 40.235 14.005 ;
        RECT 40.450 13.455 40.780 13.835 ;
        RECT 40.950 13.625 41.205 14.200 ;
        RECT 41.380 13.455 41.640 14.295 ;
        RECT 41.815 14.130 41.995 14.930 ;
        RECT 42.270 14.905 42.945 15.075 ;
        RECT 42.270 14.760 42.440 14.905 ;
        RECT 42.165 14.430 42.440 14.760 ;
        RECT 42.270 14.175 42.440 14.430 ;
        RECT 42.665 14.355 43.005 14.725 ;
        RECT 41.815 13.625 42.075 14.130 ;
        RECT 42.270 14.005 42.935 14.175 ;
        RECT 44.175 14.135 44.475 14.985 ;
        RECT 44.645 14.505 44.880 15.155 ;
        RECT 45.050 14.845 45.335 15.790 ;
        RECT 45.515 15.535 46.200 16.005 ;
        RECT 45.510 15.015 46.205 15.325 ;
        RECT 46.380 14.950 46.685 15.735 ;
        RECT 45.050 14.695 45.910 14.845 ;
        RECT 45.050 14.675 46.335 14.695 ;
        RECT 44.645 14.175 45.180 14.505 ;
        RECT 45.350 14.315 46.335 14.675 ;
        RECT 44.645 14.025 44.865 14.175 ;
        RECT 42.255 13.455 42.585 13.835 ;
        RECT 42.765 13.625 42.935 14.005 ;
        RECT 44.120 13.455 44.455 13.960 ;
        RECT 44.625 13.650 44.865 14.025 ;
        RECT 45.350 13.980 45.520 14.315 ;
        RECT 46.510 14.145 46.685 14.950 ;
        RECT 47.335 14.915 48.545 16.005 ;
        RECT 47.335 14.375 47.855 14.915 ;
        RECT 48.025 14.205 48.545 14.745 ;
        RECT 45.145 13.785 45.520 13.980 ;
        RECT 45.145 13.640 45.315 13.785 ;
        RECT 45.880 13.455 46.275 13.950 ;
        RECT 46.445 13.625 46.685 14.145 ;
        RECT 47.335 13.455 48.545 14.205 ;
        RECT 12.750 13.285 48.630 13.455 ;
      LAYER met1 ;
        RECT 12.750 48.490 48.630 48.970 ;
        RECT 21.575 48.290 21.865 48.335 ;
        RECT 26.620 48.290 26.940 48.350 ;
        RECT 21.575 48.150 26.940 48.290 ;
        RECT 21.575 48.105 21.865 48.150 ;
        RECT 26.620 48.090 26.940 48.150 ;
        RECT 32.155 48.290 32.445 48.335 ;
        RECT 33.060 48.290 33.380 48.350 ;
        RECT 32.155 48.150 33.380 48.290 ;
        RECT 32.155 48.105 32.445 48.150 ;
        RECT 33.060 48.090 33.380 48.150 ;
        RECT 39.500 48.290 39.820 48.350 ;
        RECT 40.435 48.290 40.725 48.335 ;
        RECT 39.500 48.150 40.725 48.290 ;
        RECT 39.500 48.090 39.820 48.150 ;
        RECT 40.435 48.105 40.725 48.150 ;
        RECT 23.875 47.950 24.165 47.995 ;
        RECT 31.220 47.950 31.540 48.010 ;
        RECT 38.120 47.950 38.440 48.010 ;
        RECT 23.875 47.810 31.540 47.950 ;
        RECT 23.875 47.765 24.165 47.810 ;
        RECT 31.220 47.750 31.540 47.810 ;
        RECT 32.690 47.810 38.440 47.950 ;
        RECT 27.095 47.610 27.385 47.655 ;
        RECT 20.730 47.470 27.385 47.610 ;
        RECT 18.340 47.270 18.660 47.330 ;
        RECT 20.730 47.315 20.870 47.470 ;
        RECT 27.095 47.425 27.385 47.470 ;
        RECT 20.655 47.270 20.945 47.315 ;
        RECT 18.340 47.130 20.945 47.270 ;
        RECT 18.340 47.070 18.660 47.130 ;
        RECT 20.655 47.085 20.945 47.130 ;
        RECT 22.940 47.070 23.260 47.330 ;
        RECT 23.400 47.070 23.720 47.330 ;
        RECT 24.335 47.270 24.625 47.315 ;
        RECT 32.690 47.270 32.830 47.810 ;
        RECT 38.120 47.750 38.440 47.810 ;
        RECT 24.335 47.130 32.830 47.270 ;
        RECT 33.075 47.270 33.365 47.315 ;
        RECT 33.520 47.270 33.840 47.330 ;
        RECT 33.075 47.130 33.840 47.270 ;
        RECT 24.335 47.085 24.625 47.130 ;
        RECT 33.075 47.085 33.365 47.130 ;
        RECT 33.520 47.070 33.840 47.130 ;
        RECT 36.280 47.270 36.600 47.330 ;
        RECT 37.215 47.270 37.505 47.315 ;
        RECT 36.280 47.130 37.505 47.270 ;
        RECT 36.280 47.070 36.600 47.130 ;
        RECT 37.215 47.085 37.505 47.130 ;
        RECT 41.340 47.070 41.660 47.330 ;
        RECT 44.100 47.070 44.420 47.330 ;
        RECT 45.480 47.070 45.800 47.330 ;
        RECT 46.860 47.070 47.180 47.330 ;
        RECT 25.240 46.390 25.560 46.650 ;
        RECT 30.300 46.390 30.620 46.650 ;
        RECT 33.980 46.590 34.300 46.650 ;
        RECT 36.755 46.590 37.045 46.635 ;
        RECT 33.980 46.450 37.045 46.590 ;
        RECT 33.980 46.390 34.300 46.450 ;
        RECT 36.755 46.405 37.045 46.450 ;
        RECT 39.960 46.590 40.280 46.650 ;
        RECT 43.195 46.590 43.485 46.635 ;
        RECT 39.960 46.450 43.485 46.590 ;
        RECT 39.960 46.390 40.280 46.450 ;
        RECT 43.195 46.405 43.485 46.450 ;
        RECT 43.640 46.590 43.960 46.650 ;
        RECT 44.575 46.590 44.865 46.635 ;
        RECT 43.640 46.450 44.865 46.590 ;
        RECT 43.640 46.390 43.960 46.450 ;
        RECT 44.575 46.405 44.865 46.450 ;
        RECT 45.955 46.590 46.245 46.635 ;
        RECT 46.400 46.590 46.720 46.650 ;
        RECT 45.955 46.450 46.720 46.590 ;
        RECT 45.955 46.405 46.245 46.450 ;
        RECT 46.400 46.390 46.720 46.450 ;
        RECT 12.750 45.770 48.630 46.250 ;
        RECT 18.340 45.370 18.660 45.630 ;
        RECT 22.940 45.570 23.260 45.630 ;
        RECT 32.615 45.570 32.905 45.615 ;
        RECT 33.520 45.570 33.840 45.630 ;
        RECT 22.940 45.430 28.230 45.570 ;
        RECT 22.940 45.370 23.260 45.430 ;
        RECT 25.240 45.230 25.560 45.290 ;
        RECT 26.940 45.230 27.230 45.275 ;
        RECT 25.240 45.090 27.230 45.230 ;
        RECT 28.090 45.230 28.230 45.430 ;
        RECT 32.615 45.430 33.840 45.570 ;
        RECT 32.615 45.385 32.905 45.430 ;
        RECT 33.520 45.370 33.840 45.430 ;
        RECT 33.075 45.230 33.365 45.275 ;
        RECT 28.090 45.090 33.365 45.230 ;
        RECT 25.240 45.030 25.560 45.090 ;
        RECT 26.940 45.045 27.230 45.090 ;
        RECT 33.075 45.045 33.365 45.090 ;
        RECT 33.980 45.030 34.300 45.290 ;
        RECT 23.975 44.890 24.265 44.935 ;
        RECT 26.160 44.890 26.480 44.950 ;
        RECT 23.975 44.750 26.480 44.890 ;
        RECT 23.975 44.705 24.265 44.750 ;
        RECT 26.160 44.690 26.480 44.750 ;
        RECT 34.900 44.690 35.220 44.950 ;
        RECT 35.375 44.705 35.665 44.935 ;
        RECT 36.280 44.890 36.600 44.950 ;
        RECT 37.215 44.890 37.505 44.935 ;
        RECT 36.280 44.750 37.505 44.890 ;
        RECT 20.665 44.550 20.955 44.595 ;
        RECT 23.185 44.550 23.475 44.595 ;
        RECT 24.375 44.550 24.665 44.595 ;
        RECT 20.665 44.410 24.665 44.550 ;
        RECT 20.665 44.365 20.955 44.410 ;
        RECT 23.185 44.365 23.475 44.410 ;
        RECT 24.375 44.365 24.665 44.410 ;
        RECT 25.255 44.550 25.545 44.595 ;
        RECT 25.715 44.550 26.005 44.595 ;
        RECT 25.255 44.410 26.005 44.550 ;
        RECT 25.255 44.365 25.545 44.410 ;
        RECT 25.715 44.365 26.005 44.410 ;
        RECT 26.595 44.550 26.885 44.595 ;
        RECT 27.785 44.550 28.075 44.595 ;
        RECT 30.305 44.550 30.595 44.595 ;
        RECT 26.595 44.410 30.595 44.550 ;
        RECT 26.595 44.365 26.885 44.410 ;
        RECT 27.785 44.365 28.075 44.410 ;
        RECT 30.305 44.365 30.595 44.410 ;
        RECT 31.680 44.550 32.000 44.610 ;
        RECT 35.450 44.550 35.590 44.705 ;
        RECT 36.280 44.690 36.600 44.750 ;
        RECT 37.215 44.705 37.505 44.750 ;
        RECT 38.120 44.890 38.440 44.950 ;
        RECT 39.975 44.890 40.265 44.935 ;
        RECT 38.120 44.750 40.265 44.890 ;
        RECT 38.120 44.690 38.440 44.750 ;
        RECT 39.975 44.705 40.265 44.750 ;
        RECT 40.880 44.690 41.200 44.950 ;
        RECT 41.355 44.890 41.645 44.935 ;
        RECT 44.100 44.890 44.420 44.950 ;
        RECT 41.355 44.750 44.420 44.890 ;
        RECT 41.355 44.705 41.645 44.750 ;
        RECT 44.100 44.690 44.420 44.750 ;
        RECT 46.860 44.690 47.180 44.950 ;
        RECT 31.680 44.410 35.590 44.550 ;
        RECT 35.820 44.550 36.140 44.610 ;
        RECT 38.210 44.550 38.350 44.690 ;
        RECT 35.820 44.410 38.350 44.550 ;
        RECT 21.100 44.210 21.390 44.255 ;
        RECT 22.670 44.210 22.960 44.255 ;
        RECT 24.770 44.210 25.060 44.255 ;
        RECT 21.100 44.070 25.060 44.210 ;
        RECT 21.100 44.025 21.390 44.070 ;
        RECT 22.670 44.025 22.960 44.070 ;
        RECT 24.770 44.025 25.060 44.070 ;
        RECT 23.860 43.870 24.180 43.930 ;
        RECT 25.790 43.870 25.930 44.365 ;
        RECT 31.680 44.350 32.000 44.410 ;
        RECT 35.820 44.350 36.140 44.410 ;
        RECT 42.275 44.365 42.565 44.595 ;
        RECT 26.200 44.210 26.490 44.255 ;
        RECT 28.300 44.210 28.590 44.255 ;
        RECT 29.870 44.210 30.160 44.255 ;
        RECT 26.200 44.070 30.160 44.210 ;
        RECT 26.200 44.025 26.490 44.070 ;
        RECT 28.300 44.025 28.590 44.070 ;
        RECT 29.870 44.025 30.160 44.070 ;
        RECT 30.760 44.210 31.080 44.270 ;
        RECT 36.295 44.210 36.585 44.255 ;
        RECT 30.760 44.070 36.585 44.210 ;
        RECT 30.760 44.010 31.080 44.070 ;
        RECT 36.295 44.025 36.585 44.070 ;
        RECT 37.675 44.210 37.965 44.255 ;
        RECT 40.435 44.210 40.725 44.255 ;
        RECT 37.675 44.070 40.725 44.210 ;
        RECT 37.675 44.025 37.965 44.070 ;
        RECT 40.435 44.025 40.725 44.070 ;
        RECT 41.340 44.210 41.660 44.270 ;
        RECT 42.350 44.210 42.490 44.365 ;
        RECT 41.340 44.070 42.490 44.210 ;
        RECT 44.560 44.210 44.880 44.270 ;
        RECT 45.955 44.210 46.245 44.255 ;
        RECT 44.560 44.070 46.245 44.210 ;
        RECT 41.340 44.010 41.660 44.070 ;
        RECT 44.560 44.010 44.880 44.070 ;
        RECT 45.955 44.025 46.245 44.070 ;
        RECT 34.440 43.870 34.760 43.930 ;
        RECT 23.860 43.730 34.760 43.870 ;
        RECT 23.860 43.670 24.180 43.730 ;
        RECT 34.440 43.670 34.760 43.730 ;
        RECT 37.200 43.870 37.520 43.930 ;
        RECT 39.055 43.870 39.345 43.915 ;
        RECT 37.200 43.730 39.345 43.870 ;
        RECT 37.200 43.670 37.520 43.730 ;
        RECT 39.055 43.685 39.345 43.730 ;
        RECT 43.180 43.870 43.500 43.930 ;
        RECT 45.495 43.870 45.785 43.915 ;
        RECT 43.180 43.730 45.785 43.870 ;
        RECT 43.180 43.670 43.500 43.730 ;
        RECT 45.495 43.685 45.785 43.730 ;
        RECT 12.750 43.050 48.630 43.530 ;
        RECT 26.160 42.650 26.480 42.910 ;
        RECT 31.220 42.850 31.540 42.910 ;
        RECT 33.535 42.850 33.825 42.895 ;
        RECT 36.280 42.850 36.600 42.910 ;
        RECT 31.220 42.710 33.825 42.850 ;
        RECT 31.220 42.650 31.540 42.710 ;
        RECT 33.535 42.665 33.825 42.710 ;
        RECT 34.530 42.710 39.730 42.850 ;
        RECT 14.700 42.510 14.990 42.555 ;
        RECT 16.800 42.510 17.090 42.555 ;
        RECT 18.370 42.510 18.660 42.555 ;
        RECT 34.530 42.510 34.670 42.710 ;
        RECT 36.280 42.650 36.600 42.710 ;
        RECT 14.700 42.370 18.660 42.510 ;
        RECT 14.700 42.325 14.990 42.370 ;
        RECT 16.800 42.325 17.090 42.370 ;
        RECT 18.370 42.325 18.660 42.370 ;
        RECT 29.470 42.370 34.670 42.510 ;
        RECT 34.940 42.510 35.230 42.555 ;
        RECT 37.040 42.510 37.330 42.555 ;
        RECT 38.610 42.510 38.900 42.555 ;
        RECT 34.940 42.370 38.900 42.510 ;
        RECT 29.470 42.215 29.610 42.370 ;
        RECT 34.940 42.325 35.230 42.370 ;
        RECT 37.040 42.325 37.330 42.370 ;
        RECT 38.610 42.325 38.900 42.370 ;
        RECT 15.095 42.170 15.385 42.215 ;
        RECT 16.285 42.170 16.575 42.215 ;
        RECT 18.805 42.170 19.095 42.215 ;
        RECT 15.095 42.030 19.095 42.170 ;
        RECT 15.095 41.985 15.385 42.030 ;
        RECT 16.285 41.985 16.575 42.030 ;
        RECT 18.805 41.985 19.095 42.030 ;
        RECT 29.395 41.985 29.685 42.215 ;
        RECT 34.440 41.970 34.760 42.230 ;
        RECT 35.335 42.170 35.625 42.215 ;
        RECT 36.525 42.170 36.815 42.215 ;
        RECT 39.045 42.170 39.335 42.215 ;
        RECT 35.335 42.030 39.335 42.170 ;
        RECT 35.335 41.985 35.625 42.030 ;
        RECT 36.525 41.985 36.815 42.030 ;
        RECT 39.045 41.985 39.335 42.030 ;
        RECT 14.215 41.830 14.505 41.875 ;
        RECT 23.860 41.830 24.180 41.890 ;
        RECT 14.215 41.690 24.180 41.830 ;
        RECT 14.215 41.645 14.505 41.690 ;
        RECT 23.860 41.630 24.180 41.690 ;
        RECT 24.335 41.645 24.625 41.875 ;
        RECT 28.015 41.830 28.305 41.875 ;
        RECT 30.300 41.830 30.620 41.890 ;
        RECT 28.015 41.690 30.620 41.830 ;
        RECT 28.015 41.645 28.305 41.690 ;
        RECT 15.550 41.490 15.840 41.535 ;
        RECT 16.040 41.490 16.360 41.550 ;
        RECT 24.410 41.490 24.550 41.645 ;
        RECT 30.300 41.630 30.620 41.690 ;
        RECT 30.760 41.630 31.080 41.890 ;
        RECT 31.680 41.830 32.000 41.890 ;
        RECT 33.520 41.830 33.840 41.890 ;
        RECT 31.680 41.690 33.840 41.830 ;
        RECT 31.680 41.630 32.000 41.690 ;
        RECT 33.520 41.630 33.840 41.690 ;
        RECT 33.980 41.830 34.300 41.890 ;
        RECT 34.900 41.830 35.220 41.890 ;
        RECT 33.980 41.690 35.220 41.830 ;
        RECT 33.980 41.630 34.300 41.690 ;
        RECT 34.900 41.630 35.220 41.690 ;
        RECT 35.790 41.830 36.080 41.875 ;
        RECT 37.200 41.830 37.520 41.890 ;
        RECT 35.790 41.690 37.520 41.830 ;
        RECT 39.590 41.830 39.730 42.710 ;
        RECT 41.340 42.650 41.660 42.910 ;
        RECT 44.100 42.650 44.420 42.910 ;
        RECT 42.275 41.830 42.565 41.875 ;
        RECT 39.590 41.690 42.565 41.830 ;
        RECT 35.790 41.645 36.080 41.690 ;
        RECT 37.200 41.630 37.520 41.690 ;
        RECT 42.275 41.645 42.565 41.690 ;
        RECT 43.180 41.630 43.500 41.890 ;
        RECT 44.560 41.630 44.880 41.890 ;
        RECT 46.860 41.630 47.180 41.890 ;
        RECT 15.550 41.350 16.360 41.490 ;
        RECT 15.550 41.305 15.840 41.350 ;
        RECT 16.040 41.290 16.360 41.350 ;
        RECT 21.190 41.350 24.550 41.490 ;
        RECT 28.475 41.490 28.765 41.535 ;
        RECT 36.280 41.490 36.600 41.550 ;
        RECT 28.475 41.350 36.600 41.490 ;
        RECT 21.190 41.210 21.330 41.350 ;
        RECT 28.475 41.305 28.765 41.350 ;
        RECT 36.280 41.290 36.600 41.350 ;
        RECT 21.100 40.950 21.420 41.210 ;
        RECT 21.560 40.950 21.880 41.210 ;
        RECT 30.300 41.150 30.620 41.210 ;
        RECT 32.615 41.150 32.905 41.195 ;
        RECT 30.300 41.010 32.905 41.150 ;
        RECT 30.300 40.950 30.620 41.010 ;
        RECT 32.615 40.965 32.905 41.010 ;
        RECT 45.480 40.950 45.800 41.210 ;
        RECT 45.940 40.950 46.260 41.210 ;
        RECT 12.750 40.330 48.630 40.810 ;
        RECT 13.740 40.130 14.060 40.190 ;
        RECT 14.675 40.130 14.965 40.175 ;
        RECT 13.740 39.990 14.965 40.130 ;
        RECT 13.740 39.930 14.060 39.990 ;
        RECT 14.675 39.945 14.965 39.990 ;
        RECT 16.040 39.930 16.360 40.190 ;
        RECT 17.895 40.130 18.185 40.175 ;
        RECT 21.560 40.130 21.880 40.190 ;
        RECT 17.895 39.990 21.880 40.130 ;
        RECT 17.895 39.945 18.185 39.990 ;
        RECT 21.560 39.930 21.880 39.990 ;
        RECT 23.860 40.130 24.180 40.190 ;
        RECT 26.160 40.130 26.480 40.190 ;
        RECT 23.860 39.990 26.480 40.130 ;
        RECT 23.860 39.930 24.180 39.990 ;
        RECT 26.160 39.930 26.480 39.990 ;
        RECT 27.080 40.130 27.400 40.190 ;
        RECT 30.760 40.130 31.080 40.190 ;
        RECT 43.640 40.130 43.960 40.190 ;
        RECT 27.080 39.990 31.080 40.130 ;
        RECT 27.080 39.930 27.400 39.990 ;
        RECT 30.760 39.930 31.080 39.990 ;
        RECT 37.290 39.990 43.960 40.130 ;
        RECT 35.820 39.590 36.140 39.850 ;
        RECT 15.595 39.450 15.885 39.495 ;
        RECT 21.100 39.450 21.420 39.510 ;
        RECT 15.595 39.310 21.420 39.450 ;
        RECT 15.595 39.265 15.885 39.310 ;
        RECT 21.100 39.250 21.420 39.310 ;
        RECT 30.315 39.450 30.605 39.495 ;
        RECT 30.760 39.450 31.080 39.510 ;
        RECT 37.290 39.495 37.430 39.990 ;
        RECT 43.640 39.930 43.960 39.990 ;
        RECT 45.940 39.930 46.260 40.190 ;
        RECT 39.055 39.790 39.345 39.835 ;
        RECT 40.420 39.790 40.740 39.850 ;
        RECT 39.055 39.650 40.740 39.790 ;
        RECT 39.055 39.605 39.345 39.650 ;
        RECT 40.420 39.590 40.740 39.650 ;
        RECT 40.880 39.790 41.200 39.850 ;
        RECT 46.030 39.790 46.170 39.930 ;
        RECT 40.880 39.650 46.170 39.790 ;
        RECT 40.880 39.590 41.200 39.650 ;
        RECT 30.315 39.310 31.080 39.450 ;
        RECT 30.315 39.265 30.605 39.310 ;
        RECT 30.760 39.250 31.080 39.310 ;
        RECT 37.215 39.265 37.505 39.495 ;
        RECT 39.960 39.250 40.280 39.510 ;
        RECT 42.350 39.495 42.490 39.650 ;
        RECT 41.355 39.265 41.645 39.495 ;
        RECT 42.275 39.265 42.565 39.495 ;
        RECT 18.355 38.925 18.645 39.155 ;
        RECT 19.275 39.110 19.565 39.155 ;
        RECT 19.720 39.110 20.040 39.170 ;
        RECT 19.275 38.970 20.040 39.110 ;
        RECT 19.275 38.925 19.565 38.970 ;
        RECT 16.500 38.770 16.820 38.830 ;
        RECT 18.430 38.770 18.570 38.925 ;
        RECT 19.720 38.910 20.040 38.970 ;
        RECT 33.995 39.110 34.285 39.155 ;
        RECT 34.440 39.110 34.760 39.170 ;
        RECT 33.995 38.970 34.760 39.110 ;
        RECT 33.995 38.925 34.285 38.970 ;
        RECT 34.440 38.910 34.760 38.970 ;
        RECT 36.755 39.110 37.045 39.155 ;
        RECT 40.050 39.110 40.190 39.250 ;
        RECT 36.755 38.970 40.190 39.110 ;
        RECT 41.430 39.110 41.570 39.265 ;
        RECT 43.640 39.250 43.960 39.510 ;
        RECT 45.020 39.250 45.340 39.510 ;
        RECT 45.955 39.450 46.245 39.495 ;
        RECT 46.400 39.450 46.720 39.510 ;
        RECT 45.955 39.310 46.720 39.450 ;
        RECT 45.955 39.265 46.245 39.310 ;
        RECT 46.400 39.250 46.720 39.310 ;
        RECT 42.735 39.110 43.025 39.155 ;
        RECT 41.430 38.970 43.025 39.110 ;
        RECT 36.755 38.925 37.045 38.970 ;
        RECT 42.735 38.925 43.025 38.970 ;
        RECT 36.280 38.770 36.600 38.830 ;
        RECT 40.880 38.770 41.200 38.830 ;
        RECT 16.500 38.630 36.600 38.770 ;
        RECT 16.500 38.570 16.820 38.630 ;
        RECT 36.280 38.570 36.600 38.630 ;
        RECT 37.290 38.630 41.200 38.770 ;
        RECT 30.775 38.430 31.065 38.475 ;
        RECT 31.220 38.430 31.540 38.490 ;
        RECT 37.290 38.475 37.430 38.630 ;
        RECT 40.880 38.570 41.200 38.630 ;
        RECT 30.775 38.290 31.540 38.430 ;
        RECT 30.775 38.245 31.065 38.290 ;
        RECT 31.220 38.230 31.540 38.290 ;
        RECT 37.215 38.245 37.505 38.475 ;
        RECT 38.120 38.230 38.440 38.490 ;
        RECT 12.750 37.610 48.630 38.090 ;
        RECT 27.080 37.410 27.400 37.470 ;
        RECT 18.430 37.270 27.400 37.410 ;
        RECT 16.500 36.530 16.820 36.790 ;
        RECT 17.435 36.730 17.725 36.775 ;
        RECT 18.430 36.730 18.570 37.270 ;
        RECT 27.080 37.210 27.400 37.270 ;
        RECT 33.075 37.410 33.365 37.455 ;
        RECT 33.520 37.410 33.840 37.470 ;
        RECT 33.075 37.270 33.840 37.410 ;
        RECT 33.075 37.225 33.365 37.270 ;
        RECT 33.520 37.210 33.840 37.270 ;
        RECT 43.195 37.410 43.485 37.455 ;
        RECT 45.020 37.410 45.340 37.470 ;
        RECT 43.195 37.270 45.340 37.410 ;
        RECT 43.195 37.225 43.485 37.270 ;
        RECT 45.020 37.210 45.340 37.270 ;
        RECT 18.840 37.070 19.130 37.115 ;
        RECT 20.940 37.070 21.230 37.115 ;
        RECT 22.510 37.070 22.800 37.115 ;
        RECT 18.840 36.930 22.800 37.070 ;
        RECT 18.840 36.885 19.130 36.930 ;
        RECT 20.940 36.885 21.230 36.930 ;
        RECT 22.510 36.885 22.800 36.930 ;
        RECT 25.255 36.885 25.545 37.115 ;
        RECT 26.660 37.070 26.950 37.115 ;
        RECT 28.760 37.070 29.050 37.115 ;
        RECT 30.330 37.070 30.620 37.115 ;
        RECT 26.660 36.930 30.620 37.070 ;
        RECT 26.660 36.885 26.950 36.930 ;
        RECT 28.760 36.885 29.050 36.930 ;
        RECT 30.330 36.885 30.620 36.930 ;
        RECT 17.435 36.590 18.570 36.730 ;
        RECT 19.235 36.730 19.525 36.775 ;
        RECT 20.425 36.730 20.715 36.775 ;
        RECT 22.945 36.730 23.235 36.775 ;
        RECT 19.235 36.590 23.235 36.730 ;
        RECT 17.435 36.545 17.725 36.590 ;
        RECT 19.235 36.545 19.525 36.590 ;
        RECT 20.425 36.545 20.715 36.590 ;
        RECT 22.945 36.545 23.235 36.590 ;
        RECT 18.355 36.390 18.645 36.435 ;
        RECT 21.100 36.390 21.420 36.450 ;
        RECT 23.860 36.390 24.180 36.450 ;
        RECT 18.355 36.250 24.180 36.390 ;
        RECT 25.330 36.390 25.470 36.885 ;
        RECT 34.900 36.870 35.220 37.130 ;
        RECT 41.800 37.070 42.120 37.130 ;
        RECT 46.400 37.070 46.720 37.130 ;
        RECT 39.590 36.930 46.720 37.070 ;
        RECT 26.160 36.530 26.480 36.790 ;
        RECT 39.590 36.775 39.730 36.930 ;
        RECT 41.800 36.870 42.120 36.930 ;
        RECT 46.400 36.870 46.720 36.930 ;
        RECT 27.055 36.730 27.345 36.775 ;
        RECT 28.245 36.730 28.535 36.775 ;
        RECT 30.765 36.730 31.055 36.775 ;
        RECT 27.055 36.590 31.055 36.730 ;
        RECT 27.055 36.545 27.345 36.590 ;
        RECT 28.245 36.545 28.535 36.590 ;
        RECT 30.765 36.545 31.055 36.590 ;
        RECT 39.515 36.545 39.805 36.775 ;
        RECT 39.975 36.730 40.265 36.775 ;
        RECT 42.720 36.730 43.040 36.790 ;
        RECT 39.975 36.590 43.040 36.730 ;
        RECT 39.975 36.545 40.265 36.590 ;
        RECT 42.720 36.530 43.040 36.590 ;
        RECT 34.440 36.390 34.760 36.450 ;
        RECT 25.330 36.250 35.590 36.390 ;
        RECT 18.355 36.205 18.645 36.250 ;
        RECT 21.100 36.190 21.420 36.250 ;
        RECT 23.860 36.190 24.180 36.250 ;
        RECT 34.440 36.190 34.760 36.250 ;
        RECT 35.450 36.110 35.590 36.250 ;
        RECT 39.055 36.205 39.345 36.435 ;
        RECT 40.435 36.205 40.725 36.435 ;
        RECT 40.880 36.390 41.200 36.450 ;
        RECT 41.355 36.390 41.645 36.435 ;
        RECT 40.880 36.250 41.645 36.390 ;
        RECT 19.720 36.095 20.040 36.110 ;
        RECT 19.690 36.050 20.040 36.095 ;
        RECT 27.510 36.050 27.800 36.095 ;
        RECT 33.980 36.050 34.300 36.110 ;
        RECT 19.285 35.910 27.310 36.050 ;
        RECT 19.690 35.865 20.040 35.910 ;
        RECT 19.720 35.850 20.040 35.865 ;
        RECT 14.200 35.510 14.520 35.770 ;
        RECT 16.055 35.710 16.345 35.755 ;
        RECT 18.800 35.710 19.120 35.770 ;
        RECT 16.055 35.570 19.120 35.710 ;
        RECT 27.170 35.710 27.310 35.910 ;
        RECT 27.510 35.910 34.300 36.050 ;
        RECT 27.510 35.865 27.800 35.910 ;
        RECT 33.980 35.850 34.300 35.910 ;
        RECT 35.360 36.050 35.680 36.110 ;
        RECT 36.755 36.050 37.045 36.095 ;
        RECT 35.360 35.910 37.045 36.050 ;
        RECT 39.130 36.050 39.270 36.205 ;
        RECT 40.510 36.050 40.650 36.205 ;
        RECT 40.880 36.190 41.200 36.250 ;
        RECT 41.355 36.205 41.645 36.250 ;
        RECT 42.275 36.390 42.565 36.435 ;
        RECT 43.640 36.390 43.960 36.450 ;
        RECT 42.275 36.250 43.960 36.390 ;
        RECT 42.275 36.205 42.565 36.250 ;
        RECT 43.640 36.190 43.960 36.250 ;
        RECT 44.100 36.190 44.420 36.450 ;
        RECT 45.480 36.190 45.800 36.450 ;
        RECT 45.940 36.390 46.260 36.450 ;
        RECT 46.415 36.390 46.705 36.435 ;
        RECT 45.940 36.250 46.705 36.390 ;
        RECT 45.940 36.190 46.260 36.250 ;
        RECT 46.415 36.205 46.705 36.250 ;
        RECT 41.815 36.050 42.105 36.095 ;
        RECT 39.130 35.910 39.730 36.050 ;
        RECT 40.510 35.910 42.105 36.050 ;
        RECT 35.360 35.850 35.680 35.910 ;
        RECT 36.755 35.865 37.045 35.910 ;
        RECT 33.520 35.710 33.840 35.770 ;
        RECT 34.455 35.710 34.745 35.755 ;
        RECT 27.170 35.570 34.745 35.710 ;
        RECT 16.055 35.525 16.345 35.570 ;
        RECT 18.800 35.510 19.120 35.570 ;
        RECT 33.520 35.510 33.840 35.570 ;
        RECT 34.455 35.525 34.745 35.570 ;
        RECT 38.135 35.710 38.425 35.755 ;
        RECT 39.040 35.710 39.360 35.770 ;
        RECT 38.135 35.570 39.360 35.710 ;
        RECT 39.590 35.710 39.730 35.910 ;
        RECT 41.815 35.865 42.105 35.910 ;
        RECT 44.190 35.710 44.330 36.190 ;
        RECT 39.590 35.570 44.330 35.710 ;
        RECT 38.135 35.525 38.425 35.570 ;
        RECT 39.040 35.510 39.360 35.570 ;
        RECT 12.750 34.890 48.630 35.370 ;
        RECT 33.980 34.490 34.300 34.750 ;
        RECT 36.280 34.690 36.600 34.750 ;
        RECT 40.895 34.690 41.185 34.735 ;
        RECT 36.280 34.550 41.185 34.690 ;
        RECT 36.280 34.490 36.600 34.550 ;
        RECT 40.895 34.505 41.185 34.550 ;
        RECT 45.955 34.505 46.245 34.735 ;
        RECT 14.200 34.350 14.520 34.410 ;
        RECT 19.780 34.350 20.070 34.395 ;
        RECT 14.200 34.210 20.070 34.350 ;
        RECT 14.200 34.150 14.520 34.210 ;
        RECT 19.780 34.165 20.070 34.210 ;
        RECT 24.780 34.150 25.100 34.410 ;
        RECT 46.030 34.350 46.170 34.505 ;
        RECT 44.650 34.210 46.170 34.350 ;
        RECT 44.650 34.070 44.790 34.210 ;
        RECT 21.100 33.810 21.420 34.070 ;
        RECT 39.040 33.810 39.360 34.070 ;
        RECT 39.960 33.810 40.280 34.070 ;
        RECT 44.560 33.810 44.880 34.070 ;
        RECT 45.495 34.010 45.785 34.055 ;
        RECT 45.940 34.010 46.260 34.070 ;
        RECT 45.495 33.870 46.260 34.010 ;
        RECT 45.495 33.825 45.785 33.870 ;
        RECT 45.940 33.810 46.260 33.870 ;
        RECT 46.860 33.810 47.180 34.070 ;
        RECT 16.525 33.670 16.815 33.715 ;
        RECT 19.045 33.670 19.335 33.715 ;
        RECT 20.235 33.670 20.525 33.715 ;
        RECT 16.525 33.530 20.525 33.670 ;
        RECT 16.525 33.485 16.815 33.530 ;
        RECT 19.045 33.485 19.335 33.530 ;
        RECT 20.235 33.485 20.525 33.530 ;
        RECT 31.220 33.670 31.540 33.730 ;
        RECT 36.755 33.670 37.045 33.715 ;
        RECT 31.220 33.530 37.045 33.670 ;
        RECT 31.220 33.470 31.540 33.530 ;
        RECT 36.755 33.485 37.045 33.530 ;
        RECT 16.960 33.330 17.250 33.375 ;
        RECT 18.530 33.330 18.820 33.375 ;
        RECT 20.630 33.330 20.920 33.375 ;
        RECT 16.960 33.190 20.920 33.330 ;
        RECT 16.960 33.145 17.250 33.190 ;
        RECT 18.530 33.145 18.820 33.190 ;
        RECT 20.630 33.145 20.920 33.190 ;
        RECT 14.200 32.790 14.520 33.050 ;
        RECT 30.760 32.990 31.080 33.050 ;
        RECT 31.235 32.990 31.525 33.035 ;
        RECT 30.760 32.850 31.525 32.990 ;
        RECT 30.760 32.790 31.080 32.850 ;
        RECT 31.235 32.805 31.525 32.850 ;
        RECT 35.820 32.990 36.140 33.050 ;
        RECT 39.055 32.990 39.345 33.035 ;
        RECT 35.820 32.850 39.345 32.990 ;
        RECT 35.820 32.790 36.140 32.850 ;
        RECT 39.055 32.805 39.345 32.850 ;
        RECT 42.260 32.990 42.580 33.050 ;
        RECT 45.495 32.990 45.785 33.035 ;
        RECT 42.260 32.850 45.785 32.990 ;
        RECT 42.260 32.790 42.580 32.850 ;
        RECT 45.495 32.805 45.785 32.850 ;
        RECT 12.750 32.170 48.630 32.650 ;
        RECT 18.800 31.770 19.120 32.030 ;
        RECT 27.080 31.770 27.400 32.030 ;
        RECT 27.540 31.970 27.860 32.030 ;
        RECT 29.395 31.970 29.685 32.015 ;
        RECT 27.540 31.830 29.685 31.970 ;
        RECT 27.540 31.770 27.860 31.830 ;
        RECT 29.395 31.785 29.685 31.830 ;
        RECT 38.120 31.770 38.440 32.030 ;
        RECT 45.480 31.970 45.800 32.030 ;
        RECT 46.415 31.970 46.705 32.015 ;
        RECT 45.480 31.830 46.705 31.970 ;
        RECT 45.480 31.770 45.800 31.830 ;
        RECT 46.415 31.785 46.705 31.830 ;
        RECT 28.475 31.630 28.765 31.675 ;
        RECT 31.680 31.630 32.000 31.690 ;
        RECT 35.820 31.630 36.140 31.690 ;
        RECT 28.475 31.490 32.000 31.630 ;
        RECT 28.475 31.445 28.765 31.490 ;
        RECT 14.200 31.290 14.520 31.350 ;
        RECT 15.595 31.290 15.885 31.335 ;
        RECT 28.550 31.290 28.690 31.445 ;
        RECT 31.680 31.430 32.000 31.490 ;
        RECT 34.530 31.490 36.140 31.630 ;
        RECT 14.200 31.150 15.885 31.290 ;
        RECT 14.200 31.090 14.520 31.150 ;
        RECT 15.595 31.105 15.885 31.150 ;
        RECT 27.170 31.150 28.690 31.290 ;
        RECT 28.935 31.290 29.225 31.335 ;
        RECT 34.530 31.290 34.670 31.490 ;
        RECT 35.820 31.430 36.140 31.490 ;
        RECT 44.100 31.430 44.420 31.690 ;
        RECT 28.935 31.150 34.670 31.290 ;
        RECT 22.020 30.750 22.340 31.010 ;
        RECT 27.170 30.995 27.310 31.150 ;
        RECT 28.935 31.105 29.225 31.150 ;
        RECT 34.900 31.090 35.220 31.350 ;
        RECT 44.190 31.290 44.330 31.430 ;
        RECT 37.750 31.150 44.330 31.290 ;
        RECT 26.175 30.765 26.465 30.995 ;
        RECT 27.095 30.765 27.385 30.995 ;
        RECT 26.250 30.610 26.390 30.765 ;
        RECT 27.540 30.750 27.860 31.010 ;
        RECT 29.855 30.950 30.145 30.995 ;
        RECT 30.300 30.950 30.620 31.010 ;
        RECT 29.855 30.810 30.620 30.950 ;
        RECT 29.855 30.765 30.145 30.810 ;
        RECT 30.300 30.750 30.620 30.810 ;
        RECT 31.220 30.750 31.540 31.010 ;
        RECT 37.750 30.995 37.890 31.150 ;
        RECT 37.675 30.765 37.965 30.995 ;
        RECT 38.595 30.950 38.885 30.995 ;
        RECT 40.435 30.950 40.725 30.995 ;
        RECT 40.880 30.950 41.200 31.010 ;
        RECT 41.430 30.995 41.570 31.150 ;
        RECT 38.595 30.810 41.200 30.950 ;
        RECT 38.595 30.765 38.885 30.810 ;
        RECT 40.435 30.765 40.725 30.810 ;
        RECT 40.880 30.750 41.200 30.810 ;
        RECT 41.355 30.765 41.645 30.995 ;
        RECT 41.800 30.750 42.120 31.010 ;
        RECT 43.195 30.765 43.485 30.995 ;
        RECT 31.695 30.610 31.985 30.655 ;
        RECT 26.250 30.470 31.985 30.610 ;
        RECT 31.695 30.425 31.985 30.470 ;
        RECT 39.975 30.610 40.265 30.655 ;
        RECT 42.260 30.610 42.580 30.670 ;
        RECT 43.270 30.610 43.410 30.765 ;
        RECT 44.100 30.750 44.420 31.010 ;
        RECT 44.560 30.950 44.880 31.010 ;
        RECT 45.495 30.950 45.785 30.995 ;
        RECT 44.560 30.810 45.785 30.950 ;
        RECT 44.560 30.750 44.880 30.810 ;
        RECT 45.495 30.765 45.785 30.810 ;
        RECT 45.020 30.610 45.340 30.670 ;
        RECT 39.975 30.470 42.580 30.610 ;
        RECT 39.975 30.425 40.265 30.470 ;
        RECT 42.260 30.410 42.580 30.470 ;
        RECT 42.810 30.470 45.340 30.610 ;
        RECT 19.260 30.070 19.580 30.330 ;
        RECT 36.755 30.270 37.045 30.315 ;
        RECT 37.660 30.270 37.980 30.330 ;
        RECT 36.755 30.130 37.980 30.270 ;
        RECT 36.755 30.085 37.045 30.130 ;
        RECT 37.660 30.070 37.980 30.130 ;
        RECT 40.420 30.270 40.740 30.330 ;
        RECT 42.810 30.315 42.950 30.470 ;
        RECT 45.020 30.410 45.340 30.470 ;
        RECT 40.895 30.270 41.185 30.315 ;
        RECT 40.420 30.130 41.185 30.270 ;
        RECT 40.420 30.070 40.740 30.130 ;
        RECT 40.895 30.085 41.185 30.130 ;
        RECT 42.735 30.085 43.025 30.315 ;
        RECT 12.750 29.450 48.630 29.930 ;
        RECT 13.740 29.250 14.060 29.310 ;
        RECT 14.675 29.250 14.965 29.295 ;
        RECT 13.740 29.110 14.965 29.250 ;
        RECT 13.740 29.050 14.060 29.110 ;
        RECT 14.675 29.065 14.965 29.110 ;
        RECT 18.355 29.250 18.645 29.295 ;
        RECT 19.260 29.250 19.580 29.310 ;
        RECT 18.355 29.110 19.580 29.250 ;
        RECT 18.355 29.065 18.645 29.110 ;
        RECT 19.260 29.050 19.580 29.110 ;
        RECT 27.540 29.250 27.860 29.310 ;
        RECT 34.440 29.250 34.760 29.310 ;
        RECT 27.540 29.110 34.760 29.250 ;
        RECT 27.540 29.050 27.860 29.110 ;
        RECT 34.440 29.050 34.760 29.110 ;
        RECT 44.100 29.250 44.420 29.310 ;
        RECT 46.415 29.250 46.705 29.295 ;
        RECT 44.100 29.110 46.705 29.250 ;
        RECT 44.100 29.050 44.420 29.110 ;
        RECT 46.415 29.065 46.705 29.110 ;
        RECT 21.990 28.910 22.280 28.955 ;
        RECT 25.700 28.910 26.020 28.970 ;
        RECT 27.080 28.910 27.400 28.970 ;
        RECT 42.260 28.910 42.580 28.970 ;
        RECT 21.990 28.770 27.400 28.910 ;
        RECT 21.990 28.725 22.280 28.770 ;
        RECT 25.700 28.710 26.020 28.770 ;
        RECT 27.080 28.710 27.400 28.770 ;
        RECT 40.050 28.770 42.580 28.910 ;
        RECT 14.200 28.570 14.520 28.630 ;
        RECT 15.595 28.570 15.885 28.615 ;
        RECT 14.200 28.430 15.885 28.570 ;
        RECT 14.200 28.370 14.520 28.430 ;
        RECT 15.595 28.385 15.885 28.430 ;
        RECT 29.855 28.570 30.145 28.615 ;
        RECT 32.155 28.570 32.445 28.615 ;
        RECT 29.855 28.430 32.445 28.570 ;
        RECT 29.855 28.385 30.145 28.430 ;
        RECT 32.155 28.385 32.445 28.430 ;
        RECT 38.120 28.570 38.440 28.630 ;
        RECT 40.050 28.615 40.190 28.770 ;
        RECT 42.260 28.710 42.580 28.770 ;
        RECT 39.515 28.570 39.805 28.615 ;
        RECT 38.120 28.430 39.805 28.570 ;
        RECT 38.120 28.370 38.440 28.430 ;
        RECT 39.515 28.385 39.805 28.430 ;
        RECT 39.975 28.385 40.265 28.615 ;
        RECT 40.420 28.370 40.740 28.630 ;
        RECT 43.195 28.570 43.485 28.615 ;
        RECT 43.640 28.570 43.960 28.630 ;
        RECT 43.195 28.430 43.960 28.570 ;
        RECT 43.195 28.385 43.485 28.430 ;
        RECT 43.640 28.370 43.960 28.430 ;
        RECT 44.100 28.370 44.420 28.630 ;
        RECT 45.495 28.570 45.785 28.615 ;
        RECT 45.940 28.570 46.260 28.630 ;
        RECT 45.495 28.430 46.260 28.570 ;
        RECT 45.495 28.385 45.785 28.430 ;
        RECT 45.940 28.370 46.260 28.430 ;
        RECT 18.815 28.230 19.105 28.275 ;
        RECT 19.260 28.230 19.580 28.290 ;
        RECT 18.815 28.090 19.580 28.230 ;
        RECT 18.815 28.045 19.105 28.090 ;
        RECT 19.260 28.030 19.580 28.090 ;
        RECT 19.720 28.030 20.040 28.290 ;
        RECT 20.655 28.045 20.945 28.275 ;
        RECT 21.535 28.230 21.825 28.275 ;
        RECT 22.725 28.230 23.015 28.275 ;
        RECT 25.245 28.230 25.535 28.275 ;
        RECT 21.535 28.090 25.535 28.230 ;
        RECT 21.535 28.045 21.825 28.090 ;
        RECT 22.725 28.045 23.015 28.090 ;
        RECT 25.245 28.045 25.535 28.090 ;
        RECT 30.315 28.045 30.605 28.275 ;
        RECT 31.235 28.230 31.525 28.275 ;
        RECT 33.520 28.230 33.840 28.290 ;
        RECT 31.235 28.090 33.840 28.230 ;
        RECT 31.235 28.045 31.525 28.090 ;
        RECT 14.200 27.890 14.520 27.950 ;
        RECT 20.730 27.890 20.870 28.045 ;
        RECT 14.200 27.750 20.870 27.890 ;
        RECT 21.140 27.890 21.430 27.935 ;
        RECT 23.240 27.890 23.530 27.935 ;
        RECT 24.810 27.890 25.100 27.935 ;
        RECT 21.140 27.750 25.100 27.890 ;
        RECT 14.200 27.690 14.520 27.750 ;
        RECT 21.140 27.705 21.430 27.750 ;
        RECT 23.240 27.705 23.530 27.750 ;
        RECT 24.810 27.705 25.100 27.750 ;
        RECT 27.080 27.890 27.400 27.950 ;
        RECT 28.015 27.890 28.305 27.935 ;
        RECT 27.080 27.750 28.305 27.890 ;
        RECT 30.390 27.890 30.530 28.045 ;
        RECT 33.520 28.030 33.840 28.090 ;
        RECT 33.980 28.230 34.300 28.290 ;
        RECT 34.915 28.230 35.205 28.275 ;
        RECT 33.980 28.090 35.205 28.230 ;
        RECT 33.980 28.030 34.300 28.090 ;
        RECT 34.915 28.045 35.205 28.090 ;
        RECT 40.895 28.230 41.185 28.275 ;
        RECT 44.560 28.230 44.880 28.290 ;
        RECT 40.895 28.090 44.880 28.230 ;
        RECT 40.895 28.045 41.185 28.090 ;
        RECT 44.560 28.030 44.880 28.090 ;
        RECT 35.820 27.890 36.140 27.950 ;
        RECT 41.815 27.890 42.105 27.935 ;
        RECT 30.390 27.750 42.105 27.890 ;
        RECT 27.080 27.690 27.400 27.750 ;
        RECT 28.015 27.705 28.305 27.750 ;
        RECT 35.820 27.690 36.140 27.750 ;
        RECT 41.815 27.705 42.105 27.750 ;
        RECT 16.500 27.350 16.820 27.610 ;
        RECT 12.750 26.730 48.630 27.210 ;
        RECT 21.115 26.530 21.405 26.575 ;
        RECT 22.020 26.530 22.340 26.590 ;
        RECT 21.115 26.390 22.340 26.530 ;
        RECT 21.115 26.345 21.405 26.390 ;
        RECT 22.020 26.330 22.340 26.390 ;
        RECT 35.835 26.530 36.125 26.575 ;
        RECT 36.740 26.530 37.060 26.590 ;
        RECT 35.835 26.390 37.060 26.530 ;
        RECT 35.835 26.345 36.125 26.390 ;
        RECT 36.740 26.330 37.060 26.390 ;
        RECT 42.720 26.530 43.040 26.590 ;
        RECT 43.655 26.530 43.945 26.575 ;
        RECT 42.720 26.390 43.945 26.530 ;
        RECT 42.720 26.330 43.040 26.390 ;
        RECT 43.655 26.345 43.945 26.390 ;
        RECT 14.700 26.190 14.990 26.235 ;
        RECT 16.800 26.190 17.090 26.235 ;
        RECT 18.370 26.190 18.660 26.235 ;
        RECT 14.700 26.050 18.660 26.190 ;
        RECT 14.700 26.005 14.990 26.050 ;
        RECT 16.800 26.005 17.090 26.050 ;
        RECT 18.370 26.005 18.660 26.050 ;
        RECT 26.660 26.190 26.950 26.235 ;
        RECT 28.760 26.190 29.050 26.235 ;
        RECT 30.330 26.190 30.620 26.235 ;
        RECT 26.660 26.050 30.620 26.190 ;
        RECT 26.660 26.005 26.950 26.050 ;
        RECT 28.760 26.005 29.050 26.050 ;
        RECT 30.330 26.005 30.620 26.050 ;
        RECT 35.360 25.990 35.680 26.250 ;
        RECT 14.200 25.650 14.520 25.910 ;
        RECT 15.095 25.850 15.385 25.895 ;
        RECT 16.285 25.850 16.575 25.895 ;
        RECT 18.805 25.850 19.095 25.895 ;
        RECT 15.095 25.710 19.095 25.850 ;
        RECT 15.095 25.665 15.385 25.710 ;
        RECT 16.285 25.665 16.575 25.710 ;
        RECT 18.805 25.665 19.095 25.710 ;
        RECT 27.055 25.850 27.345 25.895 ;
        RECT 28.245 25.850 28.535 25.895 ;
        RECT 30.765 25.850 31.055 25.895 ;
        RECT 27.055 25.710 31.055 25.850 ;
        RECT 27.055 25.665 27.345 25.710 ;
        RECT 28.245 25.665 28.535 25.710 ;
        RECT 30.765 25.665 31.055 25.710 ;
        RECT 33.535 25.850 33.825 25.895 ;
        RECT 34.440 25.850 34.760 25.910 ;
        RECT 33.535 25.710 34.760 25.850 ;
        RECT 33.535 25.665 33.825 25.710 ;
        RECT 34.440 25.650 34.760 25.710 ;
        RECT 42.260 25.850 42.580 25.910 ;
        RECT 42.260 25.710 46.170 25.850 ;
        RECT 42.260 25.650 42.580 25.710 ;
        RECT 14.290 25.510 14.430 25.650 ;
        RECT 21.100 25.510 21.420 25.570 ;
        RECT 26.175 25.510 26.465 25.555 ;
        RECT 14.290 25.370 26.465 25.510 ;
        RECT 21.100 25.310 21.420 25.370 ;
        RECT 26.175 25.325 26.465 25.370 ;
        RECT 27.510 25.325 27.800 25.555 ;
        RECT 15.550 25.170 15.840 25.215 ;
        RECT 16.500 25.170 16.820 25.230 ;
        RECT 15.550 25.030 16.820 25.170 ;
        RECT 15.550 24.985 15.840 25.030 ;
        RECT 16.500 24.970 16.820 25.030 ;
        RECT 26.250 24.830 26.390 25.325 ;
        RECT 27.080 25.170 27.400 25.230 ;
        RECT 27.630 25.170 27.770 25.325 ;
        RECT 39.960 25.310 40.280 25.570 ;
        RECT 42.720 25.510 43.040 25.570 ;
        RECT 44.575 25.510 44.865 25.555 ;
        RECT 42.720 25.370 44.865 25.510 ;
        RECT 42.720 25.310 43.040 25.370 ;
        RECT 44.575 25.325 44.865 25.370 ;
        RECT 45.020 25.310 45.340 25.570 ;
        RECT 45.480 25.310 45.800 25.570 ;
        RECT 46.030 25.555 46.170 25.710 ;
        RECT 45.955 25.325 46.245 25.555 ;
        RECT 27.080 25.030 27.770 25.170 ;
        RECT 27.080 24.970 27.400 25.030 ;
        RECT 31.220 24.830 31.540 24.890 ;
        RECT 26.250 24.690 31.540 24.830 ;
        RECT 31.220 24.630 31.540 24.690 ;
        RECT 33.075 24.830 33.365 24.875 ;
        RECT 33.980 24.830 34.300 24.890 ;
        RECT 33.075 24.690 34.300 24.830 ;
        RECT 33.075 24.645 33.365 24.690 ;
        RECT 33.980 24.630 34.300 24.690 ;
        RECT 40.880 24.830 41.200 24.890 ;
        RECT 43.195 24.830 43.485 24.875 ;
        RECT 40.880 24.690 43.485 24.830 ;
        RECT 40.880 24.630 41.200 24.690 ;
        RECT 43.195 24.645 43.485 24.690 ;
        RECT 12.750 24.010 48.630 24.490 ;
        RECT 40.880 23.610 41.200 23.870 ;
        RECT 44.560 23.610 44.880 23.870 ;
        RECT 35.820 23.470 36.140 23.530 ;
        RECT 30.850 23.330 36.140 23.470 ;
        RECT 15.595 23.130 15.885 23.175 ;
        RECT 22.020 23.130 22.340 23.190 ;
        RECT 15.595 22.990 22.340 23.130 ;
        RECT 15.595 22.945 15.885 22.990 ;
        RECT 22.020 22.930 22.340 22.990 ;
        RECT 24.795 23.130 25.085 23.175 ;
        RECT 27.095 23.130 27.385 23.175 ;
        RECT 24.795 22.990 27.385 23.130 ;
        RECT 24.795 22.945 25.085 22.990 ;
        RECT 27.095 22.945 27.385 22.990 ;
        RECT 14.200 22.790 14.520 22.850 ;
        RECT 16.975 22.790 17.265 22.835 ;
        RECT 14.200 22.650 17.265 22.790 ;
        RECT 14.200 22.590 14.520 22.650 ;
        RECT 16.975 22.605 17.265 22.650 ;
        RECT 21.560 22.590 21.880 22.850 ;
        RECT 25.700 22.590 26.020 22.850 ;
        RECT 26.635 22.790 26.925 22.835 ;
        RECT 30.850 22.790 30.990 23.330 ;
        RECT 35.820 23.270 36.140 23.330 ;
        RECT 45.020 23.470 45.340 23.530 ;
        RECT 46.875 23.470 47.165 23.515 ;
        RECT 45.020 23.330 47.165 23.470 ;
        RECT 45.020 23.270 45.340 23.330 ;
        RECT 46.875 23.285 47.165 23.330 ;
        RECT 31.220 22.930 31.540 23.190 ;
        RECT 32.570 23.130 32.860 23.175 ;
        RECT 36.740 23.130 37.060 23.190 ;
        RECT 32.570 22.990 36.510 23.130 ;
        RECT 32.570 22.945 32.860 22.990 ;
        RECT 26.635 22.650 30.990 22.790 ;
        RECT 32.115 22.790 32.405 22.835 ;
        RECT 33.305 22.790 33.595 22.835 ;
        RECT 35.825 22.790 36.115 22.835 ;
        RECT 32.115 22.650 36.115 22.790 ;
        RECT 26.635 22.605 26.925 22.650 ;
        RECT 32.115 22.605 32.405 22.650 ;
        RECT 33.305 22.605 33.595 22.650 ;
        RECT 35.825 22.605 36.115 22.650 ;
        RECT 13.740 22.450 14.060 22.510 ;
        RECT 14.675 22.450 14.965 22.495 ;
        RECT 13.740 22.310 14.965 22.450 ;
        RECT 13.740 22.250 14.060 22.310 ;
        RECT 14.675 22.265 14.965 22.310 ;
        RECT 19.260 22.450 19.580 22.510 ;
        RECT 31.720 22.450 32.010 22.495 ;
        RECT 33.820 22.450 34.110 22.495 ;
        RECT 35.390 22.450 35.680 22.495 ;
        RECT 19.260 22.310 31.450 22.450 ;
        RECT 19.260 22.250 19.580 22.310 ;
        RECT 18.800 22.110 19.120 22.170 ;
        RECT 20.195 22.110 20.485 22.155 ;
        RECT 18.800 21.970 20.485 22.110 ;
        RECT 18.800 21.910 19.120 21.970 ;
        RECT 20.195 21.925 20.485 21.970 ;
        RECT 28.935 22.110 29.225 22.155 ;
        RECT 30.300 22.110 30.620 22.170 ;
        RECT 28.935 21.970 30.620 22.110 ;
        RECT 31.310 22.110 31.450 22.310 ;
        RECT 31.720 22.310 35.680 22.450 ;
        RECT 36.370 22.450 36.510 22.990 ;
        RECT 36.740 22.990 42.030 23.130 ;
        RECT 36.740 22.930 37.060 22.990 ;
        RECT 37.660 22.790 37.980 22.850 ;
        RECT 41.890 22.835 42.030 22.990 ;
        RECT 43.180 22.930 43.500 23.190 ;
        RECT 44.560 23.130 44.880 23.190 ;
        RECT 45.495 23.130 45.785 23.175 ;
        RECT 44.560 22.990 45.785 23.130 ;
        RECT 44.560 22.930 44.880 22.990 ;
        RECT 45.495 22.945 45.785 22.990 ;
        RECT 41.355 22.790 41.645 22.835 ;
        RECT 37.660 22.650 41.645 22.790 ;
        RECT 37.660 22.590 37.980 22.650 ;
        RECT 41.355 22.605 41.645 22.650 ;
        RECT 41.815 22.605 42.105 22.835 ;
        RECT 42.720 22.790 43.040 22.850 ;
        RECT 45.940 22.790 46.260 22.850 ;
        RECT 42.720 22.650 46.260 22.790 ;
        RECT 42.720 22.590 43.040 22.650 ;
        RECT 45.940 22.590 46.260 22.650 ;
        RECT 39.055 22.450 39.345 22.495 ;
        RECT 36.370 22.310 39.345 22.450 ;
        RECT 31.720 22.265 32.010 22.310 ;
        RECT 33.820 22.265 34.110 22.310 ;
        RECT 35.390 22.265 35.680 22.310 ;
        RECT 39.055 22.265 39.345 22.310 ;
        RECT 44.115 22.450 44.405 22.495 ;
        RECT 46.860 22.450 47.180 22.510 ;
        RECT 44.115 22.310 47.180 22.450 ;
        RECT 44.115 22.265 44.405 22.310 ;
        RECT 46.860 22.250 47.180 22.310 ;
        RECT 37.660 22.110 37.980 22.170 ;
        RECT 31.310 21.970 37.980 22.110 ;
        RECT 28.935 21.925 29.225 21.970 ;
        RECT 30.300 21.910 30.620 21.970 ;
        RECT 37.660 21.910 37.980 21.970 ;
        RECT 38.135 22.110 38.425 22.155 ;
        RECT 39.960 22.110 40.280 22.170 ;
        RECT 38.135 21.970 40.280 22.110 ;
        RECT 38.135 21.925 38.425 21.970 ;
        RECT 39.960 21.910 40.280 21.970 ;
        RECT 43.640 22.110 43.960 22.170 ;
        RECT 45.495 22.110 45.785 22.155 ;
        RECT 43.640 21.970 45.785 22.110 ;
        RECT 43.640 21.910 43.960 21.970 ;
        RECT 45.495 21.925 45.785 21.970 ;
        RECT 12.750 21.290 48.630 21.770 ;
        RECT 14.200 20.890 14.520 21.150 ;
        RECT 31.220 21.090 31.540 21.150 ;
        RECT 32.615 21.090 32.905 21.135 ;
        RECT 31.220 20.950 32.905 21.090 ;
        RECT 31.220 20.890 31.540 20.950 ;
        RECT 32.615 20.905 32.905 20.950 ;
        RECT 40.435 21.090 40.725 21.135 ;
        RECT 42.720 21.090 43.040 21.150 ;
        RECT 40.435 20.950 43.040 21.090 ;
        RECT 40.435 20.905 40.725 20.950 ;
        RECT 42.720 20.890 43.040 20.950 ;
        RECT 43.655 21.090 43.945 21.135 ;
        RECT 44.100 21.090 44.420 21.150 ;
        RECT 43.655 20.950 44.420 21.090 ;
        RECT 43.655 20.905 43.945 20.950 ;
        RECT 44.100 20.890 44.420 20.950 ;
        RECT 16.960 20.750 17.250 20.795 ;
        RECT 18.530 20.750 18.820 20.795 ;
        RECT 20.630 20.750 20.920 20.795 ;
        RECT 16.960 20.610 20.920 20.750 ;
        RECT 16.960 20.565 17.250 20.610 ;
        RECT 18.530 20.565 18.820 20.610 ;
        RECT 20.630 20.565 20.920 20.610 ;
        RECT 37.675 20.750 37.965 20.795 ;
        RECT 43.180 20.750 43.500 20.810 ;
        RECT 37.675 20.610 43.500 20.750 ;
        RECT 37.675 20.565 37.965 20.610 ;
        RECT 43.180 20.550 43.500 20.610 ;
        RECT 16.525 20.410 16.815 20.455 ;
        RECT 19.045 20.410 19.335 20.455 ;
        RECT 20.235 20.410 20.525 20.455 ;
        RECT 16.525 20.270 20.525 20.410 ;
        RECT 16.525 20.225 16.815 20.270 ;
        RECT 19.045 20.225 19.335 20.270 ;
        RECT 20.235 20.225 20.525 20.270 ;
        RECT 21.100 20.210 21.420 20.470 ;
        RECT 46.400 20.410 46.720 20.470 ;
        RECT 36.830 20.270 46.720 20.410 ;
        RECT 26.175 20.070 26.465 20.115 ;
        RECT 30.760 20.070 31.080 20.130 ;
        RECT 36.830 20.115 36.970 20.270 ;
        RECT 46.400 20.210 46.720 20.270 ;
        RECT 26.175 19.930 31.080 20.070 ;
        RECT 26.175 19.885 26.465 19.930 ;
        RECT 30.760 19.870 31.080 19.930 ;
        RECT 36.755 19.885 37.045 20.115 ;
        RECT 38.120 19.870 38.440 20.130 ;
        RECT 39.500 19.870 39.820 20.130 ;
        RECT 40.880 19.870 41.200 20.130 ;
        RECT 42.275 19.885 42.565 20.115 ;
        RECT 43.195 20.070 43.485 20.115 ;
        RECT 43.640 20.070 43.960 20.130 ;
        RECT 43.195 19.930 43.960 20.070 ;
        RECT 43.195 19.885 43.485 19.930 ;
        RECT 16.960 19.730 17.280 19.790 ;
        RECT 19.780 19.730 20.070 19.775 ;
        RECT 42.350 19.730 42.490 19.885 ;
        RECT 43.640 19.870 43.960 19.930 ;
        RECT 44.560 19.870 44.880 20.130 ;
        RECT 45.940 19.870 46.260 20.130 ;
        RECT 46.860 19.870 47.180 20.130 ;
        RECT 44.650 19.730 44.790 19.870 ;
        RECT 16.960 19.590 20.070 19.730 ;
        RECT 16.960 19.530 17.280 19.590 ;
        RECT 19.780 19.545 20.070 19.590 ;
        RECT 39.130 19.590 44.790 19.730 ;
        RECT 39.130 19.435 39.270 19.590 ;
        RECT 39.055 19.205 39.345 19.435 ;
        RECT 41.815 19.390 42.105 19.435 ;
        RECT 42.260 19.390 42.580 19.450 ;
        RECT 41.815 19.250 42.580 19.390 ;
        RECT 41.815 19.205 42.105 19.250 ;
        RECT 42.260 19.190 42.580 19.250 ;
        RECT 42.720 19.190 43.040 19.450 ;
        RECT 12.750 18.570 48.630 19.050 ;
        RECT 16.960 18.170 17.280 18.430 ;
        RECT 18.800 18.170 19.120 18.430 ;
        RECT 19.260 18.170 19.580 18.430 ;
        RECT 21.560 18.370 21.880 18.430 ;
        RECT 23.860 18.370 24.180 18.430 ;
        RECT 26.175 18.370 26.465 18.415 ;
        RECT 21.560 18.230 26.465 18.370 ;
        RECT 21.560 18.170 21.880 18.230 ;
        RECT 23.860 18.170 24.180 18.230 ;
        RECT 26.175 18.185 26.465 18.230 ;
        RECT 30.300 18.170 30.620 18.430 ;
        RECT 35.820 18.170 36.140 18.430 ;
        RECT 45.480 18.370 45.800 18.430 ;
        RECT 45.955 18.370 46.245 18.415 ;
        RECT 45.480 18.230 46.245 18.370 ;
        RECT 45.480 18.170 45.800 18.230 ;
        RECT 45.955 18.185 46.245 18.230 ;
        RECT 14.200 17.690 14.520 17.750 ;
        RECT 15.595 17.690 15.885 17.735 ;
        RECT 14.200 17.550 15.885 17.690 ;
        RECT 30.390 17.690 30.530 18.170 ;
        RECT 31.220 18.030 31.540 18.090 ;
        RECT 31.220 17.890 33.290 18.030 ;
        RECT 31.220 17.830 31.540 17.890 ;
        RECT 33.150 17.735 33.290 17.890 ;
        RECT 31.740 17.690 32.030 17.735 ;
        RECT 30.390 17.550 32.030 17.690 ;
        RECT 14.200 17.490 14.520 17.550 ;
        RECT 15.595 17.505 15.885 17.550 ;
        RECT 31.740 17.505 32.030 17.550 ;
        RECT 33.075 17.505 33.365 17.735 ;
        RECT 35.375 17.690 35.665 17.735 ;
        RECT 39.055 17.690 39.345 17.735 ;
        RECT 35.375 17.550 39.345 17.690 ;
        RECT 35.375 17.505 35.665 17.550 ;
        RECT 39.055 17.505 39.345 17.550 ;
        RECT 42.720 17.690 43.040 17.750 ;
        RECT 45.035 17.690 45.325 17.735 ;
        RECT 42.720 17.550 45.325 17.690 ;
        RECT 42.720 17.490 43.040 17.550 ;
        RECT 45.035 17.505 45.325 17.550 ;
        RECT 20.195 17.350 20.485 17.395 ;
        RECT 25.700 17.350 26.020 17.410 ;
        RECT 20.195 17.210 26.020 17.350 ;
        RECT 20.195 17.165 20.485 17.210 ;
        RECT 25.700 17.150 26.020 17.210 ;
        RECT 28.485 17.350 28.775 17.395 ;
        RECT 31.005 17.350 31.295 17.395 ;
        RECT 32.195 17.350 32.485 17.395 ;
        RECT 28.485 17.210 32.485 17.350 ;
        RECT 28.485 17.165 28.775 17.210 ;
        RECT 31.005 17.165 31.295 17.210 ;
        RECT 32.195 17.165 32.485 17.210 ;
        RECT 36.740 17.150 37.060 17.410 ;
        RECT 37.200 17.350 37.520 17.410 ;
        RECT 41.815 17.350 42.105 17.395 ;
        RECT 37.200 17.210 42.105 17.350 ;
        RECT 37.200 17.150 37.520 17.210 ;
        RECT 41.815 17.165 42.105 17.210 ;
        RECT 42.260 17.350 42.580 17.410 ;
        RECT 43.655 17.350 43.945 17.395 ;
        RECT 42.260 17.210 43.945 17.350 ;
        RECT 42.260 17.150 42.580 17.210 ;
        RECT 43.655 17.165 43.945 17.210 ;
        RECT 44.115 17.350 44.405 17.395 ;
        RECT 46.860 17.350 47.180 17.410 ;
        RECT 44.115 17.210 47.180 17.350 ;
        RECT 44.115 17.165 44.405 17.210 ;
        RECT 46.860 17.150 47.180 17.210 ;
        RECT 11.440 17.010 11.760 17.070 ;
        RECT 14.675 17.010 14.965 17.055 ;
        RECT 11.440 16.870 14.965 17.010 ;
        RECT 11.440 16.810 11.760 16.870 ;
        RECT 14.675 16.825 14.965 16.870 ;
        RECT 28.920 17.010 29.210 17.055 ;
        RECT 30.490 17.010 30.780 17.055 ;
        RECT 32.590 17.010 32.880 17.055 ;
        RECT 28.920 16.870 32.880 17.010 ;
        RECT 28.920 16.825 29.210 16.870 ;
        RECT 30.490 16.825 30.780 16.870 ;
        RECT 32.590 16.825 32.880 16.870 ;
        RECT 31.220 16.670 31.540 16.730 ;
        RECT 33.535 16.670 33.825 16.715 ;
        RECT 31.220 16.530 33.825 16.670 ;
        RECT 31.220 16.470 31.540 16.530 ;
        RECT 33.535 16.485 33.825 16.530 ;
        RECT 12.750 15.850 48.630 16.330 ;
        RECT 33.980 15.650 34.300 15.710 ;
        RECT 28.090 15.510 34.300 15.650 ;
        RECT 23.860 14.430 24.180 14.690 ;
        RECT 28.090 14.675 28.230 15.510 ;
        RECT 33.980 15.450 34.300 15.510 ;
        RECT 41.815 15.650 42.105 15.695 ;
        RECT 43.640 15.650 43.960 15.710 ;
        RECT 41.815 15.510 43.960 15.650 ;
        RECT 41.815 15.465 42.105 15.510 ;
        RECT 43.640 15.450 43.960 15.510 ;
        RECT 45.940 15.650 46.260 15.710 ;
        RECT 46.415 15.650 46.705 15.695 ;
        RECT 45.940 15.510 46.705 15.650 ;
        RECT 45.940 15.450 46.260 15.510 ;
        RECT 46.415 15.465 46.705 15.510 ;
        RECT 28.960 15.310 29.250 15.355 ;
        RECT 31.060 15.310 31.350 15.355 ;
        RECT 32.630 15.310 32.920 15.355 ;
        RECT 28.960 15.170 32.920 15.310 ;
        RECT 28.960 15.125 29.250 15.170 ;
        RECT 31.060 15.125 31.350 15.170 ;
        RECT 32.630 15.125 32.920 15.170 ;
        RECT 35.375 15.310 35.665 15.355 ;
        RECT 37.200 15.310 37.520 15.370 ;
        RECT 35.375 15.170 37.520 15.310 ;
        RECT 35.375 15.125 35.665 15.170 ;
        RECT 37.200 15.110 37.520 15.170 ;
        RECT 43.180 15.310 43.500 15.370 ;
        RECT 45.495 15.310 45.785 15.355 ;
        RECT 43.180 15.170 45.785 15.310 ;
        RECT 43.180 15.110 43.500 15.170 ;
        RECT 45.495 15.125 45.785 15.170 ;
        RECT 29.355 14.970 29.645 15.015 ;
        RECT 30.545 14.970 30.835 15.015 ;
        RECT 33.065 14.970 33.355 15.015 ;
        RECT 29.355 14.830 33.355 14.970 ;
        RECT 29.355 14.785 29.645 14.830 ;
        RECT 30.545 14.785 30.835 14.830 ;
        RECT 33.065 14.785 33.355 14.830 ;
        RECT 42.260 14.970 42.580 15.030 ;
        RECT 44.115 14.970 44.405 15.015 ;
        RECT 42.260 14.830 44.405 14.970 ;
        RECT 42.260 14.770 42.580 14.830 ;
        RECT 44.115 14.785 44.405 14.830 ;
        RECT 28.015 14.445 28.305 14.675 ;
        RECT 28.475 14.630 28.765 14.675 ;
        RECT 28.920 14.630 29.240 14.690 ;
        RECT 28.475 14.490 29.240 14.630 ;
        RECT 28.475 14.445 28.765 14.490 ;
        RECT 28.920 14.430 29.240 14.490 ;
        RECT 37.200 14.430 37.520 14.690 ;
        RECT 39.960 14.430 40.280 14.690 ;
        RECT 42.720 14.430 43.040 14.690 ;
        RECT 29.810 14.290 30.100 14.335 ;
        RECT 31.220 14.290 31.540 14.350 ;
        RECT 29.810 14.150 31.540 14.290 ;
        RECT 29.810 14.105 30.100 14.150 ;
        RECT 31.220 14.090 31.540 14.150 ;
        RECT 33.610 14.150 36.510 14.290 ;
        RECT 33.610 14.010 33.750 14.150 ;
        RECT 24.795 13.950 25.085 13.995 ;
        RECT 26.620 13.950 26.940 14.010 ;
        RECT 24.795 13.810 26.940 13.950 ;
        RECT 24.795 13.765 25.085 13.810 ;
        RECT 26.620 13.750 26.940 13.810 ;
        RECT 27.095 13.950 27.385 13.995 ;
        RECT 29.380 13.950 29.700 14.010 ;
        RECT 27.095 13.810 29.700 13.950 ;
        RECT 27.095 13.765 27.385 13.810 ;
        RECT 29.380 13.750 29.700 13.810 ;
        RECT 33.520 13.750 33.840 14.010 ;
        RECT 36.370 13.995 36.510 14.150 ;
        RECT 36.295 13.765 36.585 13.995 ;
        RECT 39.500 13.950 39.820 14.010 ;
        RECT 40.895 13.950 41.185 13.995 ;
        RECT 39.500 13.810 41.185 13.950 ;
        RECT 39.500 13.750 39.820 13.810 ;
        RECT 40.895 13.765 41.185 13.810 ;
        RECT 12.750 13.130 48.630 13.610 ;
      LAYER met2 ;
        RECT 26.640 56.255 26.920 60.255 ;
        RECT 29.860 56.255 30.140 60.255 ;
        RECT 33.080 56.255 33.360 60.255 ;
        RECT 36.300 56.255 36.580 60.255 ;
        RECT 39.520 56.255 39.800 60.255 ;
        RECT 26.710 48.380 26.850 56.255 ;
        RECT 29.930 49.820 30.070 56.255 ;
        RECT 29.930 49.680 30.990 49.820 ;
        RECT 28.300 48.545 29.840 48.915 ;
        RECT 26.650 48.060 26.910 48.380 ;
        RECT 18.370 47.040 18.630 47.360 ;
        RECT 22.970 47.040 23.230 47.360 ;
        RECT 23.430 47.040 23.690 47.360 ;
        RECT 18.430 45.660 18.570 47.040 ;
        RECT 23.030 45.660 23.170 47.040 ;
        RECT 18.370 45.340 18.630 45.660 ;
        RECT 22.970 45.340 23.230 45.660 ;
        RECT 23.490 45.175 23.630 47.040 ;
        RECT 25.270 46.360 25.530 46.680 ;
        RECT 30.330 46.360 30.590 46.680 ;
        RECT 25.330 45.320 25.470 46.360 ;
        RECT 23.420 44.805 23.700 45.175 ;
        RECT 25.270 45.000 25.530 45.320 ;
        RECT 26.190 44.660 26.450 44.980 ;
        RECT 27.560 44.805 27.840 45.175 ;
        RECT 23.890 43.640 24.150 43.960 ;
        RECT 23.950 41.920 24.090 43.640 ;
        RECT 24.800 43.445 25.080 43.815 ;
        RECT 23.890 41.600 24.150 41.920 ;
        RECT 16.070 41.260 16.330 41.580 ;
        RECT 13.760 40.045 14.040 40.415 ;
        RECT 16.130 40.220 16.270 41.260 ;
        RECT 21.130 40.920 21.390 41.240 ;
        RECT 21.590 40.920 21.850 41.240 ;
        RECT 13.770 39.900 14.030 40.045 ;
        RECT 16.070 39.900 16.330 40.220 ;
        RECT 21.190 39.540 21.330 40.920 ;
        RECT 21.650 40.220 21.790 40.920 ;
        RECT 23.950 40.220 24.090 41.600 ;
        RECT 21.590 39.900 21.850 40.220 ;
        RECT 23.890 39.900 24.150 40.220 ;
        RECT 21.130 39.220 21.390 39.540 ;
        RECT 19.750 38.880 20.010 39.200 ;
        RECT 16.530 38.540 16.790 38.860 ;
        RECT 16.590 36.820 16.730 38.540 ;
        RECT 16.530 36.500 16.790 36.820 ;
        RECT 19.810 36.140 19.950 38.880 ;
        RECT 23.950 36.480 24.090 39.900 ;
        RECT 21.130 36.160 21.390 36.480 ;
        RECT 23.890 36.160 24.150 36.480 ;
        RECT 19.750 35.820 20.010 36.140 ;
        RECT 14.230 35.480 14.490 35.800 ;
        RECT 18.830 35.480 19.090 35.800 ;
        RECT 14.290 34.440 14.430 35.480 ;
        RECT 14.230 34.120 14.490 34.440 ;
        RECT 13.760 33.245 14.040 33.615 ;
        RECT 13.830 29.340 13.970 33.245 ;
        RECT 14.230 32.760 14.490 33.080 ;
        RECT 14.290 31.380 14.430 32.760 ;
        RECT 18.890 32.060 19.030 35.480 ;
        RECT 18.830 31.740 19.090 32.060 ;
        RECT 14.230 31.060 14.490 31.380 ;
        RECT 13.770 29.020 14.030 29.340 ;
        RECT 14.290 28.660 14.430 31.060 ;
        RECT 19.290 30.040 19.550 30.360 ;
        RECT 19.350 29.340 19.490 30.040 ;
        RECT 19.290 29.020 19.550 29.340 ;
        RECT 14.230 28.340 14.490 28.660 ;
        RECT 19.810 28.320 19.950 35.820 ;
        RECT 21.190 34.100 21.330 36.160 ;
        RECT 24.870 34.440 25.010 43.445 ;
        RECT 26.250 42.940 26.390 44.660 ;
        RECT 26.190 42.620 26.450 42.940 ;
        RECT 26.190 39.900 26.450 40.220 ;
        RECT 27.110 39.900 27.370 40.220 ;
        RECT 26.250 36.820 26.390 39.900 ;
        RECT 27.170 37.500 27.310 39.900 ;
        RECT 27.110 37.180 27.370 37.500 ;
        RECT 26.190 36.500 26.450 36.820 ;
        RECT 24.810 34.120 25.070 34.440 ;
        RECT 21.130 33.780 21.390 34.100 ;
        RECT 27.170 32.060 27.310 37.180 ;
        RECT 27.630 32.060 27.770 44.805 ;
        RECT 28.300 43.105 29.840 43.475 ;
        RECT 30.390 41.920 30.530 46.360 ;
        RECT 30.850 44.300 30.990 49.680 ;
        RECT 33.150 48.380 33.290 56.255 ;
        RECT 33.090 48.060 33.350 48.380 ;
        RECT 31.250 47.720 31.510 48.040 ;
        RECT 30.790 43.980 31.050 44.300 ;
        RECT 31.310 42.940 31.450 47.720 ;
        RECT 36.370 47.360 36.510 56.255 ;
        RECT 39.590 48.380 39.730 56.255 ;
        RECT 46.880 53.645 47.160 54.015 ;
        RECT 44.120 50.245 44.400 50.615 ;
        RECT 39.530 48.060 39.790 48.380 ;
        RECT 38.150 47.720 38.410 48.040 ;
        RECT 33.550 47.040 33.810 47.360 ;
        RECT 36.310 47.040 36.570 47.360 ;
        RECT 31.600 45.825 33.140 46.195 ;
        RECT 33.610 45.660 33.750 47.040 ;
        RECT 34.010 46.360 34.270 46.680 ;
        RECT 33.550 45.340 33.810 45.660 ;
        RECT 34.070 45.320 34.210 46.360 ;
        RECT 34.010 45.000 34.270 45.320 ;
        RECT 38.210 44.980 38.350 47.720 ;
        RECT 44.190 47.360 44.330 50.245 ;
        RECT 46.950 47.360 47.090 53.645 ;
        RECT 41.370 47.040 41.630 47.360 ;
        RECT 44.130 47.040 44.390 47.360 ;
        RECT 45.510 47.215 45.770 47.360 ;
        RECT 39.990 46.360 40.250 46.680 ;
        RECT 34.930 44.660 35.190 44.980 ;
        RECT 36.310 44.660 36.570 44.980 ;
        RECT 38.150 44.660 38.410 44.980 ;
        RECT 31.710 44.320 31.970 44.640 ;
        RECT 31.250 42.620 31.510 42.940 ;
        RECT 31.770 41.920 31.910 44.320 ;
        RECT 34.470 43.640 34.730 43.960 ;
        RECT 34.530 42.260 34.670 43.640 ;
        RECT 34.470 41.940 34.730 42.260 ;
        RECT 34.990 41.920 35.130 44.660 ;
        RECT 35.850 44.320 36.110 44.640 ;
        RECT 30.330 41.600 30.590 41.920 ;
        RECT 30.790 41.600 31.050 41.920 ;
        RECT 31.710 41.600 31.970 41.920 ;
        RECT 33.550 41.600 33.810 41.920 ;
        RECT 34.010 41.600 34.270 41.920 ;
        RECT 34.930 41.600 35.190 41.920 ;
        RECT 30.330 40.920 30.590 41.240 ;
        RECT 28.300 37.665 29.840 38.035 ;
        RECT 28.300 32.225 29.840 32.595 ;
        RECT 27.110 31.740 27.370 32.060 ;
        RECT 27.570 31.740 27.830 32.060 ;
        RECT 22.050 30.720 22.310 31.040 ;
        RECT 19.290 28.000 19.550 28.320 ;
        RECT 19.750 28.000 20.010 28.320 ;
        RECT 14.230 27.660 14.490 27.980 ;
        RECT 13.760 26.445 14.040 26.815 ;
        RECT 13.830 22.540 13.970 26.445 ;
        RECT 14.290 25.940 14.430 27.660 ;
        RECT 16.530 27.320 16.790 27.640 ;
        RECT 14.230 25.620 14.490 25.940 ;
        RECT 16.590 25.260 16.730 27.320 ;
        RECT 16.530 24.940 16.790 25.260 ;
        RECT 14.230 22.560 14.490 22.880 ;
        RECT 13.770 22.220 14.030 22.540 ;
        RECT 14.290 21.180 14.430 22.560 ;
        RECT 19.350 22.540 19.490 28.000 ;
        RECT 22.110 26.620 22.250 30.720 ;
        RECT 27.170 29.000 27.310 31.740 ;
        RECT 30.390 31.040 30.530 40.920 ;
        RECT 30.850 40.220 30.990 41.600 ;
        RECT 31.600 40.385 33.140 40.755 ;
        RECT 30.790 39.900 31.050 40.220 ;
        RECT 30.790 39.220 31.050 39.540 ;
        RECT 30.850 33.080 30.990 39.220 ;
        RECT 31.250 38.200 31.510 38.520 ;
        RECT 31.310 34.180 31.450 38.200 ;
        RECT 33.610 37.500 33.750 41.600 ;
        RECT 33.550 37.180 33.810 37.500 ;
        RECT 34.070 36.900 34.210 41.600 ;
        RECT 35.910 39.880 36.050 44.320 ;
        RECT 36.370 42.940 36.510 44.660 ;
        RECT 37.230 43.640 37.490 43.960 ;
        RECT 36.310 42.620 36.570 42.940 ;
        RECT 36.370 42.340 36.510 42.620 ;
        RECT 36.370 42.200 36.970 42.340 ;
        RECT 36.310 41.260 36.570 41.580 ;
        RECT 35.850 39.560 36.110 39.880 ;
        RECT 34.470 38.880 34.730 39.200 ;
        RECT 33.610 36.760 34.210 36.900 ;
        RECT 33.610 35.800 33.750 36.760 ;
        RECT 34.530 36.480 34.670 38.880 ;
        RECT 34.930 36.840 35.190 37.160 ;
        RECT 34.470 36.160 34.730 36.480 ;
        RECT 34.010 35.820 34.270 36.140 ;
        RECT 33.550 35.480 33.810 35.800 ;
        RECT 31.600 34.945 33.140 35.315 ;
        RECT 31.310 34.040 31.910 34.180 ;
        RECT 31.250 33.440 31.510 33.760 ;
        RECT 30.790 32.760 31.050 33.080 ;
        RECT 27.570 30.720 27.830 31.040 ;
        RECT 30.330 30.720 30.590 31.040 ;
        RECT 27.630 29.340 27.770 30.720 ;
        RECT 27.570 29.020 27.830 29.340 ;
        RECT 25.730 28.680 25.990 29.000 ;
        RECT 27.110 28.680 27.370 29.000 ;
        RECT 22.050 26.300 22.310 26.620 ;
        RECT 21.130 25.280 21.390 25.600 ;
        RECT 19.290 22.220 19.550 22.540 ;
        RECT 18.830 21.880 19.090 22.200 ;
        RECT 14.230 20.860 14.490 21.180 ;
        RECT 14.290 17.780 14.430 20.860 ;
        RECT 16.990 19.500 17.250 19.820 ;
        RECT 17.050 18.460 17.190 19.500 ;
        RECT 18.890 18.460 19.030 21.880 ;
        RECT 19.350 18.460 19.490 22.220 ;
        RECT 21.190 20.500 21.330 25.280 ;
        RECT 22.110 23.220 22.250 26.300 ;
        RECT 22.050 22.900 22.310 23.220 ;
        RECT 25.790 22.880 25.930 28.680 ;
        RECT 27.110 27.660 27.370 27.980 ;
        RECT 27.170 25.260 27.310 27.660 ;
        RECT 28.300 26.785 29.840 27.155 ;
        RECT 27.110 24.940 27.370 25.260 ;
        RECT 21.590 22.560 21.850 22.880 ;
        RECT 25.730 22.560 25.990 22.880 ;
        RECT 21.130 20.180 21.390 20.500 ;
        RECT 21.650 18.460 21.790 22.560 ;
        RECT 16.990 18.140 17.250 18.460 ;
        RECT 18.830 18.140 19.090 18.460 ;
        RECT 19.290 18.140 19.550 18.460 ;
        RECT 21.590 18.140 21.850 18.460 ;
        RECT 23.890 18.140 24.150 18.460 ;
        RECT 14.230 17.460 14.490 17.780 ;
        RECT 11.460 16.925 11.740 17.295 ;
        RECT 11.470 16.780 11.730 16.925 ;
        RECT 23.950 14.720 24.090 18.140 ;
        RECT 25.790 17.440 25.930 22.560 ;
        RECT 30.330 21.880 30.590 22.200 ;
        RECT 28.300 21.345 29.840 21.715 ;
        RECT 30.390 18.460 30.530 21.880 ;
        RECT 30.850 20.160 30.990 32.760 ;
        RECT 31.310 31.040 31.450 33.440 ;
        RECT 31.770 31.720 31.910 34.040 ;
        RECT 31.710 31.400 31.970 31.720 ;
        RECT 31.250 30.720 31.510 31.040 ;
        RECT 31.600 29.505 33.140 29.875 ;
        RECT 33.610 28.320 33.750 35.480 ;
        RECT 34.070 34.780 34.210 35.820 ;
        RECT 34.010 34.460 34.270 34.780 ;
        RECT 34.990 31.380 35.130 36.840 ;
        RECT 35.390 35.820 35.650 36.140 ;
        RECT 34.930 31.060 35.190 31.380 ;
        RECT 34.470 29.250 34.730 29.340 ;
        RECT 34.990 29.250 35.130 31.060 ;
        RECT 34.470 29.110 35.130 29.250 ;
        RECT 34.470 29.020 34.730 29.110 ;
        RECT 33.550 28.000 33.810 28.320 ;
        RECT 34.010 28.000 34.270 28.320 ;
        RECT 34.070 24.920 34.210 28.000 ;
        RECT 34.990 26.020 35.130 29.110 ;
        RECT 35.450 26.280 35.590 35.820 ;
        RECT 35.910 33.080 36.050 39.560 ;
        RECT 36.370 38.860 36.510 41.260 ;
        RECT 36.310 38.540 36.570 38.860 ;
        RECT 36.370 34.780 36.510 38.540 ;
        RECT 36.310 34.460 36.570 34.780 ;
        RECT 35.850 32.760 36.110 33.080 ;
        RECT 35.910 31.720 36.050 32.760 ;
        RECT 35.850 31.400 36.110 31.720 ;
        RECT 35.850 27.660 36.110 27.980 ;
        RECT 34.530 25.940 35.130 26.020 ;
        RECT 35.390 25.960 35.650 26.280 ;
        RECT 34.470 25.880 35.130 25.940 ;
        RECT 34.470 25.620 34.730 25.880 ;
        RECT 31.250 24.600 31.510 24.920 ;
        RECT 34.010 24.600 34.270 24.920 ;
        RECT 31.310 23.220 31.450 24.600 ;
        RECT 31.600 24.065 33.140 24.435 ;
        RECT 31.250 22.900 31.510 23.220 ;
        RECT 31.310 21.180 31.450 22.900 ;
        RECT 31.250 20.860 31.510 21.180 ;
        RECT 30.790 19.840 31.050 20.160 ;
        RECT 30.330 18.140 30.590 18.460 ;
        RECT 31.310 18.120 31.450 20.860 ;
        RECT 31.600 18.625 33.140 18.995 ;
        RECT 31.250 17.860 31.510 18.120 ;
        RECT 30.390 17.800 31.510 17.860 ;
        RECT 30.390 17.720 31.450 17.800 ;
        RECT 25.730 17.120 25.990 17.440 ;
        RECT 28.300 15.905 29.840 16.275 ;
        RECT 23.890 14.400 24.150 14.720 ;
        RECT 28.950 14.630 29.210 14.720 ;
        RECT 30.390 14.630 30.530 17.720 ;
        RECT 31.250 16.440 31.510 16.760 ;
        RECT 28.950 14.490 30.530 14.630 ;
        RECT 28.950 14.400 29.210 14.490 ;
        RECT 31.310 14.380 31.450 16.440 ;
        RECT 34.070 15.740 34.210 24.600 ;
        RECT 35.910 23.560 36.050 27.660 ;
        RECT 36.830 26.620 36.970 42.200 ;
        RECT 37.290 41.920 37.430 43.640 ;
        RECT 37.230 41.600 37.490 41.920 ;
        RECT 40.050 39.540 40.190 46.360 ;
        RECT 40.900 44.890 41.180 45.175 ;
        RECT 40.510 44.805 41.180 44.890 ;
        RECT 40.510 44.750 41.170 44.805 ;
        RECT 40.510 39.880 40.650 44.750 ;
        RECT 40.910 44.660 41.170 44.750 ;
        RECT 41.430 44.300 41.570 47.040 ;
        RECT 45.500 46.845 45.780 47.215 ;
        RECT 46.890 47.040 47.150 47.360 ;
        RECT 43.670 46.360 43.930 46.680 ;
        RECT 46.430 46.360 46.690 46.680 ;
        RECT 41.370 43.980 41.630 44.300 ;
        RECT 41.430 42.940 41.570 43.980 ;
        RECT 43.210 43.640 43.470 43.960 ;
        RECT 41.370 42.620 41.630 42.940 ;
        RECT 43.270 41.920 43.410 43.640 ;
        RECT 43.210 41.600 43.470 41.920 ;
        RECT 43.730 40.220 43.870 46.360 ;
        RECT 44.130 44.660 44.390 44.980 ;
        RECT 44.190 42.940 44.330 44.660 ;
        RECT 44.590 43.980 44.850 44.300 ;
        RECT 44.130 42.620 44.390 42.940 ;
        RECT 44.650 42.340 44.790 43.980 ;
        RECT 44.190 42.200 44.790 42.340 ;
        RECT 43.670 39.900 43.930 40.220 ;
        RECT 40.450 39.560 40.710 39.880 ;
        RECT 40.910 39.560 41.170 39.880 ;
        RECT 39.990 39.220 40.250 39.540 ;
        RECT 38.150 38.200 38.410 38.520 ;
        RECT 38.210 32.060 38.350 38.200 ;
        RECT 39.070 35.480 39.330 35.800 ;
        RECT 39.130 34.100 39.270 35.480 ;
        RECT 40.050 34.100 40.190 39.220 ;
        RECT 40.970 38.860 41.110 39.560 ;
        RECT 43.730 39.540 43.870 39.900 ;
        RECT 43.670 39.220 43.930 39.540 ;
        RECT 40.910 38.540 41.170 38.860 ;
        RECT 40.970 36.480 41.110 38.540 ;
        RECT 41.830 36.840 42.090 37.160 ;
        RECT 40.910 36.160 41.170 36.480 ;
        RECT 39.070 33.780 39.330 34.100 ;
        RECT 39.990 33.780 40.250 34.100 ;
        RECT 38.150 31.740 38.410 32.060 ;
        RECT 37.690 30.040 37.950 30.360 ;
        RECT 36.770 26.300 37.030 26.620 ;
        RECT 35.850 23.240 36.110 23.560 ;
        RECT 35.910 18.460 36.050 23.240 ;
        RECT 36.830 23.220 36.970 26.300 ;
        RECT 36.770 22.900 37.030 23.220 ;
        RECT 35.850 18.140 36.110 18.460 ;
        RECT 36.830 17.440 36.970 22.900 ;
        RECT 37.750 22.880 37.890 30.040 ;
        RECT 38.210 28.660 38.350 31.740 ;
        RECT 41.890 31.460 42.030 36.840 ;
        RECT 42.750 36.500 43.010 36.820 ;
        RECT 42.290 32.760 42.550 33.080 ;
        RECT 40.970 31.320 42.030 31.460 ;
        RECT 40.970 31.040 41.110 31.320 ;
        RECT 40.910 30.720 41.170 31.040 ;
        RECT 41.830 30.720 42.090 31.040 ;
        RECT 40.450 30.040 40.710 30.360 ;
        RECT 41.890 30.215 42.030 30.720 ;
        RECT 42.350 30.700 42.490 32.760 ;
        RECT 42.290 30.380 42.550 30.700 ;
        RECT 40.510 28.660 40.650 30.040 ;
        RECT 41.820 29.845 42.100 30.215 ;
        RECT 42.350 29.000 42.490 30.380 ;
        RECT 42.290 28.680 42.550 29.000 ;
        RECT 38.150 28.340 38.410 28.660 ;
        RECT 40.450 28.340 40.710 28.660 ;
        RECT 39.520 26.445 39.800 26.815 ;
        RECT 37.690 22.560 37.950 22.880 ;
        RECT 37.750 22.200 37.890 22.560 ;
        RECT 37.690 21.880 37.950 22.200 ;
        RECT 39.590 20.160 39.730 26.445 ;
        RECT 42.350 25.940 42.490 28.680 ;
        RECT 42.810 26.620 42.950 36.500 ;
        RECT 43.730 36.480 43.870 39.220 ;
        RECT 44.190 36.480 44.330 42.200 ;
        RECT 44.590 41.600 44.850 41.920 ;
        RECT 44.650 37.015 44.790 41.600 ;
        RECT 45.510 40.920 45.770 41.240 ;
        RECT 45.970 40.920 46.230 41.240 ;
        RECT 45.050 39.220 45.310 39.540 ;
        RECT 45.110 37.500 45.250 39.220 ;
        RECT 45.050 37.180 45.310 37.500 ;
        RECT 44.580 36.645 44.860 37.015 ;
        RECT 45.570 36.900 45.710 40.920 ;
        RECT 46.030 40.220 46.170 40.920 ;
        RECT 45.970 39.900 46.230 40.220 ;
        RECT 46.490 39.540 46.630 46.360 ;
        RECT 46.890 44.660 47.150 44.980 ;
        RECT 46.950 43.815 47.090 44.660 ;
        RECT 46.880 43.445 47.160 43.815 ;
        RECT 46.890 41.600 47.150 41.920 ;
        RECT 46.950 40.415 47.090 41.600 ;
        RECT 46.880 40.045 47.160 40.415 ;
        RECT 46.430 39.220 46.690 39.540 ;
        RECT 46.490 37.160 46.630 39.220 ;
        RECT 45.570 36.760 46.170 36.900 ;
        RECT 46.430 36.840 46.690 37.160 ;
        RECT 46.030 36.480 46.170 36.760 ;
        RECT 43.670 36.160 43.930 36.480 ;
        RECT 44.130 36.160 44.390 36.480 ;
        RECT 45.510 36.160 45.770 36.480 ;
        RECT 45.970 36.160 46.230 36.480 ;
        RECT 44.190 31.720 44.330 36.160 ;
        RECT 44.590 33.780 44.850 34.100 ;
        RECT 44.130 31.400 44.390 31.720 ;
        RECT 44.650 31.040 44.790 33.780 ;
        RECT 45.570 32.060 45.710 36.160 ;
        RECT 46.030 34.100 46.170 36.160 ;
        RECT 45.970 33.780 46.230 34.100 ;
        RECT 46.890 33.780 47.150 34.100 ;
        RECT 46.950 33.615 47.090 33.780 ;
        RECT 46.880 33.245 47.160 33.615 ;
        RECT 45.510 31.740 45.770 32.060 ;
        RECT 44.130 30.720 44.390 31.040 ;
        RECT 44.590 30.720 44.850 31.040 ;
        RECT 44.190 29.340 44.330 30.720 ;
        RECT 45.050 30.380 45.310 30.700 ;
        RECT 44.130 29.020 44.390 29.340 ;
        RECT 43.670 28.340 43.930 28.660 ;
        RECT 44.130 28.340 44.390 28.660 ;
        RECT 42.750 26.300 43.010 26.620 ;
        RECT 42.290 25.620 42.550 25.940 ;
        RECT 39.990 25.280 40.250 25.600 ;
        RECT 42.750 25.280 43.010 25.600 ;
        RECT 40.050 22.200 40.190 25.280 ;
        RECT 40.910 24.600 41.170 24.920 ;
        RECT 40.970 23.900 41.110 24.600 ;
        RECT 40.910 23.580 41.170 23.900 ;
        RECT 42.810 22.880 42.950 25.280 ;
        RECT 43.200 23.045 43.480 23.415 ;
        RECT 43.210 22.900 43.470 23.045 ;
        RECT 42.750 22.560 43.010 22.880 ;
        RECT 39.990 21.880 40.250 22.200 ;
        RECT 38.150 19.840 38.410 20.160 ;
        RECT 39.530 19.840 39.790 20.160 ;
        RECT 36.770 17.120 37.030 17.440 ;
        RECT 37.230 17.120 37.490 17.440 ;
        RECT 34.010 15.420 34.270 15.740 ;
        RECT 37.290 15.400 37.430 17.120 ;
        RECT 38.210 16.615 38.350 19.840 ;
        RECT 38.140 16.245 38.420 16.615 ;
        RECT 37.230 15.080 37.490 15.400 ;
        RECT 37.290 14.720 37.430 15.080 ;
        RECT 40.050 14.720 40.190 21.880 ;
        RECT 42.810 21.180 42.950 22.560 ;
        RECT 43.730 22.200 43.870 28.340 ;
        RECT 43.670 21.880 43.930 22.200 ;
        RECT 42.750 20.860 43.010 21.180 ;
        RECT 43.210 20.520 43.470 20.840 ;
        RECT 40.910 20.015 41.170 20.160 ;
        RECT 40.900 19.645 41.180 20.015 ;
        RECT 42.290 19.160 42.550 19.480 ;
        RECT 42.750 19.160 43.010 19.480 ;
        RECT 42.350 17.440 42.490 19.160 ;
        RECT 42.810 17.780 42.950 19.160 ;
        RECT 42.750 17.460 43.010 17.780 ;
        RECT 42.290 17.120 42.550 17.440 ;
        RECT 42.350 15.060 42.490 17.120 ;
        RECT 43.270 15.400 43.410 20.520 ;
        RECT 43.730 20.160 43.870 21.880 ;
        RECT 44.190 21.180 44.330 28.340 ;
        RECT 44.590 28.000 44.850 28.320 ;
        RECT 44.650 23.900 44.790 28.000 ;
        RECT 45.110 25.600 45.250 30.380 ;
        RECT 45.970 28.340 46.230 28.660 ;
        RECT 45.050 25.280 45.310 25.600 ;
        RECT 45.510 25.280 45.770 25.600 ;
        RECT 44.590 23.580 44.850 23.900 ;
        RECT 45.110 23.560 45.250 25.280 ;
        RECT 45.050 23.240 45.310 23.560 ;
        RECT 44.590 22.900 44.850 23.220 ;
        RECT 44.130 20.860 44.390 21.180 ;
        RECT 44.650 20.160 44.790 22.900 ;
        RECT 43.670 19.840 43.930 20.160 ;
        RECT 44.590 19.840 44.850 20.160 ;
        RECT 43.730 15.740 43.870 19.840 ;
        RECT 45.570 18.460 45.710 25.280 ;
        RECT 46.030 22.880 46.170 28.340 ;
        RECT 45.970 22.560 46.230 22.880 ;
        RECT 46.890 22.220 47.150 22.540 ;
        RECT 46.430 20.180 46.690 20.500 ;
        RECT 45.970 19.840 46.230 20.160 ;
        RECT 45.510 18.140 45.770 18.460 ;
        RECT 46.030 15.740 46.170 19.840 ;
        RECT 43.670 15.420 43.930 15.740 ;
        RECT 45.970 15.420 46.230 15.740 ;
        RECT 43.210 15.080 43.470 15.400 ;
        RECT 42.290 14.740 42.550 15.060 ;
        RECT 37.230 14.400 37.490 14.720 ;
        RECT 39.990 14.400 40.250 14.720 ;
        RECT 42.750 14.400 43.010 14.720 ;
        RECT 31.250 14.060 31.510 14.380 ;
        RECT 26.650 13.720 26.910 14.040 ;
        RECT 29.410 13.720 29.670 14.040 ;
        RECT 33.550 13.720 33.810 14.040 ;
        RECT 39.530 13.720 39.790 14.040 ;
        RECT 26.710 6.490 26.850 13.720 ;
        RECT 29.470 8.340 29.610 13.720 ;
        RECT 31.600 13.185 33.140 13.555 ;
        RECT 33.610 8.340 33.750 13.720 ;
        RECT 29.470 8.200 30.070 8.340 ;
        RECT 29.930 6.490 30.070 8.200 ;
        RECT 33.150 8.200 33.750 8.340 ;
        RECT 33.150 6.490 33.290 8.200 ;
        RECT 39.590 6.490 39.730 13.720 ;
        RECT 42.810 13.215 42.950 14.400 ;
        RECT 42.740 12.845 43.020 13.215 ;
        RECT 46.490 9.815 46.630 20.180 ;
        RECT 46.950 20.160 47.090 22.220 ;
        RECT 46.890 19.840 47.150 20.160 ;
        RECT 46.950 17.440 47.090 19.840 ;
        RECT 46.890 17.120 47.150 17.440 ;
        RECT 46.420 9.445 46.700 9.815 ;
        RECT 26.640 2.490 26.920 6.490 ;
        RECT 29.860 2.490 30.140 6.490 ;
        RECT 33.080 2.490 33.360 6.490 ;
        RECT 39.520 2.490 39.800 6.490 ;
      LAYER met3 ;
        RECT 46.855 53.980 47.185 53.995 ;
        RECT 50.275 53.980 54.275 54.130 ;
        RECT 46.855 53.680 54.275 53.980 ;
        RECT 46.855 53.665 47.185 53.680 ;
        RECT 50.275 53.530 54.275 53.680 ;
        RECT 44.095 50.580 44.425 50.595 ;
        RECT 50.275 50.580 54.275 50.730 ;
        RECT 44.095 50.280 54.275 50.580 ;
        RECT 44.095 50.265 44.425 50.280 ;
        RECT 50.275 50.130 54.275 50.280 ;
        RECT 28.280 48.565 29.860 48.895 ;
        RECT 45.475 47.180 45.805 47.195 ;
        RECT 50.275 47.180 54.275 47.330 ;
        RECT 45.475 46.880 54.275 47.180 ;
        RECT 45.475 46.865 45.805 46.880 ;
        RECT 50.275 46.730 54.275 46.880 ;
        RECT 31.580 45.845 33.160 46.175 ;
        RECT 23.395 45.140 23.725 45.155 ;
        RECT 27.535 45.140 27.865 45.155 ;
        RECT 40.875 45.140 41.205 45.155 ;
        RECT 23.395 44.840 41.205 45.140 ;
        RECT 23.395 44.825 23.725 44.840 ;
        RECT 27.535 44.825 27.865 44.840 ;
        RECT 40.875 44.825 41.205 44.840 ;
        RECT 7.230 43.780 11.230 43.930 ;
        RECT 24.775 43.780 25.105 43.795 ;
        RECT 7.230 43.480 25.105 43.780 ;
        RECT 7.230 43.330 11.230 43.480 ;
        RECT 24.775 43.465 25.105 43.480 ;
        RECT 46.855 43.780 47.185 43.795 ;
        RECT 50.275 43.780 54.275 43.930 ;
        RECT 46.855 43.480 54.275 43.780 ;
        RECT 46.855 43.465 47.185 43.480 ;
        RECT 28.280 43.125 29.860 43.455 ;
        RECT 50.275 43.330 54.275 43.480 ;
        RECT 7.230 40.380 11.230 40.530 ;
        RECT 31.580 40.405 33.160 40.735 ;
        RECT 13.735 40.380 14.065 40.395 ;
        RECT 7.230 40.080 14.065 40.380 ;
        RECT 7.230 39.930 11.230 40.080 ;
        RECT 13.735 40.065 14.065 40.080 ;
        RECT 46.855 40.380 47.185 40.395 ;
        RECT 50.275 40.380 54.275 40.530 ;
        RECT 46.855 40.080 54.275 40.380 ;
        RECT 46.855 40.065 47.185 40.080 ;
        RECT 50.275 39.930 54.275 40.080 ;
        RECT 28.280 37.685 29.860 38.015 ;
        RECT 44.555 36.980 44.885 36.995 ;
        RECT 50.275 36.980 54.275 37.130 ;
        RECT 44.555 36.680 54.275 36.980 ;
        RECT 44.555 36.665 44.885 36.680 ;
        RECT 50.275 36.530 54.275 36.680 ;
        RECT 31.580 34.965 33.160 35.295 ;
        RECT 7.230 33.580 11.230 33.730 ;
        RECT 13.735 33.580 14.065 33.595 ;
        RECT 7.230 33.280 14.065 33.580 ;
        RECT 7.230 33.130 11.230 33.280 ;
        RECT 13.735 33.265 14.065 33.280 ;
        RECT 46.855 33.580 47.185 33.595 ;
        RECT 50.275 33.580 54.275 33.730 ;
        RECT 46.855 33.280 54.275 33.580 ;
        RECT 46.855 33.265 47.185 33.280 ;
        RECT 50.275 33.130 54.275 33.280 ;
        RECT 28.280 32.245 29.860 32.575 ;
        RECT 41.795 30.180 42.125 30.195 ;
        RECT 50.275 30.180 54.275 30.330 ;
        RECT 41.795 29.880 54.275 30.180 ;
        RECT 41.795 29.865 42.125 29.880 ;
        RECT 31.580 29.525 33.160 29.855 ;
        RECT 50.275 29.730 54.275 29.880 ;
        RECT 7.230 26.780 11.230 26.930 ;
        RECT 28.280 26.805 29.860 27.135 ;
        RECT 13.735 26.780 14.065 26.795 ;
        RECT 7.230 26.480 14.065 26.780 ;
        RECT 7.230 26.330 11.230 26.480 ;
        RECT 13.735 26.465 14.065 26.480 ;
        RECT 39.495 26.780 39.825 26.795 ;
        RECT 50.275 26.780 54.275 26.930 ;
        RECT 39.495 26.480 54.275 26.780 ;
        RECT 39.495 26.465 39.825 26.480 ;
        RECT 50.275 26.330 54.275 26.480 ;
        RECT 31.580 24.085 33.160 24.415 ;
        RECT 43.175 23.380 43.505 23.395 ;
        RECT 50.275 23.380 54.275 23.530 ;
        RECT 43.175 23.080 54.275 23.380 ;
        RECT 43.175 23.065 43.505 23.080 ;
        RECT 50.275 22.930 54.275 23.080 ;
        RECT 28.280 21.365 29.860 21.695 ;
        RECT 40.875 19.980 41.205 19.995 ;
        RECT 50.275 19.980 54.275 20.130 ;
        RECT 40.875 19.680 54.275 19.980 ;
        RECT 40.875 19.665 41.205 19.680 ;
        RECT 50.275 19.530 54.275 19.680 ;
        RECT 31.580 18.645 33.160 18.975 ;
        RECT 11.435 17.260 11.765 17.275 ;
        RECT 11.220 16.945 11.765 17.260 ;
        RECT 11.220 16.730 11.520 16.945 ;
        RECT 7.230 16.280 11.520 16.730 ;
        RECT 38.115 16.580 38.445 16.595 ;
        RECT 50.275 16.580 54.275 16.730 ;
        RECT 38.115 16.280 54.275 16.580 ;
        RECT 7.230 16.130 11.230 16.280 ;
        RECT 38.115 16.265 38.445 16.280 ;
        RECT 28.280 15.925 29.860 16.255 ;
        RECT 50.275 16.130 54.275 16.280 ;
        RECT 31.580 13.205 33.160 13.535 ;
        RECT 42.715 13.180 43.045 13.195 ;
        RECT 50.275 13.180 54.275 13.330 ;
        RECT 42.715 12.880 54.275 13.180 ;
        RECT 42.715 12.865 43.045 12.880 ;
        RECT 50.275 12.730 54.275 12.880 ;
        RECT 46.395 9.780 46.725 9.795 ;
        RECT 50.275 9.780 54.275 9.930 ;
        RECT 46.395 9.480 54.275 9.780 ;
        RECT 46.395 9.465 46.725 9.480 ;
        RECT 50.275 9.330 54.275 9.480 ;
      LAYER met4 ;
        RECT 64.090 225.055 64.145 225.385 ;
        RECT 66.455 224.965 66.550 225.295 ;
        RECT 69.305 225.135 69.310 225.465 ;
        RECT 69.610 225.135 69.635 225.465 ;
        RECT 71.995 224.895 72.070 225.225 ;
        RECT 74.785 224.945 74.830 225.275 ;
        RECT 77.515 224.760 77.590 225.085 ;
        RECT 80.295 224.925 80.350 225.255 ;
        RECT 83.025 224.760 83.110 225.085 ;
        RECT 85.795 224.915 85.870 225.245 ;
        RECT 88.535 224.915 88.630 225.245 ;
        RECT 91.350 224.835 91.390 225.165 ;
        RECT 94.125 224.815 94.150 225.145 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 77.515 224.755 77.845 224.760 ;
        RECT 83.025 224.755 83.355 224.760 ;
        RECT 6.000 197.560 6.140 199.160 ;
        RECT 28.270 13.130 29.870 48.970 ;
        RECT 31.570 13.130 33.170 48.970 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

