VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 110.585 217.835 111.395 217.975 ;
        RECT 110.395 217.665 111.395 217.835 ;
        RECT 110.585 216.605 111.395 217.665 ;
        RECT 110.585 216.455 111.395 216.595 ;
        RECT 110.395 216.285 111.395 216.455 ;
        RECT 110.585 211.085 111.395 216.285 ;
        RECT 110.585 210.935 111.395 211.075 ;
        RECT 110.395 210.765 111.395 210.935 ;
        RECT 110.585 207.405 111.395 210.765 ;
        RECT 110.425 207.140 110.535 207.260 ;
        RECT 110.585 206.795 111.265 206.935 ;
        RECT 110.395 206.625 111.265 206.795 ;
        RECT 110.585 206.450 111.265 206.625 ;
        RECT 110.585 205.105 111.495 206.450 ;
        RECT 110.670 204.655 111.455 205.085 ;
        RECT 110.425 204.380 110.535 204.500 ;
        RECT 110.585 202.830 111.495 204.175 ;
        RECT 110.585 202.655 111.265 202.830 ;
        RECT 110.395 202.485 111.265 202.655 ;
        RECT 110.585 202.345 111.265 202.485 ;
        RECT 110.585 202.195 111.265 202.335 ;
        RECT 110.395 202.025 111.265 202.195 ;
        RECT 110.585 198.820 111.265 202.025 ;
        RECT 110.585 197.910 111.485 198.820 ;
        RECT 110.585 196.375 111.265 197.910 ;
        RECT 110.585 195.025 111.495 196.375 ;
        RECT 110.585 193.630 111.495 194.975 ;
        RECT 110.585 193.455 111.265 193.630 ;
        RECT 110.395 193.285 111.265 193.455 ;
        RECT 110.585 193.145 111.265 193.285 ;
        RECT 110.430 192.825 110.540 192.985 ;
        RECT 110.670 191.775 111.455 192.205 ;
        RECT 110.430 191.445 110.540 191.605 ;
        RECT 110.585 190.695 111.265 190.835 ;
        RECT 110.395 190.525 111.265 190.695 ;
        RECT 110.585 190.350 111.265 190.525 ;
        RECT 110.585 189.005 111.495 190.350 ;
        RECT 110.585 187.945 111.365 188.995 ;
        RECT 110.395 187.775 111.365 187.945 ;
        RECT 110.585 187.625 111.365 187.775 ;
        RECT 110.430 187.305 110.540 187.465 ;
        RECT 110.585 186.555 111.265 186.695 ;
        RECT 110.395 186.385 111.265 186.555 ;
        RECT 110.585 184.875 111.265 186.385 ;
        RECT 110.585 183.945 111.495 184.875 ;
        RECT 110.425 183.680 110.535 183.800 ;
        RECT 110.585 182.415 111.395 183.475 ;
        RECT 110.395 182.245 111.395 182.415 ;
        RECT 110.585 182.105 111.395 182.245 ;
      LAYER nwell ;
        RECT 111.785 181.910 114.615 218.170 ;
      LAYER pwell ;
        RECT 115.005 217.835 115.815 217.975 ;
        RECT 116.025 217.835 116.835 217.975 ;
        RECT 115.005 217.665 116.835 217.835 ;
        RECT 115.005 216.605 115.815 217.665 ;
        RECT 116.025 216.605 116.835 217.665 ;
        RECT 114.905 215.250 115.815 216.595 ;
        RECT 115.135 215.075 115.815 215.250 ;
        RECT 116.025 215.205 116.935 216.555 ;
        RECT 115.135 214.905 116.005 215.075 ;
        RECT 115.135 214.765 115.815 214.905 ;
        RECT 115.860 214.445 115.970 214.605 ;
        RECT 114.905 213.420 115.815 213.835 ;
        RECT 116.025 213.670 116.705 215.205 ;
        RECT 114.905 213.250 116.005 213.420 ;
        RECT 114.905 212.905 115.815 213.250 ;
        RECT 115.135 209.935 115.815 212.905 ;
        RECT 116.025 212.760 116.925 213.670 ;
        RECT 115.005 209.555 115.815 209.695 ;
        RECT 116.025 209.555 116.705 212.760 ;
        RECT 115.005 209.385 116.705 209.555 ;
        RECT 115.005 206.025 115.815 209.385 ;
        RECT 116.025 209.245 116.705 209.385 ;
        RECT 116.025 209.095 116.835 209.235 ;
        RECT 115.835 208.925 116.835 209.095 ;
        RECT 115.005 205.875 115.815 206.015 ;
        RECT 115.005 205.705 116.005 205.875 ;
        RECT 115.005 204.645 115.815 205.705 ;
        RECT 116.025 205.565 116.835 208.925 ;
        RECT 115.865 205.300 115.975 205.420 ;
        RECT 116.110 204.655 116.895 205.085 ;
        RECT 114.905 203.245 115.815 204.595 ;
        RECT 116.025 204.495 116.705 204.635 ;
        RECT 115.835 204.325 116.705 204.495 ;
        RECT 115.135 201.710 115.815 203.245 ;
        RECT 114.915 200.800 115.815 201.710 ;
        RECT 115.135 197.595 115.815 200.800 ;
        RECT 115.135 197.425 116.005 197.595 ;
        RECT 115.135 197.285 115.815 197.425 ;
        RECT 114.905 196.860 115.815 197.275 ;
        RECT 114.905 196.690 116.005 196.860 ;
        RECT 114.905 196.345 115.815 196.690 ;
        RECT 115.135 193.375 115.815 196.345 ;
        RECT 116.025 195.530 116.705 204.325 ;
        RECT 116.025 195.295 116.835 195.435 ;
        RECT 115.835 195.125 116.835 195.295 ;
        RECT 116.025 194.065 116.835 195.125 ;
        RECT 116.025 193.915 116.805 194.055 ;
        RECT 115.835 193.745 116.805 193.915 ;
        RECT 115.860 192.825 115.970 192.985 ;
        RECT 116.025 192.685 116.805 193.745 ;
        RECT 116.025 192.535 116.805 192.675 ;
        RECT 115.835 192.365 116.805 192.535 ;
        RECT 114.945 191.775 115.730 192.205 ;
        RECT 114.905 190.740 115.815 191.660 ;
        RECT 116.025 191.305 116.805 192.365 ;
        RECT 116.025 191.155 116.805 191.295 ;
        RECT 115.835 190.985 116.805 191.155 ;
        RECT 115.135 188.395 115.815 190.740 ;
        RECT 116.025 189.925 116.805 190.985 ;
        RECT 116.025 189.775 116.805 189.915 ;
        RECT 115.835 189.605 116.805 189.775 ;
        RECT 116.025 188.545 116.805 189.605 ;
        RECT 115.135 188.225 116.005 188.395 ;
        RECT 115.135 188.195 115.815 188.225 ;
        RECT 115.860 187.765 115.970 187.925 ;
        RECT 116.025 187.480 116.935 188.515 ;
        RECT 115.835 187.310 116.935 187.480 ;
        RECT 116.025 187.165 116.935 187.310 ;
        RECT 114.905 184.715 115.815 187.155 ;
        RECT 116.025 187.015 116.935 187.075 ;
        RECT 115.835 186.845 116.935 187.015 ;
        RECT 114.905 184.545 116.005 184.715 ;
        RECT 114.905 184.405 115.815 184.545 ;
        RECT 115.860 184.085 115.970 184.245 ;
        RECT 116.025 183.625 116.935 186.845 ;
        RECT 115.005 182.415 115.815 183.475 ;
        RECT 116.025 182.415 116.835 183.475 ;
        RECT 115.005 182.245 116.835 182.415 ;
        RECT 115.005 182.105 115.815 182.245 ;
        RECT 116.025 182.105 116.835 182.245 ;
      LAYER nwell ;
        RECT 117.225 181.910 120.055 218.170 ;
      LAYER pwell ;
        RECT 120.445 217.835 121.255 217.975 ;
        RECT 121.465 217.835 122.275 217.975 ;
        RECT 120.445 217.665 122.275 217.835 ;
        RECT 120.445 216.605 121.255 217.665 ;
        RECT 121.465 216.605 122.275 217.665 ;
        RECT 120.345 215.250 121.255 216.595 ;
        RECT 121.465 216.455 122.145 216.595 ;
        RECT 121.275 216.285 122.145 216.455 ;
        RECT 120.575 215.075 121.255 215.250 ;
        RECT 120.575 214.905 121.445 215.075 ;
        RECT 120.575 214.765 121.255 214.905 ;
        RECT 121.300 214.445 121.410 214.605 ;
        RECT 120.575 213.695 121.255 213.725 ;
        RECT 120.575 213.525 121.445 213.695 ;
        RECT 120.575 211.180 121.255 213.525 ;
        RECT 120.345 210.260 121.255 211.180 ;
        RECT 121.465 213.080 122.145 216.285 ;
        RECT 121.465 212.170 122.365 213.080 ;
        RECT 121.465 210.635 122.145 212.170 ;
        RECT 121.300 209.845 121.410 210.005 ;
        RECT 121.465 209.285 122.375 210.635 ;
        RECT 120.575 209.095 121.255 209.125 ;
        RECT 121.465 209.095 122.275 209.235 ;
        RECT 120.575 208.925 122.275 209.095 ;
        RECT 120.575 206.580 121.255 208.925 ;
        RECT 120.345 205.660 121.255 206.580 ;
        RECT 121.465 205.565 122.275 208.925 ;
        RECT 120.575 202.355 121.255 205.325 ;
        RECT 121.305 205.300 121.415 205.420 ;
        RECT 121.550 204.655 122.335 205.085 ;
        RECT 121.465 204.495 122.145 204.635 ;
        RECT 121.275 204.325 122.145 204.495 ;
        RECT 120.345 202.010 121.255 202.355 ;
        RECT 120.345 201.840 121.445 202.010 ;
        RECT 120.345 201.425 121.255 201.840 ;
        RECT 120.445 201.275 121.255 201.415 ;
        RECT 120.445 201.105 121.445 201.275 ;
        RECT 121.465 201.120 122.145 204.325 ;
        RECT 120.445 199.585 121.255 201.105 ;
        RECT 121.465 200.210 122.365 201.120 ;
        RECT 120.575 199.435 121.255 199.575 ;
        RECT 120.575 199.265 121.445 199.435 ;
        RECT 120.575 196.060 121.255 199.265 ;
        RECT 121.465 198.675 122.145 200.210 ;
        RECT 121.465 197.325 122.375 198.675 ;
        RECT 121.465 197.130 122.145 197.275 ;
        RECT 121.275 196.960 122.145 197.130 ;
        RECT 120.355 195.150 121.255 196.060 ;
        RECT 120.575 193.615 121.255 195.150 ;
        RECT 121.465 195.430 122.145 196.960 ;
        RECT 121.465 194.065 122.375 195.430 ;
        RECT 121.465 193.915 122.275 194.055 ;
        RECT 121.275 193.745 122.275 193.915 ;
        RECT 120.345 192.265 121.255 193.615 ;
        RECT 120.385 191.775 121.170 192.205 ;
        RECT 120.345 191.340 121.255 191.755 ;
        RECT 120.345 191.170 121.445 191.340 ;
        RECT 121.465 191.305 122.275 193.745 ;
        RECT 120.345 190.825 121.255 191.170 ;
        RECT 121.305 191.040 121.415 191.160 ;
        RECT 120.575 187.855 121.255 190.825 ;
        RECT 121.465 190.695 122.145 190.725 ;
        RECT 121.275 190.525 122.145 190.695 ;
        RECT 121.465 188.180 122.145 190.525 ;
        RECT 120.475 187.475 121.255 187.615 ;
        RECT 120.475 187.305 121.445 187.475 ;
        RECT 120.475 186.245 121.255 187.305 ;
        RECT 121.465 187.260 122.375 188.180 ;
        RECT 121.465 187.015 122.375 187.075 ;
        RECT 121.275 186.845 122.375 187.015 ;
        RECT 120.345 185.290 121.255 186.235 ;
        RECT 120.545 183.800 121.225 185.290 ;
        RECT 121.465 184.075 122.375 186.845 ;
        RECT 120.545 183.630 121.445 183.800 ;
        RECT 120.545 183.485 121.225 183.630 ;
        RECT 120.445 182.415 121.255 183.475 ;
        RECT 121.465 182.415 122.275 183.475 ;
        RECT 120.445 182.245 122.275 182.415 ;
        RECT 120.445 182.105 121.255 182.245 ;
        RECT 121.465 182.105 122.275 182.245 ;
      LAYER nwell ;
        RECT 122.665 181.910 125.495 218.170 ;
      LAYER pwell ;
        RECT 125.885 217.835 126.695 217.975 ;
        RECT 126.905 217.835 127.715 217.975 ;
        RECT 125.885 217.665 127.715 217.835 ;
        RECT 125.885 216.605 126.695 217.665 ;
        RECT 126.905 216.605 127.715 217.665 ;
        RECT 125.785 215.250 126.695 216.595 ;
        RECT 126.905 216.455 127.715 216.595 ;
        RECT 126.715 216.285 127.715 216.455 ;
        RECT 126.015 215.075 126.695 215.250 ;
        RECT 126.905 215.225 127.715 216.285 ;
        RECT 126.905 215.075 127.585 215.105 ;
        RECT 126.015 214.905 127.585 215.075 ;
        RECT 126.015 214.765 126.695 214.905 ;
        RECT 126.745 214.500 126.855 214.620 ;
        RECT 125.785 213.880 126.695 214.295 ;
        RECT 125.785 213.710 126.885 213.880 ;
        RECT 125.785 213.365 126.695 213.710 ;
        RECT 126.015 210.395 126.695 213.365 ;
        RECT 126.905 212.560 127.585 214.905 ;
        RECT 126.905 211.640 127.815 212.560 ;
        RECT 126.905 210.520 127.815 211.440 ;
        RECT 126.015 210.015 126.695 210.155 ;
        RECT 126.015 209.845 126.885 210.015 ;
        RECT 126.015 206.640 126.695 209.845 ;
        RECT 126.905 208.175 127.585 210.520 ;
        RECT 126.715 208.005 127.585 208.175 ;
        RECT 126.905 207.975 127.585 208.005 ;
        RECT 126.905 207.715 127.715 207.855 ;
        RECT 126.715 207.545 127.715 207.715 ;
        RECT 125.795 205.730 126.695 206.640 ;
        RECT 126.015 204.195 126.695 205.730 ;
        RECT 126.905 205.105 127.715 207.545 ;
        RECT 126.990 204.655 127.775 205.085 ;
        RECT 125.785 202.845 126.695 204.195 ;
        RECT 126.905 203.580 127.815 204.615 ;
        RECT 126.715 203.410 127.815 203.580 ;
        RECT 126.905 203.265 127.815 203.410 ;
        RECT 125.785 202.380 126.695 202.795 ;
        RECT 125.785 202.210 126.885 202.380 ;
        RECT 125.785 201.865 126.695 202.210 ;
        RECT 126.015 198.895 126.695 201.865 ;
        RECT 126.905 199.435 127.815 203.185 ;
        RECT 126.715 199.265 127.815 199.435 ;
        RECT 126.905 199.125 127.815 199.265 ;
        RECT 125.785 197.640 126.695 198.560 ;
        RECT 126.015 195.295 126.695 197.640 ;
        RECT 126.905 198.100 127.815 199.020 ;
        RECT 126.905 195.755 127.585 198.100 ;
        RECT 126.715 195.585 127.585 195.755 ;
        RECT 126.905 195.555 127.585 195.585 ;
        RECT 126.905 195.295 127.715 195.435 ;
        RECT 126.015 195.125 127.715 195.295 ;
        RECT 126.015 195.095 126.695 195.125 ;
        RECT 125.885 194.835 126.695 194.975 ;
        RECT 125.885 194.665 126.885 194.835 ;
        RECT 125.885 192.225 126.695 194.665 ;
        RECT 126.905 194.065 127.715 195.125 ;
        RECT 126.905 193.105 127.815 194.055 ;
        RECT 125.825 191.775 126.610 192.205 ;
        RECT 125.785 188.860 126.695 191.465 ;
        RECT 126.935 190.700 127.615 193.105 ;
        RECT 126.715 190.530 127.615 190.700 ;
        RECT 126.935 190.385 127.615 190.530 ;
        RECT 126.905 190.230 127.815 190.375 ;
        RECT 126.715 190.060 127.815 190.230 ;
        RECT 126.905 189.025 127.815 190.060 ;
        RECT 125.785 188.845 126.885 188.860 ;
        RECT 126.905 188.845 127.685 188.995 ;
        RECT 125.785 188.690 127.685 188.845 ;
        RECT 125.785 188.545 126.695 188.690 ;
        RECT 126.715 188.675 127.685 188.690 ;
        RECT 126.740 188.225 126.850 188.385 ;
        RECT 126.905 187.625 127.685 188.675 ;
        RECT 125.785 184.255 126.695 187.475 ;
        RECT 126.905 184.255 127.815 187.475 ;
        RECT 125.785 184.085 127.815 184.255 ;
        RECT 125.785 184.025 126.695 184.085 ;
        RECT 126.905 184.025 127.815 184.085 ;
        RECT 126.745 183.680 126.855 183.800 ;
        RECT 125.885 182.415 126.695 183.475 ;
        RECT 126.905 182.415 127.715 183.475 ;
        RECT 125.885 182.245 127.715 182.415 ;
        RECT 125.885 182.105 126.695 182.245 ;
        RECT 126.905 182.105 127.715 182.245 ;
      LAYER nwell ;
        RECT 128.105 181.910 130.935 218.170 ;
      LAYER pwell ;
        RECT 131.325 217.835 132.135 217.975 ;
        RECT 132.345 217.835 133.155 217.975 ;
        RECT 131.325 217.665 133.155 217.835 ;
        RECT 131.325 216.605 132.135 217.665 ;
        RECT 132.345 216.605 133.155 217.665 ;
        RECT 131.225 215.205 132.135 216.555 ;
        RECT 132.345 216.180 133.255 216.595 ;
        RECT 132.155 216.010 133.255 216.180 ;
        RECT 131.455 213.670 132.135 215.205 ;
        RECT 131.235 212.760 132.135 213.670 ;
        RECT 131.455 209.555 132.135 212.760 ;
        RECT 132.345 215.665 133.255 216.010 ;
        RECT 132.345 212.695 133.025 215.665 ;
        RECT 132.345 212.315 133.025 212.455 ;
        RECT 132.155 212.145 133.025 212.315 ;
        RECT 131.455 209.385 132.325 209.555 ;
        RECT 131.455 209.245 132.135 209.385 ;
        RECT 131.325 209.095 132.135 209.235 ;
        RECT 131.325 208.925 132.325 209.095 ;
        RECT 132.345 208.940 133.025 212.145 ;
        RECT 131.325 206.485 132.135 208.925 ;
        RECT 132.345 208.030 133.245 208.940 ;
        RECT 132.345 206.495 133.025 208.030 ;
        RECT 132.185 206.220 132.295 206.340 ;
        RECT 131.455 205.875 132.135 206.015 ;
        RECT 131.455 205.705 132.325 205.875 ;
        RECT 131.455 196.910 132.135 205.705 ;
        RECT 132.345 205.145 133.255 206.495 ;
        RECT 132.430 204.655 133.215 205.085 ;
        RECT 132.345 204.495 133.025 204.635 ;
        RECT 132.155 204.325 133.025 204.495 ;
        RECT 132.345 201.120 133.025 204.325 ;
        RECT 132.345 200.210 133.245 201.120 ;
        RECT 132.345 198.675 133.025 200.210 ;
        RECT 132.345 197.325 133.255 198.675 ;
        RECT 132.185 197.020 132.295 197.140 ;
        RECT 131.225 195.800 132.135 196.720 ;
        RECT 131.455 193.455 132.135 195.800 ;
        RECT 132.345 195.450 133.255 196.815 ;
        RECT 132.345 193.920 133.025 195.450 ;
        RECT 132.155 193.750 133.025 193.920 ;
        RECT 132.345 193.605 133.025 193.750 ;
        RECT 131.455 193.285 132.325 193.455 ;
        RECT 131.455 193.255 132.135 193.285 ;
        RECT 132.180 192.825 132.290 192.985 ;
        RECT 132.345 192.535 133.255 192.595 ;
        RECT 132.155 192.365 133.255 192.535 ;
        RECT 131.265 191.775 132.050 192.205 ;
        RECT 131.425 191.620 132.105 191.745 ;
        RECT 131.425 191.450 132.325 191.620 ;
        RECT 131.425 190.420 132.105 191.450 ;
        RECT 131.225 189.465 132.135 190.420 ;
        RECT 132.345 189.595 133.255 192.365 ;
        RECT 131.325 189.315 132.135 189.455 ;
        RECT 131.325 189.310 132.325 189.315 ;
        RECT 132.345 189.310 133.255 189.455 ;
        RECT 131.325 189.145 133.255 189.310 ;
        RECT 131.325 186.705 132.135 189.145 ;
        RECT 132.155 189.140 133.255 189.145 ;
        RECT 132.345 188.105 133.255 189.140 ;
        RECT 132.185 187.820 132.295 187.940 ;
        RECT 132.345 187.475 133.255 187.535 ;
        RECT 132.155 187.305 133.255 187.475 ;
        RECT 132.185 186.440 132.295 186.560 ;
        RECT 131.225 185.180 132.135 186.215 ;
        RECT 131.225 185.010 132.325 185.180 ;
        RECT 131.225 184.865 132.135 185.010 ;
        RECT 131.355 183.795 132.135 184.855 ;
        RECT 132.345 184.085 133.255 187.305 ;
        RECT 132.185 183.795 132.295 183.800 ;
        RECT 131.355 183.625 132.325 183.795 ;
        RECT 131.355 183.485 132.135 183.625 ;
        RECT 131.325 182.415 132.135 183.475 ;
        RECT 132.345 182.415 133.155 183.475 ;
        RECT 131.325 182.245 133.155 182.415 ;
        RECT 131.325 182.105 132.135 182.245 ;
        RECT 132.345 182.105 133.155 182.245 ;
      LAYER nwell ;
        RECT 133.545 181.910 136.375 218.170 ;
      LAYER pwell ;
        RECT 136.765 217.835 137.575 217.975 ;
        RECT 137.785 217.835 138.595 217.975 ;
        RECT 136.765 217.665 138.595 217.835 ;
        RECT 136.765 216.605 137.575 217.665 ;
        RECT 137.785 216.605 138.595 217.665 ;
        RECT 136.665 215.250 137.575 216.595 ;
        RECT 137.785 216.455 138.465 216.595 ;
        RECT 137.595 216.285 138.465 216.455 ;
        RECT 136.895 215.075 137.575 215.250 ;
        RECT 136.895 214.905 137.765 215.075 ;
        RECT 136.895 214.765 137.575 214.905 ;
        RECT 136.665 214.340 137.575 214.755 ;
        RECT 136.665 214.170 137.765 214.340 ;
        RECT 136.665 213.825 137.575 214.170 ;
        RECT 136.895 210.855 137.575 213.825 ;
        RECT 137.785 213.080 138.465 216.285 ;
        RECT 137.785 212.170 138.685 213.080 ;
        RECT 137.785 210.635 138.465 212.170 ;
        RECT 136.765 210.475 137.575 210.615 ;
        RECT 136.765 210.305 137.765 210.475 ;
        RECT 136.765 209.245 137.575 210.305 ;
        RECT 137.785 209.285 138.695 210.635 ;
        RECT 136.895 200.355 137.575 209.150 ;
        RECT 137.785 208.220 138.695 209.140 ;
        RECT 137.785 205.875 138.465 208.220 ;
        RECT 137.595 205.705 138.465 205.875 ;
        RECT 137.785 205.675 138.465 205.705 ;
        RECT 137.625 205.300 137.735 205.420 ;
        RECT 137.870 204.655 138.655 205.085 ;
        RECT 137.785 204.220 138.695 204.635 ;
        RECT 137.595 204.050 138.695 204.220 ;
        RECT 137.785 203.705 138.695 204.050 ;
        RECT 137.785 200.735 138.465 203.705 ;
        RECT 137.625 200.355 137.735 200.360 ;
        RECT 136.895 200.185 137.765 200.355 ;
        RECT 136.895 200.045 137.575 200.185 ;
        RECT 136.665 199.020 137.575 199.940 ;
        RECT 137.595 199.890 137.765 199.895 ;
        RECT 137.595 199.725 138.465 199.890 ;
        RECT 136.895 196.675 137.575 199.020 ;
        RECT 137.785 198.985 138.465 199.725 ;
        RECT 137.785 198.055 138.695 198.985 ;
        RECT 137.785 196.675 138.695 197.725 ;
        RECT 136.895 196.505 138.695 196.675 ;
        RECT 136.895 196.475 137.575 196.505 ;
        RECT 137.785 196.375 138.695 196.505 ;
        RECT 136.765 196.215 137.575 196.355 ;
        RECT 137.785 196.215 138.465 196.355 ;
        RECT 136.765 196.045 138.465 196.215 ;
        RECT 136.765 194.985 137.575 196.045 ;
        RECT 136.865 194.830 137.545 194.975 ;
        RECT 136.865 194.660 137.765 194.830 ;
        RECT 136.865 193.170 137.545 194.660 ;
        RECT 136.665 192.225 137.575 193.170 ;
        RECT 137.785 192.840 138.465 196.045 ;
        RECT 136.705 191.775 137.490 192.205 ;
        RECT 137.785 191.930 138.685 192.840 ;
        RECT 136.665 191.615 137.575 191.675 ;
        RECT 136.665 191.445 137.765 191.615 ;
        RECT 136.665 188.225 137.575 191.445 ;
        RECT 137.785 190.395 138.465 191.930 ;
        RECT 137.785 189.045 138.695 190.395 ;
        RECT 137.625 188.740 137.735 188.860 ;
        RECT 137.595 188.390 137.765 188.395 ;
        RECT 137.595 188.225 138.465 188.390 ;
        RECT 136.665 187.935 137.575 187.995 ;
        RECT 136.665 187.765 137.765 187.935 ;
        RECT 136.665 184.545 137.575 187.765 ;
        RECT 137.785 187.485 138.465 188.225 ;
        RECT 137.785 186.555 138.695 187.485 ;
        RECT 137.785 186.095 138.565 186.235 ;
        RECT 137.595 185.925 138.565 186.095 ;
        RECT 137.785 184.865 138.565 185.925 ;
        RECT 137.620 184.085 137.730 184.245 ;
        RECT 137.785 183.805 138.565 184.855 ;
        RECT 137.595 183.635 138.565 183.805 ;
        RECT 137.785 183.485 138.565 183.635 ;
        RECT 136.765 182.415 137.575 183.475 ;
        RECT 137.785 182.415 138.595 183.475 ;
        RECT 136.765 182.245 138.595 182.415 ;
        RECT 136.765 182.105 137.575 182.245 ;
        RECT 137.785 182.105 138.595 182.245 ;
      LAYER nwell ;
        RECT 138.985 181.910 141.815 218.170 ;
      LAYER pwell ;
        RECT 142.205 217.835 143.015 217.975 ;
        RECT 143.225 217.835 144.035 217.975 ;
        RECT 142.205 217.665 144.035 217.835 ;
        RECT 142.205 216.605 143.015 217.665 ;
        RECT 143.225 216.605 144.035 217.665 ;
        RECT 142.205 216.455 143.015 216.595 ;
        RECT 143.225 216.455 144.035 216.595 ;
        RECT 142.205 216.285 144.035 216.455 ;
        RECT 142.205 212.925 143.015 216.285 ;
        RECT 143.065 212.660 143.175 212.780 ;
        RECT 142.105 211.065 143.015 212.415 ;
        RECT 143.225 211.085 144.035 216.285 ;
        RECT 142.335 209.530 143.015 211.065 ;
        RECT 143.070 210.765 143.180 210.925 ;
        RECT 143.225 210.015 143.905 210.155 ;
        RECT 143.035 209.845 143.905 210.015 ;
        RECT 142.115 208.620 143.015 209.530 ;
        RECT 142.335 205.415 143.015 208.620 ;
        RECT 143.225 209.670 143.905 209.845 ;
        RECT 143.225 208.325 144.135 209.670 ;
        RECT 143.225 205.415 144.135 208.185 ;
        RECT 142.335 205.245 144.135 205.415 ;
        RECT 142.335 205.105 143.015 205.245 ;
        RECT 143.225 205.185 144.135 205.245 ;
        RECT 142.335 204.955 143.015 205.095 ;
        RECT 142.335 204.785 143.205 204.955 ;
        RECT 142.335 201.580 143.015 204.785 ;
        RECT 143.310 204.655 144.095 205.085 ;
        RECT 143.070 204.325 143.180 204.485 ;
        RECT 143.225 203.575 143.905 203.605 ;
        RECT 143.035 203.405 143.905 203.575 ;
        RECT 142.115 200.670 143.015 201.580 ;
        RECT 142.335 199.135 143.015 200.670 ;
        RECT 143.225 201.060 143.905 203.405 ;
        RECT 143.225 200.140 144.135 201.060 ;
        RECT 143.070 199.725 143.180 199.885 ;
        RECT 142.105 197.785 143.015 199.135 ;
        RECT 143.225 197.770 144.135 199.115 ;
        RECT 143.225 197.595 143.905 197.770 ;
        RECT 143.035 197.425 143.905 197.595 ;
        RECT 142.105 196.495 143.015 197.425 ;
        RECT 143.225 197.285 143.905 197.425 ;
        RECT 143.225 197.135 143.905 197.165 ;
        RECT 143.035 196.965 143.905 197.135 ;
        RECT 142.335 195.755 143.015 196.495 ;
        RECT 142.335 195.590 143.205 195.755 ;
        RECT 143.035 195.585 143.205 195.590 ;
        RECT 142.335 195.295 143.015 195.435 ;
        RECT 142.335 195.125 143.205 195.295 ;
        RECT 142.335 194.950 143.015 195.125 ;
        RECT 142.105 193.605 143.015 194.950 ;
        RECT 143.225 194.620 143.905 196.965 ;
        RECT 143.225 193.700 144.135 194.620 ;
        RECT 142.105 193.455 143.015 193.585 ;
        RECT 142.105 193.445 143.205 193.455 ;
        RECT 143.225 193.445 144.005 193.595 ;
        RECT 142.105 193.285 144.005 193.445 ;
        RECT 142.105 192.235 143.015 193.285 ;
        RECT 143.035 193.275 144.005 193.285 ;
        RECT 143.225 192.225 144.005 193.275 ;
        RECT 142.145 191.775 142.930 192.205 ;
        RECT 143.310 191.775 144.095 192.205 ;
        RECT 142.105 191.615 143.015 191.675 ;
        RECT 142.105 191.445 143.205 191.615 ;
        RECT 142.105 188.675 143.015 191.445 ;
        RECT 143.225 189.490 144.135 190.835 ;
        RECT 143.225 189.315 143.905 189.490 ;
        RECT 143.035 189.145 143.905 189.315 ;
        RECT 143.225 189.005 143.905 189.145 ;
        RECT 143.225 188.855 144.035 188.995 ;
        RECT 143.035 188.685 144.035 188.855 ;
        RECT 142.335 188.395 143.015 188.425 ;
        RECT 142.335 188.225 143.205 188.395 ;
        RECT 142.335 185.880 143.015 188.225 ;
        RECT 143.225 187.625 144.035 188.685 ;
        RECT 143.225 186.555 144.005 187.615 ;
        RECT 143.035 186.385 144.005 186.555 ;
        RECT 143.225 186.245 144.005 186.385 ;
        RECT 142.105 184.960 143.015 185.880 ;
        RECT 143.225 185.175 144.005 186.235 ;
        RECT 143.035 185.005 144.005 185.175 ;
        RECT 143.225 184.865 144.005 185.005 ;
        RECT 142.235 183.805 143.015 184.855 ;
        RECT 143.225 183.805 144.005 184.855 ;
        RECT 142.235 183.635 144.005 183.805 ;
        RECT 142.235 183.485 143.015 183.635 ;
        RECT 143.225 183.485 144.005 183.635 ;
        RECT 142.205 182.415 143.015 183.475 ;
        RECT 143.225 182.415 144.035 183.475 ;
        RECT 142.205 182.245 144.035 182.415 ;
        RECT 142.205 182.105 143.015 182.245 ;
        RECT 143.225 182.105 144.035 182.245 ;
      LAYER nwell ;
        RECT 144.425 181.910 146.030 218.170 ;
      LAYER pwell ;
        RECT 100.770 163.670 106.870 173.460 ;
        RECT 100.770 163.640 106.880 163.670 ;
        RECT 100.970 163.240 102.130 163.640 ;
        RECT 104.090 161.560 106.880 163.640 ;
      LAYER nwell ;
        RECT 101.980 159.450 106.820 161.560 ;
        RECT 108.100 161.220 118.290 173.470 ;
      LAYER pwell ;
        RECT 119.810 163.700 125.910 173.490 ;
        RECT 119.810 163.670 125.920 163.700 ;
        RECT 120.010 163.270 121.170 163.670 ;
        RECT 123.130 161.590 125.920 163.670 ;
      LAYER nwell ;
        RECT 121.020 159.480 125.860 161.590 ;
        RECT 127.140 161.250 137.330 173.500 ;
      LAYER pwell ;
        RECT 138.760 163.740 144.860 173.530 ;
        RECT 138.760 163.710 144.870 163.740 ;
        RECT 138.960 163.310 140.120 163.710 ;
        RECT 142.080 161.630 144.870 163.710 ;
      LAYER nwell ;
        RECT 139.970 159.520 144.810 161.630 ;
        RECT 146.090 161.290 156.280 173.540 ;
      LAYER pwell ;
        RECT 100.770 148.680 106.870 158.470 ;
        RECT 100.770 148.650 106.880 148.680 ;
        RECT 100.970 148.250 102.130 148.650 ;
        RECT 104.090 146.570 106.880 148.650 ;
      LAYER nwell ;
        RECT 101.980 144.460 106.820 146.570 ;
        RECT 108.100 146.230 118.290 158.480 ;
      LAYER pwell ;
        RECT 119.810 148.680 125.910 158.470 ;
        RECT 119.810 148.650 125.920 148.680 ;
        RECT 120.010 148.250 121.170 148.650 ;
        RECT 123.130 146.570 125.920 148.650 ;
      LAYER nwell ;
        RECT 121.020 144.460 125.860 146.570 ;
        RECT 127.140 146.230 137.330 158.480 ;
      LAYER pwell ;
        RECT 138.810 148.680 144.910 158.470 ;
        RECT 138.810 148.650 144.920 148.680 ;
        RECT 139.010 148.250 140.170 148.650 ;
        RECT 142.130 146.570 144.920 148.650 ;
      LAYER nwell ;
        RECT 140.020 144.460 144.860 146.570 ;
        RECT 146.140 146.230 156.330 158.480 ;
      LAYER pwell ;
        RECT 100.770 133.700 106.870 143.490 ;
        RECT 100.770 133.670 106.880 133.700 ;
        RECT 100.970 133.270 102.130 133.670 ;
        RECT 104.090 131.590 106.880 133.670 ;
      LAYER nwell ;
        RECT 101.980 129.480 106.820 131.590 ;
        RECT 108.100 131.250 118.290 143.500 ;
      LAYER pwell ;
        RECT 119.760 133.660 125.860 143.450 ;
        RECT 119.760 133.630 125.870 133.660 ;
        RECT 119.960 133.230 121.120 133.630 ;
        RECT 123.080 131.550 125.870 133.630 ;
      LAYER nwell ;
        RECT 120.970 129.440 125.810 131.550 ;
        RECT 127.090 131.210 137.280 143.460 ;
      LAYER pwell ;
        RECT 138.760 133.660 144.860 143.450 ;
        RECT 138.760 133.630 144.870 133.660 ;
        RECT 138.960 133.230 140.120 133.630 ;
        RECT 142.080 131.550 144.870 133.630 ;
      LAYER nwell ;
        RECT 139.970 129.440 144.810 131.550 ;
        RECT 146.090 131.210 156.280 143.460 ;
      LAYER pwell ;
        RECT 100.770 118.670 106.870 128.460 ;
        RECT 100.770 118.640 106.880 118.670 ;
        RECT 100.970 118.240 102.130 118.640 ;
        RECT 104.090 116.560 106.880 118.640 ;
      LAYER nwell ;
        RECT 101.980 114.450 106.820 116.560 ;
        RECT 108.100 116.220 118.290 128.470 ;
      LAYER pwell ;
        RECT 119.760 118.640 125.860 128.430 ;
        RECT 119.760 118.610 125.870 118.640 ;
        RECT 119.960 118.210 121.120 118.610 ;
        RECT 123.080 116.530 125.870 118.610 ;
      LAYER nwell ;
        RECT 120.970 114.420 125.810 116.530 ;
        RECT 127.090 116.190 137.280 128.440 ;
      LAYER pwell ;
        RECT 138.760 118.640 144.860 128.430 ;
        RECT 138.760 118.610 144.870 118.640 ;
        RECT 138.960 118.210 140.120 118.610 ;
        RECT 142.080 116.530 144.870 118.610 ;
      LAYER nwell ;
        RECT 139.970 114.420 144.810 116.530 ;
        RECT 146.090 116.190 156.280 128.440 ;
      LAYER pwell ;
        RECT 100.770 103.680 106.870 113.470 ;
        RECT 100.770 103.650 106.880 103.680 ;
        RECT 100.970 103.250 102.130 103.650 ;
        RECT 104.090 101.570 106.880 103.650 ;
      LAYER nwell ;
        RECT 101.980 99.460 106.820 101.570 ;
        RECT 108.100 101.230 118.290 113.480 ;
      LAYER pwell ;
        RECT 119.760 103.660 125.860 113.450 ;
        RECT 119.760 103.630 125.870 103.660 ;
        RECT 119.960 103.230 121.120 103.630 ;
        RECT 123.080 101.550 125.870 103.630 ;
      LAYER nwell ;
        RECT 120.970 99.440 125.810 101.550 ;
        RECT 127.090 101.210 137.280 113.460 ;
      LAYER pwell ;
        RECT 138.810 103.660 144.910 113.450 ;
        RECT 138.810 103.630 144.920 103.660 ;
        RECT 139.010 103.230 140.170 103.630 ;
        RECT 142.130 101.550 144.920 103.630 ;
      LAYER nwell ;
        RECT 140.020 99.440 144.860 101.550 ;
        RECT 146.140 101.210 156.330 113.460 ;
      LAYER pwell ;
        RECT 102.490 96.920 156.930 98.930 ;
        RECT 102.490 95.440 144.950 96.920 ;
      LAYER li1 ;
        RECT 110.395 217.895 110.565 217.980 ;
        RECT 113.115 217.895 113.285 217.980 ;
        RECT 115.835 217.895 116.005 217.980 ;
        RECT 118.555 217.895 118.725 217.980 ;
        RECT 121.275 217.895 121.445 217.980 ;
        RECT 123.995 217.895 124.165 217.980 ;
        RECT 126.715 217.895 126.885 217.980 ;
        RECT 129.435 217.895 129.605 217.980 ;
        RECT 132.155 217.895 132.325 217.980 ;
        RECT 134.875 217.895 135.045 217.980 ;
        RECT 137.595 217.895 137.765 217.980 ;
        RECT 140.315 217.895 140.485 217.980 ;
        RECT 143.035 217.895 143.205 217.980 ;
        RECT 145.755 217.895 145.925 217.980 ;
        RECT 110.395 217.375 111.855 217.895 ;
        RECT 110.395 216.685 111.315 217.375 ;
        RECT 112.025 217.205 114.375 217.895 ;
        RECT 114.545 217.375 117.295 217.895 ;
        RECT 111.485 216.685 114.915 217.205 ;
        RECT 115.085 216.685 116.755 217.375 ;
        RECT 117.465 217.205 119.815 217.895 ;
        RECT 119.985 217.375 122.735 217.895 ;
        RECT 116.925 216.685 120.355 217.205 ;
        RECT 120.525 216.685 122.195 217.375 ;
        RECT 122.905 217.205 125.255 217.895 ;
        RECT 125.425 217.375 128.175 217.895 ;
        RECT 122.365 216.685 125.795 217.205 ;
        RECT 125.965 216.685 127.635 217.375 ;
        RECT 128.345 217.205 130.695 217.895 ;
        RECT 130.865 217.375 133.615 217.895 ;
        RECT 127.805 216.685 131.235 217.205 ;
        RECT 131.405 216.685 133.075 217.375 ;
        RECT 133.785 217.205 136.135 217.895 ;
        RECT 136.305 217.375 139.055 217.895 ;
        RECT 133.245 216.685 136.675 217.205 ;
        RECT 136.845 216.685 138.515 217.375 ;
        RECT 139.225 217.205 141.575 217.895 ;
        RECT 141.745 217.375 144.495 217.895 ;
        RECT 138.685 216.685 142.115 217.205 ;
        RECT 142.285 216.685 143.955 217.375 ;
        RECT 144.665 217.205 145.925 217.895 ;
        RECT 144.125 216.685 145.925 217.205 ;
        RECT 110.395 216.515 110.565 216.685 ;
        RECT 113.115 216.515 113.285 216.685 ;
        RECT 110.395 214.930 111.110 216.515 ;
        RECT 112.680 216.510 113.285 216.515 ;
        RECT 115.835 216.510 116.005 216.685 ;
        RECT 112.680 216.250 114.435 216.510 ;
        RECT 114.995 216.250 116.005 216.510 ;
        RECT 116.660 216.465 117.495 216.515 ;
        RECT 112.680 215.650 113.285 216.250 ;
        RECT 113.455 215.905 115.665 216.075 ;
        RECT 113.455 215.820 114.360 215.905 ;
        RECT 115.090 215.820 115.665 215.905 ;
        RECT 115.835 215.965 116.005 216.250 ;
        RECT 116.225 216.455 117.495 216.465 ;
        RECT 118.555 216.510 118.725 216.685 ;
        RECT 121.275 216.510 121.445 216.685 ;
        RECT 123.995 216.510 124.165 216.685 ;
        RECT 126.715 216.515 126.885 216.685 ;
        RECT 129.435 216.515 129.605 216.685 ;
        RECT 126.715 216.510 128.175 216.515 ;
        RECT 116.225 216.345 118.340 216.455 ;
        RECT 116.225 216.290 116.785 216.345 ;
        RECT 117.365 216.300 118.340 216.345 ;
        RECT 116.225 216.135 116.745 216.290 ;
        RECT 115.835 215.795 116.615 215.965 ;
        RECT 114.595 215.650 114.925 215.735 ;
        RECT 115.835 215.650 116.005 215.795 ;
        RECT 112.680 215.320 114.045 215.650 ;
        RECT 114.215 215.480 115.285 215.650 ;
        RECT 110.395 214.590 111.940 214.930 ;
        RECT 110.395 211.170 111.110 214.590 ;
        RECT 112.680 213.245 113.285 215.320 ;
        RECT 114.215 215.105 114.385 215.480 ;
        RECT 113.455 214.935 114.385 215.105 ;
        RECT 114.565 214.845 114.935 215.200 ;
        RECT 115.115 215.105 115.285 215.480 ;
        RECT 115.455 215.320 116.005 215.650 ;
        RECT 116.915 215.625 117.245 216.175 ;
        RECT 117.415 216.125 118.340 216.300 ;
        RECT 118.555 216.250 119.875 216.510 ;
        RECT 120.435 216.250 121.445 216.510 ;
        RECT 121.705 216.255 122.165 216.425 ;
        RECT 118.555 215.955 118.725 216.250 ;
        RECT 121.275 216.085 121.445 216.250 ;
        RECT 117.545 215.785 118.725 215.955 ;
        RECT 118.895 215.905 121.105 216.075 ;
        RECT 118.895 215.820 119.800 215.905 ;
        RECT 120.530 215.820 121.105 215.905 ;
        RECT 115.115 214.935 115.665 215.105 ;
        RECT 115.835 215.035 116.005 215.320 ;
        RECT 116.220 215.615 117.245 215.625 ;
        RECT 118.555 215.650 118.725 215.785 ;
        RECT 121.275 215.755 121.825 216.085 ;
        RECT 121.995 215.990 122.165 216.255 ;
        RECT 122.335 216.160 122.985 216.510 ;
        RECT 123.155 216.255 123.825 216.425 ;
        RECT 123.155 215.990 123.325 216.255 ;
        RECT 123.995 216.250 125.315 216.510 ;
        RECT 125.875 216.250 128.175 216.510 ;
        RECT 123.995 216.085 124.165 216.250 ;
        RECT 121.995 215.760 123.325 215.990 ;
        RECT 123.495 215.755 124.165 216.085 ;
        RECT 124.335 215.905 126.545 216.075 ;
        RECT 124.335 215.820 125.240 215.905 ;
        RECT 125.970 215.820 126.545 215.905 ;
        RECT 126.715 215.995 128.175 216.250 ;
        RECT 120.035 215.650 120.365 215.735 ;
        RECT 121.275 215.650 121.445 215.755 ;
        RECT 116.220 215.425 118.385 215.615 ;
        RECT 116.220 215.295 116.745 215.425 ;
        RECT 117.450 215.275 118.385 215.425 ;
        RECT 118.555 215.320 119.485 215.650 ;
        RECT 119.655 215.480 120.725 215.650 ;
        RECT 115.835 214.825 116.535 215.035 ;
        RECT 113.455 213.580 115.665 213.750 ;
        RECT 113.455 213.415 114.425 213.580 ;
        RECT 115.095 213.495 115.665 213.580 ;
        RECT 114.595 213.325 114.925 213.410 ;
        RECT 115.835 213.325 116.005 214.825 ;
        RECT 116.915 214.550 117.245 215.255 ;
        RECT 117.450 214.720 117.825 215.275 ;
        RECT 118.555 215.045 118.725 215.320 ;
        RECT 119.655 215.105 119.825 215.480 ;
        RECT 118.055 214.730 118.725 215.045 ;
        RECT 118.895 214.935 119.825 215.105 ;
        RECT 120.005 214.845 120.375 215.200 ;
        RECT 120.555 215.105 120.725 215.480 ;
        RECT 120.895 215.320 121.445 215.650 ;
        RECT 123.995 215.650 124.165 215.755 ;
        RECT 125.475 215.650 125.805 215.735 ;
        RECT 126.715 215.650 127.635 215.995 ;
        RECT 128.345 215.955 129.605 216.515 ;
        RECT 130.665 216.465 131.500 216.515 ;
        RECT 130.665 216.455 131.935 216.465 ;
        RECT 129.820 216.345 131.935 216.455 ;
        RECT 129.820 216.300 130.795 216.345 ;
        RECT 129.820 216.125 130.745 216.300 ;
        RECT 131.375 216.290 131.935 216.345 ;
        RECT 128.345 215.825 130.615 215.955 ;
        RECT 121.705 215.400 123.825 215.585 ;
        RECT 121.275 215.145 121.445 215.320 ;
        RECT 123.995 215.320 124.925 215.650 ;
        RECT 125.095 215.480 126.165 215.650 ;
        RECT 120.555 214.935 121.105 215.105 ;
        RECT 121.275 214.895 121.905 215.145 ;
        RECT 122.075 214.950 123.025 215.230 ;
        RECT 123.995 215.160 124.165 215.320 ;
        RECT 123.535 214.895 124.165 215.160 ;
        RECT 125.095 215.105 125.265 215.480 ;
        RECT 124.335 214.935 125.265 215.105 ;
        RECT 116.285 214.380 118.255 214.550 ;
        RECT 116.285 213.765 116.455 214.380 ;
        RECT 116.625 213.890 117.915 214.210 ;
        RECT 116.625 213.745 116.955 213.890 ;
        RECT 112.680 213.110 114.425 213.245 ;
        RECT 114.595 213.155 115.265 213.325 ;
        RECT 111.430 213.075 114.425 213.110 ;
        RECT 111.430 212.760 113.285 213.075 ;
        RECT 114.595 212.905 114.925 212.930 ;
        RECT 112.680 211.170 113.285 212.760 ;
        RECT 110.395 210.995 110.565 211.170 ;
        RECT 113.115 210.995 113.285 211.170 ;
        RECT 110.395 209.345 111.855 210.995 ;
        RECT 112.025 210.705 113.285 210.995 ;
        RECT 113.455 212.735 114.925 212.905 ;
        RECT 113.455 211.045 113.625 212.735 ;
        RECT 115.095 212.570 115.265 213.155 ;
        RECT 115.435 213.010 116.005 213.325 ;
        RECT 116.285 213.360 116.455 213.595 ;
        RECT 117.165 213.530 117.885 213.720 ;
        RECT 118.085 213.665 118.255 214.380 ;
        RECT 118.055 213.360 118.385 213.440 ;
        RECT 116.285 213.190 118.385 213.360 ;
        RECT 115.435 212.995 116.505 213.010 ;
        RECT 115.835 212.640 116.505 212.995 ;
        RECT 116.685 212.730 116.985 213.190 ;
        RECT 118.555 213.185 118.725 214.730 ;
        RECT 118.895 213.355 119.575 213.640 ;
        RECT 118.555 213.020 119.185 213.185 ;
        RECT 117.165 212.850 117.495 213.020 ;
        RECT 117.755 212.915 119.185 213.020 ;
        RECT 117.755 212.850 118.725 212.915 ;
        RECT 115.095 212.565 115.665 212.570 ;
        RECT 113.795 212.395 115.665 212.565 ;
        RECT 113.795 211.440 113.965 212.395 ;
        RECT 114.135 212.055 115.105 212.225 ;
        RECT 114.135 211.405 114.305 212.055 ;
        RECT 115.300 212.040 115.665 212.395 ;
        RECT 115.325 211.850 115.495 211.855 ;
        RECT 114.505 211.575 115.665 211.850 ;
        RECT 114.135 211.215 115.665 211.405 ;
        RECT 113.455 210.875 114.480 211.045 ;
        RECT 115.835 211.035 116.005 212.640 ;
        RECT 116.685 212.530 117.015 212.730 ;
        RECT 117.235 212.680 117.495 212.850 ;
        RECT 117.235 212.510 118.280 212.680 ;
        RECT 117.235 212.320 117.405 212.510 ;
        RECT 116.285 212.150 117.405 212.320 ;
        RECT 116.285 211.645 116.455 212.150 ;
        RECT 117.575 211.980 117.940 212.340 ;
        RECT 116.655 211.810 117.940 211.980 ;
        RECT 116.655 211.455 116.875 211.810 ;
        RECT 116.285 211.285 116.455 211.450 ;
        RECT 117.045 211.400 117.640 211.640 ;
        RECT 118.110 211.575 118.280 212.510 ;
        RECT 116.285 211.230 116.725 211.285 ;
        RECT 117.830 211.230 118.385 211.365 ;
        RECT 116.285 211.115 118.385 211.230 ;
        RECT 118.555 211.125 118.725 212.850 ;
        RECT 119.355 212.895 119.575 213.355 ;
        RECT 119.745 213.065 120.305 213.755 ;
        RECT 120.475 213.355 121.105 213.640 ;
        RECT 120.475 212.895 120.645 213.355 ;
        RECT 121.275 213.200 121.445 214.895 ;
        RECT 122.035 214.725 123.400 214.780 ;
        RECT 121.725 214.610 123.825 214.725 ;
        RECT 121.725 214.555 122.165 214.610 ;
        RECT 121.725 214.390 121.895 214.555 ;
        RECT 123.270 214.475 123.825 214.610 ;
        RECT 121.725 213.690 121.895 214.195 ;
        RECT 122.095 214.030 122.315 214.385 ;
        RECT 122.485 214.200 123.080 214.440 ;
        RECT 122.095 213.860 123.380 214.030 ;
        RECT 121.725 213.520 122.845 213.690 ;
        RECT 122.675 213.330 122.845 213.520 ;
        RECT 123.015 213.500 123.380 213.860 ;
        RECT 123.550 213.330 123.720 214.265 ;
        RECT 121.275 213.185 121.945 213.200 ;
        RECT 120.815 212.915 121.945 213.185 ;
        RECT 119.355 212.685 120.645 212.895 ;
        RECT 121.275 212.830 121.945 212.915 ;
        RECT 122.125 213.110 122.455 213.310 ;
        RECT 122.675 213.160 123.720 213.330 ;
        RECT 123.995 213.705 124.165 214.895 ;
        RECT 125.445 214.845 125.815 215.200 ;
        RECT 125.995 215.105 126.165 215.480 ;
        RECT 126.335 215.320 127.635 215.650 ;
        RECT 126.715 215.305 127.635 215.320 ;
        RECT 127.805 215.785 130.615 215.825 ;
        RECT 127.805 215.305 129.605 215.785 ;
        RECT 130.915 215.625 131.245 216.175 ;
        RECT 131.415 216.135 131.935 216.290 ;
        RECT 132.155 216.085 132.325 216.685 ;
        RECT 134.875 216.510 135.045 216.685 ;
        RECT 137.595 216.510 137.765 216.685 ;
        RECT 140.315 216.515 140.485 216.685 ;
        RECT 143.035 216.515 143.205 216.685 ;
        RECT 145.755 216.515 145.925 216.685 ;
        RECT 132.495 216.340 134.705 216.510 ;
        RECT 132.495 216.255 133.065 216.340 ;
        RECT 133.735 216.175 134.705 216.340 ;
        RECT 134.875 216.250 136.195 216.510 ;
        RECT 136.755 216.250 137.765 216.510 ;
        RECT 138.025 216.255 138.485 216.425 ;
        RECT 133.235 216.085 133.565 216.170 ;
        RECT 132.155 215.965 132.725 216.085 ;
        RECT 131.545 215.795 132.725 215.965 ;
        RECT 132.155 215.755 132.725 215.795 ;
        RECT 132.895 215.915 133.565 216.085 ;
        RECT 134.875 216.005 135.045 216.250 ;
        RECT 137.595 216.085 137.765 216.250 ;
        RECT 130.915 215.615 131.940 215.625 ;
        RECT 125.995 214.935 126.545 215.105 ;
        RECT 126.715 214.565 126.885 215.305 ;
        RECT 127.055 214.735 127.685 215.020 ;
        RECT 126.715 214.295 127.345 214.565 ;
        RECT 124.335 214.040 126.545 214.210 ;
        RECT 124.335 213.875 125.305 214.040 ;
        RECT 125.975 213.955 126.545 214.040 ;
        RECT 125.475 213.785 125.805 213.870 ;
        RECT 126.715 213.785 126.885 214.295 ;
        RECT 127.515 214.275 127.685 214.735 ;
        RECT 127.855 214.445 128.415 215.135 ;
        RECT 129.435 215.045 129.605 215.305 ;
        RECT 129.775 215.425 131.940 215.615 ;
        RECT 129.775 215.275 130.710 215.425 ;
        RECT 131.415 215.295 131.940 215.425 ;
        RECT 128.585 214.735 129.265 215.020 ;
        RECT 128.585 214.275 128.805 214.735 ;
        RECT 129.435 214.730 130.105 215.045 ;
        RECT 129.435 214.565 129.605 214.730 ;
        RECT 130.335 214.720 130.710 215.275 ;
        RECT 128.975 214.295 129.605 214.565 ;
        RECT 130.915 214.550 131.245 215.255 ;
        RECT 132.155 215.035 132.325 215.755 ;
        RECT 132.895 215.330 133.065 215.915 ;
        RECT 133.735 215.835 135.045 216.005 ;
        RECT 133.235 215.665 133.565 215.690 ;
        RECT 133.235 215.495 134.705 215.665 ;
        RECT 131.625 214.825 132.325 215.035 ;
        RECT 127.515 214.065 128.805 214.275 ;
        RECT 123.995 213.535 125.305 213.705 ;
        RECT 125.475 213.615 126.145 213.785 ;
        RECT 118.895 212.115 121.105 212.515 ;
        RECT 118.895 211.645 119.575 211.925 ;
        RECT 119.355 211.250 119.575 211.645 ;
        RECT 119.745 211.420 120.305 212.115 ;
        RECT 120.475 211.645 121.105 211.925 ;
        RECT 120.475 211.250 120.645 211.645 ;
        RECT 116.595 211.060 117.960 211.115 ;
        RECT 112.025 210.535 114.045 210.705 ;
        RECT 112.025 209.615 113.285 210.535 ;
        RECT 113.635 210.125 114.045 210.300 ;
        RECT 114.290 210.295 114.480 210.875 ;
        RECT 114.855 210.305 115.025 211.015 ;
        RECT 115.300 210.945 116.005 211.035 ;
        RECT 118.555 210.945 119.185 211.125 ;
        RECT 115.300 210.695 116.465 210.945 ;
        RECT 115.300 210.525 116.005 210.695 ;
        RECT 116.635 210.610 117.585 210.890 ;
        RECT 118.095 210.800 119.185 210.945 ;
        RECT 119.355 210.800 120.645 211.250 ;
        RECT 121.275 211.125 121.445 212.830 ;
        RECT 122.125 212.650 122.425 213.110 ;
        RECT 122.675 212.990 122.935 213.160 ;
        RECT 123.995 212.990 124.165 213.535 ;
        RECT 125.475 213.365 125.805 213.390 ;
        RECT 122.605 212.820 122.935 212.990 ;
        RECT 123.195 212.820 124.165 212.990 ;
        RECT 121.725 212.480 123.825 212.650 ;
        RECT 121.725 212.245 121.895 212.480 ;
        RECT 123.495 212.400 123.825 212.480 ;
        RECT 122.605 212.120 123.325 212.310 ;
        RECT 121.725 211.460 121.895 212.075 ;
        RECT 122.065 211.950 122.395 212.095 ;
        RECT 122.065 211.630 123.355 211.950 ;
        RECT 123.525 211.460 123.695 212.175 ;
        RECT 121.725 211.290 123.695 211.460 ;
        RECT 120.815 211.015 121.445 211.125 ;
        RECT 120.815 210.805 121.975 211.015 ;
        RECT 120.815 210.800 121.445 210.805 ;
        RECT 118.095 210.680 118.725 210.800 ;
        RECT 120.035 210.695 120.365 210.800 ;
        RECT 114.855 210.125 115.630 210.305 ;
        RECT 113.635 210.060 115.630 210.125 ;
        RECT 115.835 210.085 116.005 210.525 ;
        RECT 116.265 210.255 118.385 210.440 ;
        RECT 118.555 210.085 118.725 210.680 ;
        RECT 118.895 210.525 119.865 210.630 ;
        RECT 120.535 210.525 121.105 210.630 ;
        RECT 118.895 210.245 121.105 210.525 ;
        RECT 113.635 209.785 115.025 210.060 ;
        RECT 115.835 209.755 116.385 210.085 ;
        RECT 116.555 209.850 117.885 210.080 ;
        RECT 115.835 209.615 116.005 209.755 ;
        RECT 110.395 207.485 111.335 209.345 ;
        RECT 112.025 209.175 114.375 209.615 ;
        RECT 111.505 207.795 114.375 209.175 ;
        RECT 114.545 209.155 116.005 209.615 ;
        RECT 116.555 209.585 116.725 209.850 ;
        RECT 116.265 209.415 116.725 209.585 ;
        RECT 116.895 209.330 117.545 209.680 ;
        RECT 117.715 209.585 117.885 209.850 ;
        RECT 118.055 209.755 118.725 210.085 ;
        RECT 117.715 209.415 118.385 209.585 ;
        RECT 118.555 209.155 118.725 209.755 ;
        RECT 121.275 210.045 121.445 210.800 ;
        RECT 122.355 210.585 122.685 211.290 ;
        RECT 123.995 211.165 124.165 212.820 ;
        RECT 124.335 213.195 125.805 213.365 ;
        RECT 124.335 211.505 124.505 213.195 ;
        RECT 125.975 213.030 126.145 213.615 ;
        RECT 126.315 213.455 126.885 213.785 ;
        RECT 127.055 213.495 129.265 213.895 ;
        RECT 125.975 213.025 126.545 213.030 ;
        RECT 124.675 212.855 126.545 213.025 ;
        RECT 124.675 211.900 124.845 212.855 ;
        RECT 125.015 212.515 125.985 212.685 ;
        RECT 125.015 211.865 125.185 212.515 ;
        RECT 126.180 212.500 126.545 212.855 ;
        RECT 126.715 212.505 126.885 213.455 ;
        RECT 127.055 213.025 127.685 213.305 ;
        RECT 127.515 212.630 127.685 213.025 ;
        RECT 127.855 212.800 128.415 213.495 ;
        RECT 128.585 213.025 129.265 213.305 ;
        RECT 128.585 212.630 128.805 213.025 ;
        RECT 126.205 212.310 126.375 212.315 ;
        RECT 125.385 212.035 126.545 212.310 ;
        RECT 126.715 212.180 127.345 212.505 ;
        RECT 127.515 212.180 128.805 212.630 ;
        RECT 129.435 213.020 129.605 214.295 ;
        RECT 129.905 214.380 131.875 214.550 ;
        RECT 129.905 213.665 130.075 214.380 ;
        RECT 130.245 213.890 131.535 214.210 ;
        RECT 131.205 213.745 131.535 213.890 ;
        RECT 131.705 213.765 131.875 214.380 ;
        RECT 132.155 213.795 132.325 214.825 ;
        RECT 132.495 215.325 133.065 215.330 ;
        RECT 132.495 215.155 134.365 215.325 ;
        RECT 132.495 214.800 132.860 215.155 ;
        RECT 133.055 214.815 134.025 214.985 ;
        RECT 132.665 214.610 132.835 214.615 ;
        RECT 132.495 214.335 133.655 214.610 ;
        RECT 133.855 214.165 134.025 214.815 ;
        RECT 134.195 214.200 134.365 215.155 ;
        RECT 132.495 213.975 134.025 214.165 ;
        RECT 134.535 213.805 134.705 215.495 ;
        RECT 130.275 213.530 130.995 213.720 ;
        RECT 129.775 213.360 130.105 213.440 ;
        RECT 131.705 213.360 131.875 213.595 ;
        RECT 129.775 213.190 131.875 213.360 ;
        RECT 132.155 213.285 132.860 213.795 ;
        RECT 129.435 212.850 130.405 213.020 ;
        RECT 130.665 212.850 130.995 213.020 ;
        RECT 129.435 212.505 129.605 212.850 ;
        RECT 130.665 212.680 130.925 212.850 ;
        RECT 131.175 212.730 131.475 213.190 ;
        RECT 132.155 213.010 132.325 213.285 ;
        RECT 133.135 213.065 133.305 213.775 ;
        RECT 128.975 212.180 129.605 212.505 ;
        RECT 125.015 211.675 126.545 211.865 ;
        RECT 124.335 211.335 125.360 211.505 ;
        RECT 126.715 211.495 126.885 212.180 ;
        RECT 127.795 212.075 128.125 212.180 ;
        RECT 127.055 211.905 127.625 212.010 ;
        RECT 128.295 211.905 129.265 212.010 ;
        RECT 127.055 211.625 129.265 211.905 ;
        RECT 122.890 210.565 123.265 211.120 ;
        RECT 123.995 211.110 124.925 211.165 ;
        RECT 123.495 210.995 124.925 211.110 ;
        RECT 123.495 210.795 124.165 210.995 ;
        RECT 121.660 210.415 122.185 210.545 ;
        RECT 122.890 210.415 123.825 210.565 ;
        RECT 121.660 210.225 123.825 210.415 ;
        RECT 121.660 210.215 122.685 210.225 ;
        RECT 121.275 209.875 122.055 210.045 ;
        RECT 121.275 209.155 121.445 209.875 ;
        RECT 121.665 209.550 122.185 209.705 ;
        RECT 122.355 209.665 122.685 210.215 ;
        RECT 123.995 210.055 124.165 210.795 ;
        RECT 124.515 210.585 124.925 210.760 ;
        RECT 125.170 210.755 125.360 211.335 ;
        RECT 125.735 210.765 125.905 211.475 ;
        RECT 126.180 210.985 126.885 211.495 ;
        RECT 127.055 211.175 129.265 211.455 ;
        RECT 127.055 211.070 127.625 211.175 ;
        RECT 128.295 211.070 129.265 211.175 ;
        RECT 126.715 210.900 126.885 210.985 ;
        RECT 127.795 210.900 128.125 211.005 ;
        RECT 129.435 210.945 129.605 212.180 ;
        RECT 129.880 212.510 130.925 212.680 ;
        RECT 131.145 212.530 131.475 212.730 ;
        RECT 131.655 212.640 132.325 213.010 ;
        RECT 132.530 212.885 133.305 213.065 ;
        RECT 133.680 213.635 134.705 213.805 ;
        RECT 134.875 215.650 135.045 215.835 ;
        RECT 135.215 215.905 137.425 216.075 ;
        RECT 135.215 215.820 136.120 215.905 ;
        RECT 136.850 215.820 137.425 215.905 ;
        RECT 137.595 215.755 138.145 216.085 ;
        RECT 138.315 215.990 138.485 216.255 ;
        RECT 138.655 216.160 139.305 216.510 ;
        RECT 139.475 216.255 140.145 216.425 ;
        RECT 139.475 215.990 139.645 216.255 ;
        RECT 140.315 216.085 141.575 216.515 ;
        RECT 138.315 215.760 139.645 215.990 ;
        RECT 139.815 215.755 141.575 216.085 ;
        RECT 136.355 215.650 136.685 215.735 ;
        RECT 137.595 215.650 137.765 215.755 ;
        RECT 134.875 215.320 135.805 215.650 ;
        RECT 135.975 215.480 137.045 215.650 ;
        RECT 134.875 214.165 135.045 215.320 ;
        RECT 135.975 215.105 136.145 215.480 ;
        RECT 135.215 214.935 136.145 215.105 ;
        RECT 136.325 214.845 136.695 215.200 ;
        RECT 136.875 215.105 137.045 215.480 ;
        RECT 137.215 215.320 137.765 215.650 ;
        RECT 138.025 215.400 140.145 215.585 ;
        RECT 137.595 215.145 137.765 215.320 ;
        RECT 136.875 214.935 137.425 215.105 ;
        RECT 137.595 214.895 138.225 215.145 ;
        RECT 138.395 214.950 139.345 215.230 ;
        RECT 140.315 215.160 141.575 215.755 ;
        RECT 139.855 214.895 141.575 215.160 ;
        RECT 135.215 214.500 137.425 214.670 ;
        RECT 135.215 214.335 136.185 214.500 ;
        RECT 136.855 214.415 137.425 214.500 ;
        RECT 136.355 214.245 136.685 214.330 ;
        RECT 137.595 214.245 137.765 214.895 ;
        RECT 138.355 214.725 139.720 214.780 ;
        RECT 138.045 214.610 140.145 214.725 ;
        RECT 138.045 214.555 138.485 214.610 ;
        RECT 138.045 214.390 138.215 214.555 ;
        RECT 139.590 214.475 140.145 214.610 ;
        RECT 140.315 214.695 141.575 214.895 ;
        RECT 141.745 214.930 143.750 216.515 ;
        RECT 141.745 214.865 144.580 214.930 ;
        RECT 134.875 213.995 136.185 214.165 ;
        RECT 136.355 214.075 137.025 214.245 ;
        RECT 133.680 213.055 133.870 213.635 ;
        RECT 134.875 213.465 135.045 213.995 ;
        RECT 136.355 213.825 136.685 213.850 ;
        RECT 134.115 213.295 135.045 213.465 ;
        RECT 134.115 212.885 134.525 213.060 ;
        RECT 132.530 212.820 134.525 212.885 ;
        RECT 129.880 211.575 130.050 212.510 ;
        RECT 130.220 211.980 130.585 212.340 ;
        RECT 130.755 212.320 130.925 212.510 ;
        RECT 130.755 212.150 131.875 212.320 ;
        RECT 130.220 211.810 131.505 211.980 ;
        RECT 130.520 211.400 131.115 211.640 ;
        RECT 131.285 211.455 131.505 211.810 ;
        RECT 131.705 211.645 131.875 212.150 ;
        RECT 132.155 211.945 132.325 212.640 ;
        RECT 133.135 212.545 134.525 212.820 ;
        RECT 132.585 212.115 133.045 212.285 ;
        RECT 132.155 211.615 132.705 211.945 ;
        RECT 132.875 211.850 133.045 212.115 ;
        RECT 133.215 212.020 133.865 212.370 ;
        RECT 134.035 212.115 134.705 212.285 ;
        RECT 134.035 211.850 134.205 212.115 ;
        RECT 134.875 211.945 135.045 213.295 ;
        RECT 132.875 211.620 134.205 211.850 ;
        RECT 134.375 211.625 135.045 211.945 ;
        RECT 135.215 213.655 136.685 213.825 ;
        RECT 135.215 211.965 135.385 213.655 ;
        RECT 136.855 213.490 137.025 214.075 ;
        RECT 137.195 213.915 137.765 214.245 ;
        RECT 136.855 213.485 137.425 213.490 ;
        RECT 135.555 213.315 137.425 213.485 ;
        RECT 135.555 212.360 135.725 213.315 ;
        RECT 135.895 212.975 136.865 213.145 ;
        RECT 135.895 212.325 136.065 212.975 ;
        RECT 137.060 212.960 137.425 213.315 ;
        RECT 137.595 213.200 137.765 213.915 ;
        RECT 138.045 213.690 138.215 214.195 ;
        RECT 138.415 214.030 138.635 214.385 ;
        RECT 138.805 214.200 139.400 214.440 ;
        RECT 138.415 213.860 139.700 214.030 ;
        RECT 138.045 213.520 139.165 213.690 ;
        RECT 138.995 213.330 139.165 213.520 ;
        RECT 139.335 213.500 139.700 213.860 ;
        RECT 139.870 213.330 140.040 214.265 ;
        RECT 137.595 212.830 138.265 213.200 ;
        RECT 138.445 213.110 138.775 213.310 ;
        RECT 138.995 213.160 140.040 213.330 ;
        RECT 137.085 212.770 137.255 212.775 ;
        RECT 136.265 212.495 137.425 212.770 ;
        RECT 135.895 212.135 137.425 212.325 ;
        RECT 135.215 211.795 136.240 211.965 ;
        RECT 137.595 211.955 137.765 212.830 ;
        RECT 138.445 212.650 138.745 213.110 ;
        RECT 138.995 212.990 139.255 213.160 ;
        RECT 140.315 213.005 142.095 214.695 ;
        RECT 142.265 214.590 144.580 214.865 ;
        RECT 142.265 213.005 143.750 214.590 ;
        RECT 145.320 213.110 145.925 216.515 ;
        RECT 140.315 212.990 140.485 213.005 ;
        RECT 138.925 212.820 139.255 212.990 ;
        RECT 139.515 212.820 140.485 212.990 ;
        RECT 138.045 212.480 140.145 212.650 ;
        RECT 138.045 212.245 138.215 212.480 ;
        RECT 139.815 212.400 140.145 212.480 ;
        RECT 138.925 212.120 139.645 212.310 ;
        RECT 134.375 211.615 135.805 211.625 ;
        RECT 129.775 211.230 130.330 211.365 ;
        RECT 131.705 211.285 131.875 211.450 ;
        RECT 131.435 211.230 131.875 211.285 ;
        RECT 129.775 211.115 131.875 211.230 ;
        RECT 130.200 211.060 131.565 211.115 ;
        RECT 132.155 211.005 132.325 211.615 ;
        RECT 134.875 211.455 135.805 211.615 ;
        RECT 132.585 211.260 134.705 211.445 ;
        RECT 132.155 210.945 132.785 211.005 ;
        RECT 129.435 210.900 130.065 210.945 ;
        RECT 125.735 210.585 126.510 210.765 ;
        RECT 124.515 210.520 126.510 210.585 ;
        RECT 126.715 210.575 127.345 210.900 ;
        RECT 124.515 210.245 125.905 210.520 ;
        RECT 122.985 209.885 124.165 210.055 ;
        RECT 121.665 209.495 122.225 209.550 ;
        RECT 122.855 209.540 123.780 209.715 ;
        RECT 122.805 209.495 123.780 209.540 ;
        RECT 121.665 209.385 123.780 209.495 ;
        RECT 123.995 209.645 124.165 209.885 ;
        RECT 124.335 209.815 125.005 209.985 ;
        RECT 121.665 209.375 122.935 209.385 ;
        RECT 122.100 209.325 122.935 209.375 ;
        RECT 123.995 209.315 124.665 209.645 ;
        RECT 124.835 209.550 125.005 209.815 ;
        RECT 125.175 209.720 125.825 210.070 ;
        RECT 125.995 209.815 126.455 209.985 ;
        RECT 125.995 209.550 126.165 209.815 ;
        RECT 126.715 209.645 126.885 210.575 ;
        RECT 127.515 210.450 128.805 210.900 ;
        RECT 128.975 210.680 130.065 210.900 ;
        RECT 128.975 210.575 129.605 210.680 ;
        RECT 130.575 210.610 131.525 210.890 ;
        RECT 131.695 210.755 132.785 210.945 ;
        RECT 132.955 210.810 133.905 211.090 ;
        RECT 134.875 211.020 135.045 211.455 ;
        RECT 134.415 210.755 135.045 211.020 ;
        RECT 131.695 210.695 132.325 210.755 ;
        RECT 127.515 210.055 127.685 210.450 ;
        RECT 127.055 209.775 127.685 210.055 ;
        RECT 124.835 209.320 126.165 209.550 ;
        RECT 126.335 209.315 126.885 209.645 ;
        RECT 127.855 209.585 128.415 210.280 ;
        RECT 128.585 210.055 128.805 210.450 ;
        RECT 129.435 210.085 129.605 210.575 ;
        RECT 129.775 210.255 131.895 210.440 ;
        RECT 132.155 210.085 132.325 210.695 ;
        RECT 132.915 210.585 134.280 210.640 ;
        RECT 132.605 210.470 134.705 210.585 ;
        RECT 132.605 210.415 133.045 210.470 ;
        RECT 132.605 210.250 132.775 210.415 ;
        RECT 134.150 210.335 134.705 210.470 ;
        RECT 134.875 210.535 135.045 210.755 ;
        RECT 135.395 211.045 135.805 211.220 ;
        RECT 136.050 211.215 136.240 211.795 ;
        RECT 136.615 211.225 136.785 211.935 ;
        RECT 137.060 211.445 137.765 211.955 ;
        RECT 136.615 211.045 137.390 211.225 ;
        RECT 135.395 210.980 137.390 211.045 ;
        RECT 137.595 211.015 137.765 211.445 ;
        RECT 138.045 211.460 138.215 212.075 ;
        RECT 138.385 211.950 138.715 212.095 ;
        RECT 138.385 211.630 139.675 211.950 ;
        RECT 139.845 211.460 140.015 212.175 ;
        RECT 138.045 211.290 140.015 211.460 ;
        RECT 140.315 211.815 140.485 212.820 ;
        RECT 141.545 212.325 142.380 212.375 ;
        RECT 141.545 212.315 142.815 212.325 ;
        RECT 140.700 212.205 142.815 212.315 ;
        RECT 140.700 212.160 141.675 212.205 ;
        RECT 140.700 211.985 141.625 212.160 ;
        RECT 142.255 212.150 142.815 212.205 ;
        RECT 140.315 211.645 141.495 211.815 ;
        RECT 135.395 210.705 136.785 210.980 ;
        RECT 137.595 210.805 138.295 211.015 ;
        RECT 137.595 210.535 137.765 210.805 ;
        RECT 138.675 210.585 139.005 211.290 ;
        RECT 139.210 210.565 139.585 211.120 ;
        RECT 140.315 211.110 140.485 211.645 ;
        RECT 141.795 211.485 142.125 212.035 ;
        RECT 142.295 211.995 142.815 212.150 ;
        RECT 143.035 211.825 143.750 213.005 ;
        RECT 144.070 212.760 145.925 213.110 ;
        RECT 142.425 211.655 143.750 211.825 ;
        RECT 141.795 211.475 142.820 211.485 ;
        RECT 140.655 211.285 142.820 211.475 ;
        RECT 140.655 211.135 141.590 211.285 ;
        RECT 142.295 211.155 142.820 211.285 ;
        RECT 143.035 211.170 143.750 211.655 ;
        RECT 145.320 211.170 145.925 212.760 ;
        RECT 139.815 210.905 140.485 211.110 ;
        RECT 139.815 210.795 140.985 210.905 ;
        RECT 140.315 210.590 140.985 210.795 ;
        RECT 128.585 209.775 129.265 210.055 ;
        RECT 129.435 209.755 130.105 210.085 ;
        RECT 130.275 209.850 131.605 210.080 ;
        RECT 123.995 209.155 124.165 209.315 ;
        RECT 114.545 207.965 117.295 209.155 ;
        RECT 111.505 207.485 114.895 207.795 ;
        RECT 110.395 206.380 110.565 207.485 ;
        RECT 110.735 206.595 111.285 206.765 ;
        RECT 110.395 206.050 110.945 206.380 ;
        RECT 111.115 206.220 111.285 206.595 ;
        RECT 111.465 206.500 111.835 206.855 ;
        RECT 112.015 206.595 112.945 206.765 ;
        RECT 112.015 206.220 112.185 206.595 ;
        RECT 113.115 206.380 114.895 207.485 ;
        RECT 111.115 206.050 112.185 206.220 ;
        RECT 112.355 206.105 114.895 206.380 ;
        RECT 115.065 207.505 117.295 207.965 ;
        RECT 117.465 208.585 118.725 209.155 ;
        RECT 118.895 208.755 119.575 209.040 ;
        RECT 117.465 208.315 119.185 208.585 ;
        RECT 115.065 206.105 116.775 207.505 ;
        RECT 117.465 207.335 118.725 208.315 ;
        RECT 119.355 208.295 119.575 208.755 ;
        RECT 119.745 208.465 120.305 209.155 ;
        RECT 120.475 208.755 121.105 209.040 ;
        RECT 120.475 208.295 120.645 208.755 ;
        RECT 121.275 208.585 122.735 209.155 ;
        RECT 120.815 208.315 122.735 208.585 ;
        RECT 119.355 208.085 120.645 208.295 ;
        RECT 118.895 207.515 121.105 207.915 ;
        RECT 112.355 206.050 113.285 206.105 ;
        RECT 110.395 205.450 110.565 206.050 ;
        RECT 111.475 205.965 111.805 206.050 ;
        RECT 113.115 205.935 113.285 206.050 ;
        RECT 115.835 205.935 116.775 206.105 ;
        RECT 110.735 205.795 111.310 205.880 ;
        RECT 112.040 205.795 112.945 205.880 ;
        RECT 110.735 205.625 112.945 205.795 ;
        RECT 113.115 205.450 114.375 205.935 ;
        RECT 110.395 205.190 111.405 205.450 ;
        RECT 111.965 205.245 114.375 205.450 ;
        RECT 114.545 205.645 116.775 205.935 ;
        RECT 116.945 206.525 118.725 207.335 ;
        RECT 118.895 207.045 119.575 207.325 ;
        RECT 119.355 206.650 119.575 207.045 ;
        RECT 119.745 206.820 120.305 207.515 ;
        RECT 121.275 207.505 122.735 208.315 ;
        RECT 122.905 208.720 124.165 209.155 ;
        RECT 124.335 208.960 126.455 209.145 ;
        RECT 122.905 208.455 124.625 208.720 ;
        RECT 125.135 208.510 126.085 208.790 ;
        RECT 126.715 208.785 126.885 209.315 ;
        RECT 127.055 209.185 129.265 209.585 ;
        RECT 129.435 209.155 129.605 209.755 ;
        RECT 130.275 209.585 130.445 209.850 ;
        RECT 129.775 209.415 130.445 209.585 ;
        RECT 130.615 209.330 131.265 209.680 ;
        RECT 131.435 209.585 131.605 209.850 ;
        RECT 131.775 209.755 132.325 210.085 ;
        RECT 131.435 209.415 131.895 209.585 ;
        RECT 132.155 209.155 132.325 209.755 ;
        RECT 132.605 209.550 132.775 210.055 ;
        RECT 132.975 209.890 133.195 210.245 ;
        RECT 133.365 210.060 133.960 210.300 ;
        RECT 132.975 209.720 134.260 209.890 ;
        RECT 132.605 209.380 133.725 209.550 ;
        RECT 133.555 209.190 133.725 209.380 ;
        RECT 133.895 209.360 134.260 209.720 ;
        RECT 134.430 209.190 134.600 210.125 ;
        RECT 127.515 208.805 128.805 209.015 ;
        RECT 126.715 208.705 127.345 208.785 ;
        RECT 126.255 208.515 127.345 208.705 ;
        RECT 126.255 208.455 126.885 208.515 ;
        RECT 120.475 207.045 121.105 207.325 ;
        RECT 120.475 206.650 120.645 207.045 ;
        RECT 116.945 206.200 119.185 206.525 ;
        RECT 119.355 206.200 120.645 206.650 ;
        RECT 121.275 206.525 122.215 207.505 ;
        RECT 122.905 207.335 124.165 208.455 ;
        RECT 124.760 208.285 126.125 208.340 ;
        RECT 124.335 208.170 126.435 208.285 ;
        RECT 124.335 208.035 124.890 208.170 ;
        RECT 125.995 208.115 126.435 208.170 ;
        RECT 120.815 206.200 122.215 206.525 ;
        RECT 116.945 205.645 118.725 206.200 ;
        RECT 120.035 206.095 120.365 206.200 ;
        RECT 118.895 205.925 119.865 206.030 ;
        RECT 120.535 205.925 121.105 206.030 ;
        RECT 118.895 205.645 121.105 205.925 ;
        RECT 121.275 205.645 122.215 206.200 ;
        RECT 122.385 206.550 124.165 207.335 ;
        RECT 124.440 206.890 124.610 207.825 ;
        RECT 125.080 207.760 125.675 208.000 ;
        RECT 126.265 207.950 126.435 208.115 ;
        RECT 125.845 207.590 126.065 207.945 ;
        RECT 126.715 207.775 126.885 208.455 ;
        RECT 127.515 208.345 127.685 208.805 ;
        RECT 127.055 208.060 127.685 208.345 ;
        RECT 127.855 207.945 128.415 208.635 ;
        RECT 128.585 208.345 128.805 208.805 ;
        RECT 129.435 208.785 130.695 209.155 ;
        RECT 128.975 208.515 130.695 208.785 ;
        RECT 128.585 208.060 129.265 208.345 ;
        RECT 129.435 207.775 130.695 208.515 ;
        RECT 130.865 209.060 132.325 209.155 ;
        RECT 130.865 208.690 132.825 209.060 ;
        RECT 133.005 208.970 133.335 209.170 ;
        RECT 133.555 209.020 134.600 209.190 ;
        RECT 134.875 209.845 136.135 210.535 ;
        RECT 136.305 210.045 137.765 210.535 ;
        RECT 137.980 210.415 138.505 210.545 ;
        RECT 139.210 210.415 140.145 210.565 ;
        RECT 137.980 210.225 140.145 210.415 ;
        RECT 137.980 210.215 139.005 210.225 ;
        RECT 136.305 210.015 138.375 210.045 ;
        RECT 136.845 209.875 138.375 210.015 ;
        RECT 134.875 209.325 136.675 209.845 ;
        RECT 136.845 209.325 137.765 209.875 ;
        RECT 137.985 209.550 138.505 209.705 ;
        RECT 138.675 209.665 139.005 210.215 ;
        RECT 140.315 210.055 140.485 210.590 ;
        RECT 141.215 210.580 141.590 211.135 ;
        RECT 141.795 210.410 142.125 211.115 ;
        RECT 143.035 210.895 143.205 211.170 ;
        RECT 142.505 210.685 143.205 210.895 ;
        RECT 139.305 209.885 140.485 210.055 ;
        RECT 137.985 209.495 138.545 209.550 ;
        RECT 139.175 209.540 140.100 209.715 ;
        RECT 139.125 209.495 140.100 209.540 ;
        RECT 137.985 209.385 140.100 209.495 ;
        RECT 137.985 209.375 139.255 209.385 ;
        RECT 138.420 209.325 139.255 209.375 ;
        RECT 134.875 209.065 135.045 209.325 ;
        RECT 137.595 209.065 137.765 209.325 ;
        RECT 130.865 207.945 132.325 208.690 ;
        RECT 133.005 208.510 133.305 208.970 ;
        RECT 133.555 208.850 133.815 209.020 ;
        RECT 134.875 208.850 135.790 209.065 ;
        RECT 133.485 208.680 133.815 208.850 ;
        RECT 134.075 208.795 135.790 208.850 ;
        RECT 134.075 208.680 135.045 208.795 ;
        RECT 132.605 208.340 134.705 208.510 ;
        RECT 132.605 208.105 132.775 208.340 ;
        RECT 134.375 208.260 134.705 208.340 ;
        RECT 133.485 207.980 134.205 208.170 ;
        RECT 134.875 208.165 135.045 208.680 ;
        RECT 135.960 208.625 136.945 209.065 ;
        RECT 137.115 208.765 137.765 209.065 ;
        RECT 137.935 208.875 140.145 209.155 ;
        RECT 137.935 208.770 138.505 208.875 ;
        RECT 139.175 208.770 140.145 208.875 ;
        RECT 140.315 208.880 140.485 209.885 ;
        RECT 140.785 210.240 142.755 210.410 ;
        RECT 140.785 209.525 140.955 210.240 ;
        RECT 141.125 209.750 142.415 210.070 ;
        RECT 142.085 209.605 142.415 209.750 ;
        RECT 142.585 209.625 142.755 210.240 ;
        RECT 143.035 209.600 143.205 210.685 ;
        RECT 143.375 209.815 143.925 209.985 ;
        RECT 141.155 209.390 141.875 209.580 ;
        RECT 140.655 209.220 140.985 209.300 ;
        RECT 142.585 209.220 142.755 209.455 ;
        RECT 140.655 209.050 142.755 209.220 ;
        RECT 143.035 209.270 143.585 209.600 ;
        RECT 143.755 209.440 143.925 209.815 ;
        RECT 144.105 209.720 144.475 210.075 ;
        RECT 144.655 209.815 145.585 209.985 ;
        RECT 144.655 209.440 144.825 209.815 ;
        RECT 145.755 209.600 145.925 211.170 ;
        RECT 143.755 209.270 144.825 209.440 ;
        RECT 144.995 209.270 145.925 209.600 ;
        RECT 135.220 208.595 136.945 208.625 ;
        RECT 137.595 208.600 137.765 208.765 ;
        RECT 140.315 208.710 141.285 208.880 ;
        RECT 141.545 208.710 141.875 208.880 ;
        RECT 138.675 208.600 139.005 208.705 ;
        RECT 140.315 208.600 140.485 208.710 ;
        RECT 135.220 208.335 137.400 208.595 ;
        RECT 124.780 207.420 126.065 207.590 ;
        RECT 124.780 207.060 125.145 207.420 ;
        RECT 126.265 207.250 126.435 207.755 ;
        RECT 125.315 207.080 126.435 207.250 ;
        RECT 125.315 206.890 125.485 207.080 ;
        RECT 124.440 206.720 125.485 206.890 ;
        RECT 125.225 206.550 125.485 206.720 ;
        RECT 125.705 206.670 126.035 206.870 ;
        RECT 126.715 206.760 128.175 207.775 ;
        RECT 122.385 206.380 124.965 206.550 ;
        RECT 125.225 206.380 125.555 206.550 ;
        RECT 122.385 205.645 124.165 206.380 ;
        RECT 125.735 206.210 126.035 206.670 ;
        RECT 126.215 206.565 128.175 206.760 ;
        RECT 128.345 206.565 131.215 207.775 ;
        RECT 131.385 206.875 132.325 207.945 ;
        RECT 132.605 207.320 132.775 207.935 ;
        RECT 132.945 207.810 133.275 207.955 ;
        RECT 132.945 207.490 134.235 207.810 ;
        RECT 134.405 207.320 134.575 208.035 ;
        RECT 132.605 207.150 134.575 207.320 ;
        RECT 134.875 207.910 135.775 208.165 ;
        RECT 134.875 207.295 135.050 207.910 ;
        RECT 135.960 207.900 136.945 208.335 ;
        RECT 137.595 208.275 138.225 208.600 ;
        RECT 137.595 208.165 137.765 208.275 ;
        RECT 137.115 207.905 137.765 208.165 ;
        RECT 135.960 207.725 136.185 207.900 ;
        RECT 135.220 207.465 136.185 207.725 ;
        RECT 131.385 206.665 132.855 206.875 ;
        RECT 131.385 206.565 132.325 206.665 ;
        RECT 126.215 206.390 127.655 206.565 ;
        RECT 128.345 206.395 129.605 206.565 ;
        RECT 124.335 206.040 126.435 206.210 ;
        RECT 124.335 205.960 124.665 206.040 ;
        RECT 114.545 205.415 116.005 205.645 ;
        RECT 111.965 205.190 114.915 205.245 ;
        RECT 110.395 205.015 110.565 205.190 ;
        RECT 113.115 205.015 114.915 205.190 ;
        RECT 110.395 204.725 111.290 205.015 ;
        RECT 111.950 204.725 114.915 205.015 ;
        RECT 115.085 205.015 116.005 205.415 ;
        RECT 118.555 205.015 118.725 205.645 ;
        RECT 115.085 204.725 116.730 205.015 ;
        RECT 117.390 204.725 118.725 205.015 ;
        RECT 119.075 205.200 120.465 205.475 ;
        RECT 119.075 205.135 121.070 205.200 ;
        RECT 119.075 204.960 119.485 205.135 ;
        RECT 110.395 204.090 110.565 204.725 ;
        RECT 113.115 204.090 113.285 204.725 ;
        RECT 115.835 204.555 116.005 204.725 ;
        RECT 118.555 204.555 119.485 204.725 ;
        RECT 114.345 204.505 115.180 204.555 ;
        RECT 114.345 204.495 115.615 204.505 ;
        RECT 113.500 204.385 115.615 204.495 ;
        RECT 113.500 204.340 114.475 204.385 ;
        RECT 113.500 204.165 114.425 204.340 ;
        RECT 115.055 204.330 115.615 204.385 ;
        RECT 110.395 203.830 111.405 204.090 ;
        RECT 111.965 203.995 113.285 204.090 ;
        RECT 111.965 203.830 114.295 203.995 ;
        RECT 110.395 203.230 110.565 203.830 ;
        RECT 113.115 203.825 114.295 203.830 ;
        RECT 110.735 203.485 112.945 203.655 ;
        RECT 110.735 203.400 111.310 203.485 ;
        RECT 112.040 203.400 112.945 203.485 ;
        RECT 111.475 203.230 111.805 203.315 ;
        RECT 113.115 203.230 113.285 203.825 ;
        RECT 114.595 203.665 114.925 204.215 ;
        RECT 115.095 204.175 115.615 204.330 ;
        RECT 115.835 204.250 116.515 204.555 ;
        RECT 115.835 204.005 116.005 204.250 ;
        RECT 116.685 204.240 117.245 204.555 ;
        RECT 118.555 204.545 118.725 204.555 ;
        RECT 117.745 204.250 118.725 204.545 ;
        RECT 119.730 204.385 119.920 204.965 ;
        RECT 115.225 203.835 116.005 204.005 ;
        RECT 114.595 203.655 115.620 203.665 ;
        RECT 113.455 203.465 115.620 203.655 ;
        RECT 113.455 203.315 114.390 203.465 ;
        RECT 115.095 203.335 115.620 203.465 ;
        RECT 115.835 203.650 116.005 203.835 ;
        RECT 116.185 203.825 118.385 204.070 ;
        RECT 116.185 203.820 117.245 203.825 ;
        RECT 115.835 203.390 116.530 203.650 ;
        RECT 110.395 202.900 110.945 203.230 ;
        RECT 111.115 203.060 112.185 203.230 ;
        RECT 110.395 201.825 110.565 202.900 ;
        RECT 111.115 202.685 111.285 203.060 ;
        RECT 110.735 202.515 111.285 202.685 ;
        RECT 111.465 202.425 111.835 202.780 ;
        RECT 112.015 202.685 112.185 203.060 ;
        RECT 112.355 203.085 113.285 203.230 ;
        RECT 112.355 202.900 113.785 203.085 ;
        RECT 113.115 202.770 113.785 202.900 ;
        RECT 112.015 202.515 112.945 202.685 ;
        RECT 110.825 201.995 111.285 202.165 ;
        RECT 110.395 201.495 110.945 201.825 ;
        RECT 111.115 201.730 111.285 201.995 ;
        RECT 111.455 201.900 112.105 202.250 ;
        RECT 112.275 201.995 112.945 202.165 ;
        RECT 112.275 201.730 112.445 201.995 ;
        RECT 113.115 201.825 113.285 202.770 ;
        RECT 114.015 202.760 114.390 203.315 ;
        RECT 114.595 202.590 114.925 203.295 ;
        RECT 115.835 203.075 116.005 203.390 ;
        RECT 116.995 203.210 117.245 203.820 ;
        RECT 118.555 203.650 118.725 204.250 ;
        RECT 117.745 203.390 118.725 203.650 ;
        RECT 115.305 202.865 116.005 203.075 ;
        RECT 116.185 202.960 118.380 203.210 ;
        RECT 115.835 202.790 116.005 202.865 ;
        RECT 111.115 201.500 112.445 201.730 ;
        RECT 112.615 201.495 113.285 201.825 ;
        RECT 113.585 202.420 115.555 202.590 ;
        RECT 113.585 201.705 113.755 202.420 ;
        RECT 113.925 201.930 115.215 202.250 ;
        RECT 114.885 201.785 115.215 201.930 ;
        RECT 115.385 201.805 115.555 202.420 ;
        RECT 115.835 202.530 116.565 202.790 ;
        RECT 115.835 201.930 116.005 202.530 ;
        RECT 116.200 202.100 116.825 202.360 ;
        RECT 113.955 201.570 114.675 201.760 ;
        RECT 115.835 201.670 116.485 201.930 ;
        RECT 110.395 200.885 110.565 201.495 ;
        RECT 110.825 201.140 112.945 201.325 ;
        RECT 113.115 201.060 113.285 201.495 ;
        RECT 113.455 201.400 113.785 201.480 ;
        RECT 115.385 201.400 115.555 201.635 ;
        RECT 113.455 201.230 115.555 201.400 ;
        RECT 110.395 200.635 111.025 200.885 ;
        RECT 111.195 200.690 112.145 200.970 ;
        RECT 113.115 200.900 114.085 201.060 ;
        RECT 112.655 200.890 114.085 200.900 ;
        RECT 114.345 200.890 114.675 201.060 ;
        RECT 112.655 200.635 113.285 200.890 ;
        RECT 114.345 200.720 114.605 200.890 ;
        RECT 114.855 200.770 115.155 201.230 ;
        RECT 115.835 201.070 116.005 201.670 ;
        RECT 116.655 201.500 116.825 202.100 ;
        RECT 116.200 201.240 116.825 201.500 ;
        RECT 115.835 201.050 116.485 201.070 ;
        RECT 110.395 198.940 110.565 200.635 ;
        RECT 111.155 200.465 112.520 200.520 ;
        RECT 110.845 200.350 112.945 200.465 ;
        RECT 110.845 200.295 111.285 200.350 ;
        RECT 110.845 200.130 111.015 200.295 ;
        RECT 112.390 200.215 112.945 200.350 ;
        RECT 110.845 199.430 111.015 199.935 ;
        RECT 111.215 199.770 111.435 200.125 ;
        RECT 111.605 199.940 112.200 200.180 ;
        RECT 111.215 199.600 112.500 199.770 ;
        RECT 110.845 199.260 111.965 199.430 ;
        RECT 111.795 199.070 111.965 199.260 ;
        RECT 112.135 199.240 112.500 199.600 ;
        RECT 112.670 199.070 112.840 200.005 ;
        RECT 110.395 198.570 111.065 198.940 ;
        RECT 111.245 198.850 111.575 199.050 ;
        RECT 111.795 198.900 112.840 199.070 ;
        RECT 113.115 198.985 113.285 200.635 ;
        RECT 113.560 200.550 114.605 200.720 ;
        RECT 114.825 200.570 115.155 200.770 ;
        RECT 115.335 200.810 116.485 201.050 ;
        RECT 115.335 200.680 116.005 200.810 ;
        RECT 113.560 199.615 113.730 200.550 ;
        RECT 113.900 200.020 114.265 200.380 ;
        RECT 114.435 200.360 114.605 200.550 ;
        RECT 114.435 200.190 115.555 200.360 ;
        RECT 113.900 199.850 115.185 200.020 ;
        RECT 114.200 199.440 114.795 199.680 ;
        RECT 114.965 199.495 115.185 199.850 ;
        RECT 115.385 199.685 115.555 200.190 ;
        RECT 115.835 200.210 116.005 200.680 ;
        RECT 116.655 200.640 116.825 201.240 ;
        RECT 116.200 200.380 116.825 200.640 ;
        RECT 115.835 199.965 116.485 200.210 ;
        RECT 113.455 199.270 114.010 199.405 ;
        RECT 115.385 199.325 115.555 199.490 ;
        RECT 115.115 199.270 115.555 199.325 ;
        RECT 113.455 199.155 115.555 199.270 ;
        RECT 115.835 199.350 116.005 199.965 ;
        RECT 116.655 199.795 116.825 200.380 ;
        RECT 116.200 199.520 116.825 199.795 ;
        RECT 113.880 199.100 115.245 199.155 ;
        RECT 115.835 199.105 116.485 199.350 ;
        RECT 115.835 198.985 116.005 199.105 ;
        RECT 110.395 196.755 110.565 198.570 ;
        RECT 111.245 198.390 111.545 198.850 ;
        RECT 111.795 198.730 112.055 198.900 ;
        RECT 113.115 198.730 113.745 198.985 ;
        RECT 111.725 198.560 112.055 198.730 ;
        RECT 112.315 198.720 113.745 198.730 ;
        RECT 112.315 198.560 113.285 198.720 ;
        RECT 114.255 198.650 115.205 198.930 ;
        RECT 115.375 198.735 116.005 198.985 ;
        RECT 116.655 198.935 116.825 199.520 ;
        RECT 110.845 198.220 112.945 198.390 ;
        RECT 110.845 197.985 111.015 198.220 ;
        RECT 112.615 198.140 112.945 198.220 ;
        RECT 113.115 198.125 113.285 198.560 ;
        RECT 115.835 198.495 116.005 198.735 ;
        RECT 116.200 198.675 116.825 198.935 ;
        RECT 113.455 198.295 115.575 198.480 ;
        RECT 115.835 198.245 116.485 198.495 ;
        RECT 115.835 198.125 116.005 198.245 ;
        RECT 111.725 197.860 112.445 198.050 ;
        RECT 110.845 197.200 111.015 197.815 ;
        RECT 111.185 197.690 111.515 197.835 ;
        RECT 111.185 197.370 112.475 197.690 ;
        RECT 112.645 197.200 112.815 197.915 ;
        RECT 110.845 197.030 112.815 197.200 ;
        RECT 113.115 197.795 113.785 198.125 ;
        RECT 113.955 197.890 115.285 198.120 ;
        RECT 110.395 196.545 111.095 196.755 ;
        RECT 110.395 195.785 110.565 196.545 ;
        RECT 111.475 196.325 111.805 197.030 ;
        RECT 112.010 196.305 112.385 196.860 ;
        RECT 113.115 196.850 113.285 197.795 ;
        RECT 113.955 197.625 114.125 197.890 ;
        RECT 113.455 197.455 114.125 197.625 ;
        RECT 114.295 197.370 114.945 197.720 ;
        RECT 115.115 197.625 115.285 197.890 ;
        RECT 115.455 197.795 116.005 198.125 ;
        RECT 116.655 198.075 116.825 198.675 ;
        RECT 116.200 197.815 116.825 198.075 ;
        RECT 115.835 197.635 116.005 197.795 ;
        RECT 115.115 197.455 115.575 197.625 ;
        RECT 115.835 197.385 116.485 197.635 ;
        RECT 113.455 197.020 115.665 197.190 ;
        RECT 113.455 196.855 114.425 197.020 ;
        RECT 115.095 196.935 115.665 197.020 ;
        RECT 112.615 196.685 113.285 196.850 ;
        RECT 114.595 196.765 114.925 196.850 ;
        RECT 115.835 196.775 116.005 197.385 ;
        RECT 116.655 197.215 116.825 197.815 ;
        RECT 116.200 196.955 116.825 197.215 ;
        RECT 116.655 196.780 116.825 196.955 ;
        RECT 116.995 196.950 117.245 202.960 ;
        RECT 118.555 202.790 118.725 203.390 ;
        RECT 117.755 202.530 118.725 202.790 ;
        RECT 117.415 202.100 118.380 202.360 ;
        RECT 118.550 202.185 118.725 202.530 ;
        RECT 118.895 204.215 119.920 204.385 ;
        RECT 120.295 204.955 121.070 205.135 ;
        RECT 121.275 205.015 121.445 205.645 ;
        RECT 123.995 205.015 124.165 205.645 ;
        RECT 120.295 204.245 120.465 204.955 ;
        RECT 121.275 204.735 122.170 205.015 ;
        RECT 120.740 204.725 122.170 204.735 ;
        RECT 122.830 204.725 124.165 205.015 ;
        RECT 124.465 205.020 124.635 205.735 ;
        RECT 124.835 205.680 125.555 205.870 ;
        RECT 126.265 205.805 126.435 206.040 ;
        RECT 125.765 205.510 126.095 205.655 ;
        RECT 124.805 205.190 126.095 205.510 ;
        RECT 126.265 205.020 126.435 205.635 ;
        RECT 124.465 204.850 126.435 205.020 ;
        RECT 126.715 205.185 127.655 206.390 ;
        RECT 127.825 205.925 129.605 206.395 ;
        RECT 132.155 205.935 132.325 206.565 ;
        RECT 133.235 206.445 133.565 207.150 ;
        RECT 134.875 207.050 135.775 207.295 ;
        RECT 133.770 206.425 134.145 206.980 ;
        RECT 134.875 206.970 135.050 207.050 ;
        RECT 134.375 206.655 135.050 206.970 ;
        RECT 135.945 206.865 136.185 207.465 ;
        RECT 134.875 206.435 135.050 206.655 ;
        RECT 135.220 206.605 136.185 206.865 ;
        RECT 132.540 206.275 133.065 206.405 ;
        RECT 133.770 206.275 134.705 206.425 ;
        RECT 132.540 206.085 134.705 206.275 ;
        RECT 134.875 206.190 135.775 206.435 ;
        RECT 132.540 206.075 133.565 206.085 ;
        RECT 127.825 205.630 130.415 205.925 ;
        RECT 127.825 205.185 129.605 205.630 ;
        RECT 130.915 205.620 131.475 205.935 ;
        RECT 131.645 205.905 132.325 205.935 ;
        RECT 131.645 205.735 132.935 205.905 ;
        RECT 131.645 205.630 132.325 205.735 ;
        RECT 129.775 205.205 131.975 205.450 ;
        RECT 126.715 205.015 126.885 205.185 ;
        RECT 129.435 205.030 129.605 205.185 ;
        RECT 130.915 205.200 131.975 205.205 ;
        RECT 129.435 205.015 130.415 205.030 ;
        RECT 120.740 204.225 121.445 204.725 ;
        RECT 123.995 204.670 124.165 204.725 ;
        RECT 121.705 204.295 122.165 204.465 ;
        RECT 118.895 202.525 119.065 204.215 ;
        RECT 121.275 204.125 121.445 204.225 ;
        RECT 119.575 203.855 121.105 204.045 ;
        RECT 119.235 202.865 119.405 203.820 ;
        RECT 119.575 203.205 119.745 203.855 ;
        RECT 121.275 203.795 121.825 204.125 ;
        RECT 121.995 204.030 122.165 204.295 ;
        RECT 122.335 204.200 122.985 204.550 ;
        RECT 123.155 204.295 123.825 204.465 ;
        RECT 123.995 204.355 124.665 204.670 ;
        RECT 123.155 204.030 123.325 204.295 ;
        RECT 123.995 204.125 124.165 204.355 ;
        RECT 124.895 204.125 125.270 204.680 ;
        RECT 125.475 204.145 125.805 204.850 ;
        RECT 126.715 204.725 127.610 205.015 ;
        RECT 128.270 204.770 130.415 205.015 ;
        RECT 128.270 204.725 129.605 204.770 ;
        RECT 126.715 204.575 126.885 204.725 ;
        RECT 126.185 204.545 126.885 204.575 ;
        RECT 126.185 204.365 127.695 204.545 ;
        RECT 126.715 204.275 127.695 204.365 ;
        RECT 121.995 203.800 123.325 204.030 ;
        RECT 123.495 203.795 124.165 204.125 ;
        RECT 119.945 203.410 121.105 203.685 ;
        RECT 120.085 203.405 120.255 203.410 ;
        RECT 119.575 203.035 120.545 203.205 ;
        RECT 120.740 202.865 121.105 203.220 ;
        RECT 119.235 202.695 121.105 202.865 ;
        RECT 120.535 202.690 121.105 202.695 ;
        RECT 121.275 203.185 121.445 203.795 ;
        RECT 121.705 203.440 123.825 203.625 ;
        RECT 123.995 203.615 124.165 203.795 ;
        RECT 124.335 203.975 125.270 204.125 ;
        RECT 125.975 203.975 126.500 204.105 ;
        RECT 124.335 203.785 126.500 203.975 ;
        RECT 125.475 203.775 126.500 203.785 ;
        RECT 123.995 203.445 125.175 203.615 ;
        RECT 121.275 202.935 121.905 203.185 ;
        RECT 122.075 202.990 123.025 203.270 ;
        RECT 123.995 203.200 124.165 203.445 ;
        RECT 123.535 202.935 124.165 203.200 ;
        RECT 124.380 203.100 125.305 203.275 ;
        RECT 125.475 203.225 125.805 203.775 ;
        RECT 126.715 203.605 126.885 204.275 ;
        RECT 127.875 204.205 128.125 204.555 ;
        RECT 129.435 204.545 129.605 204.725 ;
        RECT 130.915 204.590 131.165 205.200 ;
        RECT 132.155 205.030 132.325 205.630 ;
        RECT 132.545 205.410 133.065 205.565 ;
        RECT 133.235 205.525 133.565 206.075 ;
        RECT 134.875 205.915 135.050 206.190 ;
        RECT 135.945 206.005 136.185 206.605 ;
        RECT 133.865 205.745 135.050 205.915 ;
        RECT 135.220 205.745 136.185 206.005 ;
        RECT 134.875 205.575 135.050 205.745 ;
        RECT 132.545 205.355 133.105 205.410 ;
        RECT 133.735 205.400 134.660 205.575 ;
        RECT 133.685 205.355 134.660 205.400 ;
        RECT 132.545 205.245 134.660 205.355 ;
        RECT 134.875 205.330 135.775 205.575 ;
        RECT 132.545 205.235 133.815 205.245 ;
        RECT 132.980 205.185 133.815 205.235 ;
        RECT 131.630 205.015 132.325 205.030 ;
        RECT 134.875 205.015 135.050 205.330 ;
        RECT 135.945 205.160 136.185 205.745 ;
        RECT 131.630 204.770 133.050 205.015 ;
        RECT 132.155 204.725 133.050 204.770 ;
        RECT 133.710 204.730 135.050 205.015 ;
        RECT 135.220 204.900 136.185 205.160 ;
        RECT 133.710 204.725 135.775 204.730 ;
        RECT 128.295 204.215 129.605 204.545 ;
        RECT 129.780 204.340 131.975 204.590 ;
        RECT 129.435 204.170 129.605 204.215 ;
        RECT 127.055 204.035 127.695 204.105 ;
        RECT 127.055 203.865 128.465 204.035 ;
        RECT 127.055 203.775 127.695 203.865 ;
        RECT 126.105 203.435 127.695 203.605 ;
        RECT 126.715 203.365 127.695 203.435 ;
        RECT 125.975 203.110 126.495 203.265 ;
        RECT 124.380 203.055 125.355 203.100 ;
        RECT 125.935 203.055 126.495 203.110 ;
        RECT 124.380 202.945 126.495 203.055 ;
        RECT 118.895 202.355 120.365 202.525 ;
        RECT 120.035 202.330 120.365 202.355 ;
        RECT 117.415 201.500 117.655 202.100 ;
        RECT 118.550 202.015 119.865 202.185 ;
        RECT 120.535 202.105 120.705 202.690 ;
        RECT 121.275 202.265 121.445 202.935 ;
        RECT 122.035 202.765 123.400 202.820 ;
        RECT 121.725 202.650 123.825 202.765 ;
        RECT 121.725 202.595 122.165 202.650 ;
        RECT 121.725 202.430 121.895 202.595 ;
        RECT 123.270 202.515 123.825 202.650 ;
        RECT 118.550 201.930 118.725 202.015 ;
        RECT 117.825 201.670 118.725 201.930 ;
        RECT 120.035 201.935 120.705 202.105 ;
        RECT 120.875 201.935 121.445 202.265 ;
        RECT 120.035 201.850 120.365 201.935 ;
        RECT 117.415 201.240 118.380 201.500 ;
        RECT 118.550 201.335 118.725 201.670 ;
        RECT 118.895 201.680 119.865 201.845 ;
        RECT 120.535 201.680 121.105 201.765 ;
        RECT 118.895 201.510 121.105 201.680 ;
        RECT 121.275 201.335 121.445 201.935 ;
        RECT 121.725 201.730 121.895 202.235 ;
        RECT 122.095 202.070 122.315 202.425 ;
        RECT 122.485 202.240 123.080 202.480 ;
        RECT 122.095 201.900 123.380 202.070 ;
        RECT 121.725 201.560 122.845 201.730 ;
        RECT 122.675 201.370 122.845 201.560 ;
        RECT 123.015 201.540 123.380 201.900 ;
        RECT 123.550 201.370 123.720 202.305 ;
        RECT 117.415 200.640 117.655 201.240 ;
        RECT 118.550 201.070 119.815 201.335 ;
        RECT 117.825 200.810 119.815 201.070 ;
        RECT 117.415 200.380 118.380 200.640 ;
        RECT 118.550 200.415 119.815 200.810 ;
        RECT 119.985 201.240 121.445 201.335 ;
        RECT 119.985 200.870 121.945 201.240 ;
        RECT 122.125 201.150 122.455 201.350 ;
        RECT 122.675 201.200 123.720 201.370 ;
        RECT 123.995 202.205 124.165 202.935 ;
        RECT 125.225 202.935 126.495 202.945 ;
        RECT 125.225 202.885 126.060 202.935 ;
        RECT 124.335 202.540 126.545 202.710 ;
        RECT 124.335 202.375 125.305 202.540 ;
        RECT 125.975 202.455 126.545 202.540 ;
        RECT 126.715 202.575 126.885 203.365 ;
        RECT 127.875 203.345 128.125 203.695 ;
        RECT 128.295 203.685 128.465 203.865 ;
        RECT 129.435 203.910 130.405 204.170 ;
        RECT 128.295 203.355 129.250 203.685 ;
        RECT 129.435 203.310 129.610 203.910 ;
        RECT 129.780 203.480 130.745 203.740 ;
        RECT 127.055 202.745 127.705 203.075 ;
        RECT 125.475 202.285 125.805 202.370 ;
        RECT 126.715 202.285 127.345 202.575 ;
        RECT 123.995 202.035 125.305 202.205 ;
        RECT 125.475 202.115 126.145 202.285 ;
        RECT 119.985 200.585 121.445 200.870 ;
        RECT 122.125 200.690 122.425 201.150 ;
        RECT 122.675 201.030 122.935 201.200 ;
        RECT 123.995 201.030 124.165 202.035 ;
        RECT 125.475 201.865 125.805 201.890 ;
        RECT 122.605 200.860 122.935 201.030 ;
        RECT 123.195 200.860 124.165 201.030 ;
        RECT 117.415 199.780 117.655 200.380 ;
        RECT 118.550 200.210 120.335 200.415 ;
        RECT 117.825 199.950 120.335 200.210 ;
        RECT 117.415 199.520 118.380 199.780 ;
        RECT 118.550 199.665 120.335 199.950 ;
        RECT 120.505 199.665 121.445 200.585 ;
        RECT 121.725 200.520 123.825 200.690 ;
        RECT 121.725 200.285 121.895 200.520 ;
        RECT 123.495 200.440 123.825 200.520 ;
        RECT 122.605 200.160 123.325 200.350 ;
        RECT 117.415 198.935 117.655 199.520 ;
        RECT 118.550 199.350 118.725 199.665 ;
        RECT 117.825 199.105 118.725 199.350 ;
        RECT 118.895 199.235 119.565 199.405 ;
        RECT 118.550 199.065 118.725 199.105 ;
        RECT 117.415 198.675 118.380 198.935 ;
        RECT 118.550 198.735 119.225 199.065 ;
        RECT 119.395 198.970 119.565 199.235 ;
        RECT 119.735 199.140 120.385 199.490 ;
        RECT 120.555 199.235 121.015 199.405 ;
        RECT 120.555 198.970 120.725 199.235 ;
        RECT 121.275 199.065 121.445 199.665 ;
        RECT 121.725 199.500 121.895 200.115 ;
        RECT 122.065 199.990 122.395 200.135 ;
        RECT 122.065 199.670 123.355 199.990 ;
        RECT 123.525 199.500 123.695 200.215 ;
        RECT 121.725 199.330 123.695 199.500 ;
        RECT 123.995 199.665 124.165 200.860 ;
        RECT 124.335 201.695 125.805 201.865 ;
        RECT 124.335 200.005 124.505 201.695 ;
        RECT 125.975 201.530 126.145 202.115 ;
        RECT 126.315 202.245 127.345 202.285 ;
        RECT 126.315 201.955 126.885 202.245 ;
        RECT 127.535 202.030 127.705 202.745 ;
        RECT 127.875 202.605 128.125 203.115 ;
        RECT 129.435 203.055 130.335 203.310 ;
        RECT 128.315 203.050 130.335 203.055 ;
        RECT 128.315 202.725 129.610 203.050 ;
        RECT 130.505 202.880 130.745 203.480 ;
        RECT 129.435 202.450 129.610 202.725 ;
        RECT 129.780 202.620 130.745 202.880 ;
        RECT 125.975 201.525 126.545 201.530 ;
        RECT 124.675 201.355 126.545 201.525 ;
        RECT 124.675 200.400 124.845 201.355 ;
        RECT 125.015 201.015 125.985 201.185 ;
        RECT 125.015 200.365 125.185 201.015 ;
        RECT 126.180 201.000 126.545 201.355 ;
        RECT 126.715 201.500 126.885 201.955 ;
        RECT 127.055 201.700 127.705 202.030 ;
        RECT 127.875 202.025 129.190 202.395 ;
        RECT 129.435 202.190 130.335 202.450 ;
        RECT 126.715 201.170 127.345 201.500 ;
        RECT 125.525 200.810 125.695 200.815 ;
        RECT 125.385 200.535 126.545 200.810 ;
        RECT 125.015 200.175 126.545 200.365 ;
        RECT 126.715 200.005 126.885 201.170 ;
        RECT 127.535 200.945 127.705 201.700 ;
        RECT 127.875 201.525 129.190 201.855 ;
        RECT 129.435 201.590 129.610 202.190 ;
        RECT 130.505 202.020 130.745 202.620 ;
        RECT 129.780 201.760 130.745 202.020 ;
        RECT 129.435 201.330 130.335 201.590 ;
        RECT 127.875 200.985 129.190 201.315 ;
        RECT 127.215 200.775 127.705 200.945 ;
        RECT 127.070 200.275 127.705 200.605 ;
        RECT 127.875 200.395 128.085 200.815 ;
        RECT 129.435 200.730 129.610 201.330 ;
        RECT 130.505 201.160 130.745 201.760 ;
        RECT 129.780 200.900 130.745 201.160 ;
        RECT 128.255 200.465 129.265 200.715 ;
        RECT 129.435 200.485 130.335 200.730 ;
        RECT 127.515 200.225 127.705 200.275 ;
        RECT 128.255 200.225 128.545 200.465 ;
        RECT 129.435 200.295 129.610 200.485 ;
        RECT 130.505 200.315 130.745 200.900 ;
        RECT 124.335 199.835 125.360 200.005 ;
        RECT 126.715 199.995 127.345 200.005 ;
        RECT 123.995 199.495 124.925 199.665 ;
        RECT 119.395 198.740 120.725 198.970 ;
        RECT 120.895 199.055 121.445 199.065 ;
        RECT 120.895 198.845 121.975 199.055 ;
        RECT 120.895 198.735 121.445 198.845 ;
        RECT 117.415 198.075 117.655 198.675 ;
        RECT 118.550 198.490 118.725 198.735 ;
        RECT 117.825 198.245 118.725 198.490 ;
        RECT 118.895 198.380 121.015 198.565 ;
        RECT 118.550 198.140 118.725 198.245 ;
        RECT 117.415 197.815 118.380 198.075 ;
        RECT 118.550 197.875 119.185 198.140 ;
        RECT 119.695 197.930 120.645 198.210 ;
        RECT 121.275 198.125 121.445 198.735 ;
        RECT 122.355 198.625 122.685 199.330 ;
        RECT 122.890 198.605 123.265 199.160 ;
        RECT 123.995 199.150 124.165 199.495 ;
        RECT 123.495 198.835 124.165 199.150 ;
        RECT 121.660 198.455 122.185 198.585 ;
        RECT 122.890 198.455 123.825 198.605 ;
        RECT 121.660 198.265 123.825 198.455 ;
        RECT 121.660 198.255 122.685 198.265 ;
        RECT 120.815 198.085 121.445 198.125 ;
        RECT 120.815 197.915 122.055 198.085 ;
        RECT 120.815 197.875 121.445 197.915 ;
        RECT 117.415 197.215 117.655 197.815 ;
        RECT 118.550 197.630 118.725 197.875 ;
        RECT 119.320 197.705 120.685 197.760 ;
        RECT 117.825 197.385 118.725 197.630 ;
        RECT 118.895 197.590 120.995 197.705 ;
        RECT 118.895 197.455 119.450 197.590 ;
        RECT 120.555 197.535 120.995 197.590 ;
        RECT 117.415 196.955 118.380 197.215 ;
        RECT 117.415 196.780 117.640 196.955 ;
        RECT 115.835 196.765 116.485 196.775 ;
        RECT 112.615 196.535 114.425 196.685 ;
        RECT 114.595 196.595 115.265 196.765 ;
        RECT 113.115 196.515 114.425 196.535 ;
        RECT 110.780 196.155 111.305 196.285 ;
        RECT 112.010 196.155 112.945 196.305 ;
        RECT 110.780 195.965 112.945 196.155 ;
        RECT 110.780 195.955 111.805 195.965 ;
        RECT 110.395 195.615 111.175 195.785 ;
        RECT 110.395 194.890 110.565 195.615 ;
        RECT 110.785 195.290 111.305 195.445 ;
        RECT 111.475 195.405 111.805 195.955 ;
        RECT 113.115 195.795 113.285 196.515 ;
        RECT 114.595 196.345 114.925 196.370 ;
        RECT 112.105 195.625 113.285 195.795 ;
        RECT 110.785 195.235 111.345 195.290 ;
        RECT 111.975 195.280 112.900 195.455 ;
        RECT 111.925 195.235 112.900 195.280 ;
        RECT 110.785 195.125 112.900 195.235 ;
        RECT 110.785 195.115 112.055 195.125 ;
        RECT 111.220 195.065 112.055 195.115 ;
        RECT 113.115 194.890 113.285 195.625 ;
        RECT 110.395 194.630 111.405 194.890 ;
        RECT 111.965 194.630 113.285 194.890 ;
        RECT 110.395 194.030 110.565 194.630 ;
        RECT 110.735 194.285 112.945 194.455 ;
        RECT 110.735 194.200 111.310 194.285 ;
        RECT 112.040 194.200 112.945 194.285 ;
        RECT 113.115 194.145 113.285 194.630 ;
        RECT 113.455 196.175 114.925 196.345 ;
        RECT 113.455 194.485 113.625 196.175 ;
        RECT 115.095 196.010 115.265 196.595 ;
        RECT 115.435 196.515 116.485 196.765 ;
        RECT 115.435 196.435 116.005 196.515 ;
        RECT 115.095 196.005 115.665 196.010 ;
        RECT 113.795 195.835 115.665 196.005 ;
        RECT 113.795 194.880 113.965 195.835 ;
        RECT 114.135 195.495 115.105 195.665 ;
        RECT 114.135 194.845 114.305 195.495 ;
        RECT 115.300 195.480 115.665 195.835 ;
        RECT 115.835 195.915 116.005 196.435 ;
        RECT 116.655 196.345 117.640 196.780 ;
        RECT 118.550 196.770 118.725 197.385 ;
        RECT 117.825 196.515 118.725 196.770 ;
        RECT 116.200 196.085 118.380 196.345 ;
        RECT 116.655 196.055 118.380 196.085 ;
        RECT 115.835 195.615 116.485 195.915 ;
        RECT 116.655 195.615 117.640 196.055 ;
        RECT 118.555 195.970 118.725 196.515 ;
        RECT 119.000 196.310 119.170 197.245 ;
        RECT 119.640 197.180 120.235 197.420 ;
        RECT 120.825 197.370 120.995 197.535 ;
        RECT 120.405 197.010 120.625 197.365 ;
        RECT 121.275 197.185 121.445 197.875 ;
        RECT 121.665 197.590 122.185 197.745 ;
        RECT 122.355 197.705 122.685 198.255 ;
        RECT 123.995 198.095 124.165 198.835 ;
        RECT 124.515 199.085 124.925 199.260 ;
        RECT 125.170 199.255 125.360 199.835 ;
        RECT 125.735 199.265 125.905 199.975 ;
        RECT 126.180 199.835 127.345 199.995 ;
        RECT 127.515 199.965 128.545 200.225 ;
        RECT 128.715 199.965 129.610 200.295 ;
        RECT 129.780 200.055 130.745 200.315 ;
        RECT 127.515 199.855 128.085 199.965 ;
        RECT 126.180 199.485 126.885 199.835 ;
        RECT 127.875 199.645 128.085 199.855 ;
        RECT 129.435 199.870 129.610 199.965 ;
        RECT 125.735 199.085 126.510 199.265 ;
        RECT 124.515 199.020 126.510 199.085 ;
        RECT 124.515 198.745 125.905 199.020 ;
        RECT 124.335 198.295 126.545 198.575 ;
        RECT 124.335 198.190 125.305 198.295 ;
        RECT 125.975 198.190 126.545 198.295 ;
        RECT 126.715 198.480 126.885 199.485 ;
        RECT 127.055 199.475 127.685 199.545 ;
        RECT 128.255 199.475 129.265 199.730 ;
        RECT 127.055 199.205 129.265 199.475 ;
        RECT 129.435 199.625 130.335 199.870 ;
        RECT 127.055 198.755 129.265 199.035 ;
        RECT 127.055 198.650 127.625 198.755 ;
        RECT 128.295 198.650 129.265 198.755 ;
        RECT 129.435 199.010 129.610 199.625 ;
        RECT 130.505 199.455 130.745 200.055 ;
        RECT 129.780 199.195 130.745 199.455 ;
        RECT 129.435 198.765 130.335 199.010 ;
        RECT 127.795 198.480 128.125 198.585 ;
        RECT 129.435 198.480 129.610 198.765 ;
        RECT 130.505 198.595 130.745 199.195 ;
        RECT 126.715 198.155 127.345 198.480 ;
        RECT 122.985 198.020 124.165 198.095 ;
        RECT 125.475 198.020 125.805 198.125 ;
        RECT 126.715 198.020 126.885 198.155 ;
        RECT 122.985 197.925 124.625 198.020 ;
        RECT 121.665 197.535 122.225 197.590 ;
        RECT 122.855 197.580 123.780 197.755 ;
        RECT 122.805 197.535 123.780 197.580 ;
        RECT 121.665 197.425 123.780 197.535 ;
        RECT 123.995 197.695 124.625 197.925 ;
        RECT 121.665 197.415 122.935 197.425 ;
        RECT 122.100 197.365 122.935 197.415 ;
        RECT 119.340 196.840 120.625 197.010 ;
        RECT 119.340 196.480 119.705 196.840 ;
        RECT 120.825 196.670 120.995 197.175 ;
        RECT 119.875 196.500 120.995 196.670 ;
        RECT 121.275 196.855 121.950 197.185 ;
        RECT 122.805 197.130 122.975 197.135 ;
        RECT 119.875 196.310 120.045 196.500 ;
        RECT 119.000 196.140 120.045 196.310 ;
        RECT 119.785 195.970 120.045 196.140 ;
        RECT 120.265 196.090 120.595 196.290 ;
        RECT 121.275 196.180 121.445 196.855 ;
        RECT 122.125 196.830 122.975 197.130 ;
        RECT 123.145 196.935 123.805 197.105 ;
        RECT 121.640 196.660 122.015 196.685 ;
        RECT 123.145 196.660 123.375 196.935 ;
        RECT 123.995 196.765 124.165 197.695 ;
        RECT 124.795 197.570 126.085 198.020 ;
        RECT 126.255 197.695 126.885 198.020 ;
        RECT 124.795 197.175 125.015 197.570 ;
        RECT 124.335 196.895 125.015 197.175 ;
        RECT 121.640 196.445 123.375 196.660 ;
        RECT 118.555 195.885 119.525 195.970 ;
        RECT 117.810 195.800 119.525 195.885 ;
        RECT 119.785 195.800 120.115 195.970 ;
        RECT 117.810 195.615 118.725 195.800 ;
        RECT 120.295 195.630 120.595 196.090 ;
        RECT 120.775 195.810 121.445 196.180 ;
        RECT 122.165 196.425 123.375 196.445 ;
        RECT 123.545 196.435 124.165 196.765 ;
        RECT 125.185 196.705 125.745 197.400 ;
        RECT 125.915 197.175 126.085 197.570 ;
        RECT 125.915 196.895 126.545 197.175 ;
        RECT 121.630 195.995 121.970 196.165 ;
        RECT 122.165 196.105 122.495 196.425 ;
        RECT 115.835 195.355 116.005 195.615 ;
        RECT 118.555 195.355 118.725 195.615 ;
        RECT 118.895 195.460 120.995 195.630 ;
        RECT 118.895 195.380 119.225 195.460 ;
        RECT 114.645 195.290 114.815 195.295 ;
        RECT 114.505 195.015 115.665 195.290 ;
        RECT 114.135 194.655 115.665 194.845 ;
        RECT 115.835 194.835 117.295 195.355 ;
        RECT 113.455 194.315 114.480 194.485 ;
        RECT 115.835 194.475 116.755 194.835 ;
        RECT 117.465 194.665 118.725 195.355 ;
        RECT 111.475 194.030 111.805 194.115 ;
        RECT 113.115 194.030 114.045 194.145 ;
        RECT 110.395 193.700 110.945 194.030 ;
        RECT 111.115 193.860 112.185 194.030 ;
        RECT 110.395 192.135 110.565 193.700 ;
        RECT 111.115 193.485 111.285 193.860 ;
        RECT 110.735 193.315 111.285 193.485 ;
        RECT 111.465 193.225 111.835 193.580 ;
        RECT 112.015 193.485 112.185 193.860 ;
        RECT 112.355 193.975 114.045 194.030 ;
        RECT 112.355 193.700 113.285 193.975 ;
        RECT 112.015 193.315 112.945 193.485 ;
        RECT 113.115 192.135 113.285 193.700 ;
        RECT 113.635 193.565 114.045 193.740 ;
        RECT 114.290 193.735 114.480 194.315 ;
        RECT 114.855 193.745 115.025 194.455 ;
        RECT 115.300 194.145 116.755 194.475 ;
        RECT 116.925 194.145 118.725 194.665 ;
        RECT 119.025 194.440 119.195 195.155 ;
        RECT 119.395 195.100 120.115 195.290 ;
        RECT 120.825 195.225 120.995 195.460 ;
        RECT 121.275 195.405 121.445 195.810 ;
        RECT 121.775 195.935 121.970 195.995 ;
        RECT 122.665 195.950 123.780 196.235 ;
        RECT 122.665 195.935 122.835 195.950 ;
        RECT 121.775 195.765 122.835 195.935 ;
        RECT 123.995 195.905 124.165 196.435 ;
        RECT 124.335 196.305 126.545 196.705 ;
        RECT 126.715 196.365 126.885 197.695 ;
        RECT 127.515 198.030 128.805 198.480 ;
        RECT 128.975 198.155 129.610 198.480 ;
        RECT 129.780 198.335 130.745 198.595 ;
        RECT 127.515 197.635 127.685 198.030 ;
        RECT 127.055 197.355 127.685 197.635 ;
        RECT 127.855 197.165 128.415 197.860 ;
        RECT 128.585 197.635 128.805 198.030 ;
        RECT 129.435 198.150 129.610 198.155 ;
        RECT 130.520 198.160 130.745 198.335 ;
        RECT 130.915 198.330 131.165 204.340 ;
        RECT 132.155 204.170 132.325 204.725 ;
        RECT 132.585 204.295 133.045 204.465 ;
        RECT 131.595 204.125 132.325 204.170 ;
        RECT 131.595 203.910 132.705 204.125 ;
        RECT 132.155 203.795 132.705 203.910 ;
        RECT 132.875 204.030 133.045 204.295 ;
        RECT 133.215 204.200 133.865 204.550 ;
        RECT 134.875 204.470 135.775 204.725 ;
        RECT 134.035 204.295 134.705 204.465 ;
        RECT 134.035 204.030 134.205 204.295 ;
        RECT 134.875 204.125 135.050 204.470 ;
        RECT 135.945 204.300 136.185 204.900 ;
        RECT 132.875 203.800 134.205 204.030 ;
        RECT 134.375 203.870 135.050 204.125 ;
        RECT 135.220 204.040 136.185 204.300 ;
        RECT 134.375 203.795 135.775 203.870 ;
        RECT 131.335 203.480 131.960 203.740 ;
        RECT 131.335 202.880 131.505 203.480 ;
        RECT 132.155 203.310 132.325 203.795 ;
        RECT 132.585 203.440 134.705 203.625 ;
        RECT 134.875 203.610 135.775 203.795 ;
        RECT 131.675 203.185 132.325 203.310 ;
        RECT 131.675 203.050 132.785 203.185 ;
        RECT 132.155 202.935 132.785 203.050 ;
        RECT 132.955 202.990 133.905 203.270 ;
        RECT 134.875 203.200 135.050 203.610 ;
        RECT 135.945 203.440 136.185 204.040 ;
        RECT 134.415 203.010 135.050 203.200 ;
        RECT 135.220 203.180 136.185 203.440 ;
        RECT 134.415 202.935 135.775 203.010 ;
        RECT 131.335 202.620 131.960 202.880 ;
        RECT 131.335 202.020 131.505 202.620 ;
        RECT 132.155 202.450 132.325 202.935 ;
        RECT 132.915 202.765 134.280 202.820 ;
        RECT 131.675 202.190 132.325 202.450 ;
        RECT 132.605 202.650 134.705 202.765 ;
        RECT 132.605 202.595 133.045 202.650 ;
        RECT 132.605 202.430 132.775 202.595 ;
        RECT 134.150 202.515 134.705 202.650 ;
        RECT 134.875 202.750 135.775 202.935 ;
        RECT 131.335 201.760 131.960 202.020 ;
        RECT 131.335 201.175 131.505 201.760 ;
        RECT 132.155 201.590 132.325 202.190 ;
        RECT 131.675 201.345 132.325 201.590 ;
        RECT 132.605 201.730 132.775 202.235 ;
        RECT 132.975 202.070 133.195 202.425 ;
        RECT 133.365 202.240 133.960 202.480 ;
        RECT 132.975 201.900 134.260 202.070 ;
        RECT 132.605 201.560 133.725 201.730 ;
        RECT 133.555 201.370 133.725 201.560 ;
        RECT 133.895 201.540 134.260 201.900 ;
        RECT 134.430 201.370 134.600 202.305 ;
        RECT 132.155 201.240 132.325 201.345 ;
        RECT 131.335 200.900 131.960 201.175 ;
        RECT 131.335 200.315 131.505 200.900 ;
        RECT 132.155 200.870 132.825 201.240 ;
        RECT 133.005 201.150 133.335 201.350 ;
        RECT 133.555 201.200 134.600 201.370 ;
        RECT 134.875 202.150 135.050 202.750 ;
        RECT 135.945 202.580 136.185 203.180 ;
        RECT 135.220 202.320 136.185 202.580 ;
        RECT 134.875 201.890 135.845 202.150 ;
        RECT 134.875 201.290 135.045 201.890 ;
        RECT 136.355 201.720 136.605 207.730 ;
        RECT 136.775 207.725 136.945 207.900 ;
        RECT 136.775 207.465 137.400 207.725 ;
        RECT 136.775 206.865 136.945 207.465 ;
        RECT 137.595 207.295 137.765 207.905 ;
        RECT 138.395 208.150 139.685 208.600 ;
        RECT 139.855 208.275 140.485 208.600 ;
        RECT 141.545 208.540 141.805 208.710 ;
        RECT 142.055 208.590 142.355 209.050 ;
        RECT 143.035 208.870 143.205 209.270 ;
        RECT 144.115 209.185 144.445 209.270 ;
        RECT 138.395 207.755 138.565 208.150 ;
        RECT 137.935 207.475 138.565 207.755 ;
        RECT 137.115 207.045 137.765 207.295 ;
        RECT 138.735 207.285 139.295 207.980 ;
        RECT 139.465 207.755 139.685 208.150 ;
        RECT 139.465 207.475 140.145 207.755 ;
        RECT 136.775 206.605 137.400 206.865 ;
        RECT 136.775 206.005 136.945 206.605 ;
        RECT 137.595 206.485 137.765 207.045 ;
        RECT 137.935 206.885 140.145 207.285 ;
        RECT 140.315 206.805 140.485 208.275 ;
        RECT 140.760 208.370 141.805 208.540 ;
        RECT 142.025 208.390 142.355 208.590 ;
        RECT 142.535 208.670 143.205 208.870 ;
        RECT 143.375 209.015 143.950 209.100 ;
        RECT 144.680 209.015 145.585 209.100 ;
        RECT 143.375 208.845 145.585 209.015 ;
        RECT 145.755 208.670 145.925 209.270 ;
        RECT 142.535 208.500 144.045 208.670 ;
        RECT 143.035 208.410 144.045 208.500 ;
        RECT 144.605 208.410 145.925 208.670 ;
        RECT 140.760 207.435 140.930 208.370 ;
        RECT 141.100 207.840 141.465 208.200 ;
        RECT 141.635 208.180 141.805 208.370 ;
        RECT 141.635 208.010 142.755 208.180 ;
        RECT 141.100 207.670 142.385 207.840 ;
        RECT 141.400 207.260 141.995 207.500 ;
        RECT 142.165 207.315 142.385 207.670 ;
        RECT 142.585 207.505 142.755 208.010 ;
        RECT 140.655 207.090 141.210 207.225 ;
        RECT 142.585 207.145 142.755 207.310 ;
        RECT 142.315 207.090 142.755 207.145 ;
        RECT 140.655 206.975 142.755 207.090 ;
        RECT 143.035 207.175 143.205 208.410 ;
        RECT 143.375 208.065 144.785 208.235 ;
        RECT 145.755 208.225 145.925 208.410 ;
        RECT 143.375 207.745 143.945 208.065 ;
        RECT 143.375 207.345 143.945 207.575 ;
        RECT 144.115 207.490 144.445 207.895 ;
        RECT 144.615 207.715 144.785 208.065 ;
        RECT 144.955 207.895 145.925 208.225 ;
        RECT 144.615 207.465 145.585 207.715 ;
        RECT 141.080 206.920 142.445 206.975 ;
        RECT 143.035 206.805 143.605 207.175 ;
        RECT 138.395 206.505 139.685 206.715 ;
        RECT 137.595 206.435 138.225 206.485 ;
        RECT 137.115 206.215 138.225 206.435 ;
        RECT 137.115 206.185 137.765 206.215 ;
        RECT 136.775 205.745 137.400 206.005 ;
        RECT 136.775 205.160 136.945 205.745 ;
        RECT 137.595 205.575 137.765 206.185 ;
        RECT 138.395 206.045 138.565 206.505 ;
        RECT 137.935 205.760 138.565 206.045 ;
        RECT 138.735 205.645 139.295 206.335 ;
        RECT 139.465 206.045 139.685 206.505 ;
        RECT 140.315 206.540 140.945 206.805 ;
        RECT 142.575 206.755 143.605 206.805 ;
        RECT 140.315 206.485 140.485 206.540 ;
        RECT 139.855 206.215 140.485 206.485 ;
        RECT 141.455 206.470 142.405 206.750 ;
        RECT 142.575 206.555 143.205 206.755 ;
        RECT 143.775 206.585 143.945 207.345 ;
        RECT 144.115 207.025 145.245 207.275 ;
        RECT 139.465 205.760 140.145 206.045 ;
        RECT 140.315 205.945 140.485 206.215 ;
        RECT 140.655 206.115 142.775 206.300 ;
        RECT 143.035 206.245 143.205 206.555 ;
        RECT 143.375 206.415 143.945 206.585 ;
        RECT 144.115 206.625 145.245 206.825 ;
        RECT 144.115 206.580 144.445 206.625 ;
        RECT 145.415 206.455 145.585 207.465 ;
        RECT 143.035 205.945 143.945 206.245 ;
        RECT 144.115 206.005 144.395 206.395 ;
        RECT 144.565 206.285 145.585 206.455 ;
        RECT 137.115 205.330 137.765 205.575 ;
        RECT 136.775 204.885 137.400 205.160 ;
        RECT 137.595 205.015 137.765 205.330 ;
        RECT 140.315 205.615 140.985 205.945 ;
        RECT 141.155 205.710 142.485 205.940 ;
        RECT 140.315 205.015 140.485 205.615 ;
        RECT 141.155 205.445 141.325 205.710 ;
        RECT 140.655 205.275 141.325 205.445 ;
        RECT 141.495 205.190 142.145 205.540 ;
        RECT 142.315 205.445 142.485 205.710 ;
        RECT 142.655 205.795 143.945 205.945 ;
        RECT 144.565 205.835 144.735 206.285 ;
        RECT 145.755 206.115 145.925 207.895 ;
        RECT 142.655 205.615 143.205 205.795 ;
        RECT 144.115 205.665 144.735 205.835 ;
        RECT 144.905 205.800 145.925 206.115 ;
        RECT 142.315 205.275 142.775 205.445 ;
        RECT 136.775 204.300 136.945 204.885 ;
        RECT 137.595 204.725 138.490 205.015 ;
        RECT 139.150 204.725 140.485 205.015 ;
        RECT 143.035 205.015 143.205 205.615 ;
        RECT 143.385 205.495 143.945 205.625 ;
        RECT 144.955 205.495 145.585 205.625 ;
        RECT 143.385 205.185 145.585 205.495 ;
        RECT 145.755 205.015 145.925 205.800 ;
        RECT 140.655 204.755 141.325 204.925 ;
        RECT 137.595 204.715 137.765 204.725 ;
        RECT 137.115 204.470 137.765 204.715 ;
        RECT 140.315 204.585 140.485 204.725 ;
        RECT 136.775 204.040 137.400 204.300 ;
        RECT 137.595 204.125 137.765 204.470 ;
        RECT 137.935 204.380 140.145 204.550 ;
        RECT 137.935 204.295 138.505 204.380 ;
        RECT 139.175 204.215 140.145 204.380 ;
        RECT 140.315 204.255 140.985 204.585 ;
        RECT 141.155 204.490 141.325 204.755 ;
        RECT 141.495 204.660 142.145 205.010 ;
        RECT 142.315 204.755 142.775 204.925 ;
        RECT 142.315 204.490 142.485 204.755 ;
        RECT 143.035 204.725 143.930 205.015 ;
        RECT 144.590 204.725 145.925 205.015 ;
        RECT 143.035 204.585 143.205 204.725 ;
        RECT 141.155 204.260 142.485 204.490 ;
        RECT 142.655 204.255 143.205 204.585 ;
        RECT 138.675 204.125 139.005 204.210 ;
        RECT 136.775 203.440 136.945 204.040 ;
        RECT 137.595 203.870 138.165 204.125 ;
        RECT 137.115 203.795 138.165 203.870 ;
        RECT 138.335 203.955 139.005 204.125 ;
        RECT 140.315 204.045 140.485 204.255 ;
        RECT 137.115 203.610 137.765 203.795 ;
        RECT 136.775 203.180 137.400 203.440 ;
        RECT 136.775 202.580 136.945 203.180 ;
        RECT 137.595 203.010 137.765 203.610 ;
        RECT 138.335 203.370 138.505 203.955 ;
        RECT 139.175 203.875 140.485 204.045 ;
        RECT 140.655 203.900 142.775 204.085 ;
        RECT 138.675 203.705 139.005 203.730 ;
        RECT 138.675 203.535 140.145 203.705 ;
        RECT 137.115 202.750 137.765 203.010 ;
        RECT 137.935 203.365 138.505 203.370 ;
        RECT 137.935 203.195 139.805 203.365 ;
        RECT 137.935 202.840 138.300 203.195 ;
        RECT 138.495 202.855 139.465 203.025 ;
        RECT 136.775 202.320 137.400 202.580 ;
        RECT 137.595 202.150 137.765 202.750 ;
        RECT 138.785 202.650 138.955 202.655 ;
        RECT 137.935 202.375 139.095 202.650 ;
        RECT 139.295 202.205 139.465 202.855 ;
        RECT 139.635 202.240 139.805 203.195 ;
        RECT 137.035 201.890 137.765 202.150 ;
        RECT 137.935 202.015 139.465 202.205 ;
        RECT 137.595 201.835 137.765 201.890 ;
        RECT 139.975 201.845 140.145 203.535 ;
        RECT 135.220 201.470 137.415 201.720 ;
        RECT 132.155 200.730 132.325 200.870 ;
        RECT 131.675 200.485 132.325 200.730 ;
        RECT 133.005 200.690 133.305 201.150 ;
        RECT 133.555 201.030 133.815 201.200 ;
        RECT 134.875 201.030 135.855 201.290 ;
        RECT 133.485 200.860 133.815 201.030 ;
        RECT 134.075 200.860 135.045 201.030 ;
        RECT 131.335 200.055 131.960 200.315 ;
        RECT 131.335 199.455 131.505 200.055 ;
        RECT 132.155 199.875 132.325 200.485 ;
        RECT 132.605 200.520 134.705 200.690 ;
        RECT 132.605 200.285 132.775 200.520 ;
        RECT 134.375 200.440 134.705 200.520 ;
        RECT 134.875 200.430 135.045 200.860 ;
        RECT 136.355 200.860 136.605 201.470 ;
        RECT 137.595 201.325 138.300 201.835 ;
        RECT 137.595 201.290 137.765 201.325 ;
        RECT 137.070 201.030 137.765 201.290 ;
        RECT 138.575 201.105 138.745 201.815 ;
        RECT 136.355 200.855 137.415 200.860 ;
        RECT 135.215 200.610 137.415 200.855 ;
        RECT 133.485 200.160 134.205 200.350 ;
        RECT 131.675 199.625 132.325 199.875 ;
        RECT 131.335 199.195 131.960 199.455 ;
        RECT 131.335 198.595 131.505 199.195 ;
        RECT 132.155 199.055 132.325 199.625 ;
        RECT 132.605 199.500 132.775 200.115 ;
        RECT 132.945 199.990 133.275 200.135 ;
        RECT 132.945 199.670 134.235 199.990 ;
        RECT 134.405 199.500 134.575 200.215 ;
        RECT 132.605 199.330 134.575 199.500 ;
        RECT 134.875 200.135 135.855 200.430 ;
        RECT 134.875 199.400 135.045 200.135 ;
        RECT 136.355 200.125 136.915 200.440 ;
        RECT 137.595 200.430 137.765 201.030 ;
        RECT 137.970 200.925 138.745 201.105 ;
        RECT 139.120 201.675 140.145 201.845 ;
        RECT 140.315 203.660 140.485 203.875 ;
        RECT 140.315 203.395 140.945 203.660 ;
        RECT 141.455 203.450 142.405 203.730 ;
        RECT 143.035 203.645 143.205 204.255 ;
        RECT 142.575 203.395 143.205 203.645 ;
        RECT 139.120 201.095 139.310 201.675 ;
        RECT 140.315 201.505 140.485 203.395 ;
        RECT 141.080 203.225 142.445 203.280 ;
        RECT 140.655 203.110 142.755 203.225 ;
        RECT 140.655 202.975 141.210 203.110 ;
        RECT 142.315 203.055 142.755 203.110 ;
        RECT 140.760 201.830 140.930 202.765 ;
        RECT 141.400 202.700 141.995 202.940 ;
        RECT 142.585 202.890 142.755 203.055 ;
        RECT 143.035 203.065 143.205 203.395 ;
        RECT 143.375 203.235 144.005 203.520 ;
        RECT 142.165 202.530 142.385 202.885 ;
        RECT 143.035 202.795 143.665 203.065 ;
        RECT 141.100 202.360 142.385 202.530 ;
        RECT 141.100 202.000 141.465 202.360 ;
        RECT 142.585 202.190 142.755 202.695 ;
        RECT 141.635 202.020 142.755 202.190 ;
        RECT 141.635 201.830 141.805 202.020 ;
        RECT 140.760 201.660 141.805 201.830 ;
        RECT 139.555 201.490 140.485 201.505 ;
        RECT 141.545 201.490 141.805 201.660 ;
        RECT 142.025 201.610 142.355 201.810 ;
        RECT 143.035 201.700 143.205 202.795 ;
        RECT 143.835 202.775 144.005 203.235 ;
        RECT 144.175 202.945 144.735 203.635 ;
        RECT 144.905 203.235 145.585 203.520 ;
        RECT 144.905 202.775 145.125 203.235 ;
        RECT 145.755 203.065 145.925 204.725 ;
        RECT 145.295 202.795 145.925 203.065 ;
        RECT 143.835 202.565 145.125 202.775 ;
        RECT 143.375 201.995 145.585 202.395 ;
        RECT 139.555 201.335 141.285 201.490 ;
        RECT 140.315 201.320 141.285 201.335 ;
        RECT 141.545 201.320 141.875 201.490 ;
        RECT 139.555 200.925 139.965 201.100 ;
        RECT 137.970 200.860 139.965 200.925 ;
        RECT 138.575 200.585 139.965 200.860 ;
        RECT 137.085 200.125 137.765 200.430 ;
        RECT 135.215 199.675 137.425 199.955 ;
        RECT 135.215 199.570 136.185 199.675 ;
        RECT 136.855 199.570 137.425 199.675 ;
        RECT 137.595 199.790 137.765 200.125 ;
        RECT 137.595 199.550 138.275 199.790 ;
        RECT 136.355 199.400 136.685 199.505 ;
        RECT 137.595 199.400 137.765 199.550 ;
        RECT 138.445 199.540 139.005 199.895 ;
        RECT 132.155 199.015 132.855 199.055 ;
        RECT 131.675 198.845 132.855 199.015 ;
        RECT 131.675 198.765 132.325 198.845 ;
        RECT 131.335 198.335 131.960 198.595 ;
        RECT 131.335 198.160 131.505 198.335 ;
        RECT 129.435 197.895 130.335 198.150 ;
        RECT 128.585 197.355 129.265 197.635 ;
        RECT 129.435 197.265 129.605 197.895 ;
        RECT 130.520 197.725 131.505 198.160 ;
        RECT 132.155 198.155 132.325 198.765 ;
        RECT 133.235 198.625 133.565 199.330 ;
        RECT 133.770 198.605 134.145 199.160 ;
        RECT 134.875 199.150 135.505 199.400 ;
        RECT 134.375 199.075 135.505 199.150 ;
        RECT 134.375 198.835 135.045 199.075 ;
        RECT 132.540 198.455 133.065 198.585 ;
        RECT 133.770 198.455 134.705 198.605 ;
        RECT 132.540 198.265 134.705 198.455 ;
        RECT 132.540 198.255 133.565 198.265 ;
        RECT 131.675 198.085 132.325 198.155 ;
        RECT 131.675 197.915 132.935 198.085 ;
        RECT 131.675 197.895 132.325 197.915 ;
        RECT 129.780 197.465 131.960 197.725 ;
        RECT 129.780 197.435 131.505 197.465 ;
        RECT 127.055 196.765 129.265 197.165 ;
        RECT 129.435 196.995 130.350 197.265 ;
        RECT 130.520 196.995 131.505 197.435 ;
        RECT 132.155 197.295 132.325 197.895 ;
        RECT 132.545 197.590 133.065 197.745 ;
        RECT 133.235 197.705 133.565 198.255 ;
        RECT 134.875 198.095 135.045 198.835 ;
        RECT 135.675 198.950 136.965 199.400 ;
        RECT 137.135 199.075 137.765 199.400 ;
        RECT 139.175 199.380 139.520 199.770 ;
        RECT 140.315 199.610 140.485 201.320 ;
        RECT 142.055 201.150 142.355 201.610 ;
        RECT 142.535 201.330 143.205 201.700 ;
        RECT 143.375 201.525 144.005 201.805 ;
        RECT 140.655 200.980 142.755 201.150 ;
        RECT 140.655 200.900 140.985 200.980 ;
        RECT 140.785 199.960 140.955 200.675 ;
        RECT 141.155 200.620 141.875 200.810 ;
        RECT 142.585 200.745 142.755 200.980 ;
        RECT 143.035 201.005 143.205 201.330 ;
        RECT 143.835 201.130 144.005 201.525 ;
        RECT 144.175 201.300 144.735 201.995 ;
        RECT 144.905 201.525 145.585 201.805 ;
        RECT 144.905 201.130 145.125 201.525 ;
        RECT 143.035 200.680 143.665 201.005 ;
        RECT 143.835 200.680 145.125 201.130 ;
        RECT 145.755 201.005 145.925 202.795 ;
        RECT 145.295 200.680 145.925 201.005 ;
        RECT 142.085 200.450 142.415 200.595 ;
        RECT 141.125 200.130 142.415 200.450 ;
        RECT 142.585 199.960 142.755 200.575 ;
        RECT 140.785 199.790 142.755 199.960 ;
        RECT 139.175 199.370 139.345 199.380 ;
        RECT 137.945 199.200 139.345 199.370 ;
        RECT 137.945 199.090 138.275 199.200 ;
        RECT 135.675 198.555 135.895 198.950 ;
        RECT 135.215 198.275 135.895 198.555 ;
        RECT 133.865 197.925 135.045 198.095 ;
        RECT 136.065 198.085 136.625 198.780 ;
        RECT 136.795 198.555 136.965 198.950 ;
        RECT 137.595 198.860 137.765 199.075 ;
        RECT 137.595 198.645 138.275 198.860 ;
        RECT 138.445 198.765 139.005 199.030 ;
        RECT 136.795 198.275 137.425 198.555 ;
        RECT 132.545 197.535 133.105 197.590 ;
        RECT 133.735 197.580 134.660 197.755 ;
        RECT 133.685 197.535 134.660 197.580 ;
        RECT 132.545 197.425 134.660 197.535 ;
        RECT 132.545 197.415 133.815 197.425 ;
        RECT 132.980 197.365 133.815 197.415 ;
        RECT 131.675 196.995 132.325 197.295 ;
        RECT 127.515 196.385 128.805 196.595 ;
        RECT 124.795 195.925 126.085 196.135 ;
        RECT 120.325 194.930 120.655 195.075 ;
        RECT 119.365 194.610 120.655 194.930 ;
        RECT 120.825 194.440 120.995 195.055 ;
        RECT 119.025 194.270 120.995 194.440 ;
        RECT 121.275 195.005 121.940 195.405 ;
        RECT 122.305 195.375 122.835 195.765 ;
        RECT 121.275 194.415 121.445 195.005 ;
        RECT 122.305 194.945 122.685 195.375 ;
        RECT 123.005 195.080 123.315 195.775 ;
        RECT 123.995 195.770 124.625 195.905 ;
        RECT 123.525 195.635 124.625 195.770 ;
        RECT 123.525 195.085 124.165 195.635 ;
        RECT 124.795 195.465 125.015 195.925 ;
        RECT 124.335 195.180 125.015 195.465 ;
        RECT 121.615 194.775 122.135 194.835 ;
        RECT 122.940 194.775 123.725 194.905 ;
        RECT 121.615 194.600 123.725 194.775 ;
        RECT 123.995 194.895 124.165 195.085 ;
        RECT 125.185 195.065 125.745 195.755 ;
        RECT 125.915 195.465 126.085 195.925 ;
        RECT 126.715 196.095 127.345 196.365 ;
        RECT 126.715 195.905 126.885 196.095 ;
        RECT 127.515 195.925 127.685 196.385 ;
        RECT 126.255 195.635 126.885 195.905 ;
        RECT 127.055 195.640 127.685 195.925 ;
        RECT 125.915 195.180 126.545 195.465 ;
        RECT 126.715 195.355 126.885 195.635 ;
        RECT 127.855 195.525 128.415 196.215 ;
        RECT 128.585 195.925 128.805 196.385 ;
        RECT 129.435 196.365 129.605 196.995 ;
        RECT 132.155 196.735 132.325 196.995 ;
        RECT 134.875 197.285 135.045 197.925 ;
        RECT 135.215 197.685 137.425 198.085 ;
        RECT 137.595 197.595 137.765 198.645 ;
        RECT 139.175 198.515 139.345 199.200 ;
        RECT 140.315 199.295 140.985 199.610 ;
        RECT 140.315 198.895 140.485 199.295 ;
        RECT 141.215 199.065 141.590 199.620 ;
        RECT 141.795 199.085 142.125 199.790 ;
        RECT 143.035 199.515 143.205 200.680 ;
        RECT 144.115 200.575 144.445 200.680 ;
        RECT 143.375 200.405 143.945 200.510 ;
        RECT 144.615 200.405 145.585 200.510 ;
        RECT 143.375 200.125 145.585 200.405 ;
        RECT 142.505 199.305 143.205 199.515 ;
        RECT 139.515 198.565 140.485 198.895 ;
        RECT 140.655 198.915 141.590 199.065 ;
        RECT 142.295 198.915 142.820 199.045 ;
        RECT 140.655 198.725 142.820 198.915 ;
        RECT 137.935 198.175 138.505 198.475 ;
        RECT 138.675 198.345 139.345 198.515 ;
        RECT 140.315 198.555 140.485 198.565 ;
        RECT 141.795 198.715 142.820 198.725 ;
        RECT 143.035 199.030 143.205 199.305 ;
        RECT 145.755 199.030 145.925 200.680 ;
        RECT 143.035 198.770 144.045 199.030 ;
        RECT 144.605 198.770 145.925 199.030 ;
        RECT 139.525 198.175 140.145 198.395 ;
        RECT 137.935 197.860 140.145 198.175 ;
        RECT 140.315 198.385 141.495 198.555 ;
        RECT 140.315 197.595 140.485 198.385 ;
        RECT 140.700 198.040 141.625 198.215 ;
        RECT 141.795 198.165 142.125 198.715 ;
        RECT 143.035 198.545 143.205 198.770 ;
        RECT 142.425 198.375 143.205 198.545 ;
        RECT 142.295 198.050 142.815 198.205 ;
        RECT 140.700 197.995 141.675 198.040 ;
        RECT 142.255 197.995 142.815 198.050 ;
        RECT 140.700 197.885 142.815 197.995 ;
        RECT 141.545 197.875 142.815 197.885 ;
        RECT 143.035 198.170 143.205 198.375 ;
        RECT 143.375 198.425 145.585 198.595 ;
        RECT 143.375 198.340 143.950 198.425 ;
        RECT 144.680 198.340 145.585 198.425 ;
        RECT 144.115 198.170 144.445 198.255 ;
        RECT 145.755 198.170 145.925 198.770 ;
        RECT 141.545 197.825 142.380 197.875 ;
        RECT 143.035 197.840 143.585 198.170 ;
        RECT 143.755 198.000 144.825 198.170 ;
        RECT 135.675 197.305 136.965 197.515 ;
        RECT 134.875 197.015 135.505 197.285 ;
        RECT 134.875 196.735 135.045 197.015 ;
        RECT 135.675 196.845 135.895 197.305 ;
        RECT 128.975 196.180 129.605 196.365 ;
        RECT 129.775 196.455 131.985 196.735 ;
        RECT 129.775 196.350 130.745 196.455 ;
        RECT 131.415 196.350 131.985 196.455 ;
        RECT 132.155 196.465 132.960 196.735 ;
        RECT 133.920 196.465 135.045 196.735 ;
        RECT 135.215 196.560 135.895 196.845 ;
        RECT 130.915 196.180 131.245 196.285 ;
        RECT 132.155 196.180 132.325 196.465 ;
        RECT 128.975 196.095 130.065 196.180 ;
        RECT 128.585 195.640 129.265 195.925 ;
        RECT 129.435 195.855 130.065 196.095 ;
        RECT 129.435 195.355 129.605 195.855 ;
        RECT 126.715 194.895 128.175 195.355 ;
        RECT 123.995 194.415 125.255 194.895 ;
        RECT 115.300 193.965 116.005 194.145 ;
        RECT 114.855 193.565 115.630 193.745 ;
        RECT 113.635 193.500 115.630 193.565 ;
        RECT 115.835 193.535 116.005 193.965 ;
        RECT 118.555 194.090 118.725 194.145 ;
        RECT 116.175 193.715 116.725 193.885 ;
        RECT 113.635 193.225 115.025 193.500 ;
        RECT 115.835 193.205 116.385 193.535 ;
        RECT 116.555 193.390 116.725 193.715 ;
        RECT 116.905 193.625 117.275 193.955 ;
        RECT 117.455 193.715 118.385 193.885 ;
        RECT 118.555 193.775 119.225 194.090 ;
        RECT 117.455 193.390 117.625 193.715 ;
        RECT 118.555 193.535 118.725 193.775 ;
        RECT 119.455 193.545 119.830 194.100 ;
        RECT 120.035 193.565 120.365 194.270 ;
        RECT 121.275 194.145 122.080 194.415 ;
        RECT 123.040 194.145 125.255 194.415 ;
        RECT 121.275 193.995 121.445 194.145 ;
        RECT 120.745 193.975 121.445 193.995 ;
        RECT 123.995 193.975 125.255 194.145 ;
        RECT 120.745 193.785 122.735 193.975 ;
        RECT 116.555 193.220 117.625 193.390 ;
        RECT 115.835 192.155 116.005 193.205 ;
        RECT 116.980 193.105 117.310 193.220 ;
        RECT 117.795 193.205 118.725 193.535 ;
        RECT 118.895 193.395 119.830 193.545 ;
        RECT 120.535 193.395 121.060 193.525 ;
        RECT 118.895 193.205 121.060 193.395 ;
        RECT 118.555 193.035 118.725 193.205 ;
        RECT 120.035 193.195 121.060 193.205 ;
        RECT 116.175 192.935 116.680 193.025 ;
        RECT 117.480 192.935 118.385 193.035 ;
        RECT 116.175 192.765 118.385 192.935 ;
        RECT 118.555 192.865 119.735 193.035 ;
        RECT 116.175 192.335 116.725 192.505 ;
        RECT 115.835 192.135 116.385 192.155 ;
        RECT 110.395 191.845 111.290 192.135 ;
        RECT 111.950 191.845 114.450 192.135 ;
        RECT 115.110 191.845 116.385 192.135 ;
        RECT 110.395 190.280 110.565 191.845 ;
        RECT 113.115 191.120 113.285 191.845 ;
        RECT 115.835 191.825 116.385 191.845 ;
        RECT 116.555 192.010 116.725 192.335 ;
        RECT 116.905 192.245 117.275 192.575 ;
        RECT 117.455 192.335 118.385 192.505 ;
        RECT 117.455 192.010 117.625 192.335 ;
        RECT 118.555 192.155 118.725 192.865 ;
        RECT 118.940 192.520 119.865 192.695 ;
        RECT 120.035 192.645 120.365 193.195 ;
        RECT 121.275 193.025 122.735 193.785 ;
        RECT 120.665 192.855 122.735 193.025 ;
        RECT 121.275 192.765 122.735 192.855 ;
        RECT 122.905 193.515 125.255 193.975 ;
        RECT 125.425 194.835 128.175 194.895 ;
        RECT 125.425 194.145 127.635 194.835 ;
        RECT 128.345 194.665 129.605 195.355 ;
        RECT 130.235 195.730 131.525 196.180 ;
        RECT 131.695 195.875 132.325 196.180 ;
        RECT 132.495 196.105 134.605 196.280 ;
        RECT 132.495 196.045 133.015 196.105 ;
        RECT 133.820 195.975 134.605 196.105 ;
        RECT 134.875 196.275 135.045 196.465 ;
        RECT 136.065 196.445 136.625 197.135 ;
        RECT 136.795 196.845 136.965 197.305 ;
        RECT 137.595 197.385 138.585 197.595 ;
        RECT 139.175 197.385 140.485 197.595 ;
        RECT 137.595 197.285 137.765 197.385 ;
        RECT 137.135 197.015 137.765 197.285 ;
        RECT 136.795 196.560 137.425 196.845 ;
        RECT 137.595 196.715 137.765 197.015 ;
        RECT 137.935 196.965 140.145 197.215 ;
        RECT 137.935 196.885 138.565 196.965 ;
        RECT 139.165 196.885 140.145 196.965 ;
        RECT 140.315 196.915 140.485 197.385 ;
        RECT 140.655 197.305 142.865 197.620 ;
        RECT 140.655 197.085 141.275 197.305 ;
        RECT 141.455 196.965 142.125 197.135 ;
        RECT 142.295 197.005 142.865 197.305 ;
        RECT 137.595 196.485 138.585 196.715 ;
        RECT 137.595 196.275 137.765 196.485 ;
        RECT 138.755 196.465 139.005 196.795 ;
        RECT 140.315 196.715 141.285 196.915 ;
        RECT 139.175 196.585 141.285 196.715 ;
        RECT 139.175 196.485 140.485 196.585 ;
        RECT 131.695 195.855 132.820 195.875 ;
        RECT 130.235 195.335 130.455 195.730 ;
        RECT 129.775 195.055 130.455 195.335 ;
        RECT 130.625 194.865 131.185 195.560 ;
        RECT 131.355 195.335 131.525 195.730 ;
        RECT 132.155 195.475 132.820 195.855 ;
        RECT 133.185 195.505 133.565 195.935 ;
        RECT 131.355 195.055 131.985 195.335 ;
        RECT 127.805 194.145 129.605 194.665 ;
        RECT 129.775 194.465 131.985 194.865 ;
        RECT 125.425 193.685 126.885 194.145 ;
        RECT 129.435 194.065 129.605 194.145 ;
        RECT 130.235 194.085 131.525 194.295 ;
        RECT 127.215 193.805 129.265 193.975 ;
        RECT 127.215 193.700 127.560 193.805 ;
        RECT 128.295 193.700 129.265 193.805 ;
        RECT 129.435 193.795 130.065 194.065 ;
        RECT 120.535 192.530 121.055 192.685 ;
        RECT 118.940 192.475 119.915 192.520 ;
        RECT 120.495 192.475 121.055 192.530 ;
        RECT 118.940 192.365 121.055 192.475 ;
        RECT 119.785 192.355 121.055 192.365 ;
        RECT 119.785 192.305 120.620 192.355 ;
        RECT 116.555 191.840 117.625 192.010 ;
        RECT 117.795 192.135 118.725 192.155 ;
        RECT 121.275 192.135 122.215 192.765 ;
        RECT 122.905 192.595 125.775 193.515 ;
        RECT 117.795 191.845 119.890 192.135 ;
        RECT 120.550 191.845 122.215 192.135 ;
        RECT 113.455 191.395 115.665 191.675 ;
        RECT 113.455 191.290 114.425 191.395 ;
        RECT 115.095 191.290 115.665 191.395 ;
        RECT 114.595 191.120 114.925 191.225 ;
        RECT 115.835 191.120 116.005 191.825 ;
        RECT 116.980 191.725 117.310 191.840 ;
        RECT 117.795 191.825 118.725 191.845 ;
        RECT 116.175 191.555 116.680 191.645 ;
        RECT 117.480 191.555 118.385 191.655 ;
        RECT 116.175 191.385 118.385 191.555 ;
        RECT 113.115 190.795 113.745 191.120 ;
        RECT 110.735 190.495 111.285 190.665 ;
        RECT 110.395 189.950 110.945 190.280 ;
        RECT 111.115 190.120 111.285 190.495 ;
        RECT 111.465 190.400 111.835 190.755 ;
        RECT 112.015 190.495 112.945 190.665 ;
        RECT 112.015 190.120 112.185 190.495 ;
        RECT 113.115 190.280 113.285 190.795 ;
        RECT 111.115 189.950 112.185 190.120 ;
        RECT 112.355 189.950 113.285 190.280 ;
        RECT 113.915 190.670 115.205 191.120 ;
        RECT 115.375 190.795 116.005 191.120 ;
        RECT 116.175 190.955 116.725 191.125 ;
        RECT 113.915 190.275 114.135 190.670 ;
        RECT 113.455 189.995 114.135 190.275 ;
        RECT 110.395 189.350 110.565 189.950 ;
        RECT 111.475 189.865 111.805 189.950 ;
        RECT 110.735 189.695 111.310 189.780 ;
        RECT 112.040 189.695 112.945 189.780 ;
        RECT 110.735 189.525 112.945 189.695 ;
        RECT 113.115 189.350 113.285 189.950 ;
        RECT 114.305 189.805 114.865 190.500 ;
        RECT 115.035 190.275 115.205 190.670 ;
        RECT 115.835 190.775 116.005 190.795 ;
        RECT 115.835 190.445 116.385 190.775 ;
        RECT 116.555 190.630 116.725 190.955 ;
        RECT 116.905 190.865 117.275 191.195 ;
        RECT 118.555 191.165 118.725 191.825 ;
        RECT 118.895 191.500 121.105 191.670 ;
        RECT 118.895 191.335 119.865 191.500 ;
        RECT 120.535 191.415 121.105 191.500 ;
        RECT 121.275 191.385 122.215 191.845 ;
        RECT 122.385 192.305 125.775 192.595 ;
        RECT 125.945 193.510 126.885 193.685 ;
        RECT 127.795 193.530 128.125 193.635 ;
        RECT 125.945 193.130 127.285 193.510 ;
        RECT 127.455 193.360 128.465 193.530 ;
        RECT 129.435 193.490 129.605 193.795 ;
        RECT 130.235 193.625 130.455 194.085 ;
        RECT 125.945 192.620 126.885 193.130 ;
        RECT 127.455 192.960 127.625 193.360 ;
        RECT 127.105 192.790 127.625 192.960 ;
        RECT 127.795 192.810 128.125 193.190 ;
        RECT 128.295 193.040 128.465 193.360 ;
        RECT 128.635 193.210 129.605 193.490 ;
        RECT 129.775 193.340 130.455 193.625 ;
        RECT 130.625 193.225 131.185 193.915 ;
        RECT 131.355 193.625 131.525 194.085 ;
        RECT 132.155 194.065 132.325 195.475 ;
        RECT 133.185 195.115 133.715 195.505 ;
        RECT 132.655 194.945 133.715 195.115 ;
        RECT 133.885 195.105 134.195 195.800 ;
        RECT 134.875 195.795 136.135 196.275 ;
        RECT 134.405 195.585 136.135 195.795 ;
        RECT 136.305 195.845 137.765 196.275 ;
        RECT 138.025 196.015 138.485 196.185 ;
        RECT 136.305 195.755 138.145 195.845 ;
        RECT 134.405 195.110 136.675 195.585 ;
        RECT 132.655 194.885 132.850 194.945 ;
        RECT 132.510 194.715 132.850 194.885 ;
        RECT 133.545 194.930 133.715 194.945 ;
        RECT 134.875 195.065 136.675 195.110 ;
        RECT 136.845 195.515 138.145 195.755 ;
        RECT 138.315 195.750 138.485 196.015 ;
        RECT 138.655 195.920 139.305 196.270 ;
        RECT 139.475 196.015 140.145 196.185 ;
        RECT 139.475 195.750 139.645 196.015 ;
        RECT 140.315 195.845 140.485 196.485 ;
        RECT 141.455 196.280 141.625 196.965 ;
        RECT 143.035 196.835 143.205 197.840 ;
        RECT 143.755 197.625 143.925 198.000 ;
        RECT 143.375 197.455 143.925 197.625 ;
        RECT 144.105 197.365 144.475 197.720 ;
        RECT 144.655 197.625 144.825 198.000 ;
        RECT 144.995 197.840 145.925 198.170 ;
        RECT 144.655 197.455 145.585 197.625 ;
        RECT 141.795 196.450 142.355 196.715 ;
        RECT 142.525 196.625 143.205 196.835 ;
        RECT 143.375 196.795 144.005 197.080 ;
        RECT 142.525 196.620 143.665 196.625 ;
        RECT 142.525 196.280 142.855 196.390 ;
        RECT 141.455 196.110 142.855 196.280 ;
        RECT 143.035 196.355 143.665 196.620 ;
        RECT 141.455 196.100 141.625 196.110 ;
        RECT 138.315 195.520 139.645 195.750 ;
        RECT 139.815 195.515 140.485 195.845 ;
        RECT 141.280 195.710 141.625 196.100 ;
        RECT 141.795 195.585 142.355 195.940 ;
        RECT 143.035 195.930 143.205 196.355 ;
        RECT 143.835 196.335 144.005 196.795 ;
        RECT 144.175 196.505 144.735 197.195 ;
        RECT 144.905 196.795 145.585 197.080 ;
        RECT 144.905 196.335 145.125 196.795 ;
        RECT 145.755 196.625 145.925 197.840 ;
        RECT 145.295 196.355 145.925 196.625 ;
        RECT 143.835 196.125 145.125 196.335 ;
        RECT 142.525 195.690 143.205 195.930 ;
        RECT 136.845 195.065 137.765 195.515 ;
        RECT 138.025 195.160 140.145 195.345 ;
        RECT 133.045 194.455 133.375 194.775 ;
        RECT 133.545 194.645 134.660 194.930 ;
        RECT 133.045 194.435 134.255 194.455 ;
        RECT 134.875 194.445 135.045 195.065 ;
        RECT 137.595 194.905 137.765 195.065 ;
        RECT 132.520 194.220 134.255 194.435 ;
        RECT 132.520 194.195 132.895 194.220 ;
        RECT 131.695 194.025 132.325 194.065 ;
        RECT 131.695 193.795 132.830 194.025 ;
        RECT 132.155 193.695 132.830 193.795 ;
        RECT 133.005 193.750 133.855 194.050 ;
        RECT 134.025 193.945 134.255 194.220 ;
        RECT 134.425 194.115 135.045 194.445 ;
        RECT 134.025 193.775 134.685 193.945 ;
        RECT 133.005 193.745 133.175 193.750 ;
        RECT 131.355 193.340 131.985 193.625 ;
        RECT 128.295 192.870 128.755 193.040 ;
        RECT 125.945 192.305 127.285 192.620 ;
        RECT 122.385 192.135 124.165 192.305 ;
        RECT 126.715 192.290 127.285 192.305 ;
        RECT 126.715 192.135 126.885 192.290 ;
        RECT 122.385 191.845 125.330 192.135 ;
        RECT 125.990 191.845 126.885 192.135 ;
        RECT 127.455 192.115 127.625 192.790 ;
        RECT 127.105 191.945 127.625 192.115 ;
        RECT 127.795 191.900 128.415 192.640 ;
        RECT 122.385 191.385 124.165 191.845 ;
        RECT 126.715 191.745 126.885 191.845 ;
        RECT 120.035 191.245 120.365 191.330 ;
        RECT 121.275 191.245 121.445 191.385 ;
        RECT 117.455 190.955 118.385 191.125 ;
        RECT 118.555 190.995 119.865 191.165 ;
        RECT 120.035 191.075 120.705 191.245 ;
        RECT 117.455 190.630 117.625 190.955 ;
        RECT 118.555 190.775 118.725 190.995 ;
        RECT 120.035 190.825 120.365 190.850 ;
        RECT 116.555 190.460 117.625 190.630 ;
        RECT 115.035 189.995 115.665 190.275 ;
        RECT 113.455 189.405 115.665 189.805 ;
        RECT 110.395 189.090 111.405 189.350 ;
        RECT 111.965 189.090 113.285 189.350 ;
        RECT 115.835 189.395 116.005 190.445 ;
        RECT 116.980 190.345 117.310 190.460 ;
        RECT 117.795 190.445 118.725 190.775 ;
        RECT 116.175 190.175 116.680 190.265 ;
        RECT 117.480 190.175 118.385 190.275 ;
        RECT 116.175 190.005 118.385 190.175 ;
        RECT 116.175 189.575 116.725 189.745 ;
        RECT 110.395 188.475 110.565 189.090 ;
        RECT 113.115 189.005 113.285 189.090 ;
        RECT 113.915 189.025 115.205 189.235 ;
        RECT 110.735 188.735 112.945 188.915 ;
        RECT 110.735 188.655 111.240 188.735 ;
        RECT 112.040 188.645 112.945 188.735 ;
        RECT 113.115 188.735 113.745 189.005 ;
        RECT 110.395 188.145 110.945 188.475 ;
        RECT 111.540 188.460 111.870 188.565 ;
        RECT 113.115 188.475 113.285 188.735 ;
        RECT 113.915 188.565 114.135 189.025 ;
        RECT 111.115 188.290 112.185 188.460 ;
        RECT 110.395 186.610 110.565 188.145 ;
        RECT 111.115 187.965 111.285 188.290 ;
        RECT 110.735 187.795 111.285 187.965 ;
        RECT 111.465 187.725 111.835 188.065 ;
        RECT 112.015 187.965 112.185 188.290 ;
        RECT 112.355 188.145 113.285 188.475 ;
        RECT 113.455 188.280 114.135 188.565 ;
        RECT 114.305 188.165 114.865 188.855 ;
        RECT 115.035 188.565 115.205 189.025 ;
        RECT 115.835 189.065 116.385 189.395 ;
        RECT 116.555 189.250 116.725 189.575 ;
        RECT 116.905 189.485 117.275 189.815 ;
        RECT 117.455 189.575 118.385 189.745 ;
        RECT 117.455 189.250 117.625 189.575 ;
        RECT 118.555 189.395 118.725 190.445 ;
        RECT 116.555 189.080 117.625 189.250 ;
        RECT 115.835 189.005 116.005 189.065 ;
        RECT 115.375 188.735 116.005 189.005 ;
        RECT 116.980 188.965 117.310 189.080 ;
        RECT 117.795 189.065 118.725 189.395 ;
        RECT 115.035 188.280 115.665 188.565 ;
        RECT 115.835 188.445 116.005 188.735 ;
        RECT 116.175 188.795 116.680 188.885 ;
        RECT 117.480 188.795 118.385 188.895 ;
        RECT 116.175 188.625 118.385 188.795 ;
        RECT 118.555 188.625 118.725 189.065 ;
        RECT 118.895 190.655 120.365 190.825 ;
        RECT 118.895 188.965 119.065 190.655 ;
        RECT 120.535 190.490 120.705 191.075 ;
        RECT 120.875 190.915 121.445 191.245 ;
        RECT 120.535 190.485 121.105 190.490 ;
        RECT 119.235 190.315 121.105 190.485 ;
        RECT 119.235 189.360 119.405 190.315 ;
        RECT 119.575 189.975 120.545 190.145 ;
        RECT 119.575 189.325 119.745 189.975 ;
        RECT 120.740 189.960 121.105 190.315 ;
        RECT 121.275 190.185 121.445 190.915 ;
        RECT 121.615 190.355 122.245 190.640 ;
        RECT 121.275 189.915 121.905 190.185 ;
        RECT 120.765 189.770 120.935 189.775 ;
        RECT 119.945 189.495 121.105 189.770 ;
        RECT 119.575 189.135 121.105 189.325 ;
        RECT 118.895 188.795 119.920 188.965 ;
        RECT 121.275 188.955 121.445 189.915 ;
        RECT 122.075 189.895 122.245 190.355 ;
        RECT 122.415 190.065 122.975 190.755 ;
        RECT 123.145 190.355 123.825 190.640 ;
        RECT 123.995 190.385 124.165 191.385 ;
        RECT 124.805 191.375 126.145 191.500 ;
        RECT 124.375 191.330 126.145 191.375 ;
        RECT 126.715 191.415 127.385 191.745 ;
        RECT 128.585 191.730 128.755 192.870 ;
        RECT 126.715 191.345 126.885 191.415 ;
        RECT 124.375 191.045 124.975 191.330 ;
        RECT 125.145 190.915 125.805 191.160 ;
        RECT 124.385 190.615 124.975 190.865 ;
        RECT 125.975 190.845 126.145 191.330 ;
        RECT 126.315 191.015 126.885 191.345 ;
        RECT 127.795 191.220 128.125 191.630 ;
        RECT 128.295 191.410 128.755 191.730 ;
        RECT 123.145 189.895 123.365 190.355 ;
        RECT 123.995 190.185 124.635 190.385 ;
        RECT 123.535 190.055 124.635 190.185 ;
        RECT 123.535 189.915 124.165 190.055 ;
        RECT 122.075 189.685 123.365 189.895 ;
        RECT 121.615 189.115 123.825 189.515 ;
        RECT 123.995 189.385 124.165 189.915 ;
        RECT 124.805 189.825 124.975 190.615 ;
        RECT 125.145 190.435 125.805 190.700 ;
        RECT 125.975 190.515 126.485 190.845 ;
        RECT 126.715 190.805 126.885 191.015 ;
        RECT 127.105 191.215 128.125 191.220 ;
        RECT 127.105 190.975 128.720 191.215 ;
        RECT 128.925 190.990 129.215 193.040 ;
        RECT 129.435 192.135 129.605 193.210 ;
        RECT 132.155 192.135 132.325 193.695 ;
        RECT 134.875 193.065 135.045 194.115 ;
        RECT 135.265 193.235 135.555 194.890 ;
        RECT 135.725 194.570 136.185 194.890 ;
        RECT 135.725 193.470 135.895 194.570 ;
        RECT 136.355 194.540 136.925 194.890 ;
        RECT 137.595 194.885 138.225 194.905 ;
        RECT 137.095 194.655 138.225 194.885 ;
        RECT 138.395 194.710 139.345 194.990 ;
        RECT 140.315 194.920 140.485 195.515 ;
        RECT 140.655 195.095 141.585 195.265 ;
        RECT 139.855 194.880 140.485 194.920 ;
        RECT 139.855 194.655 141.245 194.880 ;
        RECT 137.095 194.555 137.765 194.655 ;
        RECT 136.065 193.660 136.685 194.370 ;
        RECT 136.855 194.185 137.375 194.355 ;
        RECT 135.725 193.300 136.185 193.470 ;
        RECT 134.875 192.785 135.845 193.065 ;
        RECT 136.015 192.915 136.185 193.300 ;
        RECT 136.355 193.085 136.685 193.490 ;
        RECT 136.855 193.485 137.025 194.185 ;
        RECT 137.595 193.985 137.765 194.555 ;
        RECT 140.315 194.550 141.245 194.655 ;
        RECT 141.415 194.720 141.585 195.095 ;
        RECT 141.765 195.000 142.135 195.355 ;
        RECT 142.315 195.095 142.865 195.265 ;
        RECT 142.315 194.720 142.485 195.095 ;
        RECT 143.035 194.880 143.205 195.690 ;
        RECT 143.375 195.555 145.585 195.955 ;
        RECT 143.375 195.085 144.005 195.365 ;
        RECT 141.415 194.550 142.485 194.720 ;
        RECT 142.655 194.565 143.205 194.880 ;
        RECT 143.835 194.690 144.005 195.085 ;
        RECT 144.175 194.860 144.735 195.555 ;
        RECT 144.905 195.085 145.585 195.365 ;
        RECT 144.905 194.690 145.125 195.085 ;
        RECT 142.655 194.550 143.665 194.565 ;
        RECT 138.355 194.485 139.720 194.540 ;
        RECT 138.045 194.370 140.145 194.485 ;
        RECT 138.045 194.315 138.485 194.370 ;
        RECT 138.045 194.150 138.215 194.315 ;
        RECT 139.590 194.235 140.145 194.370 ;
        RECT 137.195 193.655 137.765 193.985 ;
        RECT 136.855 193.315 137.375 193.485 ;
        RECT 136.855 192.915 137.025 193.315 ;
        RECT 137.595 193.145 137.765 193.655 ;
        RECT 138.045 193.450 138.215 193.955 ;
        RECT 138.415 193.790 138.635 194.145 ;
        RECT 138.805 193.960 139.400 194.200 ;
        RECT 138.415 193.620 139.700 193.790 ;
        RECT 138.045 193.280 139.165 193.450 ;
        RECT 132.505 192.285 134.705 192.595 ;
        RECT 132.505 192.155 133.065 192.285 ;
        RECT 134.075 192.155 134.705 192.285 ;
        RECT 129.435 191.845 130.770 192.135 ;
        RECT 131.430 191.985 132.325 192.135 ;
        RECT 134.875 192.135 135.045 192.785 ;
        RECT 136.015 192.745 137.025 192.915 ;
        RECT 137.195 192.960 137.765 193.145 ;
        RECT 138.995 193.090 139.165 193.280 ;
        RECT 139.335 193.260 139.700 193.620 ;
        RECT 139.870 193.090 140.040 194.025 ;
        RECT 137.195 192.765 138.265 192.960 ;
        RECT 136.355 192.645 136.685 192.745 ;
        RECT 137.595 192.590 138.265 192.765 ;
        RECT 138.445 192.870 138.775 193.070 ;
        RECT 138.995 192.920 140.040 193.090 ;
        RECT 140.315 193.950 140.485 194.550 ;
        RECT 141.795 194.465 142.125 194.550 ;
        RECT 140.655 194.295 141.560 194.380 ;
        RECT 142.290 194.295 142.865 194.380 ;
        RECT 140.655 194.125 142.865 194.295 ;
        RECT 143.035 194.240 143.665 194.550 ;
        RECT 143.835 194.240 145.125 194.690 ;
        RECT 145.755 194.565 145.925 196.355 ;
        RECT 145.295 194.240 145.925 194.565 ;
        RECT 143.035 193.950 143.205 194.240 ;
        RECT 144.115 194.135 144.445 194.240 ;
        RECT 140.315 193.690 141.635 193.950 ;
        RECT 142.195 193.690 143.205 193.950 ;
        RECT 140.315 193.475 140.485 193.690 ;
        RECT 140.315 193.245 141.625 193.475 ;
        RECT 135.215 192.475 136.185 192.575 ;
        RECT 136.920 192.475 137.265 192.575 ;
        RECT 135.215 192.305 137.265 192.475 ;
        RECT 137.595 192.135 137.765 192.590 ;
        RECT 138.445 192.410 138.745 192.870 ;
        RECT 138.995 192.750 139.255 192.920 ;
        RECT 140.315 192.750 140.485 193.245 ;
        RECT 141.795 193.165 142.045 193.495 ;
        RECT 143.035 193.475 143.205 193.690 ;
        RECT 143.375 193.965 143.945 194.070 ;
        RECT 144.615 193.965 145.585 194.070 ;
        RECT 143.375 193.685 145.585 193.965 ;
        RECT 142.215 193.245 143.205 193.475 ;
        RECT 143.375 193.255 143.925 193.425 ;
        RECT 143.035 193.075 143.205 193.245 ;
        RECT 138.925 192.580 139.255 192.750 ;
        RECT 139.515 192.580 140.485 192.750 ;
        RECT 140.655 192.995 141.635 193.075 ;
        RECT 142.235 192.995 142.865 193.075 ;
        RECT 140.655 192.745 142.865 192.995 ;
        RECT 143.035 192.745 143.585 193.075 ;
        RECT 143.755 192.930 143.925 193.255 ;
        RECT 144.105 193.155 144.475 193.495 ;
        RECT 144.655 193.255 145.585 193.435 ;
        RECT 144.655 192.930 144.825 193.255 ;
        RECT 145.755 193.075 145.925 194.240 ;
        RECT 143.755 192.760 144.825 192.930 ;
        RECT 140.315 192.575 140.485 192.580 ;
        RECT 143.035 192.575 143.205 192.745 ;
        RECT 144.180 192.655 144.510 192.760 ;
        RECT 144.995 192.745 145.925 193.075 ;
        RECT 131.430 191.845 133.065 191.985 ;
        RECT 133.235 191.945 133.855 192.115 ;
        RECT 134.875 191.980 136.210 192.135 ;
        RECT 129.435 190.805 129.605 191.845 ;
        RECT 125.145 189.955 125.805 190.240 ;
        RECT 124.385 189.575 124.975 189.825 ;
        RECT 125.145 189.565 125.805 189.780 ;
        RECT 125.475 189.475 125.805 189.565 ;
        RECT 123.995 189.135 125.305 189.385 ;
        RECT 125.975 189.305 126.145 190.515 ;
        RECT 126.715 190.465 127.385 190.805 ;
        RECT 127.555 190.465 128.125 190.805 ;
        RECT 128.360 190.465 129.605 190.805 ;
        RECT 129.825 190.485 130.115 191.675 ;
        RECT 130.285 191.330 130.745 191.655 ;
        RECT 130.915 191.330 131.245 191.675 ;
        RECT 131.415 191.405 131.935 191.660 ;
        RECT 132.155 191.535 133.065 191.845 ;
        RECT 130.285 190.655 130.455 191.330 ;
        RECT 130.625 190.965 131.245 191.160 ;
        RECT 130.285 190.485 130.745 190.655 ;
        RECT 126.715 190.275 126.885 190.465 ;
        RECT 129.435 190.315 129.605 190.465 ;
        RECT 126.715 190.035 127.695 190.275 ;
        RECT 126.715 189.465 126.885 190.035 ;
        RECT 127.875 189.945 128.125 190.295 ;
        RECT 128.295 189.955 129.250 190.285 ;
        RECT 129.435 190.035 130.405 190.315 ;
        RECT 130.575 190.165 130.745 190.485 ;
        RECT 130.915 190.335 131.245 190.965 ;
        RECT 131.415 190.735 131.585 191.405 ;
        RECT 132.155 191.235 132.325 191.535 ;
        RECT 133.235 191.385 133.515 191.775 ;
        RECT 133.685 191.495 133.855 191.945 ;
        RECT 134.025 191.845 136.210 191.980 ;
        RECT 136.870 191.845 137.765 192.135 ;
        RECT 138.045 192.240 140.145 192.410 ;
        RECT 138.045 192.005 138.215 192.240 ;
        RECT 139.815 192.160 140.145 192.240 ;
        RECT 140.315 192.365 141.625 192.575 ;
        RECT 142.215 192.365 143.205 192.575 ;
        RECT 140.315 192.135 140.485 192.365 ;
        RECT 143.035 192.135 143.205 192.365 ;
        RECT 143.375 192.485 143.880 192.565 ;
        RECT 144.680 192.485 145.585 192.575 ;
        RECT 143.375 192.305 145.585 192.485 ;
        RECT 145.755 192.135 145.925 192.745 ;
        RECT 138.925 191.880 139.645 192.070 ;
        RECT 134.025 191.665 135.045 191.845 ;
        RECT 131.755 191.025 132.325 191.235 ;
        RECT 132.495 191.195 133.065 191.365 ;
        RECT 133.685 191.325 134.705 191.495 ;
        RECT 131.755 190.905 132.725 191.025 ;
        RECT 131.415 190.565 131.935 190.735 ;
        RECT 132.155 190.605 132.725 190.905 ;
        RECT 131.415 190.165 131.585 190.565 ;
        RECT 132.155 190.395 132.325 190.605 ;
        RECT 132.895 190.435 133.065 191.195 ;
        RECT 133.235 191.155 133.565 191.200 ;
        RECT 133.235 190.955 134.365 191.155 ;
        RECT 133.235 190.505 134.365 190.755 ;
        RECT 127.055 189.775 127.695 189.865 ;
        RECT 128.295 189.775 128.465 189.955 ;
        RECT 127.055 189.605 128.465 189.775 ;
        RECT 127.055 189.535 127.695 189.605 ;
        RECT 125.475 189.135 126.145 189.305 ;
        RECT 126.315 189.365 126.885 189.465 ;
        RECT 126.315 189.135 127.695 189.365 ;
        RECT 118.555 188.455 119.485 188.625 ;
        RECT 115.835 188.175 116.815 188.445 ;
        RECT 112.015 187.785 112.945 187.965 ;
        RECT 113.115 187.065 113.285 188.145 ;
        RECT 115.835 187.505 116.005 188.175 ;
        RECT 116.995 188.105 117.245 188.455 ;
        RECT 118.555 188.445 118.725 188.455 ;
        RECT 117.415 188.115 118.725 188.445 ;
        RECT 116.175 187.935 116.815 188.005 ;
        RECT 116.175 187.765 117.585 187.935 ;
        RECT 116.175 187.675 116.815 187.765 ;
        RECT 115.835 187.265 116.815 187.505 ;
        RECT 113.115 186.735 114.005 187.065 ;
        RECT 114.305 186.845 114.845 187.075 ;
        RECT 114.645 186.745 114.845 186.845 ;
        RECT 115.015 186.735 115.665 187.075 ;
        RECT 110.395 186.275 111.070 186.610 ;
        RECT 110.395 184.850 110.565 186.275 ;
        RECT 111.245 186.255 112.095 186.555 ;
        RECT 112.265 186.355 112.925 186.525 ;
        RECT 110.760 186.085 111.135 186.105 ;
        RECT 112.265 186.085 112.495 186.355 ;
        RECT 113.115 186.185 113.285 186.735 ;
        RECT 113.530 186.435 114.825 186.555 ;
        RECT 113.530 186.340 114.845 186.435 ;
        RECT 110.760 185.865 112.495 186.085 ;
        RECT 111.285 185.850 112.495 185.865 ;
        RECT 112.665 185.855 113.285 186.185 ;
        RECT 110.750 185.415 111.090 185.585 ;
        RECT 111.285 185.550 111.615 185.850 ;
        RECT 110.895 185.380 111.090 185.415 ;
        RECT 111.785 185.395 112.900 185.680 ;
        RECT 113.115 185.645 113.285 185.855 ;
        RECT 113.455 185.815 114.445 186.145 ;
        RECT 114.645 186.105 114.845 186.340 ;
        RECT 115.015 186.225 115.205 186.735 ;
        RECT 115.835 186.565 116.005 187.265 ;
        RECT 116.995 187.245 117.245 187.595 ;
        RECT 117.415 187.585 117.585 187.765 ;
        RECT 117.415 187.255 118.370 187.585 ;
        RECT 118.555 187.095 118.725 188.115 ;
        RECT 119.075 188.045 119.485 188.220 ;
        RECT 119.730 188.215 119.920 188.795 ;
        RECT 120.295 188.225 120.465 188.935 ;
        RECT 120.740 188.445 121.445 188.955 ;
        RECT 121.615 188.645 122.245 188.925 ;
        RECT 120.295 188.045 121.070 188.225 ;
        RECT 119.075 187.980 121.070 188.045 ;
        RECT 121.275 188.125 121.445 188.445 ;
        RECT 122.075 188.250 122.245 188.645 ;
        RECT 122.415 188.420 122.975 189.115 ;
        RECT 123.145 188.645 123.825 188.925 ;
        RECT 123.145 188.250 123.365 188.645 ;
        RECT 119.075 187.705 120.465 187.980 ;
        RECT 121.275 187.800 121.905 188.125 ;
        RECT 122.075 187.800 123.365 188.250 ;
        RECT 123.995 188.125 124.165 189.135 ;
        RECT 125.475 188.995 125.805 189.135 ;
        RECT 126.715 189.095 127.695 189.135 ;
        RECT 124.375 188.825 125.225 188.965 ;
        RECT 125.990 188.825 126.500 188.965 ;
        RECT 124.375 188.635 126.500 188.825 ;
        RECT 123.535 187.800 124.165 188.125 ;
        RECT 118.895 187.275 119.825 187.445 ;
        RECT 116.370 186.820 118.385 187.075 ;
        RECT 116.370 186.715 116.745 186.820 ;
        RECT 117.400 186.735 118.385 186.820 ;
        RECT 118.555 186.765 119.485 187.095 ;
        RECT 119.655 186.950 119.825 187.275 ;
        RECT 120.005 187.185 120.375 187.515 ;
        RECT 120.555 187.275 121.105 187.445 ;
        RECT 120.555 186.950 120.725 187.275 ;
        RECT 121.275 187.095 121.445 187.800 ;
        RECT 122.355 187.695 122.685 187.800 ;
        RECT 121.615 187.525 122.185 187.630 ;
        RECT 122.855 187.525 123.825 187.630 ;
        RECT 121.615 187.245 123.825 187.525 ;
        RECT 123.995 187.320 124.165 187.800 ;
        RECT 126.715 188.475 126.885 189.095 ;
        RECT 127.875 189.085 128.125 189.435 ;
        RECT 129.435 189.425 129.605 190.035 ;
        RECT 130.575 189.995 131.585 190.165 ;
        RECT 131.755 190.015 132.325 190.395 ;
        RECT 132.495 190.205 133.065 190.435 ;
        RECT 134.535 190.315 134.705 191.325 ;
        RECT 130.915 189.890 131.245 189.995 ;
        RECT 129.775 189.720 130.745 189.825 ;
        RECT 131.480 189.720 131.825 189.825 ;
        RECT 129.775 189.550 131.825 189.720 ;
        RECT 128.295 189.375 129.605 189.425 ;
        RECT 132.155 189.375 132.325 190.015 ;
        RECT 132.495 189.715 133.065 190.035 ;
        RECT 133.235 189.885 133.565 190.290 ;
        RECT 133.735 190.065 134.705 190.315 ;
        RECT 134.875 191.165 135.045 191.665 ;
        RECT 135.215 191.420 137.230 191.675 ;
        RECT 135.215 191.335 136.200 191.420 ;
        RECT 136.855 191.315 137.230 191.420 ;
        RECT 136.355 191.165 136.685 191.250 ;
        RECT 134.875 190.755 135.475 191.165 ;
        RECT 135.645 190.900 136.685 191.165 ;
        RECT 137.595 191.050 137.765 191.845 ;
        RECT 138.045 191.220 138.215 191.835 ;
        RECT 138.385 191.710 138.715 191.855 ;
        RECT 138.385 191.390 139.675 191.710 ;
        RECT 139.845 191.220 140.015 191.935 ;
        RECT 138.045 191.050 140.015 191.220 ;
        RECT 140.315 191.845 141.650 192.135 ;
        RECT 142.310 191.845 143.930 192.135 ;
        RECT 144.590 191.845 145.925 192.135 ;
        RECT 140.315 191.060 140.485 191.845 ;
        RECT 140.655 191.365 142.855 191.675 ;
        RECT 140.655 191.235 141.285 191.365 ;
        RECT 142.295 191.235 142.855 191.365 ;
        RECT 133.735 189.715 133.905 190.065 ;
        RECT 134.875 190.010 135.045 190.755 ;
        RECT 134.875 189.885 135.465 190.010 ;
        RECT 132.495 189.545 133.905 189.715 ;
        RECT 134.075 189.680 135.465 189.885 ;
        RECT 135.645 189.890 135.815 190.900 ;
        RECT 136.855 190.880 137.765 191.050 ;
        RECT 137.595 190.775 137.765 190.880 ;
        RECT 135.985 190.230 136.155 190.685 ;
        RECT 136.355 190.400 136.685 190.730 ;
        RECT 136.855 190.430 137.230 190.600 ;
        RECT 137.595 190.565 138.295 190.775 ;
        RECT 136.855 190.230 137.025 190.430 ;
        RECT 135.985 190.060 137.025 190.230 ;
        RECT 135.645 189.720 137.425 189.890 ;
        RECT 137.595 189.805 137.765 190.565 ;
        RECT 138.675 190.345 139.005 191.050 ;
        RECT 139.210 190.325 139.585 190.880 ;
        RECT 140.315 190.870 141.335 191.060 ;
        RECT 139.815 190.745 141.335 190.870 ;
        RECT 141.505 191.025 142.125 191.195 ;
        RECT 143.035 191.065 143.205 191.845 ;
        RECT 139.815 190.555 140.485 190.745 ;
        RECT 141.505 190.575 141.675 191.025 ;
        RECT 137.980 190.175 138.505 190.305 ;
        RECT 139.210 190.175 140.145 190.325 ;
        RECT 137.980 189.985 140.145 190.175 ;
        RECT 137.980 189.975 139.005 189.985 ;
        RECT 134.075 189.555 135.045 189.680 ;
        RECT 128.295 189.095 130.695 189.375 ;
        RECT 127.055 188.655 127.605 188.825 ;
        RECT 126.715 188.145 127.265 188.475 ;
        RECT 127.435 188.330 127.605 188.655 ;
        RECT 127.785 188.555 128.155 188.895 ;
        RECT 128.335 188.655 129.265 188.835 ;
        RECT 128.335 188.330 128.505 188.655 ;
        RECT 129.435 188.475 130.695 189.095 ;
        RECT 127.435 188.160 128.505 188.330 ;
        RECT 119.655 186.780 120.725 186.950 ;
        RECT 115.375 186.450 116.005 186.565 ;
        RECT 116.915 186.565 117.245 186.650 ;
        RECT 118.555 186.565 118.725 186.765 ;
        RECT 119.970 186.665 120.300 186.780 ;
        RECT 120.895 186.765 121.445 187.095 ;
        RECT 115.375 186.395 116.745 186.450 ;
        RECT 115.835 186.280 116.745 186.395 ;
        RECT 116.915 186.300 117.955 186.565 ;
        RECT 111.785 185.380 111.955 185.395 ;
        RECT 110.895 185.210 111.955 185.380 ;
        RECT 110.395 184.455 111.060 184.850 ;
        RECT 111.425 184.820 111.955 185.210 ;
        RECT 110.395 183.395 110.565 184.455 ;
        RECT 111.425 184.395 111.805 184.820 ;
        RECT 112.125 184.525 112.435 185.220 ;
        RECT 113.115 185.215 114.060 185.645 ;
        RECT 112.645 184.935 114.060 185.215 ;
        RECT 114.230 185.280 114.445 185.815 ;
        RECT 114.615 185.465 114.845 185.935 ;
        RECT 115.015 185.895 115.285 186.225 ;
        RECT 115.400 185.760 115.665 185.765 ;
        RECT 115.395 185.755 115.665 185.760 ;
        RECT 115.385 185.750 115.665 185.755 ;
        RECT 115.380 185.745 115.665 185.750 ;
        RECT 115.370 185.740 115.665 185.745 ;
        RECT 115.365 185.730 115.665 185.740 ;
        RECT 115.355 185.720 115.665 185.730 ;
        RECT 115.345 185.705 115.665 185.720 ;
        RECT 115.015 185.405 115.665 185.705 ;
        RECT 115.015 185.280 115.205 185.405 ;
        RECT 114.230 184.995 115.205 185.280 ;
        RECT 115.835 185.165 116.005 186.280 ;
        RECT 116.370 185.830 116.745 186.000 ;
        RECT 116.575 185.630 116.745 185.830 ;
        RECT 116.915 185.800 117.245 186.130 ;
        RECT 117.445 185.630 117.615 186.085 ;
        RECT 116.575 185.460 117.615 185.630 ;
        RECT 117.785 185.290 117.955 186.300 ;
        RECT 118.125 186.155 118.725 186.565 ;
        RECT 118.895 186.495 119.800 186.595 ;
        RECT 120.600 186.495 121.105 186.585 ;
        RECT 118.895 186.325 121.105 186.495 ;
        RECT 121.275 186.465 121.445 186.765 ;
        RECT 121.625 186.765 123.825 187.075 ;
        RECT 121.625 186.635 122.185 186.765 ;
        RECT 123.195 186.635 123.825 186.765 ;
        RECT 123.995 186.990 125.265 187.320 ;
        RECT 118.555 185.675 118.725 186.155 ;
        RECT 118.895 185.985 120.945 186.155 ;
        RECT 118.895 185.885 119.865 185.985 ;
        RECT 120.600 185.885 120.945 185.985 ;
        RECT 121.275 186.015 122.185 186.465 ;
        RECT 122.355 186.425 122.975 186.595 ;
        RECT 123.995 186.460 124.165 186.990 ;
        RECT 125.515 186.890 125.725 187.535 ;
        RECT 125.895 187.050 126.530 187.380 ;
        RECT 120.035 185.715 120.365 185.815 ;
        RECT 118.555 185.410 119.525 185.675 ;
        RECT 115.375 184.995 116.005 185.165 ;
        RECT 116.175 185.120 117.955 185.290 ;
        RECT 112.645 184.530 113.285 184.935 ;
        RECT 114.890 184.765 115.665 184.825 ;
        RECT 110.735 184.220 111.255 184.285 ;
        RECT 112.060 184.220 112.845 184.350 ;
        RECT 110.735 184.045 112.845 184.220 ;
        RECT 113.115 183.395 113.285 184.530 ;
        RECT 113.455 184.485 115.665 184.765 ;
        RECT 115.835 184.390 116.005 184.995 ;
        RECT 116.175 184.560 116.825 184.890 ;
        RECT 115.835 184.220 116.475 184.390 ;
        RECT 115.835 183.395 116.005 184.220 ;
        RECT 116.655 184.050 116.825 184.560 ;
        RECT 116.995 184.380 117.205 184.950 ;
        RECT 117.375 184.910 117.955 185.120 ;
        RECT 118.135 185.395 119.525 185.410 ;
        RECT 119.695 185.545 120.705 185.715 ;
        RECT 121.275 185.695 121.445 186.015 ;
        RECT 122.355 185.865 122.635 186.255 ;
        RECT 122.805 185.975 122.975 186.425 ;
        RECT 123.145 186.145 124.165 186.460 ;
        RECT 124.335 186.190 125.345 186.515 ;
        RECT 123.995 186.020 124.165 186.145 ;
        RECT 118.135 185.080 118.725 185.395 ;
        RECT 117.375 184.585 118.385 184.910 ;
        RECT 116.190 183.720 116.825 184.050 ;
        RECT 116.995 183.565 117.205 184.210 ;
        RECT 118.555 184.110 118.725 185.080 ;
        RECT 117.455 183.780 118.725 184.110 ;
        RECT 118.555 183.395 118.725 183.780 ;
        RECT 118.945 183.570 119.235 185.225 ;
        RECT 119.695 185.160 119.865 185.545 ;
        RECT 119.405 184.990 119.865 185.160 ;
        RECT 119.405 183.890 119.575 184.990 ;
        RECT 120.035 184.970 120.365 185.375 ;
        RECT 120.535 185.145 120.705 185.545 ;
        RECT 120.875 185.505 121.445 185.695 ;
        RECT 121.615 185.675 122.185 185.845 ;
        RECT 122.805 185.805 123.825 185.975 ;
        RECT 120.875 185.315 121.845 185.505 ;
        RECT 120.535 184.975 121.055 185.145 ;
        RECT 121.275 185.085 121.845 185.315 ;
        RECT 119.745 184.090 120.365 184.800 ;
        RECT 120.535 184.275 120.705 184.975 ;
        RECT 121.275 184.805 121.445 185.085 ;
        RECT 122.015 184.915 122.185 185.675 ;
        RECT 122.355 185.635 122.685 185.680 ;
        RECT 122.355 185.435 123.485 185.635 ;
        RECT 122.355 184.985 123.485 185.235 ;
        RECT 120.875 184.475 121.445 184.805 ;
        RECT 121.615 184.685 122.185 184.915 ;
        RECT 123.655 184.795 123.825 185.805 ;
        RECT 120.535 184.105 121.055 184.275 ;
        RECT 119.405 183.570 119.865 183.890 ;
        RECT 120.035 183.570 120.605 183.920 ;
        RECT 121.275 183.905 121.445 184.475 ;
        RECT 121.615 184.195 122.185 184.515 ;
        RECT 122.355 184.365 122.685 184.770 ;
        RECT 122.855 184.545 123.825 184.795 ;
        RECT 123.995 185.690 124.585 186.020 ;
        RECT 124.765 185.980 125.345 186.190 ;
        RECT 125.515 186.150 125.725 186.720 ;
        RECT 125.895 186.540 126.065 187.050 ;
        RECT 126.715 186.880 126.885 188.145 ;
        RECT 127.860 188.055 128.190 188.160 ;
        RECT 128.675 188.145 130.695 188.475 ;
        RECT 130.865 189.355 132.325 189.375 ;
        RECT 130.865 189.115 133.135 189.355 ;
        RECT 130.865 188.445 132.325 189.115 ;
        RECT 133.315 189.025 133.565 189.375 ;
        RECT 133.735 189.035 134.690 189.365 ;
        RECT 132.495 188.855 133.135 188.945 ;
        RECT 133.735 188.855 133.905 189.035 ;
        RECT 132.495 188.685 133.905 188.855 ;
        RECT 134.875 188.710 135.045 189.555 ;
        RECT 135.645 189.510 136.225 189.720 ;
        RECT 137.595 189.635 138.375 189.805 ;
        RECT 135.215 189.185 136.225 189.510 ;
        RECT 136.395 188.980 136.605 189.550 ;
        RECT 136.775 189.160 137.425 189.490 ;
        RECT 132.495 188.615 133.135 188.685 ;
        RECT 130.865 188.175 133.135 188.445 ;
        RECT 130.865 188.165 132.325 188.175 ;
        RECT 133.315 188.165 133.565 188.515 ;
        RECT 134.875 188.505 136.145 188.710 ;
        RECT 133.735 188.380 136.145 188.505 ;
        RECT 133.735 188.175 135.045 188.380 ;
        RECT 129.435 187.995 130.695 188.145 ;
        RECT 127.055 187.885 127.560 187.965 ;
        RECT 128.360 187.885 129.265 187.975 ;
        RECT 127.055 187.705 129.265 187.885 ;
        RECT 127.070 187.050 127.705 187.380 ;
        RECT 126.245 186.710 127.355 186.880 ;
        RECT 125.895 186.210 126.545 186.540 ;
        RECT 124.765 185.810 126.545 185.980 ;
        RECT 123.995 184.945 124.165 185.690 ;
        RECT 122.855 184.195 123.025 184.545 ;
        RECT 123.995 184.535 124.595 184.945 ;
        RECT 124.765 184.800 124.935 185.810 ;
        RECT 125.105 185.470 126.145 185.640 ;
        RECT 125.105 185.015 125.275 185.470 ;
        RECT 125.475 184.970 125.805 185.300 ;
        RECT 125.975 185.270 126.145 185.470 ;
        RECT 125.975 185.100 126.350 185.270 ;
        RECT 126.715 184.820 126.885 186.710 ;
        RECT 127.535 186.540 127.705 187.050 ;
        RECT 127.875 186.890 128.085 187.535 ;
        RECT 129.435 187.320 131.215 187.995 ;
        RECT 128.335 186.990 131.215 187.320 ;
        RECT 129.435 186.785 131.215 186.990 ;
        RECT 131.385 186.910 132.325 188.165 ;
        RECT 132.690 187.280 134.705 187.535 ;
        RECT 132.690 187.175 133.065 187.280 ;
        RECT 133.720 187.195 134.705 187.280 ;
        RECT 134.875 187.485 135.045 188.175 ;
        RECT 136.395 188.165 136.605 188.810 ;
        RECT 136.775 188.650 136.945 189.160 ;
        RECT 137.595 188.990 137.765 189.635 ;
        RECT 137.985 189.310 138.505 189.465 ;
        RECT 138.675 189.425 139.005 189.975 ;
        RECT 140.315 189.815 140.485 190.555 ;
        RECT 139.305 189.645 140.485 189.815 ;
        RECT 137.985 189.255 138.545 189.310 ;
        RECT 139.175 189.300 140.100 189.475 ;
        RECT 139.125 189.255 140.100 189.300 ;
        RECT 137.985 189.145 140.100 189.255 ;
        RECT 137.985 189.135 139.255 189.145 ;
        RECT 138.420 189.085 139.255 189.135 ;
        RECT 137.125 188.820 137.765 188.990 ;
        RECT 136.775 188.320 137.410 188.650 ;
        RECT 137.595 188.290 137.765 188.820 ;
        RECT 140.315 188.965 140.485 189.645 ;
        RECT 140.655 190.405 141.675 190.575 ;
        RECT 141.845 190.465 142.125 190.855 ;
        RECT 142.295 190.750 143.205 191.065 ;
        RECT 145.755 190.750 145.925 191.845 ;
        RECT 142.295 190.615 144.045 190.750 ;
        RECT 143.035 190.490 144.045 190.615 ;
        RECT 144.605 190.490 145.925 190.750 ;
        RECT 140.655 189.395 140.825 190.405 ;
        RECT 141.795 190.235 142.125 190.280 ;
        RECT 140.995 190.035 142.125 190.235 ;
        RECT 142.295 190.275 142.865 190.445 ;
        RECT 140.995 189.585 142.125 189.835 ;
        RECT 142.295 189.515 142.465 190.275 ;
        RECT 143.035 190.105 143.205 190.490 ;
        RECT 142.635 189.890 143.205 190.105 ;
        RECT 143.375 190.145 145.585 190.315 ;
        RECT 143.375 190.060 143.950 190.145 ;
        RECT 144.680 190.060 145.585 190.145 ;
        RECT 144.115 189.890 144.445 189.975 ;
        RECT 145.755 189.890 145.925 190.490 ;
        RECT 142.635 189.685 143.585 189.890 ;
        RECT 143.035 189.560 143.585 189.685 ;
        RECT 143.755 189.720 144.825 189.890 ;
        RECT 140.655 189.145 141.625 189.395 ;
        RECT 140.315 188.635 141.285 188.965 ;
        RECT 141.455 188.795 141.625 189.145 ;
        RECT 141.795 188.965 142.125 189.370 ;
        RECT 142.295 189.285 142.865 189.515 ;
        RECT 142.295 188.795 142.865 189.115 ;
        RECT 137.595 188.050 138.275 188.290 ;
        RECT 135.215 187.740 137.230 187.995 ;
        RECT 135.215 187.655 136.200 187.740 ;
        RECT 136.855 187.635 137.230 187.740 ;
        RECT 136.355 187.485 136.685 187.570 ;
        RECT 133.235 187.025 133.565 187.110 ;
        RECT 134.875 187.075 135.475 187.485 ;
        RECT 135.645 187.220 136.685 187.485 ;
        RECT 137.595 187.370 137.765 188.050 ;
        RECT 138.445 188.040 139.005 188.395 ;
        RECT 139.175 187.880 139.520 188.270 ;
        RECT 140.315 187.885 140.485 188.635 ;
        RECT 141.455 188.625 142.865 188.795 ;
        RECT 143.035 188.915 143.205 189.560 ;
        RECT 143.755 189.345 143.925 189.720 ;
        RECT 143.375 189.175 143.925 189.345 ;
        RECT 144.105 189.085 144.475 189.440 ;
        RECT 144.655 189.345 144.825 189.720 ;
        RECT 144.995 189.560 145.925 189.890 ;
        RECT 144.655 189.175 145.585 189.345 ;
        RECT 145.755 188.915 145.925 189.560 ;
        RECT 140.655 188.055 141.335 188.340 ;
        RECT 139.175 187.870 139.345 187.880 ;
        RECT 137.945 187.700 139.345 187.870 ;
        RECT 137.945 187.590 138.275 187.700 ;
        RECT 136.855 187.360 137.765 187.370 ;
        RECT 134.875 187.025 135.045 187.075 ;
        RECT 131.385 186.785 133.065 186.910 ;
        RECT 127.055 186.210 127.705 186.540 ;
        RECT 127.875 186.150 128.085 186.720 ;
        RECT 128.255 186.190 129.265 186.515 ;
        RECT 128.255 185.980 128.835 186.190 ;
        RECT 129.435 186.145 129.605 186.785 ;
        RECT 132.155 186.740 133.065 186.785 ;
        RECT 133.235 186.760 134.275 187.025 ;
        RECT 129.435 186.020 130.745 186.145 ;
        RECT 127.055 185.810 128.835 185.980 ;
        RECT 127.455 185.470 128.495 185.640 ;
        RECT 127.455 185.270 127.625 185.470 ;
        RECT 127.250 185.100 127.625 185.270 ;
        RECT 127.795 184.970 128.125 185.300 ;
        RECT 128.325 185.015 128.495 185.470 ;
        RECT 124.765 184.535 125.805 184.800 ;
        RECT 125.975 184.650 127.625 184.820 ;
        RECT 128.665 184.800 128.835 185.810 ;
        RECT 129.015 185.815 130.745 186.020 ;
        RECT 129.015 185.690 129.605 185.815 ;
        RECT 130.915 185.805 131.165 186.155 ;
        RECT 132.155 186.145 132.325 186.740 ;
        RECT 132.690 186.290 133.065 186.460 ;
        RECT 131.345 185.875 132.325 186.145 ;
        RECT 132.895 186.090 133.065 186.290 ;
        RECT 133.235 186.260 133.565 186.590 ;
        RECT 133.765 186.090 133.935 186.545 ;
        RECT 132.895 185.920 133.935 186.090 ;
        RECT 129.435 184.945 129.605 185.690 ;
        RECT 131.345 185.635 131.985 185.705 ;
        RECT 130.575 185.465 131.985 185.635 ;
        RECT 130.575 185.285 130.745 185.465 ;
        RECT 131.345 185.375 131.985 185.465 ;
        RECT 129.790 184.955 130.745 185.285 ;
        RECT 130.915 184.945 131.165 185.295 ;
        RECT 132.155 185.205 132.325 185.875 ;
        RECT 134.105 185.750 134.275 186.760 ;
        RECT 134.445 186.615 135.045 187.025 ;
        RECT 134.875 186.330 135.045 186.615 ;
        RECT 134.875 186.000 135.465 186.330 ;
        RECT 135.645 186.210 135.815 187.220 ;
        RECT 136.855 187.200 138.275 187.360 ;
        RECT 138.445 187.265 139.005 187.530 ;
        RECT 137.595 187.145 138.275 187.200 ;
        RECT 135.985 186.550 136.155 187.005 ;
        RECT 136.355 186.720 136.685 187.050 ;
        RECT 136.855 186.750 137.230 186.920 ;
        RECT 136.855 186.550 137.025 186.750 ;
        RECT 135.985 186.380 137.025 186.550 ;
        RECT 135.645 186.040 137.425 186.210 ;
        RECT 134.875 185.870 135.045 186.000 ;
        RECT 132.495 185.580 134.275 185.750 ;
        RECT 131.345 184.965 132.325 185.205 ;
        RECT 132.495 185.020 133.145 185.350 ;
        RECT 123.995 184.365 124.165 184.535 ;
        RECT 125.475 184.450 125.805 184.535 ;
        RECT 121.615 184.025 123.025 184.195 ;
        RECT 123.195 184.035 124.165 184.365 ;
        RECT 120.775 183.575 121.445 183.905 ;
        RECT 121.275 183.395 121.445 183.575 ;
        RECT 123.995 183.395 124.165 184.035 ;
        RECT 124.335 184.280 125.320 184.365 ;
        RECT 125.975 184.280 126.350 184.385 ;
        RECT 124.335 184.255 126.350 184.280 ;
        RECT 124.335 184.085 126.375 184.255 ;
        RECT 124.335 184.025 126.350 184.085 ;
        RECT 126.715 183.395 126.885 184.650 ;
        RECT 127.795 184.535 128.835 184.800 ;
        RECT 129.005 184.535 129.605 184.945 ;
        RECT 132.155 184.850 132.325 184.965 ;
        RECT 127.795 184.450 128.125 184.535 ;
        RECT 127.250 184.280 127.625 184.385 ;
        RECT 128.280 184.280 129.265 184.365 ;
        RECT 127.250 184.025 129.265 184.280 ;
        RECT 129.435 184.335 129.605 184.535 ;
        RECT 129.775 184.605 131.985 184.775 ;
        RECT 129.775 184.505 130.680 184.605 ;
        RECT 131.480 184.515 131.985 184.605 ;
        RECT 132.155 184.680 132.795 184.850 ;
        RECT 129.435 184.005 130.365 184.335 ;
        RECT 130.850 184.320 131.180 184.435 ;
        RECT 132.155 184.335 132.325 184.680 ;
        RECT 132.975 184.510 133.145 185.020 ;
        RECT 133.315 184.840 133.525 185.410 ;
        RECT 133.695 185.370 134.275 185.580 ;
        RECT 134.455 185.540 135.045 185.870 ;
        RECT 135.645 185.830 136.225 186.040 ;
        RECT 133.695 185.045 134.705 185.370 ;
        RECT 134.875 185.030 135.045 185.540 ;
        RECT 135.215 185.505 136.225 185.830 ;
        RECT 136.395 185.300 136.605 185.870 ;
        RECT 136.775 185.480 137.425 185.810 ;
        RECT 137.595 185.715 137.765 187.145 ;
        RECT 139.175 187.015 139.345 187.700 ;
        RECT 140.315 187.615 140.945 187.885 ;
        RECT 140.315 187.395 140.485 187.615 ;
        RECT 139.515 187.065 140.485 187.395 ;
        RECT 141.115 187.595 141.335 188.055 ;
        RECT 141.505 187.765 142.065 188.455 ;
        RECT 143.035 188.395 144.495 188.915 ;
        RECT 142.235 188.055 142.865 188.340 ;
        RECT 142.235 187.595 142.405 188.055 ;
        RECT 143.035 187.885 143.955 188.395 ;
        RECT 144.665 188.225 145.925 188.915 ;
        RECT 142.575 187.705 143.955 187.885 ;
        RECT 144.125 187.705 145.925 188.225 ;
        RECT 142.575 187.615 143.205 187.705 ;
        RECT 141.115 187.385 142.405 187.595 ;
        RECT 137.935 186.675 138.505 186.975 ;
        RECT 138.675 186.845 139.345 187.015 ;
        RECT 139.525 186.675 140.145 186.895 ;
        RECT 137.935 186.360 140.145 186.675 ;
        RECT 137.935 185.895 138.485 186.065 ;
        RECT 134.875 184.700 136.145 185.030 ;
        RECT 130.535 184.150 131.605 184.320 ;
        RECT 129.435 183.395 129.605 184.005 ;
        RECT 130.535 183.825 130.705 184.150 ;
        RECT 129.775 183.655 130.705 183.825 ;
        RECT 130.885 183.585 131.255 183.915 ;
        RECT 131.435 183.825 131.605 184.150 ;
        RECT 131.775 184.005 132.325 184.335 ;
        RECT 132.510 184.180 133.145 184.510 ;
        RECT 133.315 184.025 133.525 184.670 ;
        RECT 134.875 184.570 135.045 184.700 ;
        RECT 133.775 184.240 135.045 184.570 ;
        RECT 136.395 184.485 136.605 185.130 ;
        RECT 136.775 184.970 136.945 185.480 ;
        RECT 137.595 185.385 138.145 185.715 ;
        RECT 138.315 185.570 138.485 185.895 ;
        RECT 138.665 185.805 139.035 186.135 ;
        RECT 139.215 185.895 140.145 186.065 ;
        RECT 139.215 185.570 139.385 185.895 ;
        RECT 140.315 185.825 140.485 187.065 ;
        RECT 140.655 186.815 142.865 187.215 ;
        RECT 143.035 187.095 143.205 187.615 ;
        RECT 143.375 187.365 145.585 187.535 ;
        RECT 143.375 187.275 143.880 187.365 ;
        RECT 144.680 187.265 145.585 187.365 ;
        RECT 140.655 186.345 141.335 186.625 ;
        RECT 141.115 185.950 141.335 186.345 ;
        RECT 141.505 186.120 142.065 186.815 ;
        RECT 143.035 186.765 143.585 187.095 ;
        RECT 144.180 187.080 144.510 187.195 ;
        RECT 145.755 187.095 145.925 187.705 ;
        RECT 143.755 186.910 144.825 187.080 ;
        RECT 142.235 186.345 142.865 186.625 ;
        RECT 142.235 185.950 142.405 186.345 ;
        RECT 140.315 185.715 140.945 185.825 ;
        RECT 138.315 185.400 139.385 185.570 ;
        RECT 139.555 185.500 140.945 185.715 ;
        RECT 141.115 185.500 142.405 185.950 ;
        RECT 143.035 185.825 143.205 186.765 ;
        RECT 143.755 186.585 143.925 186.910 ;
        RECT 143.375 186.415 143.925 186.585 ;
        RECT 144.105 186.345 144.475 186.675 ;
        RECT 144.655 186.585 144.825 186.910 ;
        RECT 144.995 186.765 145.925 187.095 ;
        RECT 144.655 186.415 145.585 186.585 ;
        RECT 143.375 185.985 145.585 186.155 ;
        RECT 143.375 185.895 143.880 185.985 ;
        RECT 144.680 185.885 145.585 185.985 ;
        RECT 142.575 185.715 143.205 185.825 ;
        RECT 142.575 185.500 143.585 185.715 ;
        RECT 144.180 185.700 144.510 185.815 ;
        RECT 145.755 185.715 145.925 186.765 ;
        RECT 137.595 185.310 137.765 185.385 ;
        RECT 137.125 185.140 137.765 185.310 ;
        RECT 138.740 185.285 139.070 185.400 ;
        RECT 139.555 185.385 140.485 185.500 ;
        RECT 141.795 185.395 142.125 185.500 ;
        RECT 136.775 184.640 137.410 184.970 ;
        RECT 131.435 183.655 131.985 183.825 ;
        RECT 132.155 183.395 132.325 184.005 ;
        RECT 134.875 183.395 135.045 184.240 ;
        RECT 137.595 184.335 137.765 185.140 ;
        RECT 137.935 185.115 138.440 185.205 ;
        RECT 139.240 185.115 140.145 185.215 ;
        RECT 137.935 184.945 140.145 185.115 ;
        RECT 137.935 184.595 140.145 184.775 ;
        RECT 137.935 184.515 138.440 184.595 ;
        RECT 139.240 184.505 140.145 184.595 ;
        RECT 137.595 184.005 138.145 184.335 ;
        RECT 138.740 184.320 139.070 184.425 ;
        RECT 140.315 184.335 140.485 185.385 ;
        RECT 143.035 185.385 143.585 185.500 ;
        RECT 143.755 185.530 144.825 185.700 ;
        RECT 140.655 185.225 141.625 185.330 ;
        RECT 142.295 185.225 142.865 185.330 ;
        RECT 140.655 184.945 142.865 185.225 ;
        RECT 140.655 184.595 142.865 184.775 ;
        RECT 140.655 184.505 141.560 184.595 ;
        RECT 142.360 184.515 142.865 184.595 ;
        RECT 138.315 184.150 139.385 184.320 ;
        RECT 137.595 183.395 137.765 184.005 ;
        RECT 138.315 183.825 138.485 184.150 ;
        RECT 137.935 183.655 138.485 183.825 ;
        RECT 138.665 183.585 139.035 183.925 ;
        RECT 139.215 183.825 139.385 184.150 ;
        RECT 139.555 184.005 141.245 184.335 ;
        RECT 141.730 184.320 142.060 184.425 ;
        RECT 143.035 184.335 143.205 185.385 ;
        RECT 143.755 185.205 143.925 185.530 ;
        RECT 143.375 185.035 143.925 185.205 ;
        RECT 144.105 184.965 144.475 185.295 ;
        RECT 144.655 185.205 144.825 185.530 ;
        RECT 144.995 185.385 145.925 185.715 ;
        RECT 144.655 185.035 145.585 185.205 ;
        RECT 143.375 184.595 145.585 184.775 ;
        RECT 143.375 184.515 143.880 184.595 ;
        RECT 144.680 184.505 145.585 184.595 ;
        RECT 141.415 184.150 142.485 184.320 ;
        RECT 139.215 183.645 140.145 183.825 ;
        RECT 140.315 183.395 140.485 184.005 ;
        RECT 141.415 183.825 141.585 184.150 ;
        RECT 140.655 183.645 141.585 183.825 ;
        RECT 141.765 183.585 142.135 183.925 ;
        RECT 142.315 183.825 142.485 184.150 ;
        RECT 142.655 184.005 143.585 184.335 ;
        RECT 144.180 184.320 144.510 184.425 ;
        RECT 145.755 184.335 145.925 185.385 ;
        RECT 143.755 184.150 144.825 184.320 ;
        RECT 142.315 183.655 142.865 183.825 ;
        RECT 143.035 183.395 143.205 184.005 ;
        RECT 143.755 183.825 143.925 184.150 ;
        RECT 143.375 183.655 143.925 183.825 ;
        RECT 144.105 183.585 144.475 183.925 ;
        RECT 144.655 183.825 144.825 184.150 ;
        RECT 144.995 184.005 145.925 184.335 ;
        RECT 144.655 183.645 145.585 183.825 ;
        RECT 145.755 183.395 145.925 184.005 ;
        RECT 110.395 182.705 111.315 183.395 ;
        RECT 111.485 182.875 114.915 183.395 ;
        RECT 110.395 182.185 111.855 182.705 ;
        RECT 112.025 182.185 114.375 182.875 ;
        RECT 115.085 182.705 116.755 183.395 ;
        RECT 116.925 182.875 120.355 183.395 ;
        RECT 114.545 182.185 117.295 182.705 ;
        RECT 117.465 182.185 119.815 182.875 ;
        RECT 120.525 182.705 122.195 183.395 ;
        RECT 122.365 182.875 125.795 183.395 ;
        RECT 119.985 182.185 122.735 182.705 ;
        RECT 122.905 182.185 125.255 182.875 ;
        RECT 125.965 182.705 127.635 183.395 ;
        RECT 127.805 182.875 131.235 183.395 ;
        RECT 125.425 182.185 128.175 182.705 ;
        RECT 128.345 182.185 130.695 182.875 ;
        RECT 131.405 182.705 133.075 183.395 ;
        RECT 133.245 182.875 136.675 183.395 ;
        RECT 130.865 182.185 133.615 182.705 ;
        RECT 133.785 182.185 136.135 182.875 ;
        RECT 136.845 182.705 138.515 183.395 ;
        RECT 138.685 182.875 142.115 183.395 ;
        RECT 136.305 182.185 139.055 182.705 ;
        RECT 139.225 182.185 141.575 182.875 ;
        RECT 142.285 182.705 143.955 183.395 ;
        RECT 144.125 182.875 145.925 183.395 ;
        RECT 141.745 182.185 144.495 182.705 ;
        RECT 144.665 182.185 145.925 182.875 ;
        RECT 110.395 182.100 110.565 182.185 ;
        RECT 113.115 182.100 113.285 182.185 ;
        RECT 115.835 182.100 116.005 182.185 ;
        RECT 118.555 182.100 118.725 182.185 ;
        RECT 121.275 182.100 121.445 182.185 ;
        RECT 123.995 182.100 124.165 182.185 ;
        RECT 126.715 182.100 126.885 182.185 ;
        RECT 129.435 182.100 129.605 182.185 ;
        RECT 132.155 182.100 132.325 182.185 ;
        RECT 134.875 182.100 135.045 182.185 ;
        RECT 137.595 182.100 137.765 182.185 ;
        RECT 140.315 182.100 140.485 182.185 ;
        RECT 143.035 182.100 143.205 182.185 ;
        RECT 145.755 182.100 145.925 182.185 ;
        RECT 138.940 173.340 144.680 173.350 ;
        RECT 119.990 173.300 125.730 173.310 ;
        RECT 100.950 173.270 106.690 173.280 ;
        RECT 100.460 173.110 106.690 173.270 ;
        RECT 100.460 170.850 101.130 173.110 ;
        RECT 101.800 172.540 105.840 172.710 ;
        RECT 101.460 171.480 101.630 172.480 ;
        RECT 106.010 171.480 106.180 172.480 ;
        RECT 101.800 171.250 105.840 171.420 ;
        RECT 106.520 170.850 106.690 173.110 ;
        RECT 100.460 170.680 106.690 170.850 ;
        RECT 100.460 167.420 101.130 170.680 ;
        RECT 101.800 170.110 105.840 170.280 ;
        RECT 101.460 168.050 101.630 170.050 ;
        RECT 106.010 168.050 106.180 170.050 ;
        RECT 101.800 167.820 105.840 167.990 ;
        RECT 106.520 167.420 106.690 170.680 ;
        RECT 100.460 167.250 106.690 167.420 ;
        RECT 100.460 163.990 101.130 167.250 ;
        RECT 101.800 166.680 105.840 166.850 ;
        RECT 101.460 164.620 101.630 166.620 ;
        RECT 106.010 164.620 106.180 166.620 ;
        RECT 101.800 164.390 105.840 164.560 ;
        RECT 106.520 163.990 106.690 167.250 ;
        RECT 100.460 163.980 106.690 163.990 ;
        RECT 108.280 173.250 118.110 173.290 ;
        RECT 108.280 173.120 118.910 173.250 ;
        RECT 108.280 170.860 108.450 173.120 ;
        RECT 109.175 172.550 117.215 172.720 ;
        RECT 108.790 171.490 108.960 172.490 ;
        RECT 117.430 171.490 117.600 172.490 ;
        RECT 109.175 171.260 117.215 171.430 ;
        RECT 117.940 170.860 118.910 173.120 ;
        RECT 108.280 170.690 118.910 170.860 ;
        RECT 108.280 167.430 108.450 170.690 ;
        RECT 109.175 170.120 117.215 170.290 ;
        RECT 108.790 168.060 108.960 170.060 ;
        RECT 117.430 168.060 117.600 170.060 ;
        RECT 109.175 167.830 117.215 168.000 ;
        RECT 117.940 167.430 118.910 170.690 ;
        RECT 108.280 167.260 118.910 167.430 ;
        RECT 108.280 164.000 108.450 167.260 ;
        RECT 109.175 166.690 117.215 166.860 ;
        RECT 108.790 164.630 108.960 166.630 ;
        RECT 117.430 164.630 117.600 166.630 ;
        RECT 109.175 164.400 117.215 164.570 ;
        RECT 117.940 164.000 118.910 167.260 ;
        RECT 100.460 163.880 106.700 163.980 ;
        RECT 100.450 163.320 106.700 163.880 ;
        RECT 100.450 163.300 105.620 163.320 ;
        RECT 100.450 163.230 104.440 163.300 ;
        RECT 100.450 161.960 102.370 163.230 ;
        RECT 103.880 163.220 104.440 163.230 ;
        RECT 104.110 162.130 104.440 163.220 ;
        RECT 104.810 162.750 105.850 162.920 ;
        RECT 104.810 162.310 105.850 162.480 ;
        RECT 106.020 162.450 106.190 162.780 ;
        RECT 104.270 161.910 104.440 162.130 ;
        RECT 106.530 161.910 106.700 163.320 ;
        RECT 104.270 161.740 106.700 161.910 ;
        RECT 108.280 163.830 118.910 164.000 ;
        RECT 119.500 173.140 125.730 173.300 ;
        RECT 119.500 170.880 120.170 173.140 ;
        RECT 120.840 172.570 124.880 172.740 ;
        RECT 120.500 171.510 120.670 172.510 ;
        RECT 125.050 171.510 125.220 172.510 ;
        RECT 120.840 171.280 124.880 171.450 ;
        RECT 125.560 170.880 125.730 173.140 ;
        RECT 119.500 170.710 125.730 170.880 ;
        RECT 119.500 167.450 120.170 170.710 ;
        RECT 120.840 170.140 124.880 170.310 ;
        RECT 120.500 168.080 120.670 170.080 ;
        RECT 125.050 168.080 125.220 170.080 ;
        RECT 120.840 167.850 124.880 168.020 ;
        RECT 125.560 167.450 125.730 170.710 ;
        RECT 119.500 167.280 125.730 167.450 ;
        RECT 119.500 164.020 120.170 167.280 ;
        RECT 120.840 166.710 124.880 166.880 ;
        RECT 120.500 164.650 120.670 166.650 ;
        RECT 125.050 164.650 125.220 166.650 ;
        RECT 120.840 164.420 124.880 164.590 ;
        RECT 125.560 164.020 125.730 167.280 ;
        RECT 119.500 164.010 125.730 164.020 ;
        RECT 127.320 173.280 137.150 173.320 ;
        RECT 127.320 173.150 137.950 173.280 ;
        RECT 127.320 170.890 127.490 173.150 ;
        RECT 128.215 172.580 136.255 172.750 ;
        RECT 127.830 171.520 128.000 172.520 ;
        RECT 136.470 171.520 136.640 172.520 ;
        RECT 128.215 171.290 136.255 171.460 ;
        RECT 136.980 170.890 137.950 173.150 ;
        RECT 127.320 170.720 137.950 170.890 ;
        RECT 127.320 167.460 127.490 170.720 ;
        RECT 128.215 170.150 136.255 170.320 ;
        RECT 127.830 168.090 128.000 170.090 ;
        RECT 136.470 168.090 136.640 170.090 ;
        RECT 128.215 167.860 136.255 168.030 ;
        RECT 136.980 167.460 137.950 170.720 ;
        RECT 127.320 167.290 137.950 167.460 ;
        RECT 127.320 164.030 127.490 167.290 ;
        RECT 128.215 166.720 136.255 166.890 ;
        RECT 127.830 164.660 128.000 166.660 ;
        RECT 136.470 164.660 136.640 166.660 ;
        RECT 128.215 164.430 136.255 164.600 ;
        RECT 136.980 164.030 137.950 167.290 ;
        RECT 119.500 163.910 125.740 164.010 ;
        RECT 108.280 161.570 108.450 163.830 ;
        RECT 109.175 163.260 117.215 163.430 ;
        RECT 108.790 162.200 108.960 163.200 ;
        RECT 117.430 162.200 117.600 163.200 ;
        RECT 109.175 161.970 117.215 162.140 ;
        RECT 117.940 161.570 118.910 163.830 ;
        RECT 119.490 163.350 125.740 163.910 ;
        RECT 119.490 163.330 124.660 163.350 ;
        RECT 119.490 163.260 123.480 163.330 ;
        RECT 119.490 161.990 121.410 163.260 ;
        RECT 122.920 163.250 123.480 163.260 ;
        RECT 123.150 162.160 123.480 163.250 ;
        RECT 123.850 162.780 124.890 162.950 ;
        RECT 123.850 162.340 124.890 162.510 ;
        RECT 125.060 162.480 125.230 162.810 ;
        RECT 123.310 161.940 123.480 162.160 ;
        RECT 125.570 161.940 125.740 163.350 ;
        RECT 123.310 161.770 125.740 161.940 ;
        RECT 127.320 163.860 137.950 164.030 ;
        RECT 138.450 173.180 144.680 173.340 ;
        RECT 138.450 170.920 139.120 173.180 ;
        RECT 139.790 172.610 143.830 172.780 ;
        RECT 139.450 171.550 139.620 172.550 ;
        RECT 144.000 171.550 144.170 172.550 ;
        RECT 139.790 171.320 143.830 171.490 ;
        RECT 144.510 170.920 144.680 173.180 ;
        RECT 138.450 170.750 144.680 170.920 ;
        RECT 138.450 167.490 139.120 170.750 ;
        RECT 139.790 170.180 143.830 170.350 ;
        RECT 139.450 168.120 139.620 170.120 ;
        RECT 144.000 168.120 144.170 170.120 ;
        RECT 139.790 167.890 143.830 168.060 ;
        RECT 144.510 167.490 144.680 170.750 ;
        RECT 138.450 167.320 144.680 167.490 ;
        RECT 138.450 164.060 139.120 167.320 ;
        RECT 139.790 166.750 143.830 166.920 ;
        RECT 139.450 164.690 139.620 166.690 ;
        RECT 144.000 164.690 144.170 166.690 ;
        RECT 139.790 164.460 143.830 164.630 ;
        RECT 144.510 164.060 144.680 167.320 ;
        RECT 138.450 164.050 144.680 164.060 ;
        RECT 146.270 173.320 156.100 173.360 ;
        RECT 146.270 173.190 156.900 173.320 ;
        RECT 146.270 170.930 146.440 173.190 ;
        RECT 147.165 172.620 155.205 172.790 ;
        RECT 146.780 171.560 146.950 172.560 ;
        RECT 155.420 171.560 155.590 172.560 ;
        RECT 147.165 171.330 155.205 171.500 ;
        RECT 155.930 170.930 156.900 173.190 ;
        RECT 146.270 170.760 156.900 170.930 ;
        RECT 146.270 167.500 146.440 170.760 ;
        RECT 147.165 170.190 155.205 170.360 ;
        RECT 146.780 168.130 146.950 170.130 ;
        RECT 155.420 168.130 155.590 170.130 ;
        RECT 147.165 167.900 155.205 168.070 ;
        RECT 155.930 167.500 156.900 170.760 ;
        RECT 146.270 167.330 156.900 167.500 ;
        RECT 146.270 164.070 146.440 167.330 ;
        RECT 147.165 166.760 155.205 166.930 ;
        RECT 146.780 164.700 146.950 166.700 ;
        RECT 155.420 164.700 155.590 166.700 ;
        RECT 147.165 164.470 155.205 164.640 ;
        RECT 155.930 164.070 156.900 167.330 ;
        RECT 138.450 163.950 144.690 164.050 ;
        RECT 127.320 161.600 127.490 163.860 ;
        RECT 128.215 163.290 136.255 163.460 ;
        RECT 127.830 162.230 128.000 163.230 ;
        RECT 136.470 162.230 136.640 163.230 ;
        RECT 128.215 162.000 136.255 162.170 ;
        RECT 136.980 161.600 137.950 163.860 ;
        RECT 138.440 163.390 144.690 163.950 ;
        RECT 138.440 163.370 143.610 163.390 ;
        RECT 138.440 163.300 142.430 163.370 ;
        RECT 138.440 162.030 140.360 163.300 ;
        RECT 141.870 163.290 142.430 163.300 ;
        RECT 142.100 162.200 142.430 163.290 ;
        RECT 142.800 162.820 143.840 162.990 ;
        RECT 142.800 162.380 143.840 162.550 ;
        RECT 144.010 162.520 144.180 162.850 ;
        RECT 142.260 161.980 142.430 162.200 ;
        RECT 144.520 161.980 144.690 163.390 ;
        RECT 142.260 161.810 144.690 161.980 ;
        RECT 146.270 163.900 156.900 164.070 ;
        RECT 146.270 161.640 146.440 163.900 ;
        RECT 147.165 163.330 155.205 163.500 ;
        RECT 146.780 162.270 146.950 163.270 ;
        RECT 155.420 162.270 155.590 163.270 ;
        RECT 147.165 162.040 155.205 162.210 ;
        RECT 155.930 161.640 156.900 163.900 ;
        RECT 146.270 161.610 156.900 161.640 ;
        RECT 127.320 161.570 137.950 161.600 ;
        RECT 108.280 161.540 118.910 161.570 ;
        RECT 108.250 161.430 118.910 161.540 ;
        RECT 127.290 161.460 137.950 161.570 ;
        RECT 146.240 161.500 156.900 161.610 ;
        RECT 106.500 161.380 118.910 161.430 ;
        RECT 125.540 161.410 137.950 161.460 ;
        RECT 144.490 161.450 156.900 161.500 ;
        RECT 102.160 161.210 118.910 161.380 ;
        RECT 102.160 159.800 102.330 161.210 ;
        RECT 102.700 160.640 105.740 160.810 ;
        RECT 102.700 160.200 105.740 160.370 ;
        RECT 105.955 160.340 106.125 160.670 ;
        RECT 106.460 160.450 118.910 161.210 ;
        RECT 121.200 161.240 137.950 161.410 ;
        RECT 106.460 160.440 118.800 160.450 ;
        RECT 106.460 160.430 112.340 160.440 ;
        RECT 106.460 160.410 107.030 160.430 ;
        RECT 108.250 160.420 112.340 160.430 ;
        RECT 106.470 159.800 106.640 160.410 ;
        RECT 102.160 159.630 106.640 159.800 ;
        RECT 121.200 159.830 121.370 161.240 ;
        RECT 121.740 160.670 124.780 160.840 ;
        RECT 121.740 160.230 124.780 160.400 ;
        RECT 124.995 160.370 125.165 160.700 ;
        RECT 125.500 160.480 137.950 161.240 ;
        RECT 140.150 161.280 156.900 161.450 ;
        RECT 125.500 160.470 137.840 160.480 ;
        RECT 125.500 160.460 131.380 160.470 ;
        RECT 125.500 160.440 126.070 160.460 ;
        RECT 127.290 160.450 131.380 160.460 ;
        RECT 125.510 159.830 125.680 160.440 ;
        RECT 121.200 159.660 125.680 159.830 ;
        RECT 140.150 159.870 140.320 161.280 ;
        RECT 140.690 160.710 143.730 160.880 ;
        RECT 140.690 160.270 143.730 160.440 ;
        RECT 143.945 160.410 144.115 160.740 ;
        RECT 144.450 160.520 156.900 161.280 ;
        RECT 144.450 160.510 156.790 160.520 ;
        RECT 144.450 160.500 150.330 160.510 ;
        RECT 144.450 160.480 145.020 160.500 ;
        RECT 146.240 160.490 150.330 160.500 ;
        RECT 144.460 159.870 144.630 160.480 ;
        RECT 140.150 159.700 144.630 159.870 ;
        RECT 100.950 158.280 106.690 158.290 ;
        RECT 100.460 158.120 106.690 158.280 ;
        RECT 100.460 155.860 101.130 158.120 ;
        RECT 101.800 157.550 105.840 157.720 ;
        RECT 101.460 156.490 101.630 157.490 ;
        RECT 106.010 156.490 106.180 157.490 ;
        RECT 101.800 156.260 105.840 156.430 ;
        RECT 106.520 155.860 106.690 158.120 ;
        RECT 100.460 155.690 106.690 155.860 ;
        RECT 100.460 152.430 101.130 155.690 ;
        RECT 101.800 155.120 105.840 155.290 ;
        RECT 101.460 153.060 101.630 155.060 ;
        RECT 106.010 153.060 106.180 155.060 ;
        RECT 101.800 152.830 105.840 153.000 ;
        RECT 106.520 152.430 106.690 155.690 ;
        RECT 100.460 152.260 106.690 152.430 ;
        RECT 100.460 149.000 101.130 152.260 ;
        RECT 101.800 151.690 105.840 151.860 ;
        RECT 101.460 149.630 101.630 151.630 ;
        RECT 106.010 149.630 106.180 151.630 ;
        RECT 101.800 149.400 105.840 149.570 ;
        RECT 106.520 149.000 106.690 152.260 ;
        RECT 100.460 148.990 106.690 149.000 ;
        RECT 108.280 158.260 118.110 158.300 ;
        RECT 119.990 158.280 125.730 158.290 ;
        RECT 108.280 158.130 118.910 158.260 ;
        RECT 108.280 155.870 108.450 158.130 ;
        RECT 109.175 157.560 117.215 157.730 ;
        RECT 108.790 156.500 108.960 157.500 ;
        RECT 117.430 156.500 117.600 157.500 ;
        RECT 109.175 156.270 117.215 156.440 ;
        RECT 117.940 155.870 118.910 158.130 ;
        RECT 108.280 155.700 118.910 155.870 ;
        RECT 108.280 152.440 108.450 155.700 ;
        RECT 109.175 155.130 117.215 155.300 ;
        RECT 108.790 153.070 108.960 155.070 ;
        RECT 117.430 153.070 117.600 155.070 ;
        RECT 109.175 152.840 117.215 153.010 ;
        RECT 117.940 152.440 118.910 155.700 ;
        RECT 108.280 152.270 118.910 152.440 ;
        RECT 108.280 149.010 108.450 152.270 ;
        RECT 109.175 151.700 117.215 151.870 ;
        RECT 108.790 149.640 108.960 151.640 ;
        RECT 117.430 149.640 117.600 151.640 ;
        RECT 109.175 149.410 117.215 149.580 ;
        RECT 117.940 149.010 118.910 152.270 ;
        RECT 100.460 148.890 106.700 148.990 ;
        RECT 100.450 148.330 106.700 148.890 ;
        RECT 100.450 148.310 105.620 148.330 ;
        RECT 100.450 148.240 104.440 148.310 ;
        RECT 100.450 146.970 102.370 148.240 ;
        RECT 103.880 148.230 104.440 148.240 ;
        RECT 104.110 147.140 104.440 148.230 ;
        RECT 104.810 147.760 105.850 147.930 ;
        RECT 104.810 147.320 105.850 147.490 ;
        RECT 106.020 147.460 106.190 147.790 ;
        RECT 104.270 146.920 104.440 147.140 ;
        RECT 106.530 146.920 106.700 148.330 ;
        RECT 104.270 146.750 106.700 146.920 ;
        RECT 108.280 148.840 118.910 149.010 ;
        RECT 119.500 158.120 125.730 158.280 ;
        RECT 119.500 155.860 120.170 158.120 ;
        RECT 120.840 157.550 124.880 157.720 ;
        RECT 120.500 156.490 120.670 157.490 ;
        RECT 125.050 156.490 125.220 157.490 ;
        RECT 120.840 156.260 124.880 156.430 ;
        RECT 125.560 155.860 125.730 158.120 ;
        RECT 119.500 155.690 125.730 155.860 ;
        RECT 119.500 152.430 120.170 155.690 ;
        RECT 120.840 155.120 124.880 155.290 ;
        RECT 120.500 153.060 120.670 155.060 ;
        RECT 125.050 153.060 125.220 155.060 ;
        RECT 120.840 152.830 124.880 153.000 ;
        RECT 125.560 152.430 125.730 155.690 ;
        RECT 119.500 152.260 125.730 152.430 ;
        RECT 119.500 149.000 120.170 152.260 ;
        RECT 120.840 151.690 124.880 151.860 ;
        RECT 120.500 149.630 120.670 151.630 ;
        RECT 125.050 149.630 125.220 151.630 ;
        RECT 120.840 149.400 124.880 149.570 ;
        RECT 125.560 149.000 125.730 152.260 ;
        RECT 119.500 148.990 125.730 149.000 ;
        RECT 127.320 158.260 137.150 158.300 ;
        RECT 138.990 158.280 144.730 158.290 ;
        RECT 127.320 158.130 137.950 158.260 ;
        RECT 127.320 155.870 127.490 158.130 ;
        RECT 128.215 157.560 136.255 157.730 ;
        RECT 127.830 156.500 128.000 157.500 ;
        RECT 136.470 156.500 136.640 157.500 ;
        RECT 128.215 156.270 136.255 156.440 ;
        RECT 136.980 155.870 137.950 158.130 ;
        RECT 127.320 155.700 137.950 155.870 ;
        RECT 127.320 152.440 127.490 155.700 ;
        RECT 128.215 155.130 136.255 155.300 ;
        RECT 127.830 153.070 128.000 155.070 ;
        RECT 136.470 153.070 136.640 155.070 ;
        RECT 128.215 152.840 136.255 153.010 ;
        RECT 136.980 152.440 137.950 155.700 ;
        RECT 127.320 152.270 137.950 152.440 ;
        RECT 127.320 149.010 127.490 152.270 ;
        RECT 128.215 151.700 136.255 151.870 ;
        RECT 127.830 149.640 128.000 151.640 ;
        RECT 136.470 149.640 136.640 151.640 ;
        RECT 128.215 149.410 136.255 149.580 ;
        RECT 136.980 149.010 137.950 152.270 ;
        RECT 119.500 148.890 125.740 148.990 ;
        RECT 108.280 146.580 108.450 148.840 ;
        RECT 109.175 148.270 117.215 148.440 ;
        RECT 108.790 147.210 108.960 148.210 ;
        RECT 117.430 147.210 117.600 148.210 ;
        RECT 109.175 146.980 117.215 147.150 ;
        RECT 117.940 146.580 118.910 148.840 ;
        RECT 119.490 148.330 125.740 148.890 ;
        RECT 119.490 148.310 124.660 148.330 ;
        RECT 119.490 148.240 123.480 148.310 ;
        RECT 119.490 146.970 121.410 148.240 ;
        RECT 122.920 148.230 123.480 148.240 ;
        RECT 123.150 147.140 123.480 148.230 ;
        RECT 123.850 147.760 124.890 147.930 ;
        RECT 123.850 147.320 124.890 147.490 ;
        RECT 125.060 147.460 125.230 147.790 ;
        RECT 123.310 146.920 123.480 147.140 ;
        RECT 125.570 146.920 125.740 148.330 ;
        RECT 123.310 146.750 125.740 146.920 ;
        RECT 127.320 148.840 137.950 149.010 ;
        RECT 138.500 158.120 144.730 158.280 ;
        RECT 138.500 155.860 139.170 158.120 ;
        RECT 139.840 157.550 143.880 157.720 ;
        RECT 139.500 156.490 139.670 157.490 ;
        RECT 144.050 156.490 144.220 157.490 ;
        RECT 139.840 156.260 143.880 156.430 ;
        RECT 144.560 155.860 144.730 158.120 ;
        RECT 138.500 155.690 144.730 155.860 ;
        RECT 138.500 152.430 139.170 155.690 ;
        RECT 139.840 155.120 143.880 155.290 ;
        RECT 139.500 153.060 139.670 155.060 ;
        RECT 144.050 153.060 144.220 155.060 ;
        RECT 139.840 152.830 143.880 153.000 ;
        RECT 144.560 152.430 144.730 155.690 ;
        RECT 138.500 152.260 144.730 152.430 ;
        RECT 138.500 149.000 139.170 152.260 ;
        RECT 139.840 151.690 143.880 151.860 ;
        RECT 139.500 149.630 139.670 151.630 ;
        RECT 144.050 149.630 144.220 151.630 ;
        RECT 139.840 149.400 143.880 149.570 ;
        RECT 144.560 149.000 144.730 152.260 ;
        RECT 138.500 148.990 144.730 149.000 ;
        RECT 146.320 158.260 156.150 158.300 ;
        RECT 146.320 158.130 156.950 158.260 ;
        RECT 146.320 155.870 146.490 158.130 ;
        RECT 147.215 157.560 155.255 157.730 ;
        RECT 146.830 156.500 147.000 157.500 ;
        RECT 155.470 156.500 155.640 157.500 ;
        RECT 147.215 156.270 155.255 156.440 ;
        RECT 155.980 155.870 156.950 158.130 ;
        RECT 146.320 155.700 156.950 155.870 ;
        RECT 146.320 152.440 146.490 155.700 ;
        RECT 147.215 155.130 155.255 155.300 ;
        RECT 146.830 153.070 147.000 155.070 ;
        RECT 155.470 153.070 155.640 155.070 ;
        RECT 147.215 152.840 155.255 153.010 ;
        RECT 155.980 152.440 156.950 155.700 ;
        RECT 146.320 152.270 156.950 152.440 ;
        RECT 146.320 149.010 146.490 152.270 ;
        RECT 147.215 151.700 155.255 151.870 ;
        RECT 146.830 149.640 147.000 151.640 ;
        RECT 155.470 149.640 155.640 151.640 ;
        RECT 147.215 149.410 155.255 149.580 ;
        RECT 155.980 149.010 156.950 152.270 ;
        RECT 138.500 148.890 144.740 148.990 ;
        RECT 108.280 146.550 118.910 146.580 ;
        RECT 127.320 146.580 127.490 148.840 ;
        RECT 128.215 148.270 136.255 148.440 ;
        RECT 127.830 147.210 128.000 148.210 ;
        RECT 136.470 147.210 136.640 148.210 ;
        RECT 128.215 146.980 136.255 147.150 ;
        RECT 136.980 146.580 137.950 148.840 ;
        RECT 138.490 148.330 144.740 148.890 ;
        RECT 138.490 148.310 143.660 148.330 ;
        RECT 138.490 148.240 142.480 148.310 ;
        RECT 138.490 146.970 140.410 148.240 ;
        RECT 141.920 148.230 142.480 148.240 ;
        RECT 142.150 147.140 142.480 148.230 ;
        RECT 142.850 147.760 143.890 147.930 ;
        RECT 142.850 147.320 143.890 147.490 ;
        RECT 144.060 147.460 144.230 147.790 ;
        RECT 142.310 146.920 142.480 147.140 ;
        RECT 144.570 146.920 144.740 148.330 ;
        RECT 142.310 146.750 144.740 146.920 ;
        RECT 146.320 148.840 156.950 149.010 ;
        RECT 127.320 146.550 137.950 146.580 ;
        RECT 146.320 146.580 146.490 148.840 ;
        RECT 147.215 148.270 155.255 148.440 ;
        RECT 146.830 147.210 147.000 148.210 ;
        RECT 155.470 147.210 155.640 148.210 ;
        RECT 147.215 146.980 155.255 147.150 ;
        RECT 155.980 146.580 156.950 148.840 ;
        RECT 146.320 146.550 156.950 146.580 ;
        RECT 108.250 146.440 118.910 146.550 ;
        RECT 127.290 146.440 137.950 146.550 ;
        RECT 146.290 146.440 156.950 146.550 ;
        RECT 106.500 146.390 118.910 146.440 ;
        RECT 125.540 146.390 137.950 146.440 ;
        RECT 144.540 146.390 156.950 146.440 ;
        RECT 102.160 146.220 118.910 146.390 ;
        RECT 102.160 144.810 102.330 146.220 ;
        RECT 102.700 145.650 105.740 145.820 ;
        RECT 102.700 145.210 105.740 145.380 ;
        RECT 105.955 145.350 106.125 145.680 ;
        RECT 106.460 145.460 118.910 146.220 ;
        RECT 121.200 146.220 137.950 146.390 ;
        RECT 106.460 145.450 118.800 145.460 ;
        RECT 106.460 145.440 112.340 145.450 ;
        RECT 106.460 145.420 107.030 145.440 ;
        RECT 108.250 145.430 112.340 145.440 ;
        RECT 106.470 144.810 106.640 145.420 ;
        RECT 102.160 144.640 106.640 144.810 ;
        RECT 121.200 144.810 121.370 146.220 ;
        RECT 121.740 145.650 124.780 145.820 ;
        RECT 121.740 145.210 124.780 145.380 ;
        RECT 124.995 145.350 125.165 145.680 ;
        RECT 125.500 145.460 137.950 146.220 ;
        RECT 140.200 146.220 156.950 146.390 ;
        RECT 125.500 145.450 137.840 145.460 ;
        RECT 125.500 145.440 131.380 145.450 ;
        RECT 125.500 145.420 126.070 145.440 ;
        RECT 127.290 145.430 131.380 145.440 ;
        RECT 125.510 144.810 125.680 145.420 ;
        RECT 121.200 144.640 125.680 144.810 ;
        RECT 140.200 144.810 140.370 146.220 ;
        RECT 140.740 145.650 143.780 145.820 ;
        RECT 140.740 145.210 143.780 145.380 ;
        RECT 143.995 145.350 144.165 145.680 ;
        RECT 144.500 145.460 156.950 146.220 ;
        RECT 144.500 145.450 156.840 145.460 ;
        RECT 144.500 145.440 150.380 145.450 ;
        RECT 144.500 145.420 145.070 145.440 ;
        RECT 146.290 145.430 150.380 145.440 ;
        RECT 144.510 144.810 144.680 145.420 ;
        RECT 140.200 144.640 144.680 144.810 ;
        RECT 100.950 143.300 106.690 143.310 ;
        RECT 100.460 143.140 106.690 143.300 ;
        RECT 100.460 140.880 101.130 143.140 ;
        RECT 101.800 142.570 105.840 142.740 ;
        RECT 101.460 141.510 101.630 142.510 ;
        RECT 106.010 141.510 106.180 142.510 ;
        RECT 101.800 141.280 105.840 141.450 ;
        RECT 106.520 140.880 106.690 143.140 ;
        RECT 100.460 140.710 106.690 140.880 ;
        RECT 100.460 137.450 101.130 140.710 ;
        RECT 101.800 140.140 105.840 140.310 ;
        RECT 101.460 138.080 101.630 140.080 ;
        RECT 106.010 138.080 106.180 140.080 ;
        RECT 101.800 137.850 105.840 138.020 ;
        RECT 106.520 137.450 106.690 140.710 ;
        RECT 100.460 137.280 106.690 137.450 ;
        RECT 100.460 134.020 101.130 137.280 ;
        RECT 101.800 136.710 105.840 136.880 ;
        RECT 101.460 134.650 101.630 136.650 ;
        RECT 106.010 134.650 106.180 136.650 ;
        RECT 101.800 134.420 105.840 134.590 ;
        RECT 106.520 134.020 106.690 137.280 ;
        RECT 100.460 134.010 106.690 134.020 ;
        RECT 108.280 143.280 118.110 143.320 ;
        RECT 108.280 143.150 118.910 143.280 ;
        RECT 119.940 143.260 125.680 143.270 ;
        RECT 108.280 140.890 108.450 143.150 ;
        RECT 109.175 142.580 117.215 142.750 ;
        RECT 108.790 141.520 108.960 142.520 ;
        RECT 117.430 141.520 117.600 142.520 ;
        RECT 109.175 141.290 117.215 141.460 ;
        RECT 117.940 140.890 118.910 143.150 ;
        RECT 108.280 140.720 118.910 140.890 ;
        RECT 108.280 137.460 108.450 140.720 ;
        RECT 109.175 140.150 117.215 140.320 ;
        RECT 108.790 138.090 108.960 140.090 ;
        RECT 117.430 138.090 117.600 140.090 ;
        RECT 109.175 137.860 117.215 138.030 ;
        RECT 117.940 137.460 118.910 140.720 ;
        RECT 108.280 137.290 118.910 137.460 ;
        RECT 108.280 134.030 108.450 137.290 ;
        RECT 109.175 136.720 117.215 136.890 ;
        RECT 108.790 134.660 108.960 136.660 ;
        RECT 117.430 134.660 117.600 136.660 ;
        RECT 109.175 134.430 117.215 134.600 ;
        RECT 117.940 134.030 118.910 137.290 ;
        RECT 100.460 133.910 106.700 134.010 ;
        RECT 100.450 133.350 106.700 133.910 ;
        RECT 100.450 133.330 105.620 133.350 ;
        RECT 100.450 133.260 104.440 133.330 ;
        RECT 100.450 131.990 102.370 133.260 ;
        RECT 103.880 133.250 104.440 133.260 ;
        RECT 104.110 132.160 104.440 133.250 ;
        RECT 104.810 132.780 105.850 132.950 ;
        RECT 104.810 132.340 105.850 132.510 ;
        RECT 106.020 132.480 106.190 132.810 ;
        RECT 104.270 131.940 104.440 132.160 ;
        RECT 106.530 131.940 106.700 133.350 ;
        RECT 104.270 131.770 106.700 131.940 ;
        RECT 108.280 133.860 118.910 134.030 ;
        RECT 119.450 143.100 125.680 143.260 ;
        RECT 119.450 140.840 120.120 143.100 ;
        RECT 120.790 142.530 124.830 142.700 ;
        RECT 120.450 141.470 120.620 142.470 ;
        RECT 125.000 141.470 125.170 142.470 ;
        RECT 120.790 141.240 124.830 141.410 ;
        RECT 125.510 140.840 125.680 143.100 ;
        RECT 119.450 140.670 125.680 140.840 ;
        RECT 119.450 137.410 120.120 140.670 ;
        RECT 120.790 140.100 124.830 140.270 ;
        RECT 120.450 138.040 120.620 140.040 ;
        RECT 125.000 138.040 125.170 140.040 ;
        RECT 120.790 137.810 124.830 137.980 ;
        RECT 125.510 137.410 125.680 140.670 ;
        RECT 119.450 137.240 125.680 137.410 ;
        RECT 119.450 133.980 120.120 137.240 ;
        RECT 120.790 136.670 124.830 136.840 ;
        RECT 120.450 134.610 120.620 136.610 ;
        RECT 125.000 134.610 125.170 136.610 ;
        RECT 120.790 134.380 124.830 134.550 ;
        RECT 125.510 133.980 125.680 137.240 ;
        RECT 119.450 133.970 125.680 133.980 ;
        RECT 127.270 143.240 137.100 143.280 ;
        RECT 138.940 143.260 144.680 143.270 ;
        RECT 127.270 143.110 137.900 143.240 ;
        RECT 127.270 140.850 127.440 143.110 ;
        RECT 128.165 142.540 136.205 142.710 ;
        RECT 127.780 141.480 127.950 142.480 ;
        RECT 136.420 141.480 136.590 142.480 ;
        RECT 128.165 141.250 136.205 141.420 ;
        RECT 136.930 140.850 137.900 143.110 ;
        RECT 127.270 140.680 137.900 140.850 ;
        RECT 127.270 137.420 127.440 140.680 ;
        RECT 128.165 140.110 136.205 140.280 ;
        RECT 127.780 138.050 127.950 140.050 ;
        RECT 136.420 138.050 136.590 140.050 ;
        RECT 128.165 137.820 136.205 137.990 ;
        RECT 136.930 137.420 137.900 140.680 ;
        RECT 127.270 137.250 137.900 137.420 ;
        RECT 127.270 133.990 127.440 137.250 ;
        RECT 128.165 136.680 136.205 136.850 ;
        RECT 127.780 134.620 127.950 136.620 ;
        RECT 136.420 134.620 136.590 136.620 ;
        RECT 128.165 134.390 136.205 134.560 ;
        RECT 136.930 133.990 137.900 137.250 ;
        RECT 119.450 133.870 125.690 133.970 ;
        RECT 108.280 131.600 108.450 133.860 ;
        RECT 109.175 133.290 117.215 133.460 ;
        RECT 108.790 132.230 108.960 133.230 ;
        RECT 117.430 132.230 117.600 133.230 ;
        RECT 109.175 132.000 117.215 132.170 ;
        RECT 117.940 131.600 118.910 133.860 ;
        RECT 119.440 133.310 125.690 133.870 ;
        RECT 119.440 133.290 124.610 133.310 ;
        RECT 119.440 133.220 123.430 133.290 ;
        RECT 119.440 131.950 121.360 133.220 ;
        RECT 122.870 133.210 123.430 133.220 ;
        RECT 123.100 132.120 123.430 133.210 ;
        RECT 123.800 132.740 124.840 132.910 ;
        RECT 123.800 132.300 124.840 132.470 ;
        RECT 125.010 132.440 125.180 132.770 ;
        RECT 123.260 131.900 123.430 132.120 ;
        RECT 125.520 131.900 125.690 133.310 ;
        RECT 123.260 131.730 125.690 131.900 ;
        RECT 127.270 133.820 137.900 133.990 ;
        RECT 138.450 143.100 144.680 143.260 ;
        RECT 138.450 140.840 139.120 143.100 ;
        RECT 139.790 142.530 143.830 142.700 ;
        RECT 139.450 141.470 139.620 142.470 ;
        RECT 144.000 141.470 144.170 142.470 ;
        RECT 139.790 141.240 143.830 141.410 ;
        RECT 144.510 140.840 144.680 143.100 ;
        RECT 138.450 140.670 144.680 140.840 ;
        RECT 138.450 137.410 139.120 140.670 ;
        RECT 139.790 140.100 143.830 140.270 ;
        RECT 139.450 138.040 139.620 140.040 ;
        RECT 144.000 138.040 144.170 140.040 ;
        RECT 139.790 137.810 143.830 137.980 ;
        RECT 144.510 137.410 144.680 140.670 ;
        RECT 138.450 137.240 144.680 137.410 ;
        RECT 138.450 133.980 139.120 137.240 ;
        RECT 139.790 136.670 143.830 136.840 ;
        RECT 139.450 134.610 139.620 136.610 ;
        RECT 144.000 134.610 144.170 136.610 ;
        RECT 139.790 134.380 143.830 134.550 ;
        RECT 144.510 133.980 144.680 137.240 ;
        RECT 138.450 133.970 144.680 133.980 ;
        RECT 146.270 143.240 156.100 143.280 ;
        RECT 146.270 143.110 156.900 143.240 ;
        RECT 146.270 140.850 146.440 143.110 ;
        RECT 147.165 142.540 155.205 142.710 ;
        RECT 146.780 141.480 146.950 142.480 ;
        RECT 155.420 141.480 155.590 142.480 ;
        RECT 147.165 141.250 155.205 141.420 ;
        RECT 155.930 140.850 156.900 143.110 ;
        RECT 146.270 140.680 156.900 140.850 ;
        RECT 146.270 137.420 146.440 140.680 ;
        RECT 147.165 140.110 155.205 140.280 ;
        RECT 146.780 138.050 146.950 140.050 ;
        RECT 155.420 138.050 155.590 140.050 ;
        RECT 147.165 137.820 155.205 137.990 ;
        RECT 155.930 137.420 156.900 140.680 ;
        RECT 146.270 137.250 156.900 137.420 ;
        RECT 146.270 133.990 146.440 137.250 ;
        RECT 147.165 136.680 155.205 136.850 ;
        RECT 146.780 134.620 146.950 136.620 ;
        RECT 155.420 134.620 155.590 136.620 ;
        RECT 147.165 134.390 155.205 134.560 ;
        RECT 155.930 133.990 156.900 137.250 ;
        RECT 138.450 133.870 144.690 133.970 ;
        RECT 108.280 131.570 118.910 131.600 ;
        RECT 108.250 131.460 118.910 131.570 ;
        RECT 127.270 131.560 127.440 133.820 ;
        RECT 128.165 133.250 136.205 133.420 ;
        RECT 127.780 132.190 127.950 133.190 ;
        RECT 136.420 132.190 136.590 133.190 ;
        RECT 128.165 131.960 136.205 132.130 ;
        RECT 136.930 131.560 137.900 133.820 ;
        RECT 138.440 133.310 144.690 133.870 ;
        RECT 138.440 133.290 143.610 133.310 ;
        RECT 138.440 133.220 142.430 133.290 ;
        RECT 138.440 131.950 140.360 133.220 ;
        RECT 141.870 133.210 142.430 133.220 ;
        RECT 142.100 132.120 142.430 133.210 ;
        RECT 142.800 132.740 143.840 132.910 ;
        RECT 142.800 132.300 143.840 132.470 ;
        RECT 144.010 132.440 144.180 132.770 ;
        RECT 142.260 131.900 142.430 132.120 ;
        RECT 144.520 131.900 144.690 133.310 ;
        RECT 142.260 131.730 144.690 131.900 ;
        RECT 146.270 133.820 156.900 133.990 ;
        RECT 127.270 131.530 137.900 131.560 ;
        RECT 146.270 131.560 146.440 133.820 ;
        RECT 147.165 133.250 155.205 133.420 ;
        RECT 146.780 132.190 146.950 133.190 ;
        RECT 155.420 132.190 155.590 133.190 ;
        RECT 147.165 131.960 155.205 132.130 ;
        RECT 155.930 131.560 156.900 133.820 ;
        RECT 146.270 131.530 156.900 131.560 ;
        RECT 106.500 131.410 118.910 131.460 ;
        RECT 127.240 131.420 137.900 131.530 ;
        RECT 146.240 131.420 156.900 131.530 ;
        RECT 102.160 131.240 118.910 131.410 ;
        RECT 125.490 131.370 137.900 131.420 ;
        RECT 144.490 131.370 156.900 131.420 ;
        RECT 102.160 129.830 102.330 131.240 ;
        RECT 102.700 130.670 105.740 130.840 ;
        RECT 102.700 130.230 105.740 130.400 ;
        RECT 105.955 130.370 106.125 130.700 ;
        RECT 106.460 130.480 118.910 131.240 ;
        RECT 121.150 131.200 137.900 131.370 ;
        RECT 106.460 130.470 118.800 130.480 ;
        RECT 106.460 130.460 112.340 130.470 ;
        RECT 106.460 130.440 107.030 130.460 ;
        RECT 108.250 130.450 112.340 130.460 ;
        RECT 106.470 129.830 106.640 130.440 ;
        RECT 102.160 129.660 106.640 129.830 ;
        RECT 121.150 129.790 121.320 131.200 ;
        RECT 121.690 130.630 124.730 130.800 ;
        RECT 121.690 130.190 124.730 130.360 ;
        RECT 124.945 130.330 125.115 130.660 ;
        RECT 125.450 130.440 137.900 131.200 ;
        RECT 140.150 131.200 156.900 131.370 ;
        RECT 125.450 130.430 137.790 130.440 ;
        RECT 125.450 130.420 131.330 130.430 ;
        RECT 125.450 130.400 126.020 130.420 ;
        RECT 127.240 130.410 131.330 130.420 ;
        RECT 125.460 129.790 125.630 130.400 ;
        RECT 121.150 129.620 125.630 129.790 ;
        RECT 140.150 129.790 140.320 131.200 ;
        RECT 140.690 130.630 143.730 130.800 ;
        RECT 140.690 130.190 143.730 130.360 ;
        RECT 143.945 130.330 144.115 130.660 ;
        RECT 144.450 130.440 156.900 131.200 ;
        RECT 144.450 130.430 156.790 130.440 ;
        RECT 144.450 130.420 150.330 130.430 ;
        RECT 144.450 130.400 145.020 130.420 ;
        RECT 146.240 130.410 150.330 130.420 ;
        RECT 144.460 129.790 144.630 130.400 ;
        RECT 140.150 129.620 144.630 129.790 ;
        RECT 100.950 128.270 106.690 128.280 ;
        RECT 100.460 128.110 106.690 128.270 ;
        RECT 100.460 125.850 101.130 128.110 ;
        RECT 101.800 127.540 105.840 127.710 ;
        RECT 101.460 126.480 101.630 127.480 ;
        RECT 106.010 126.480 106.180 127.480 ;
        RECT 101.800 126.250 105.840 126.420 ;
        RECT 106.520 125.850 106.690 128.110 ;
        RECT 100.460 125.680 106.690 125.850 ;
        RECT 100.460 122.420 101.130 125.680 ;
        RECT 101.800 125.110 105.840 125.280 ;
        RECT 101.460 123.050 101.630 125.050 ;
        RECT 106.010 123.050 106.180 125.050 ;
        RECT 101.800 122.820 105.840 122.990 ;
        RECT 106.520 122.420 106.690 125.680 ;
        RECT 100.460 122.250 106.690 122.420 ;
        RECT 100.460 118.990 101.130 122.250 ;
        RECT 101.800 121.680 105.840 121.850 ;
        RECT 101.460 119.620 101.630 121.620 ;
        RECT 106.010 119.620 106.180 121.620 ;
        RECT 101.800 119.390 105.840 119.560 ;
        RECT 106.520 118.990 106.690 122.250 ;
        RECT 100.460 118.980 106.690 118.990 ;
        RECT 108.280 128.250 118.110 128.290 ;
        RECT 108.280 128.120 118.910 128.250 ;
        RECT 119.940 128.240 125.680 128.250 ;
        RECT 108.280 125.860 108.450 128.120 ;
        RECT 109.175 127.550 117.215 127.720 ;
        RECT 108.790 126.490 108.960 127.490 ;
        RECT 117.430 126.490 117.600 127.490 ;
        RECT 109.175 126.260 117.215 126.430 ;
        RECT 117.940 125.860 118.910 128.120 ;
        RECT 108.280 125.690 118.910 125.860 ;
        RECT 108.280 122.430 108.450 125.690 ;
        RECT 109.175 125.120 117.215 125.290 ;
        RECT 108.790 123.060 108.960 125.060 ;
        RECT 117.430 123.060 117.600 125.060 ;
        RECT 109.175 122.830 117.215 123.000 ;
        RECT 117.940 122.430 118.910 125.690 ;
        RECT 108.280 122.260 118.910 122.430 ;
        RECT 108.280 119.000 108.450 122.260 ;
        RECT 109.175 121.690 117.215 121.860 ;
        RECT 108.790 119.630 108.960 121.630 ;
        RECT 117.430 119.630 117.600 121.630 ;
        RECT 109.175 119.400 117.215 119.570 ;
        RECT 117.940 119.000 118.910 122.260 ;
        RECT 100.460 118.880 106.700 118.980 ;
        RECT 100.450 118.320 106.700 118.880 ;
        RECT 100.450 118.300 105.620 118.320 ;
        RECT 100.450 118.230 104.440 118.300 ;
        RECT 100.450 116.960 102.370 118.230 ;
        RECT 103.880 118.220 104.440 118.230 ;
        RECT 104.110 117.130 104.440 118.220 ;
        RECT 104.810 117.750 105.850 117.920 ;
        RECT 104.810 117.310 105.850 117.480 ;
        RECT 106.020 117.450 106.190 117.780 ;
        RECT 104.270 116.910 104.440 117.130 ;
        RECT 106.530 116.910 106.700 118.320 ;
        RECT 104.270 116.740 106.700 116.910 ;
        RECT 108.280 118.830 118.910 119.000 ;
        RECT 119.450 128.080 125.680 128.240 ;
        RECT 119.450 125.820 120.120 128.080 ;
        RECT 120.790 127.510 124.830 127.680 ;
        RECT 120.450 126.450 120.620 127.450 ;
        RECT 125.000 126.450 125.170 127.450 ;
        RECT 120.790 126.220 124.830 126.390 ;
        RECT 125.510 125.820 125.680 128.080 ;
        RECT 119.450 125.650 125.680 125.820 ;
        RECT 119.450 122.390 120.120 125.650 ;
        RECT 120.790 125.080 124.830 125.250 ;
        RECT 120.450 123.020 120.620 125.020 ;
        RECT 125.000 123.020 125.170 125.020 ;
        RECT 120.790 122.790 124.830 122.960 ;
        RECT 125.510 122.390 125.680 125.650 ;
        RECT 119.450 122.220 125.680 122.390 ;
        RECT 119.450 118.960 120.120 122.220 ;
        RECT 120.790 121.650 124.830 121.820 ;
        RECT 120.450 119.590 120.620 121.590 ;
        RECT 125.000 119.590 125.170 121.590 ;
        RECT 120.790 119.360 124.830 119.530 ;
        RECT 125.510 118.960 125.680 122.220 ;
        RECT 119.450 118.950 125.680 118.960 ;
        RECT 127.270 128.220 137.100 128.260 ;
        RECT 138.940 128.240 144.680 128.250 ;
        RECT 127.270 128.090 137.900 128.220 ;
        RECT 127.270 125.830 127.440 128.090 ;
        RECT 128.165 127.520 136.205 127.690 ;
        RECT 127.780 126.460 127.950 127.460 ;
        RECT 136.420 126.460 136.590 127.460 ;
        RECT 128.165 126.230 136.205 126.400 ;
        RECT 136.930 125.830 137.900 128.090 ;
        RECT 127.270 125.660 137.900 125.830 ;
        RECT 127.270 122.400 127.440 125.660 ;
        RECT 128.165 125.090 136.205 125.260 ;
        RECT 127.780 123.030 127.950 125.030 ;
        RECT 136.420 123.030 136.590 125.030 ;
        RECT 128.165 122.800 136.205 122.970 ;
        RECT 136.930 122.400 137.900 125.660 ;
        RECT 127.270 122.230 137.900 122.400 ;
        RECT 127.270 118.970 127.440 122.230 ;
        RECT 128.165 121.660 136.205 121.830 ;
        RECT 127.780 119.600 127.950 121.600 ;
        RECT 136.420 119.600 136.590 121.600 ;
        RECT 128.165 119.370 136.205 119.540 ;
        RECT 136.930 118.970 137.900 122.230 ;
        RECT 119.450 118.850 125.690 118.950 ;
        RECT 108.280 116.570 108.450 118.830 ;
        RECT 109.175 118.260 117.215 118.430 ;
        RECT 108.790 117.200 108.960 118.200 ;
        RECT 117.430 117.200 117.600 118.200 ;
        RECT 109.175 116.970 117.215 117.140 ;
        RECT 117.940 116.570 118.910 118.830 ;
        RECT 119.440 118.290 125.690 118.850 ;
        RECT 119.440 118.270 124.610 118.290 ;
        RECT 119.440 118.200 123.430 118.270 ;
        RECT 119.440 116.930 121.360 118.200 ;
        RECT 122.870 118.190 123.430 118.200 ;
        RECT 123.100 117.100 123.430 118.190 ;
        RECT 123.800 117.720 124.840 117.890 ;
        RECT 123.800 117.280 124.840 117.450 ;
        RECT 125.010 117.420 125.180 117.750 ;
        RECT 123.260 116.880 123.430 117.100 ;
        RECT 125.520 116.880 125.690 118.290 ;
        RECT 123.260 116.710 125.690 116.880 ;
        RECT 127.270 118.800 137.900 118.970 ;
        RECT 138.450 128.080 144.680 128.240 ;
        RECT 138.450 125.820 139.120 128.080 ;
        RECT 139.790 127.510 143.830 127.680 ;
        RECT 139.450 126.450 139.620 127.450 ;
        RECT 144.000 126.450 144.170 127.450 ;
        RECT 139.790 126.220 143.830 126.390 ;
        RECT 144.510 125.820 144.680 128.080 ;
        RECT 138.450 125.650 144.680 125.820 ;
        RECT 138.450 122.390 139.120 125.650 ;
        RECT 139.790 125.080 143.830 125.250 ;
        RECT 139.450 123.020 139.620 125.020 ;
        RECT 144.000 123.020 144.170 125.020 ;
        RECT 139.790 122.790 143.830 122.960 ;
        RECT 144.510 122.390 144.680 125.650 ;
        RECT 138.450 122.220 144.680 122.390 ;
        RECT 138.450 118.960 139.120 122.220 ;
        RECT 139.790 121.650 143.830 121.820 ;
        RECT 139.450 119.590 139.620 121.590 ;
        RECT 144.000 119.590 144.170 121.590 ;
        RECT 139.790 119.360 143.830 119.530 ;
        RECT 144.510 118.960 144.680 122.220 ;
        RECT 138.450 118.950 144.680 118.960 ;
        RECT 146.270 128.220 156.100 128.260 ;
        RECT 146.270 128.090 156.900 128.220 ;
        RECT 146.270 125.830 146.440 128.090 ;
        RECT 147.165 127.520 155.205 127.690 ;
        RECT 146.780 126.460 146.950 127.460 ;
        RECT 155.420 126.460 155.590 127.460 ;
        RECT 147.165 126.230 155.205 126.400 ;
        RECT 155.930 125.830 156.900 128.090 ;
        RECT 146.270 125.660 156.900 125.830 ;
        RECT 146.270 122.400 146.440 125.660 ;
        RECT 147.165 125.090 155.205 125.260 ;
        RECT 146.780 123.030 146.950 125.030 ;
        RECT 155.420 123.030 155.590 125.030 ;
        RECT 147.165 122.800 155.205 122.970 ;
        RECT 155.930 122.400 156.900 125.660 ;
        RECT 146.270 122.230 156.900 122.400 ;
        RECT 146.270 118.970 146.440 122.230 ;
        RECT 147.165 121.660 155.205 121.830 ;
        RECT 146.780 119.600 146.950 121.600 ;
        RECT 155.420 119.600 155.590 121.600 ;
        RECT 147.165 119.370 155.205 119.540 ;
        RECT 155.930 118.970 156.900 122.230 ;
        RECT 138.450 118.850 144.690 118.950 ;
        RECT 108.280 116.540 118.910 116.570 ;
        RECT 108.250 116.430 118.910 116.540 ;
        RECT 127.270 116.540 127.440 118.800 ;
        RECT 128.165 118.230 136.205 118.400 ;
        RECT 127.780 117.170 127.950 118.170 ;
        RECT 136.420 117.170 136.590 118.170 ;
        RECT 128.165 116.940 136.205 117.110 ;
        RECT 136.930 116.540 137.900 118.800 ;
        RECT 138.440 118.290 144.690 118.850 ;
        RECT 138.440 118.270 143.610 118.290 ;
        RECT 138.440 118.200 142.430 118.270 ;
        RECT 138.440 116.930 140.360 118.200 ;
        RECT 141.870 118.190 142.430 118.200 ;
        RECT 142.100 117.100 142.430 118.190 ;
        RECT 142.800 117.720 143.840 117.890 ;
        RECT 142.800 117.280 143.840 117.450 ;
        RECT 144.010 117.420 144.180 117.750 ;
        RECT 142.260 116.880 142.430 117.100 ;
        RECT 144.520 116.880 144.690 118.290 ;
        RECT 142.260 116.710 144.690 116.880 ;
        RECT 146.270 118.800 156.900 118.970 ;
        RECT 127.270 116.510 137.900 116.540 ;
        RECT 146.270 116.540 146.440 118.800 ;
        RECT 147.165 118.230 155.205 118.400 ;
        RECT 146.780 117.170 146.950 118.170 ;
        RECT 155.420 117.170 155.590 118.170 ;
        RECT 147.165 116.940 155.205 117.110 ;
        RECT 155.930 116.540 156.900 118.800 ;
        RECT 146.270 116.510 156.900 116.540 ;
        RECT 106.500 116.380 118.910 116.430 ;
        RECT 127.240 116.400 137.900 116.510 ;
        RECT 146.240 116.400 156.900 116.510 ;
        RECT 102.160 116.210 118.910 116.380 ;
        RECT 125.490 116.350 137.900 116.400 ;
        RECT 144.490 116.350 156.900 116.400 ;
        RECT 102.160 114.800 102.330 116.210 ;
        RECT 102.700 115.640 105.740 115.810 ;
        RECT 102.700 115.200 105.740 115.370 ;
        RECT 105.955 115.340 106.125 115.670 ;
        RECT 106.460 115.450 118.910 116.210 ;
        RECT 121.150 116.180 137.900 116.350 ;
        RECT 106.460 115.440 118.800 115.450 ;
        RECT 106.460 115.430 112.340 115.440 ;
        RECT 106.460 115.410 107.030 115.430 ;
        RECT 108.250 115.420 112.340 115.430 ;
        RECT 106.470 114.800 106.640 115.410 ;
        RECT 102.160 114.630 106.640 114.800 ;
        RECT 121.150 114.770 121.320 116.180 ;
        RECT 121.690 115.610 124.730 115.780 ;
        RECT 121.690 115.170 124.730 115.340 ;
        RECT 124.945 115.310 125.115 115.640 ;
        RECT 125.450 115.420 137.900 116.180 ;
        RECT 140.150 116.180 156.900 116.350 ;
        RECT 125.450 115.410 137.790 115.420 ;
        RECT 125.450 115.400 131.330 115.410 ;
        RECT 125.450 115.380 126.020 115.400 ;
        RECT 127.240 115.390 131.330 115.400 ;
        RECT 125.460 114.770 125.630 115.380 ;
        RECT 121.150 114.600 125.630 114.770 ;
        RECT 140.150 114.770 140.320 116.180 ;
        RECT 140.690 115.610 143.730 115.780 ;
        RECT 140.690 115.170 143.730 115.340 ;
        RECT 143.945 115.310 144.115 115.640 ;
        RECT 144.450 115.420 156.900 116.180 ;
        RECT 144.450 115.410 156.790 115.420 ;
        RECT 144.450 115.400 150.330 115.410 ;
        RECT 144.450 115.380 145.020 115.400 ;
        RECT 146.240 115.390 150.330 115.400 ;
        RECT 144.460 114.770 144.630 115.380 ;
        RECT 140.150 114.600 144.630 114.770 ;
        RECT 100.950 113.280 106.690 113.290 ;
        RECT 100.460 113.120 106.690 113.280 ;
        RECT 100.460 110.860 101.130 113.120 ;
        RECT 101.800 112.550 105.840 112.720 ;
        RECT 101.460 111.490 101.630 112.490 ;
        RECT 106.010 111.490 106.180 112.490 ;
        RECT 101.800 111.260 105.840 111.430 ;
        RECT 106.520 110.860 106.690 113.120 ;
        RECT 100.460 110.690 106.690 110.860 ;
        RECT 100.460 107.430 101.130 110.690 ;
        RECT 101.800 110.120 105.840 110.290 ;
        RECT 101.460 108.060 101.630 110.060 ;
        RECT 106.010 108.060 106.180 110.060 ;
        RECT 101.800 107.830 105.840 108.000 ;
        RECT 106.520 107.430 106.690 110.690 ;
        RECT 100.460 107.260 106.690 107.430 ;
        RECT 100.460 104.000 101.130 107.260 ;
        RECT 101.800 106.690 105.840 106.860 ;
        RECT 101.460 104.630 101.630 106.630 ;
        RECT 106.010 104.630 106.180 106.630 ;
        RECT 101.800 104.400 105.840 104.570 ;
        RECT 106.520 104.000 106.690 107.260 ;
        RECT 100.460 103.990 106.690 104.000 ;
        RECT 108.280 113.260 118.110 113.300 ;
        RECT 119.940 113.260 125.680 113.270 ;
        RECT 108.280 113.130 118.910 113.260 ;
        RECT 108.280 110.870 108.450 113.130 ;
        RECT 109.175 112.560 117.215 112.730 ;
        RECT 108.790 111.500 108.960 112.500 ;
        RECT 117.430 111.500 117.600 112.500 ;
        RECT 109.175 111.270 117.215 111.440 ;
        RECT 117.940 110.870 118.910 113.130 ;
        RECT 108.280 110.700 118.910 110.870 ;
        RECT 108.280 107.440 108.450 110.700 ;
        RECT 109.175 110.130 117.215 110.300 ;
        RECT 108.790 108.070 108.960 110.070 ;
        RECT 117.430 108.070 117.600 110.070 ;
        RECT 109.175 107.840 117.215 108.010 ;
        RECT 117.940 107.440 118.910 110.700 ;
        RECT 108.280 107.270 118.910 107.440 ;
        RECT 108.280 104.010 108.450 107.270 ;
        RECT 109.175 106.700 117.215 106.870 ;
        RECT 108.790 104.640 108.960 106.640 ;
        RECT 117.430 104.640 117.600 106.640 ;
        RECT 109.175 104.410 117.215 104.580 ;
        RECT 117.940 104.010 118.910 107.270 ;
        RECT 100.460 103.890 106.700 103.990 ;
        RECT 100.450 103.330 106.700 103.890 ;
        RECT 100.450 103.310 105.620 103.330 ;
        RECT 100.450 103.240 104.440 103.310 ;
        RECT 100.450 101.970 102.370 103.240 ;
        RECT 103.880 103.230 104.440 103.240 ;
        RECT 104.110 102.140 104.440 103.230 ;
        RECT 104.810 102.760 105.850 102.930 ;
        RECT 104.810 102.320 105.850 102.490 ;
        RECT 106.020 102.460 106.190 102.790 ;
        RECT 100.460 98.780 101.400 101.970 ;
        RECT 104.270 101.920 104.440 102.140 ;
        RECT 106.530 101.920 106.700 103.330 ;
        RECT 104.270 101.750 106.700 101.920 ;
        RECT 108.280 103.840 118.910 104.010 ;
        RECT 119.450 113.100 125.680 113.260 ;
        RECT 119.450 110.840 120.120 113.100 ;
        RECT 120.790 112.530 124.830 112.700 ;
        RECT 120.450 111.470 120.620 112.470 ;
        RECT 125.000 111.470 125.170 112.470 ;
        RECT 120.790 111.240 124.830 111.410 ;
        RECT 125.510 110.840 125.680 113.100 ;
        RECT 119.450 110.670 125.680 110.840 ;
        RECT 119.450 107.410 120.120 110.670 ;
        RECT 120.790 110.100 124.830 110.270 ;
        RECT 120.450 108.040 120.620 110.040 ;
        RECT 125.000 108.040 125.170 110.040 ;
        RECT 120.790 107.810 124.830 107.980 ;
        RECT 125.510 107.410 125.680 110.670 ;
        RECT 119.450 107.240 125.680 107.410 ;
        RECT 119.450 103.980 120.120 107.240 ;
        RECT 120.790 106.670 124.830 106.840 ;
        RECT 120.450 104.610 120.620 106.610 ;
        RECT 125.000 104.610 125.170 106.610 ;
        RECT 120.790 104.380 124.830 104.550 ;
        RECT 125.510 103.980 125.680 107.240 ;
        RECT 119.450 103.970 125.680 103.980 ;
        RECT 127.270 113.240 137.100 113.280 ;
        RECT 138.990 113.260 144.730 113.270 ;
        RECT 127.270 113.110 137.900 113.240 ;
        RECT 127.270 110.850 127.440 113.110 ;
        RECT 128.165 112.540 136.205 112.710 ;
        RECT 127.780 111.480 127.950 112.480 ;
        RECT 136.420 111.480 136.590 112.480 ;
        RECT 128.165 111.250 136.205 111.420 ;
        RECT 136.930 110.850 137.900 113.110 ;
        RECT 127.270 110.680 137.900 110.850 ;
        RECT 127.270 107.420 127.440 110.680 ;
        RECT 128.165 110.110 136.205 110.280 ;
        RECT 127.780 108.050 127.950 110.050 ;
        RECT 136.420 108.050 136.590 110.050 ;
        RECT 128.165 107.820 136.205 107.990 ;
        RECT 136.930 107.420 137.900 110.680 ;
        RECT 127.270 107.250 137.900 107.420 ;
        RECT 127.270 103.990 127.440 107.250 ;
        RECT 128.165 106.680 136.205 106.850 ;
        RECT 127.780 104.620 127.950 106.620 ;
        RECT 136.420 104.620 136.590 106.620 ;
        RECT 128.165 104.390 136.205 104.560 ;
        RECT 136.930 103.990 137.900 107.250 ;
        RECT 119.450 103.870 125.690 103.970 ;
        RECT 108.280 101.580 108.450 103.840 ;
        RECT 109.175 103.270 117.215 103.440 ;
        RECT 108.790 102.210 108.960 103.210 ;
        RECT 117.430 102.210 117.600 103.210 ;
        RECT 109.175 101.980 117.215 102.150 ;
        RECT 117.940 101.580 118.910 103.840 ;
        RECT 119.440 103.310 125.690 103.870 ;
        RECT 119.440 103.290 124.610 103.310 ;
        RECT 119.440 103.220 123.430 103.290 ;
        RECT 119.440 101.950 121.360 103.220 ;
        RECT 122.870 103.210 123.430 103.220 ;
        RECT 123.100 102.120 123.430 103.210 ;
        RECT 123.800 102.740 124.840 102.910 ;
        RECT 123.800 102.300 124.840 102.470 ;
        RECT 125.010 102.440 125.180 102.770 ;
        RECT 123.260 101.900 123.430 102.120 ;
        RECT 125.520 101.900 125.690 103.310 ;
        RECT 123.260 101.730 125.690 101.900 ;
        RECT 127.270 103.820 137.900 103.990 ;
        RECT 138.500 113.100 144.730 113.260 ;
        RECT 138.500 110.840 139.170 113.100 ;
        RECT 139.840 112.530 143.880 112.700 ;
        RECT 139.500 111.470 139.670 112.470 ;
        RECT 144.050 111.470 144.220 112.470 ;
        RECT 139.840 111.240 143.880 111.410 ;
        RECT 144.560 110.840 144.730 113.100 ;
        RECT 138.500 110.670 144.730 110.840 ;
        RECT 138.500 107.410 139.170 110.670 ;
        RECT 139.840 110.100 143.880 110.270 ;
        RECT 139.500 108.040 139.670 110.040 ;
        RECT 144.050 108.040 144.220 110.040 ;
        RECT 139.840 107.810 143.880 107.980 ;
        RECT 144.560 107.410 144.730 110.670 ;
        RECT 138.500 107.240 144.730 107.410 ;
        RECT 138.500 103.980 139.170 107.240 ;
        RECT 139.840 106.670 143.880 106.840 ;
        RECT 139.500 104.610 139.670 106.610 ;
        RECT 144.050 104.610 144.220 106.610 ;
        RECT 139.840 104.380 143.880 104.550 ;
        RECT 144.560 103.980 144.730 107.240 ;
        RECT 138.500 103.970 144.730 103.980 ;
        RECT 146.320 113.240 156.150 113.280 ;
        RECT 146.320 113.110 156.950 113.240 ;
        RECT 146.320 110.850 146.490 113.110 ;
        RECT 147.215 112.540 155.255 112.710 ;
        RECT 146.830 111.480 147.000 112.480 ;
        RECT 155.470 111.480 155.640 112.480 ;
        RECT 147.215 111.250 155.255 111.420 ;
        RECT 155.980 110.850 156.950 113.110 ;
        RECT 146.320 110.680 156.950 110.850 ;
        RECT 146.320 107.420 146.490 110.680 ;
        RECT 147.215 110.110 155.255 110.280 ;
        RECT 146.830 108.050 147.000 110.050 ;
        RECT 155.470 108.050 155.640 110.050 ;
        RECT 147.215 107.820 155.255 107.990 ;
        RECT 155.980 107.420 156.950 110.680 ;
        RECT 146.320 107.250 156.950 107.420 ;
        RECT 146.320 103.990 146.490 107.250 ;
        RECT 147.215 106.680 155.255 106.850 ;
        RECT 146.830 104.620 147.000 106.620 ;
        RECT 155.470 104.620 155.640 106.620 ;
        RECT 147.215 104.390 155.255 104.560 ;
        RECT 155.980 103.990 156.950 107.250 ;
        RECT 138.500 103.870 144.740 103.970 ;
        RECT 108.280 101.550 118.910 101.580 ;
        RECT 108.250 101.440 118.910 101.550 ;
        RECT 127.270 101.560 127.440 103.820 ;
        RECT 128.165 103.250 136.205 103.420 ;
        RECT 127.780 102.190 127.950 103.190 ;
        RECT 136.420 102.190 136.590 103.190 ;
        RECT 128.165 101.960 136.205 102.130 ;
        RECT 136.930 101.560 137.900 103.820 ;
        RECT 138.490 103.310 144.740 103.870 ;
        RECT 138.490 103.290 143.660 103.310 ;
        RECT 138.490 103.220 142.480 103.290 ;
        RECT 138.490 101.950 140.410 103.220 ;
        RECT 141.920 103.210 142.480 103.220 ;
        RECT 142.150 102.120 142.480 103.210 ;
        RECT 142.850 102.740 143.890 102.910 ;
        RECT 142.850 102.300 143.890 102.470 ;
        RECT 144.060 102.440 144.230 102.770 ;
        RECT 142.310 101.900 142.480 102.120 ;
        RECT 144.570 101.900 144.740 103.310 ;
        RECT 142.310 101.730 144.740 101.900 ;
        RECT 146.320 103.820 156.950 103.990 ;
        RECT 127.270 101.530 137.900 101.560 ;
        RECT 146.320 101.560 146.490 103.820 ;
        RECT 147.215 103.250 155.255 103.420 ;
        RECT 146.830 102.190 147.000 103.190 ;
        RECT 155.470 102.190 155.640 103.190 ;
        RECT 147.215 101.960 155.255 102.130 ;
        RECT 155.980 101.560 156.950 103.820 ;
        RECT 146.320 101.530 156.950 101.560 ;
        RECT 106.500 101.390 118.910 101.440 ;
        RECT 127.240 101.420 137.900 101.530 ;
        RECT 146.290 101.420 156.950 101.530 ;
        RECT 102.160 101.220 118.910 101.390 ;
        RECT 125.490 101.370 137.900 101.420 ;
        RECT 144.540 101.370 156.950 101.420 ;
        RECT 102.160 99.810 102.330 101.220 ;
        RECT 102.700 100.650 105.740 100.820 ;
        RECT 102.700 100.210 105.740 100.380 ;
        RECT 105.955 100.350 106.125 100.680 ;
        RECT 106.460 100.460 118.910 101.220 ;
        RECT 121.150 101.200 137.900 101.370 ;
        RECT 106.460 100.450 118.800 100.460 ;
        RECT 106.460 100.440 112.340 100.450 ;
        RECT 106.460 100.420 107.030 100.440 ;
        RECT 108.250 100.430 112.340 100.440 ;
        RECT 106.470 99.810 106.640 100.420 ;
        RECT 102.160 99.640 106.640 99.810 ;
        RECT 121.150 99.790 121.320 101.200 ;
        RECT 121.690 100.630 124.730 100.800 ;
        RECT 121.690 100.190 124.730 100.360 ;
        RECT 124.945 100.330 125.115 100.660 ;
        RECT 125.450 100.440 137.900 101.200 ;
        RECT 140.200 101.200 156.950 101.370 ;
        RECT 125.450 100.430 137.790 100.440 ;
        RECT 125.450 100.420 131.330 100.430 ;
        RECT 125.450 100.400 126.020 100.420 ;
        RECT 127.240 100.410 131.330 100.420 ;
        RECT 125.460 99.790 125.630 100.400 ;
        RECT 121.150 99.620 125.630 99.790 ;
        RECT 140.200 99.790 140.370 101.200 ;
        RECT 140.740 100.630 143.780 100.800 ;
        RECT 140.740 100.190 143.780 100.360 ;
        RECT 143.995 100.330 144.165 100.660 ;
        RECT 144.500 100.440 156.950 101.200 ;
        RECT 144.500 100.430 156.840 100.440 ;
        RECT 144.500 100.420 150.380 100.430 ;
        RECT 144.500 100.400 145.070 100.420 ;
        RECT 146.290 100.410 150.380 100.420 ;
        RECT 144.510 99.790 144.680 100.400 ;
        RECT 140.200 99.620 144.680 99.790 ;
        RECT 100.410 98.750 102.840 98.780 ;
        RECT 100.410 98.580 156.750 98.750 ;
        RECT 100.410 97.270 102.840 98.580 ;
        RECT 103.320 97.750 105.480 98.100 ;
        RECT 106.020 97.750 108.180 98.100 ;
        RECT 108.660 97.270 108.830 98.580 ;
        RECT 109.310 97.750 111.470 98.100 ;
        RECT 112.010 97.750 114.170 98.100 ;
        RECT 114.650 97.270 114.820 98.580 ;
        RECT 115.300 97.750 117.460 98.100 ;
        RECT 118.000 97.750 120.160 98.100 ;
        RECT 120.640 97.270 120.810 98.580 ;
        RECT 121.290 97.750 123.450 98.100 ;
        RECT 123.990 97.750 126.150 98.100 ;
        RECT 126.630 97.270 126.800 98.580 ;
        RECT 127.280 97.750 129.440 98.100 ;
        RECT 129.980 97.750 132.140 98.100 ;
        RECT 132.620 97.270 132.790 98.580 ;
        RECT 133.270 97.750 135.430 98.100 ;
        RECT 135.970 97.750 138.130 98.100 ;
        RECT 138.610 97.270 138.780 98.580 ;
        RECT 139.260 97.750 141.420 98.100 ;
        RECT 141.960 97.750 144.120 98.100 ;
        RECT 144.600 97.270 144.770 98.580 ;
        RECT 145.250 97.750 147.410 98.100 ;
        RECT 147.950 97.750 150.110 98.100 ;
        RECT 150.590 97.270 150.760 98.580 ;
        RECT 151.240 97.750 153.400 98.100 ;
        RECT 153.940 97.750 156.100 98.100 ;
        RECT 156.580 97.270 156.750 98.580 ;
        RECT 100.410 97.100 156.750 97.270 ;
        RECT 100.410 95.790 102.840 97.100 ;
        RECT 103.320 96.270 105.480 96.620 ;
        RECT 106.020 96.270 108.180 96.620 ;
        RECT 108.660 95.790 108.830 97.100 ;
        RECT 109.310 96.270 111.470 96.620 ;
        RECT 112.010 96.270 114.170 96.620 ;
        RECT 114.650 95.790 114.820 97.100 ;
        RECT 115.300 96.270 117.460 96.620 ;
        RECT 118.000 96.270 120.160 96.620 ;
        RECT 120.640 95.790 120.810 97.100 ;
        RECT 121.290 96.270 123.450 96.620 ;
        RECT 123.990 96.270 126.150 96.620 ;
        RECT 126.630 95.790 126.800 97.100 ;
        RECT 127.280 96.270 129.440 96.620 ;
        RECT 129.980 96.270 132.140 96.620 ;
        RECT 132.620 95.790 132.790 97.100 ;
        RECT 133.270 96.270 135.430 96.620 ;
        RECT 135.970 96.270 138.130 96.620 ;
        RECT 138.610 95.790 138.780 97.100 ;
        RECT 139.260 96.270 141.420 96.620 ;
        RECT 141.960 96.270 144.120 96.620 ;
        RECT 144.600 95.790 144.770 97.100 ;
        RECT 100.410 95.650 144.770 95.790 ;
        RECT 102.670 95.620 144.770 95.650 ;
      LAYER met1 ;
        RECT 147.680 220.250 147.940 220.570 ;
        RECT 147.240 219.710 147.500 220.030 ;
        RECT 113.920 218.970 114.180 219.290 ;
        RECT 146.840 219.250 147.160 219.510 ;
        RECT 108.350 205.840 108.610 206.160 ;
        RECT 108.410 201.760 108.550 205.840 ;
        RECT 108.810 205.290 109.070 205.610 ;
        RECT 108.870 202.330 109.010 205.290 ;
        RECT 109.290 204.800 109.550 205.120 ;
        RECT 109.350 203.170 109.490 204.800 ;
        RECT 109.290 202.850 109.550 203.170 ;
        RECT 108.870 202.190 109.920 202.330 ;
        RECT 108.410 201.620 109.370 201.760 ;
        RECT 107.815 174.670 108.810 198.905 ;
        RECT 109.230 196.510 109.370 201.620 ;
        RECT 109.780 197.210 109.920 202.190 ;
        RECT 109.690 196.890 110.020 197.210 ;
        RECT 109.230 196.370 109.540 196.510 ;
        RECT 109.400 191.230 109.540 196.370 ;
        RECT 109.400 191.000 109.930 191.230 ;
        RECT 109.670 190.910 109.930 191.000 ;
        RECT 110.240 182.100 110.720 217.980 ;
        RECT 111.540 206.550 111.800 206.870 ;
        RECT 110.875 205.645 111.105 205.935 ;
        RECT 110.920 204.110 111.060 205.645 ;
        RECT 110.860 203.790 111.120 204.110 ;
        RECT 110.875 203.345 111.105 203.635 ;
        RECT 110.920 201.350 111.060 203.345 ;
        RECT 111.555 202.640 111.785 202.715 ;
        RECT 111.555 202.500 112.760 202.640 ;
        RECT 111.555 202.425 111.785 202.500 ;
        RECT 111.555 201.965 111.785 202.255 ;
        RECT 111.600 201.810 111.740 201.965 ;
        RECT 111.540 201.490 111.800 201.810 ;
        RECT 112.235 201.480 112.465 201.770 ;
        RECT 110.860 201.030 111.120 201.350 ;
        RECT 111.895 201.085 112.125 201.375 ;
        RECT 111.215 200.630 111.445 200.920 ;
        RECT 111.260 199.510 111.400 200.630 ;
        RECT 111.940 200.185 112.080 201.085 ;
        RECT 111.895 199.895 112.125 200.185 ;
        RECT 111.200 199.190 111.460 199.510 ;
        RECT 111.940 197.665 112.080 199.895 ;
        RECT 112.280 199.670 112.420 201.480 ;
        RECT 112.235 199.380 112.465 199.670 ;
        RECT 112.280 198.100 112.420 199.380 ;
        RECT 112.235 197.810 112.465 198.100 ;
        RECT 111.895 197.375 112.125 197.665 ;
        RECT 110.860 197.120 111.120 197.210 ;
        RECT 110.860 196.980 111.400 197.120 ;
        RECT 110.860 196.890 111.120 196.980 ;
        RECT 110.875 194.360 111.105 194.435 ;
        RECT 111.260 194.360 111.400 196.980 ;
        RECT 112.620 196.750 112.760 202.500 ;
        RECT 112.560 196.430 112.820 196.750 ;
        RECT 112.235 195.065 112.465 195.355 ;
        RECT 110.875 194.220 111.400 194.360 ;
        RECT 110.875 194.145 111.105 194.220 ;
        RECT 112.280 193.530 112.420 195.065 ;
        RECT 111.540 193.210 111.800 193.530 ;
        RECT 112.220 193.210 112.480 193.530 ;
        RECT 110.860 190.910 111.120 191.230 ;
        RECT 110.920 189.835 111.060 190.910 ;
        RECT 111.540 190.450 111.800 190.770 ;
        RECT 110.875 189.545 111.105 189.835 ;
        RECT 112.575 188.625 112.805 188.915 ;
        RECT 111.880 188.150 112.140 188.470 ;
        RECT 111.540 187.690 111.800 188.010 ;
        RECT 111.940 186.615 112.080 188.150 ;
        RECT 112.220 187.230 112.480 187.550 ;
        RECT 111.895 186.325 112.125 186.615 ;
        RECT 112.280 185.235 112.420 187.230 ;
        RECT 112.620 187.090 112.760 188.625 ;
        RECT 112.560 186.770 112.820 187.090 ;
        RECT 112.235 184.945 112.465 185.235 ;
        RECT 112.560 184.470 112.820 184.790 ;
        RECT 112.620 184.315 112.760 184.470 ;
        RECT 112.575 184.025 112.805 184.315 ;
        RECT 112.960 182.100 113.440 217.980 ;
        RECT 113.980 216.055 114.120 218.970 ;
        RECT 146.310 218.730 146.570 219.050 ;
        RECT 114.600 216.210 114.860 216.530 ;
        RECT 113.935 215.765 114.165 216.055 ;
        RECT 114.660 215.135 114.800 216.210 ;
        RECT 114.615 214.845 114.845 215.135 ;
        RECT 115.280 213.450 115.540 213.770 ;
        RECT 115.280 211.610 115.540 211.930 ;
        RECT 115.280 211.150 115.540 211.470 ;
        RECT 114.275 210.245 114.505 210.535 ;
        RECT 114.320 205.030 114.460 210.245 ;
        RECT 115.280 208.850 115.540 209.170 ;
        RECT 115.340 206.870 115.480 208.850 ;
        RECT 115.280 206.550 115.540 206.870 ;
        RECT 114.260 204.710 114.520 205.030 ;
        RECT 115.340 204.555 115.480 206.550 ;
        RECT 115.295 204.265 115.525 204.555 ;
        RECT 114.275 201.955 114.505 202.245 ;
        RECT 113.935 201.520 114.165 201.810 ;
        RECT 113.980 200.240 114.120 201.520 ;
        RECT 113.935 199.950 114.165 200.240 ;
        RECT 113.580 199.190 113.840 199.510 ;
        RECT 113.640 197.195 113.780 199.190 ;
        RECT 113.980 198.140 114.120 199.950 ;
        RECT 114.320 199.725 114.460 201.955 ;
        RECT 115.280 200.340 115.540 200.430 ;
        RECT 114.660 200.200 115.540 200.340 ;
        RECT 114.275 199.435 114.505 199.725 ;
        RECT 114.320 198.535 114.460 199.435 ;
        RECT 114.660 198.990 114.800 200.200 ;
        RECT 115.280 200.110 115.540 200.200 ;
        RECT 114.940 199.190 115.200 199.510 ;
        RECT 114.615 198.700 114.845 198.990 ;
        RECT 114.275 198.245 114.505 198.535 ;
        RECT 113.935 197.850 114.165 198.140 ;
        RECT 114.615 197.580 114.845 197.655 ;
        RECT 115.000 197.580 115.140 199.190 ;
        RECT 114.615 197.440 115.140 197.580 ;
        RECT 114.615 197.365 114.845 197.440 ;
        RECT 113.595 196.905 113.825 197.195 ;
        RECT 114.615 195.065 114.845 195.355 ;
        RECT 114.260 193.670 114.520 193.990 ;
        RECT 114.260 193.210 114.520 193.530 ;
        RECT 114.320 188.915 114.460 193.210 ;
        RECT 114.660 191.675 114.800 195.065 ;
        RECT 115.280 194.590 115.540 194.910 ;
        RECT 114.615 191.385 114.845 191.675 ;
        RECT 114.275 188.625 114.505 188.915 ;
        RECT 114.260 188.150 114.520 188.470 ;
        RECT 114.320 187.075 114.460 188.150 ;
        RECT 114.600 187.690 114.860 188.010 ;
        RECT 114.275 186.785 114.505 187.075 ;
        RECT 114.275 186.325 114.505 186.615 ;
        RECT 114.320 183.870 114.460 186.325 ;
        RECT 114.660 185.695 114.800 187.690 ;
        RECT 114.615 185.405 114.845 185.695 ;
        RECT 115.280 184.930 115.540 185.250 ;
        RECT 115.340 184.775 115.480 184.930 ;
        RECT 115.295 184.485 115.525 184.775 ;
        RECT 114.260 183.550 114.520 183.870 ;
        RECT 115.680 182.100 116.160 217.980 ;
        RECT 118.000 216.210 118.260 216.530 ;
        RECT 117.335 213.915 117.565 214.205 ;
        RECT 116.640 213.450 116.900 213.770 ;
        RECT 116.700 210.950 116.840 213.450 ;
        RECT 117.380 211.685 117.520 213.915 ;
        RECT 117.675 213.480 117.905 213.770 ;
        RECT 117.720 212.200 117.860 213.480 ;
        RECT 117.675 211.910 117.905 212.200 ;
        RECT 117.335 211.395 117.565 211.685 ;
        RECT 116.655 210.660 116.885 210.950 ;
        RECT 117.380 210.495 117.520 211.395 ;
        RECT 117.335 210.205 117.565 210.495 ;
        RECT 117.720 210.100 117.860 211.910 ;
        RECT 117.675 209.810 117.905 210.100 ;
        RECT 117.320 209.310 117.580 209.630 ;
        RECT 116.995 204.265 117.225 204.555 ;
        RECT 117.040 199.970 117.180 204.265 ;
        RECT 116.980 199.650 117.240 199.970 ;
        RECT 118.000 199.190 118.260 199.510 ;
        RECT 118.060 198.115 118.200 199.190 ;
        RECT 118.015 197.825 118.245 198.115 ;
        RECT 116.995 193.900 117.225 193.975 ;
        RECT 116.995 193.760 117.520 193.900 ;
        RECT 116.995 193.685 117.225 193.760 ;
        RECT 116.980 192.290 117.240 192.610 ;
        RECT 116.315 191.600 116.545 191.675 ;
        RECT 116.315 191.460 116.840 191.600 ;
        RECT 116.315 191.385 116.545 191.460 ;
        RECT 116.315 188.625 116.545 188.915 ;
        RECT 116.360 188.470 116.500 188.625 ;
        RECT 116.300 188.150 116.560 188.470 ;
        RECT 116.700 188.380 116.840 191.460 ;
        RECT 116.980 190.910 117.240 191.230 ;
        RECT 116.980 189.530 117.240 189.850 ;
        RECT 116.995 188.380 117.225 188.455 ;
        RECT 116.700 188.240 117.225 188.380 ;
        RECT 116.300 187.690 116.560 188.010 ;
        RECT 116.700 186.080 116.840 188.240 ;
        RECT 116.995 188.165 117.225 188.240 ;
        RECT 116.995 187.245 117.225 187.535 ;
        RECT 117.040 187.090 117.180 187.245 ;
        RECT 116.980 186.770 117.240 187.090 ;
        RECT 116.980 186.080 117.240 186.170 ;
        RECT 116.700 185.940 117.240 186.080 ;
        RECT 116.980 185.850 117.240 185.940 ;
        RECT 116.980 184.470 117.240 184.790 ;
        RECT 117.380 184.330 117.520 193.760 ;
        RECT 117.675 192.765 117.905 193.055 ;
        RECT 117.720 187.550 117.860 192.765 ;
        RECT 118.015 190.005 118.245 190.295 ;
        RECT 118.060 188.010 118.200 190.005 ;
        RECT 118.000 187.690 118.260 188.010 ;
        RECT 117.660 187.230 117.920 187.550 ;
        RECT 118.015 186.785 118.245 187.075 ;
        RECT 118.060 186.630 118.200 186.785 ;
        RECT 118.000 186.310 118.260 186.630 ;
        RECT 117.320 184.010 117.580 184.330 ;
        RECT 116.980 183.550 117.240 183.870 ;
        RECT 118.400 182.100 118.880 217.980 ;
        RECT 119.360 216.670 119.620 216.990 ;
        RECT 119.420 216.055 119.560 216.670 ;
        RECT 119.700 216.210 119.960 216.530 ;
        RECT 119.375 215.765 119.605 216.055 ;
        RECT 119.760 213.755 119.900 216.210 ;
        RECT 120.055 214.845 120.285 215.135 ;
        RECT 119.715 213.465 119.945 213.755 ;
        RECT 119.020 211.610 119.280 211.930 ;
        RECT 119.080 210.535 119.220 211.610 ;
        RECT 119.360 211.150 119.620 211.470 ;
        RECT 119.035 210.245 119.265 210.535 ;
        RECT 119.035 201.505 119.265 201.795 ;
        RECT 119.080 200.430 119.220 201.505 ;
        RECT 119.020 200.110 119.280 200.430 ;
        RECT 119.420 199.420 119.560 211.150 ;
        RECT 119.700 208.850 119.960 209.170 ;
        RECT 120.100 208.710 120.240 214.845 ;
        RECT 120.040 208.390 120.300 208.710 ;
        RECT 120.055 205.645 120.285 205.935 ;
        RECT 119.700 204.710 119.960 205.030 ;
        RECT 119.715 203.805 119.945 204.095 ;
        RECT 119.760 199.880 119.900 203.805 ;
        RECT 120.100 203.635 120.240 205.645 ;
        RECT 120.055 203.345 120.285 203.635 ;
        RECT 119.760 199.740 120.580 199.880 ;
        RECT 119.080 199.280 119.560 199.420 ;
        RECT 119.080 193.070 119.220 199.280 ;
        RECT 120.040 199.190 120.300 199.510 ;
        RECT 119.375 198.720 119.605 199.010 ;
        RECT 119.420 196.910 119.560 198.720 ;
        RECT 119.715 198.325 119.945 198.615 ;
        RECT 119.760 197.425 119.900 198.325 ;
        RECT 120.055 197.870 120.285 198.160 ;
        RECT 119.715 197.135 119.945 197.425 ;
        RECT 119.375 196.620 119.605 196.910 ;
        RECT 119.420 195.340 119.560 196.620 ;
        RECT 119.375 195.050 119.605 195.340 ;
        RECT 119.760 194.905 119.900 197.135 ;
        RECT 119.715 194.615 119.945 194.905 ;
        RECT 120.100 194.360 120.240 197.870 ;
        RECT 120.440 194.910 120.580 199.740 ;
        RECT 120.380 194.590 120.640 194.910 ;
        RECT 119.420 194.220 120.240 194.360 ;
        RECT 119.020 192.750 119.280 193.070 ;
        RECT 119.035 192.305 119.265 192.595 ;
        RECT 119.080 190.770 119.220 192.305 ;
        RECT 119.420 191.675 119.560 194.220 ;
        RECT 120.040 193.670 120.300 193.990 ;
        RECT 119.700 192.750 119.960 193.070 ;
        RECT 119.375 191.385 119.605 191.675 ;
        RECT 119.020 190.450 119.280 190.770 ;
        RECT 119.760 189.375 119.900 192.750 ;
        RECT 119.715 189.085 119.945 189.375 ;
        RECT 119.715 188.840 119.945 188.915 ;
        RECT 120.100 188.840 120.240 193.670 ;
        RECT 120.720 189.530 120.980 189.850 ;
        RECT 119.715 188.700 120.240 188.840 ;
        RECT 119.715 188.625 119.945 188.700 ;
        RECT 119.700 187.690 119.960 188.010 ;
        RECT 119.020 186.770 119.280 187.090 ;
        RECT 119.080 185.235 119.220 186.770 ;
        RECT 119.375 186.325 119.605 186.615 ;
        RECT 119.035 184.945 119.265 185.235 ;
        RECT 119.420 183.870 119.560 186.325 ;
        RECT 119.760 184.790 119.900 187.690 ;
        RECT 120.040 187.230 120.300 187.550 ;
        RECT 120.040 185.850 120.300 186.170 ;
        RECT 120.720 185.850 120.980 186.170 ;
        RECT 120.100 185.235 120.240 185.850 ;
        RECT 120.380 185.390 120.640 185.710 ;
        RECT 120.055 184.945 120.285 185.235 ;
        RECT 119.700 184.470 119.960 184.790 ;
        RECT 119.360 183.550 119.620 183.870 ;
        RECT 120.440 183.855 120.580 185.390 ;
        RECT 120.395 183.565 120.625 183.855 ;
        RECT 121.120 182.100 121.600 217.980 ;
        RECT 122.760 216.440 123.020 216.530 ;
        RECT 122.480 216.300 123.020 216.440 ;
        RECT 122.095 214.890 122.325 215.180 ;
        RECT 122.140 214.230 122.280 214.890 ;
        RECT 122.080 213.910 122.340 214.230 ;
        RECT 122.480 209.630 122.620 216.300 ;
        RECT 122.760 216.210 123.020 216.300 ;
        RECT 123.115 215.740 123.345 216.030 ;
        RECT 122.775 215.345 123.005 215.635 ;
        RECT 122.820 214.445 122.960 215.345 ;
        RECT 122.775 214.155 123.005 214.445 ;
        RECT 122.820 211.925 122.960 214.155 ;
        RECT 123.160 213.930 123.300 215.740 ;
        RECT 123.115 213.640 123.345 213.930 ;
        RECT 123.160 212.360 123.300 213.640 ;
        RECT 123.115 212.070 123.345 212.360 ;
        RECT 122.775 211.635 123.005 211.925 ;
        RECT 122.420 209.310 122.680 209.630 ;
        RECT 123.455 209.325 123.685 209.615 ;
        RECT 122.480 204.555 122.620 209.310 ;
        RECT 123.500 208.710 123.640 209.325 ;
        RECT 123.440 208.390 123.700 208.710 ;
        RECT 122.435 204.480 122.665 204.555 ;
        RECT 121.800 204.340 122.665 204.480 ;
        RECT 121.800 199.510 121.940 204.340 ;
        RECT 122.435 204.265 122.665 204.340 ;
        RECT 123.115 203.780 123.345 204.070 ;
        RECT 122.080 203.330 122.340 203.650 ;
        RECT 122.775 203.385 123.005 203.675 ;
        RECT 122.140 203.100 122.280 203.330 ;
        RECT 122.435 203.100 122.665 203.220 ;
        RECT 122.140 202.960 122.665 203.100 ;
        RECT 122.435 202.930 122.665 202.960 ;
        RECT 122.820 202.485 122.960 203.385 ;
        RECT 122.775 202.195 123.005 202.485 ;
        RECT 122.820 199.965 122.960 202.195 ;
        RECT 123.160 201.970 123.300 203.780 ;
        RECT 123.115 201.680 123.345 201.970 ;
        RECT 123.160 200.400 123.300 201.680 ;
        RECT 123.115 200.110 123.345 200.400 ;
        RECT 122.775 199.675 123.005 199.965 ;
        RECT 121.740 199.190 122.000 199.510 ;
        RECT 121.755 197.365 121.985 197.655 ;
        RECT 121.800 196.750 121.940 197.365 ;
        RECT 122.775 196.905 123.005 197.195 ;
        RECT 121.740 196.430 122.000 196.750 ;
        RECT 122.820 196.290 122.960 196.905 ;
        RECT 122.760 195.970 123.020 196.290 ;
        RECT 123.100 195.050 123.360 195.370 ;
        RECT 123.455 194.605 123.685 194.895 ;
        RECT 123.500 193.990 123.640 194.605 ;
        RECT 123.440 193.670 123.700 193.990 ;
        RECT 122.420 190.450 122.680 190.770 ;
        RECT 121.740 189.530 122.000 189.850 ;
        RECT 121.800 187.535 121.940 189.530 ;
        RECT 122.760 188.150 123.020 188.470 ;
        RECT 122.420 187.690 122.680 188.010 ;
        RECT 121.755 187.245 121.985 187.535 ;
        RECT 122.480 186.155 122.620 187.690 ;
        RECT 122.435 185.865 122.665 186.155 ;
        RECT 122.420 185.390 122.680 185.710 ;
        RECT 122.420 184.930 122.680 185.250 ;
        RECT 122.435 184.700 122.665 184.775 ;
        RECT 122.820 184.700 122.960 188.150 ;
        RECT 123.440 187.690 123.700 188.010 ;
        RECT 123.500 187.075 123.640 187.690 ;
        RECT 123.455 186.785 123.685 187.075 ;
        RECT 122.435 184.560 122.960 184.700 ;
        RECT 122.435 184.485 122.665 184.560 ;
        RECT 123.840 182.100 124.320 217.980 ;
        RECT 126.160 216.670 126.420 216.990 ;
        RECT 124.800 216.210 125.060 216.530 ;
        RECT 125.480 216.210 125.740 216.530 ;
        RECT 124.460 213.910 124.720 214.230 ;
        RECT 124.860 210.000 125.000 216.210 ;
        RECT 125.540 215.135 125.680 216.210 ;
        RECT 126.220 216.055 126.360 216.670 ;
        RECT 126.175 215.765 126.405 216.055 ;
        RECT 125.495 214.845 125.725 215.135 ;
        RECT 126.175 212.085 126.405 212.375 ;
        RECT 125.155 211.625 125.385 211.915 ;
        RECT 125.200 211.470 125.340 211.625 ;
        RECT 126.220 211.470 126.360 212.085 ;
        RECT 125.140 211.150 125.400 211.470 ;
        RECT 126.160 211.150 126.420 211.470 ;
        RECT 125.140 210.690 125.400 211.010 ;
        RECT 125.155 210.000 125.385 210.075 ;
        RECT 124.860 209.860 125.385 210.000 ;
        RECT 125.155 209.785 125.385 209.860 ;
        RECT 124.815 209.300 125.045 209.590 ;
        RECT 124.860 207.490 125.000 209.300 ;
        RECT 125.155 208.905 125.385 209.195 ;
        RECT 125.200 208.005 125.340 208.905 ;
        RECT 125.835 208.450 126.065 208.740 ;
        RECT 125.155 207.715 125.385 208.005 ;
        RECT 124.815 207.200 125.045 207.490 ;
        RECT 124.860 205.920 125.000 207.200 ;
        RECT 124.815 205.630 125.045 205.920 ;
        RECT 125.200 205.485 125.340 207.715 ;
        RECT 125.155 205.195 125.385 205.485 ;
        RECT 125.880 205.030 126.020 208.450 ;
        RECT 125.820 204.710 126.080 205.030 ;
        RECT 125.880 203.650 126.020 204.710 ;
        RECT 124.800 203.330 125.060 203.650 ;
        RECT 125.820 203.330 126.080 203.650 ;
        RECT 124.860 202.715 125.000 203.330 ;
        RECT 126.160 202.870 126.420 203.190 ;
        RECT 124.815 202.425 125.045 202.715 ;
        RECT 125.495 200.585 125.725 200.875 ;
        RECT 125.155 200.340 125.385 200.415 ;
        RECT 124.860 200.200 125.385 200.340 ;
        RECT 124.860 194.910 125.000 200.200 ;
        RECT 125.155 200.125 125.385 200.200 ;
        RECT 125.155 199.205 125.385 199.495 ;
        RECT 125.200 197.210 125.340 199.205 ;
        RECT 125.540 198.575 125.680 200.585 ;
        RECT 125.495 198.285 125.725 198.575 ;
        RECT 125.140 196.890 125.400 197.210 ;
        RECT 125.140 196.430 125.400 196.750 ;
        RECT 125.200 195.815 125.340 196.430 ;
        RECT 126.220 196.290 126.360 202.870 ;
        RECT 126.160 195.970 126.420 196.290 ;
        RECT 125.155 195.525 125.385 195.815 ;
        RECT 124.800 194.590 125.060 194.910 ;
        RECT 124.860 188.915 125.000 194.590 ;
        RECT 125.480 192.290 125.740 192.610 ;
        RECT 125.540 191.215 125.680 192.290 ;
        RECT 125.495 190.925 125.725 191.215 ;
        RECT 125.495 190.680 125.725 190.755 ;
        RECT 125.495 190.540 126.020 190.680 ;
        RECT 125.495 190.465 125.725 190.540 ;
        RECT 125.480 189.990 125.740 190.310 ;
        RECT 125.155 189.545 125.385 189.835 ;
        RECT 124.815 188.625 125.045 188.915 ;
        RECT 125.200 186.170 125.340 189.545 ;
        RECT 125.880 188.470 126.020 190.540 ;
        RECT 125.820 188.150 126.080 188.470 ;
        RECT 125.495 187.245 125.725 187.535 ;
        RECT 125.540 187.090 125.680 187.245 ;
        RECT 125.480 186.770 125.740 187.090 ;
        RECT 125.480 186.310 125.740 186.630 ;
        RECT 126.160 186.310 126.420 186.630 ;
        RECT 125.140 185.850 125.400 186.170 ;
        RECT 125.495 184.945 125.725 185.235 ;
        RECT 125.540 184.790 125.680 184.945 ;
        RECT 125.480 184.470 125.740 184.790 ;
        RECT 126.220 184.315 126.360 186.310 ;
        RECT 126.175 184.025 126.405 184.315 ;
        RECT 126.560 182.100 127.040 217.980 ;
        RECT 128.200 216.210 128.460 216.530 ;
        RECT 128.260 215.135 128.400 216.210 ;
        RECT 128.215 214.845 128.445 215.135 ;
        RECT 128.880 211.610 129.140 211.930 ;
        RECT 127.180 211.150 127.440 211.470 ;
        RECT 127.860 208.390 128.120 208.710 ;
        RECT 127.875 204.480 128.105 204.555 ;
        RECT 127.580 204.340 128.105 204.480 ;
        RECT 127.580 199.035 127.720 204.340 ;
        RECT 127.875 204.265 128.105 204.340 ;
        RECT 127.875 203.560 128.105 203.635 ;
        RECT 127.875 203.420 128.400 203.560 ;
        RECT 127.875 203.345 128.105 203.420 ;
        RECT 127.860 202.870 128.120 203.190 ;
        RECT 128.260 202.180 128.400 203.420 ;
        RECT 128.880 203.330 129.140 203.650 ;
        RECT 128.880 202.870 129.140 203.190 ;
        RECT 128.555 202.180 128.785 202.255 ;
        RECT 128.260 202.040 128.785 202.180 ;
        RECT 128.555 201.965 128.785 202.040 ;
        RECT 128.215 201.505 128.445 201.795 ;
        RECT 127.875 200.585 128.105 200.875 ;
        RECT 127.920 200.430 128.060 200.585 ;
        RECT 127.860 200.110 128.120 200.430 ;
        RECT 127.860 199.190 128.120 199.510 ;
        RECT 127.535 198.745 127.765 199.035 ;
        RECT 128.260 196.200 128.400 201.505 ;
        RECT 128.600 199.050 128.740 201.965 ;
        RECT 128.940 201.335 129.080 202.870 ;
        RECT 128.895 201.045 129.125 201.335 ;
        RECT 128.540 198.730 128.800 199.050 ;
        RECT 128.260 196.060 128.740 196.200 ;
        RECT 128.200 195.510 128.460 195.830 ;
        RECT 128.600 194.910 128.740 196.060 ;
        RECT 128.540 194.590 128.800 194.910 ;
        RECT 127.195 193.685 127.425 193.975 ;
        RECT 127.240 193.070 127.380 193.685 ;
        RECT 127.180 192.750 127.440 193.070 ;
        RECT 127.875 192.980 128.105 193.055 ;
        RECT 127.875 192.840 128.400 192.980 ;
        RECT 127.875 192.765 128.105 192.840 ;
        RECT 127.875 191.845 128.105 192.135 ;
        RECT 127.535 190.465 127.765 190.755 ;
        RECT 127.180 189.990 127.440 190.310 ;
        RECT 127.240 189.835 127.380 189.990 ;
        RECT 127.195 189.545 127.425 189.835 ;
        RECT 127.580 188.470 127.720 190.465 ;
        RECT 127.920 190.295 128.060 191.845 ;
        RECT 127.875 190.005 128.105 190.295 ;
        RECT 127.920 189.850 128.060 190.005 ;
        RECT 127.860 189.530 128.120 189.850 ;
        RECT 127.875 189.300 128.105 189.375 ;
        RECT 128.260 189.300 128.400 192.840 ;
        RECT 128.880 192.290 129.140 192.610 ;
        RECT 127.875 189.160 128.400 189.300 ;
        RECT 127.875 189.085 128.105 189.160 ;
        RECT 127.860 188.610 128.120 188.930 ;
        RECT 127.520 188.150 127.780 188.470 ;
        RECT 127.195 187.920 127.425 187.995 ;
        RECT 127.195 187.780 127.720 187.920 ;
        RECT 127.195 187.705 127.425 187.780 ;
        RECT 127.580 187.460 127.720 187.780 ;
        RECT 127.875 187.460 128.105 187.535 ;
        RECT 127.580 187.320 128.105 187.460 ;
        RECT 127.580 185.710 127.720 187.320 ;
        RECT 127.875 187.245 128.105 187.320 ;
        RECT 127.860 186.310 128.120 186.630 ;
        RECT 128.260 186.540 128.400 189.160 ;
        RECT 128.540 186.540 128.800 186.630 ;
        RECT 128.260 186.400 128.800 186.540 ;
        RECT 128.540 186.310 128.800 186.400 ;
        RECT 127.860 185.850 128.120 186.170 ;
        RECT 127.520 185.390 127.780 185.710 ;
        RECT 127.920 185.235 128.060 185.850 ;
        RECT 127.875 184.945 128.105 185.235 ;
        RECT 128.880 184.930 129.140 185.250 ;
        RECT 128.940 184.315 129.080 184.930 ;
        RECT 128.895 184.025 129.125 184.315 ;
        RECT 129.280 182.100 129.760 217.980 ;
        RECT 129.900 216.210 130.160 216.530 ;
        RECT 131.260 216.210 131.520 216.530 ;
        RECT 130.595 213.915 130.825 214.205 ;
        RECT 130.255 213.480 130.485 213.770 ;
        RECT 130.300 212.200 130.440 213.480 ;
        RECT 130.255 211.910 130.485 212.200 ;
        RECT 130.300 210.100 130.440 211.910 ;
        RECT 130.640 211.685 130.780 213.915 ;
        RECT 130.595 211.395 130.825 211.685 ;
        RECT 130.640 210.495 130.780 211.395 ;
        RECT 131.320 210.950 131.460 216.210 ;
        RECT 131.275 210.660 131.505 210.950 ;
        RECT 130.595 210.205 130.825 210.495 ;
        RECT 130.255 209.810 130.485 210.100 ;
        RECT 130.920 209.310 131.180 209.630 ;
        RECT 131.260 205.630 131.520 205.950 ;
        RECT 129.900 199.650 130.160 199.970 ;
        RECT 129.960 199.495 130.100 199.650 ;
        RECT 129.915 199.205 130.145 199.495 ;
        RECT 130.580 199.190 130.840 199.510 ;
        RECT 129.900 194.590 130.160 194.910 ;
        RECT 129.960 191.675 130.100 194.590 ;
        RECT 130.640 193.975 130.780 199.190 ;
        RECT 131.600 196.430 131.860 196.750 ;
        RECT 131.600 194.130 131.860 194.450 ;
        RECT 130.595 193.685 130.825 193.975 ;
        RECT 129.915 191.385 130.145 191.675 ;
        RECT 130.920 191.370 131.180 191.690 ;
        RECT 130.920 190.450 131.180 190.770 ;
        RECT 131.660 189.835 131.800 194.130 ;
        RECT 131.615 189.545 131.845 189.835 ;
        RECT 129.900 188.150 130.160 188.470 ;
        RECT 129.960 185.235 130.100 188.150 ;
        RECT 130.920 186.080 131.180 186.170 ;
        RECT 130.920 185.940 131.460 186.080 ;
        RECT 130.920 185.850 131.180 185.940 ;
        RECT 129.915 184.945 130.145 185.235 ;
        RECT 130.935 184.945 131.165 185.235 ;
        RECT 130.980 184.790 131.120 184.945 ;
        RECT 130.920 184.470 131.180 184.790 ;
        RECT 131.320 184.700 131.460 185.940 ;
        RECT 131.615 184.700 131.845 184.775 ;
        RECT 131.320 184.560 131.845 184.700 ;
        RECT 131.615 184.485 131.845 184.560 ;
        RECT 130.920 183.550 131.180 183.870 ;
        RECT 132.000 182.100 132.480 217.980 ;
        RECT 132.620 216.210 132.880 216.530 ;
        RECT 132.635 214.385 132.865 214.675 ;
        RECT 132.680 211.930 132.820 214.385 ;
        RECT 133.640 213.910 133.900 214.230 ;
        RECT 133.655 213.005 133.885 213.295 ;
        RECT 133.315 212.085 133.545 212.375 ;
        RECT 133.700 212.300 133.840 213.005 ;
        RECT 133.700 212.160 134.520 212.300 ;
        RECT 132.620 211.610 132.880 211.930 ;
        RECT 133.020 211.040 133.160 211.445 ;
        RECT 132.975 211.010 133.205 211.040 ;
        RECT 132.960 210.690 133.220 211.010 ;
        RECT 133.020 203.560 133.160 210.690 ;
        RECT 133.360 209.630 133.500 212.085 ;
        RECT 133.995 211.600 134.225 211.890 ;
        RECT 133.655 211.205 133.885 211.495 ;
        RECT 133.700 210.305 133.840 211.205 ;
        RECT 133.655 210.015 133.885 210.305 ;
        RECT 133.300 209.310 133.560 209.630 ;
        RECT 133.360 206.870 133.500 209.310 ;
        RECT 133.700 207.785 133.840 210.015 ;
        RECT 134.040 209.790 134.180 211.600 ;
        RECT 133.995 209.500 134.225 209.790 ;
        RECT 134.040 208.220 134.180 209.500 ;
        RECT 133.995 207.930 134.225 208.220 ;
        RECT 133.655 207.495 133.885 207.785 ;
        RECT 133.300 206.550 133.560 206.870 ;
        RECT 133.995 205.400 134.225 205.475 ;
        RECT 132.680 203.420 133.160 203.560 ;
        RECT 133.360 205.260 134.225 205.400 ;
        RECT 132.680 197.210 132.820 203.420 ;
        RECT 132.975 202.930 133.205 203.220 ;
        RECT 132.620 196.890 132.880 197.210 ;
        RECT 132.680 196.275 132.820 196.890 ;
        RECT 133.020 196.750 133.160 202.930 ;
        RECT 132.960 196.430 133.220 196.750 ;
        RECT 133.360 196.290 133.500 205.260 ;
        RECT 133.995 205.185 134.225 205.260 ;
        RECT 133.640 204.250 133.900 204.570 ;
        RECT 133.995 203.780 134.225 204.070 ;
        RECT 133.655 203.385 133.885 203.675 ;
        RECT 133.700 202.485 133.840 203.385 ;
        RECT 133.655 202.195 133.885 202.485 ;
        RECT 133.700 199.965 133.840 202.195 ;
        RECT 134.040 201.970 134.180 203.780 ;
        RECT 134.380 203.650 134.520 212.160 ;
        RECT 134.320 203.330 134.580 203.650 ;
        RECT 133.995 201.680 134.225 201.970 ;
        RECT 134.040 200.400 134.180 201.680 ;
        RECT 133.995 200.110 134.225 200.400 ;
        RECT 133.655 199.675 133.885 199.965 ;
        RECT 134.335 197.365 134.565 197.655 ;
        RECT 134.380 197.210 134.520 197.365 ;
        RECT 134.320 196.890 134.580 197.210 ;
        RECT 132.635 195.985 132.865 196.275 ;
        RECT 133.300 195.970 133.560 196.290 ;
        RECT 132.960 195.280 133.220 195.370 ;
        RECT 133.360 195.280 133.500 195.970 ;
        RECT 133.980 195.510 134.240 195.830 ;
        RECT 132.960 195.140 133.500 195.280 ;
        RECT 132.960 195.050 133.220 195.140 ;
        RECT 133.020 193.975 133.160 195.050 ;
        RECT 132.975 193.685 133.205 193.975 ;
        RECT 132.635 192.305 132.865 192.595 ;
        RECT 132.680 191.690 132.820 192.305 ;
        RECT 132.620 191.370 132.880 191.690 ;
        RECT 133.315 191.600 133.545 191.675 ;
        RECT 133.020 191.460 133.545 191.600 ;
        RECT 133.020 191.140 133.160 191.460 ;
        RECT 133.315 191.385 133.545 191.460 ;
        RECT 132.680 191.000 133.160 191.140 ;
        RECT 133.655 191.140 133.885 191.215 ;
        RECT 133.655 191.000 134.180 191.140 ;
        RECT 132.680 186.540 132.820 191.000 ;
        RECT 133.655 190.925 133.885 191.000 ;
        RECT 133.655 190.465 133.885 190.755 ;
        RECT 133.315 190.220 133.545 190.295 ;
        RECT 133.020 190.080 133.545 190.220 ;
        RECT 133.020 188.915 133.160 190.080 ;
        RECT 133.315 190.005 133.545 190.080 ;
        RECT 133.300 189.530 133.560 189.850 ;
        RECT 133.360 189.375 133.500 189.530 ;
        RECT 133.315 189.085 133.545 189.375 ;
        RECT 132.975 188.625 133.205 188.915 ;
        RECT 133.315 188.165 133.545 188.455 ;
        RECT 133.360 187.090 133.500 188.165 ;
        RECT 133.700 188.010 133.840 190.465 ;
        RECT 134.040 188.930 134.180 191.000 ;
        RECT 133.980 188.610 134.240 188.930 ;
        RECT 133.640 187.690 133.900 188.010 ;
        RECT 133.300 186.770 133.560 187.090 ;
        RECT 133.300 186.540 133.560 186.630 ;
        RECT 132.680 186.400 133.560 186.540 ;
        RECT 133.300 186.310 133.560 186.400 ;
        RECT 133.300 184.930 133.560 185.250 ;
        RECT 133.300 184.470 133.560 184.790 ;
        RECT 133.360 184.315 133.500 184.470 ;
        RECT 134.040 184.330 134.180 188.610 ;
        RECT 134.335 187.245 134.565 187.535 ;
        RECT 134.380 185.710 134.520 187.245 ;
        RECT 134.320 185.390 134.580 185.710 ;
        RECT 133.315 184.025 133.545 184.315 ;
        RECT 133.980 184.010 134.240 184.330 ;
        RECT 134.720 182.100 135.200 217.980 ;
        RECT 137.040 216.670 137.300 216.990 ;
        RECT 137.100 216.055 137.240 216.670 ;
        RECT 137.055 215.765 137.285 216.055 ;
        RECT 136.375 214.845 136.605 215.135 ;
        RECT 135.680 213.910 135.940 214.230 ;
        RECT 135.740 212.300 135.880 213.910 ;
        RECT 136.035 212.300 136.265 212.375 ;
        RECT 135.740 212.160 136.265 212.300 ;
        RECT 135.355 199.665 135.585 199.955 ;
        RECT 135.400 199.510 135.540 199.665 ;
        RECT 135.340 199.190 135.600 199.510 ;
        RECT 135.740 194.450 135.880 212.160 ;
        RECT 136.035 212.085 136.265 212.160 ;
        RECT 136.035 211.165 136.265 211.455 ;
        RECT 136.080 211.010 136.220 211.165 ;
        RECT 136.020 210.690 136.280 211.010 ;
        RECT 136.420 209.630 136.560 214.845 ;
        RECT 137.040 214.370 137.300 214.690 ;
        RECT 137.055 212.545 137.285 212.835 ;
        RECT 136.360 209.310 136.620 209.630 ;
        RECT 137.100 209.170 137.240 212.545 ;
        RECT 137.040 208.850 137.300 209.170 ;
        RECT 137.040 206.550 137.300 206.870 ;
        RECT 137.100 204.570 137.240 206.550 ;
        RECT 137.040 204.250 137.300 204.570 ;
        RECT 137.040 203.330 137.300 203.650 ;
        RECT 136.375 200.125 136.605 200.415 ;
        RECT 136.420 199.970 136.560 200.125 ;
        RECT 137.100 199.970 137.240 203.330 ;
        RECT 136.360 199.650 136.620 199.970 ;
        RECT 137.040 199.650 137.300 199.970 ;
        RECT 136.035 196.445 136.265 196.735 ;
        RECT 136.080 196.290 136.220 196.445 ;
        RECT 136.020 195.970 136.280 196.290 ;
        RECT 136.700 194.590 136.960 194.910 ;
        RECT 135.680 194.130 135.940 194.450 ;
        RECT 136.035 193.685 136.265 193.975 ;
        RECT 135.355 193.440 135.585 193.515 ;
        RECT 135.355 193.300 135.880 193.440 ;
        RECT 135.355 193.225 135.585 193.300 ;
        RECT 135.340 192.290 135.600 192.610 ;
        RECT 135.740 189.850 135.880 193.300 ;
        RECT 136.080 190.680 136.220 193.685 ;
        RECT 136.375 193.440 136.605 193.515 ;
        RECT 136.375 193.300 137.240 193.440 ;
        RECT 136.375 193.225 136.605 193.300 ;
        RECT 136.715 191.385 136.945 191.675 ;
        RECT 136.360 190.680 136.620 190.770 ;
        RECT 136.080 190.540 136.620 190.680 ;
        RECT 136.360 190.450 136.620 190.540 ;
        RECT 136.760 190.310 136.900 191.385 ;
        RECT 136.700 189.990 136.960 190.310 ;
        RECT 135.680 189.530 135.940 189.850 ;
        RECT 136.700 189.530 136.960 189.850 ;
        RECT 136.375 189.300 136.605 189.375 ;
        RECT 136.080 189.160 136.605 189.300 ;
        RECT 136.080 187.995 136.220 189.160 ;
        RECT 136.375 189.085 136.605 189.160 ;
        RECT 136.375 188.380 136.605 188.455 ;
        RECT 136.760 188.380 136.900 189.530 ;
        RECT 136.375 188.240 136.900 188.380 ;
        RECT 136.375 188.165 136.605 188.240 ;
        RECT 136.035 187.705 136.265 187.995 ;
        RECT 136.360 186.770 136.620 187.090 ;
        RECT 136.360 185.390 136.620 185.710 ;
        RECT 136.375 184.485 136.605 184.775 ;
        RECT 136.760 184.700 136.900 188.240 ;
        RECT 137.100 187.090 137.240 193.300 ;
        RECT 137.040 186.770 137.300 187.090 ;
        RECT 137.040 184.700 137.300 184.790 ;
        RECT 136.760 184.560 137.300 184.700 ;
        RECT 136.420 184.330 136.560 184.485 ;
        RECT 137.040 184.470 137.300 184.560 ;
        RECT 136.360 184.010 136.620 184.330 ;
        RECT 137.440 182.100 137.920 217.980 ;
        RECT 138.755 216.225 138.985 216.515 ;
        RECT 138.415 214.890 138.645 215.180 ;
        RECT 138.460 214.690 138.600 214.890 ;
        RECT 138.400 214.370 138.660 214.690 ;
        RECT 138.060 209.540 138.320 209.630 ;
        RECT 138.060 209.400 138.600 209.540 ;
        RECT 138.060 209.310 138.320 209.400 ;
        RECT 138.060 208.850 138.320 209.170 ;
        RECT 138.460 206.320 138.600 209.400 ;
        RECT 138.800 206.870 138.940 216.225 ;
        RECT 139.435 215.740 139.665 216.030 ;
        RECT 139.095 215.345 139.325 215.635 ;
        RECT 139.140 214.445 139.280 215.345 ;
        RECT 139.095 214.155 139.325 214.445 ;
        RECT 139.140 211.925 139.280 214.155 ;
        RECT 139.480 213.930 139.620 215.740 ;
        RECT 139.435 213.640 139.665 213.930 ;
        RECT 139.480 212.360 139.620 213.640 ;
        RECT 139.435 212.070 139.665 212.360 ;
        RECT 139.095 211.635 139.325 211.925 ;
        RECT 138.740 206.550 139.000 206.870 ;
        RECT 138.755 206.320 138.985 206.395 ;
        RECT 138.460 206.180 138.985 206.320 ;
        RECT 138.755 206.105 138.985 206.180 ;
        RECT 139.760 204.250 140.020 204.570 ;
        RECT 138.755 202.425 138.985 202.715 ;
        RECT 138.415 201.965 138.645 202.255 ;
        RECT 138.060 200.110 138.320 200.430 ;
        RECT 138.120 198.115 138.260 200.110 ;
        RECT 138.075 197.825 138.305 198.115 ;
        RECT 138.460 194.450 138.600 201.965 ;
        RECT 138.800 200.430 138.940 202.425 ;
        RECT 139.095 201.260 139.325 201.335 ;
        RECT 139.095 201.120 139.620 201.260 ;
        RECT 139.095 201.045 139.325 201.120 ;
        RECT 138.740 200.110 139.000 200.430 ;
        RECT 138.740 199.650 139.000 199.970 ;
        RECT 138.740 198.730 139.000 199.050 ;
        RECT 138.800 197.210 138.940 198.730 ;
        RECT 138.740 196.890 139.000 197.210 ;
        RECT 138.740 196.430 139.000 196.750 ;
        RECT 138.800 195.830 138.940 196.430 ;
        RECT 139.080 195.970 139.340 196.290 ;
        RECT 139.480 196.200 139.620 201.120 ;
        RECT 139.760 199.190 140.020 199.510 ;
        RECT 139.820 197.195 139.960 199.190 ;
        RECT 139.775 196.905 140.005 197.195 ;
        RECT 139.480 196.060 139.960 196.200 ;
        RECT 138.740 195.510 139.000 195.830 ;
        RECT 139.435 195.500 139.665 195.790 ;
        RECT 139.095 195.105 139.325 195.395 ;
        RECT 138.755 194.650 138.985 194.940 ;
        RECT 138.400 194.130 138.660 194.450 ;
        RECT 138.800 193.530 138.940 194.650 ;
        RECT 139.140 194.205 139.280 195.105 ;
        RECT 139.095 193.915 139.325 194.205 ;
        RECT 138.740 193.210 139.000 193.530 ;
        RECT 139.140 191.685 139.280 193.915 ;
        RECT 139.480 193.690 139.620 195.500 ;
        RECT 139.820 194.450 139.960 196.060 ;
        RECT 139.760 194.130 140.020 194.450 ;
        RECT 139.435 193.400 139.665 193.690 ;
        RECT 139.480 192.120 139.620 193.400 ;
        RECT 139.435 191.830 139.665 192.120 ;
        RECT 139.095 191.395 139.325 191.685 ;
        RECT 139.820 191.140 139.960 194.130 ;
        RECT 138.800 191.000 139.960 191.140 ;
        RECT 138.800 188.455 138.940 191.000 ;
        RECT 139.760 189.070 140.020 189.390 ;
        RECT 138.755 188.165 138.985 188.455 ;
        RECT 138.740 187.230 139.000 187.550 ;
        RECT 139.760 186.310 140.020 186.630 ;
        RECT 138.740 185.850 139.000 186.170 ;
        RECT 138.060 184.930 138.320 185.250 ;
        RECT 138.060 184.470 138.320 184.790 ;
        RECT 138.740 183.550 139.000 183.870 ;
        RECT 140.160 182.100 140.640 217.980 ;
        RECT 142.480 212.070 142.740 212.390 ;
        RECT 141.475 209.775 141.705 210.065 ;
        RECT 141.135 209.340 141.365 209.630 ;
        RECT 141.180 208.060 141.320 209.340 ;
        RECT 141.135 207.770 141.365 208.060 ;
        RECT 140.780 206.550 141.040 206.870 ;
        RECT 140.840 204.940 140.980 206.550 ;
        RECT 141.180 205.960 141.320 207.770 ;
        RECT 141.520 207.545 141.660 209.775 ;
        RECT 141.475 207.255 141.705 207.545 ;
        RECT 142.480 207.470 142.740 207.790 ;
        RECT 141.520 206.355 141.660 207.255 ;
        RECT 141.815 206.465 142.045 206.755 ;
        RECT 141.475 206.065 141.705 206.355 ;
        RECT 141.135 205.670 141.365 205.960 ;
        RECT 141.475 205.185 141.705 205.475 ;
        RECT 141.520 205.015 141.660 205.185 ;
        RECT 141.475 204.940 141.705 205.015 ;
        RECT 140.840 204.800 141.705 204.940 ;
        RECT 140.840 196.290 140.980 204.800 ;
        RECT 141.475 204.725 141.705 204.800 ;
        RECT 141.860 204.570 142.000 206.465 ;
        RECT 142.140 205.170 142.400 205.490 ;
        RECT 141.135 204.240 141.365 204.530 ;
        RECT 141.800 204.250 142.060 204.570 ;
        RECT 141.180 202.430 141.320 204.240 ;
        RECT 141.475 203.845 141.705 204.135 ;
        RECT 141.520 202.945 141.660 203.845 ;
        RECT 142.200 203.790 142.340 205.170 ;
        RECT 142.155 203.500 142.385 203.790 ;
        RECT 141.475 202.655 141.705 202.945 ;
        RECT 141.135 202.140 141.365 202.430 ;
        RECT 141.180 200.860 141.320 202.140 ;
        RECT 141.135 200.570 141.365 200.860 ;
        RECT 141.520 200.425 141.660 202.655 ;
        RECT 142.540 202.640 142.680 207.470 ;
        RECT 142.200 202.500 142.680 202.640 ;
        RECT 141.475 200.135 141.705 200.425 ;
        RECT 141.120 199.650 141.380 199.970 ;
        RECT 140.780 195.970 141.040 196.290 ;
        RECT 141.180 194.435 141.320 199.650 ;
        RECT 141.460 198.730 141.720 199.050 ;
        RECT 141.520 195.280 141.660 198.730 ;
        RECT 142.200 197.655 142.340 202.500 ;
        RECT 142.495 197.825 142.725 198.115 ;
        RECT 142.155 197.365 142.385 197.655 ;
        RECT 142.540 197.210 142.680 197.825 ;
        RECT 142.480 196.890 142.740 197.210 ;
        RECT 142.140 196.430 142.400 196.750 ;
        RECT 141.800 195.510 142.060 195.830 ;
        RECT 141.815 195.280 142.045 195.355 ;
        RECT 141.520 195.140 142.045 195.280 ;
        RECT 141.815 195.065 142.045 195.140 ;
        RECT 141.460 194.590 141.720 194.910 ;
        RECT 141.135 194.145 141.365 194.435 ;
        RECT 140.780 193.210 141.040 193.530 ;
        RECT 140.840 191.675 140.980 193.210 ;
        RECT 141.135 192.765 141.365 193.055 ;
        RECT 140.795 191.385 141.025 191.675 ;
        RECT 141.180 190.295 141.320 192.765 ;
        RECT 141.520 192.520 141.660 194.590 ;
        RECT 141.800 194.130 142.060 194.450 ;
        RECT 141.860 193.515 142.000 194.130 ;
        RECT 141.815 193.225 142.045 193.515 ;
        RECT 141.800 192.520 142.060 192.610 ;
        RECT 141.520 192.380 142.060 192.520 ;
        RECT 141.800 192.290 142.060 192.380 ;
        RECT 141.860 190.755 142.000 192.290 ;
        RECT 141.815 190.465 142.045 190.755 ;
        RECT 141.135 190.005 141.365 190.295 ;
        RECT 141.800 189.530 142.060 189.850 ;
        RECT 141.120 189.070 141.380 189.390 ;
        RECT 141.815 189.085 142.045 189.375 ;
        RECT 141.180 188.380 141.320 189.070 ;
        RECT 141.475 188.380 141.705 188.455 ;
        RECT 141.180 188.240 141.705 188.380 ;
        RECT 141.475 188.165 141.705 188.240 ;
        RECT 140.780 187.230 141.040 187.550 ;
        RECT 140.840 185.235 140.980 187.230 ;
        RECT 141.860 186.630 142.000 189.085 ;
        RECT 141.800 186.310 142.060 186.630 ;
        RECT 141.120 185.850 141.380 186.170 ;
        RECT 140.795 184.945 141.025 185.235 ;
        RECT 141.180 184.775 141.320 185.850 ;
        RECT 141.135 184.485 141.365 184.775 ;
        RECT 141.800 183.550 142.060 183.870 ;
        RECT 142.880 182.100 143.360 217.980 ;
        RECT 144.180 212.070 144.440 212.390 ;
        RECT 144.240 210.075 144.380 212.070 ;
        RECT 144.195 210.000 144.425 210.075 ;
        RECT 144.195 209.860 144.720 210.000 ;
        RECT 144.195 209.785 144.425 209.860 ;
        RECT 144.180 207.470 144.440 207.790 ;
        RECT 144.180 207.010 144.440 207.330 ;
        RECT 144.195 206.105 144.425 206.395 ;
        RECT 143.500 205.170 143.760 205.490 ;
        RECT 143.500 200.110 143.760 200.430 ;
        RECT 144.240 198.040 144.380 206.105 ;
        RECT 144.580 203.635 144.720 209.860 ;
        RECT 145.215 208.865 145.445 209.155 ;
        RECT 144.875 206.565 145.105 206.855 ;
        RECT 144.535 203.345 144.765 203.635 ;
        RECT 144.920 199.510 145.060 206.565 ;
        RECT 145.260 204.110 145.400 208.865 ;
        RECT 145.200 203.790 145.460 204.110 ;
        RECT 144.860 199.190 145.120 199.510 ;
        RECT 145.215 198.285 145.445 198.575 ;
        RECT 144.240 197.900 145.060 198.040 ;
        RECT 144.195 197.365 144.425 197.655 ;
        RECT 144.240 197.210 144.380 197.365 ;
        RECT 144.180 196.890 144.440 197.210 ;
        RECT 143.500 196.430 143.760 196.750 ;
        RECT 143.560 193.975 143.700 196.430 ;
        RECT 144.180 194.130 144.440 194.450 ;
        RECT 143.515 193.685 143.745 193.975 ;
        RECT 144.240 193.515 144.380 194.130 ;
        RECT 144.195 193.225 144.425 193.515 ;
        RECT 144.920 192.610 145.060 197.900 ;
        RECT 145.260 197.670 145.400 198.285 ;
        RECT 145.200 197.350 145.460 197.670 ;
        RECT 144.860 192.290 145.120 192.610 ;
        RECT 145.200 190.910 145.460 191.230 ;
        RECT 143.500 190.450 143.760 190.770 ;
        RECT 143.560 187.535 143.700 190.450 ;
        RECT 145.260 190.295 145.400 190.910 ;
        RECT 145.215 190.005 145.445 190.295 ;
        RECT 144.180 189.070 144.440 189.390 ;
        RECT 143.515 187.245 143.745 187.535 ;
        RECT 143.500 186.770 143.760 187.090 ;
        RECT 143.560 186.155 143.700 186.770 ;
        RECT 144.180 186.310 144.440 186.630 ;
        RECT 143.515 185.865 143.745 186.155 ;
        RECT 144.180 184.930 144.440 185.250 ;
        RECT 143.515 184.485 143.745 184.775 ;
        RECT 143.560 184.330 143.700 184.485 ;
        RECT 143.500 184.010 143.760 184.330 ;
        RECT 144.180 183.550 144.440 183.870 ;
        RECT 145.600 182.100 146.080 217.980 ;
        RECT 146.370 199.970 146.510 218.730 ;
        RECT 146.280 199.650 146.600 199.970 ;
        RECT 146.930 197.640 147.070 219.250 ;
        RECT 146.840 197.380 147.160 197.640 ;
        RECT 147.300 196.920 147.440 219.710 ;
        RECT 147.740 204.110 147.880 220.250 ;
        RECT 147.650 203.790 147.970 204.110 ;
        RECT 146.830 196.780 147.440 196.920 ;
        RECT 146.830 191.200 146.970 196.780 ;
        RECT 146.740 190.940 147.060 191.200 ;
        RECT 100.270 173.675 139.495 174.670 ;
        RECT 100.360 173.250 101.170 173.675 ;
        RECT 119.450 173.310 120.130 173.675 ;
        RECT 138.390 173.350 139.080 173.675 ;
        RECT 100.360 172.350 101.200 173.250 ;
        RECT 106.870 172.860 108.120 173.300 ;
        RECT 119.410 173.280 120.130 173.310 ;
        RECT 104.810 172.850 110.050 172.860 ;
        RECT 101.860 172.750 117.160 172.850 ;
        RECT 101.860 172.740 117.195 172.750 ;
        RECT 101.820 172.620 117.195 172.740 ;
        RECT 101.820 172.510 105.820 172.620 ;
        RECT 106.870 172.540 108.610 172.620 ;
        RECT 109.190 172.540 117.195 172.620 ;
        RECT 106.870 172.460 108.120 172.540 ;
        RECT 109.195 172.520 117.195 172.540 ;
        RECT 100.370 171.150 101.200 172.350 ;
        RECT 101.430 172.210 101.660 172.460 ;
        RECT 105.980 172.320 106.210 172.460 ;
        RECT 108.760 172.320 108.990 172.470 ;
        RECT 105.980 172.210 108.990 172.320 ;
        RECT 117.400 172.210 117.630 172.470 ;
        RECT 101.430 171.770 117.630 172.210 ;
        RECT 101.430 171.500 101.660 171.770 ;
        RECT 105.980 171.740 117.630 171.770 ;
        RECT 105.980 171.650 108.990 171.740 ;
        RECT 105.980 171.500 106.210 171.650 ;
        RECT 108.760 171.510 108.990 171.650 ;
        RECT 117.400 171.510 117.630 171.740 ;
        RECT 101.820 171.220 105.820 171.450 ;
        RECT 109.195 171.240 117.195 171.460 ;
        RECT 117.960 171.240 118.920 173.280 ;
        RECT 109.195 171.230 118.920 171.240 ;
        RECT 101.820 171.150 105.810 171.220 ;
        RECT 100.370 171.040 105.810 171.150 ;
        RECT 109.250 171.070 118.920 171.230 ;
        RECT 100.370 170.950 103.500 171.040 ;
        RECT 116.990 171.020 118.920 171.070 ;
        RECT 100.370 167.680 101.200 170.950 ;
        RECT 104.850 170.490 110.100 170.500 ;
        RECT 104.850 170.380 117.160 170.490 ;
        RECT 101.880 170.320 117.160 170.380 ;
        RECT 101.880 170.310 117.195 170.320 ;
        RECT 101.820 170.180 117.195 170.310 ;
        RECT 101.820 170.170 106.980 170.180 ;
        RECT 101.820 170.080 105.820 170.170 ;
        RECT 109.195 170.090 117.195 170.180 ;
        RECT 109.280 170.080 117.170 170.090 ;
        RECT 101.430 169.720 101.660 170.030 ;
        RECT 101.880 169.720 105.780 170.080 ;
        RECT 105.980 169.720 106.210 170.030 ;
        RECT 101.430 168.380 106.210 169.720 ;
        RECT 101.430 168.070 101.660 168.380 ;
        RECT 105.980 168.070 106.210 168.380 ;
        RECT 108.760 169.500 108.990 170.040 ;
        RECT 109.800 169.500 110.810 169.530 ;
        RECT 117.400 169.500 117.630 170.040 ;
        RECT 108.760 168.600 117.630 169.500 ;
        RECT 108.760 168.080 108.990 168.600 ;
        RECT 109.800 168.530 110.810 168.600 ;
        RECT 117.400 168.080 117.630 168.600 ;
        RECT 101.820 167.790 105.820 168.020 ;
        RECT 109.195 167.800 117.195 168.030 ;
        RECT 100.370 167.640 101.500 167.680 ;
        RECT 100.370 167.560 101.740 167.640 ;
        RECT 102.110 167.570 105.770 167.790 ;
        RECT 102.110 167.560 103.550 167.570 ;
        RECT 100.370 167.520 103.550 167.560 ;
        RECT 100.370 167.430 103.060 167.520 ;
        RECT 109.260 167.510 117.150 167.800 ;
        RECT 100.370 167.370 102.390 167.430 ;
        RECT 100.370 167.320 102.140 167.370 ;
        RECT 100.370 163.980 101.200 167.320 ;
        RECT 109.250 167.020 117.170 167.030 ;
        RECT 105.480 167.010 117.170 167.020 ;
        RECT 101.860 166.890 117.170 167.010 ;
        RECT 101.860 166.880 117.195 166.890 ;
        RECT 101.820 166.760 117.195 166.880 ;
        RECT 101.820 166.650 105.820 166.760 ;
        RECT 101.430 166.310 101.660 166.600 ;
        RECT 101.880 166.310 105.770 166.650 ;
        RECT 105.980 166.310 106.210 166.600 ;
        RECT 101.430 164.940 106.210 166.310 ;
        RECT 101.430 164.640 101.660 164.940 ;
        RECT 105.980 164.640 106.210 164.940 ;
        RECT 101.820 164.360 105.820 164.590 ;
        RECT 102.070 164.130 105.640 164.360 ;
        RECT 102.070 163.980 105.760 164.130 ;
        RECT 100.370 163.700 105.760 163.980 ;
        RECT 107.010 163.810 107.630 166.760 ;
        RECT 109.195 166.660 117.195 166.760 ;
        RECT 109.250 166.650 117.170 166.660 ;
        RECT 108.760 165.950 108.990 166.610 ;
        RECT 109.770 165.950 110.770 166.040 ;
        RECT 117.400 165.950 117.630 166.610 ;
        RECT 108.760 165.130 117.630 165.950 ;
        RECT 108.760 164.650 108.990 165.130 ;
        RECT 109.770 165.040 110.770 165.130 ;
        RECT 117.400 164.650 117.630 165.130 ;
        RECT 109.195 164.370 117.195 164.600 ;
        RECT 100.370 163.240 105.770 163.700 ;
        RECT 100.370 161.900 102.370 163.240 ;
        RECT 104.120 163.230 105.770 163.240 ;
        RECT 102.810 161.960 103.810 162.680 ;
        RECT 104.120 162.420 104.430 163.230 ;
        RECT 104.890 162.950 105.770 163.230 ;
        RECT 106.010 163.410 107.630 163.810 ;
        RECT 109.280 163.460 117.150 164.370 ;
        RECT 104.830 162.720 105.830 162.950 ;
        RECT 106.010 162.760 106.360 163.410 ;
        RECT 107.010 163.400 107.630 163.410 ;
        RECT 109.195 163.230 117.195 163.460 ;
        RECT 109.280 163.220 117.150 163.230 ;
        RECT 104.890 162.510 105.770 162.530 ;
        RECT 104.160 162.130 104.430 162.420 ;
        RECT 104.830 162.280 105.830 162.510 ;
        RECT 105.990 162.470 106.360 162.760 ;
        RECT 106.020 162.410 106.360 162.470 ;
        RECT 107.120 163.080 107.880 163.130 ;
        RECT 108.760 163.080 108.990 163.180 ;
        RECT 107.120 162.870 108.990 163.080 ;
        RECT 117.400 162.870 117.630 163.180 ;
        RECT 107.120 162.450 109.660 162.870 ;
        RECT 117.030 162.450 117.630 162.870 ;
        RECT 104.890 162.130 105.770 162.280 ;
        RECT 104.900 161.960 105.630 162.130 ;
        RECT 100.380 161.890 102.370 161.900 ;
        RECT 100.380 158.290 101.160 161.890 ;
        RECT 102.780 160.840 105.630 161.960 ;
        RECT 106.020 161.660 106.370 162.410 ;
        RECT 107.120 162.290 108.990 162.450 ;
        RECT 107.120 162.240 107.880 162.290 ;
        RECT 108.760 162.220 108.990 162.290 ;
        RECT 117.400 162.220 117.630 162.450 ;
        RECT 109.195 161.940 117.195 162.170 ;
        RECT 106.020 161.600 106.310 161.660 ;
        RECT 105.930 161.480 106.310 161.600 ;
        RECT 109.290 161.540 117.150 161.940 ;
        RECT 117.960 161.640 118.920 171.020 ;
        RECT 119.410 171.180 120.240 173.280 ;
        RECT 125.910 172.890 127.160 173.330 ;
        RECT 138.360 173.320 139.080 173.350 ;
        RECT 123.850 172.880 129.090 172.890 ;
        RECT 120.900 172.780 136.200 172.880 ;
        RECT 120.900 172.770 136.235 172.780 ;
        RECT 120.860 172.650 136.235 172.770 ;
        RECT 120.860 172.540 124.860 172.650 ;
        RECT 125.910 172.570 127.650 172.650 ;
        RECT 128.230 172.570 136.235 172.650 ;
        RECT 125.910 172.490 127.160 172.570 ;
        RECT 128.235 172.550 136.235 172.570 ;
        RECT 120.470 172.240 120.700 172.490 ;
        RECT 125.020 172.350 125.250 172.490 ;
        RECT 127.800 172.350 128.030 172.500 ;
        RECT 125.020 172.240 128.030 172.350 ;
        RECT 136.440 172.240 136.670 172.500 ;
        RECT 120.470 171.800 136.670 172.240 ;
        RECT 120.470 171.530 120.700 171.800 ;
        RECT 125.020 171.770 136.670 171.800 ;
        RECT 125.020 171.680 128.030 171.770 ;
        RECT 125.020 171.530 125.250 171.680 ;
        RECT 127.800 171.540 128.030 171.680 ;
        RECT 136.440 171.540 136.670 171.770 ;
        RECT 120.860 171.250 124.860 171.480 ;
        RECT 128.235 171.270 136.235 171.490 ;
        RECT 137.000 171.270 137.960 173.310 ;
        RECT 128.235 171.260 137.960 171.270 ;
        RECT 120.860 171.180 124.850 171.250 ;
        RECT 119.410 171.070 124.850 171.180 ;
        RECT 128.290 171.100 137.960 171.260 ;
        RECT 119.410 170.980 122.540 171.070 ;
        RECT 136.030 171.050 137.960 171.100 ;
        RECT 119.410 167.720 120.240 170.980 ;
        RECT 123.890 170.520 129.140 170.530 ;
        RECT 123.890 170.410 136.200 170.520 ;
        RECT 120.920 170.350 136.200 170.410 ;
        RECT 120.920 170.340 136.235 170.350 ;
        RECT 120.860 170.210 136.235 170.340 ;
        RECT 120.860 170.200 126.020 170.210 ;
        RECT 120.860 170.110 124.860 170.200 ;
        RECT 128.235 170.120 136.235 170.210 ;
        RECT 128.320 170.110 136.210 170.120 ;
        RECT 120.470 169.750 120.700 170.060 ;
        RECT 120.920 169.750 124.820 170.110 ;
        RECT 125.020 169.750 125.250 170.060 ;
        RECT 120.470 168.410 125.250 169.750 ;
        RECT 120.470 168.100 120.700 168.410 ;
        RECT 125.020 168.100 125.250 168.410 ;
        RECT 127.800 169.530 128.030 170.070 ;
        RECT 128.840 169.530 129.850 169.560 ;
        RECT 136.440 169.530 136.670 170.070 ;
        RECT 127.800 168.630 136.670 169.530 ;
        RECT 127.800 168.110 128.030 168.630 ;
        RECT 128.840 168.560 129.850 168.630 ;
        RECT 136.440 168.110 136.670 168.630 ;
        RECT 120.860 167.820 124.860 168.050 ;
        RECT 128.235 167.830 136.235 168.060 ;
        RECT 117.950 161.540 118.920 161.640 ;
        RECT 102.720 160.610 105.720 160.840 ;
        RECT 105.930 160.650 106.270 161.480 ;
        RECT 108.280 161.470 118.920 161.540 ;
        RECT 102.770 160.580 105.630 160.610 ;
        RECT 102.770 160.560 103.940 160.580 ;
        RECT 104.900 160.570 105.630 160.580 ;
        RECT 102.720 160.170 105.720 160.400 ;
        RECT 105.925 160.360 106.270 160.650 ;
        RECT 106.460 160.430 118.920 161.470 ;
        RECT 119.380 167.710 120.240 167.720 ;
        RECT 119.380 167.670 120.540 167.710 ;
        RECT 119.380 167.590 120.780 167.670 ;
        RECT 121.150 167.600 124.810 167.820 ;
        RECT 121.150 167.590 122.590 167.600 ;
        RECT 119.380 167.550 122.590 167.590 ;
        RECT 119.380 167.460 122.100 167.550 ;
        RECT 128.300 167.540 136.190 167.830 ;
        RECT 119.380 167.400 121.430 167.460 ;
        RECT 119.380 167.350 121.180 167.400 ;
        RECT 119.380 164.010 120.240 167.350 ;
        RECT 128.290 167.050 136.210 167.060 ;
        RECT 124.520 167.040 136.210 167.050 ;
        RECT 120.900 166.920 136.210 167.040 ;
        RECT 120.900 166.910 136.235 166.920 ;
        RECT 120.860 166.790 136.235 166.910 ;
        RECT 120.860 166.680 124.860 166.790 ;
        RECT 120.470 166.340 120.700 166.630 ;
        RECT 120.920 166.340 124.810 166.680 ;
        RECT 125.020 166.340 125.250 166.630 ;
        RECT 120.470 164.970 125.250 166.340 ;
        RECT 120.470 164.670 120.700 164.970 ;
        RECT 125.020 164.670 125.250 164.970 ;
        RECT 120.860 164.390 124.860 164.620 ;
        RECT 121.110 164.160 124.680 164.390 ;
        RECT 121.110 164.010 124.800 164.160 ;
        RECT 119.380 163.730 124.800 164.010 ;
        RECT 126.050 163.840 126.670 166.790 ;
        RECT 128.235 166.690 136.235 166.790 ;
        RECT 128.290 166.680 136.210 166.690 ;
        RECT 127.800 165.980 128.030 166.640 ;
        RECT 128.810 165.980 129.810 166.070 ;
        RECT 136.440 165.980 136.670 166.640 ;
        RECT 127.800 165.160 136.670 165.980 ;
        RECT 127.800 164.680 128.030 165.160 ;
        RECT 128.810 165.070 129.810 165.160 ;
        RECT 136.440 164.680 136.670 165.160 ;
        RECT 128.235 164.400 136.235 164.630 ;
        RECT 119.380 163.270 124.810 163.730 ;
        RECT 119.380 161.920 121.410 163.270 ;
        RECT 123.160 163.260 124.810 163.270 ;
        RECT 121.850 161.990 122.850 162.710 ;
        RECT 123.160 162.450 123.470 163.260 ;
        RECT 123.930 162.980 124.810 163.260 ;
        RECT 125.050 163.440 126.670 163.840 ;
        RECT 128.320 163.490 136.190 164.400 ;
        RECT 123.870 162.750 124.870 162.980 ;
        RECT 125.050 162.790 125.400 163.440 ;
        RECT 126.050 163.430 126.670 163.440 ;
        RECT 128.235 163.260 136.235 163.490 ;
        RECT 128.320 163.250 136.190 163.260 ;
        RECT 123.930 162.540 124.810 162.560 ;
        RECT 123.200 162.160 123.470 162.450 ;
        RECT 123.870 162.310 124.870 162.540 ;
        RECT 125.030 162.500 125.400 162.790 ;
        RECT 125.060 162.440 125.400 162.500 ;
        RECT 126.160 163.110 126.920 163.160 ;
        RECT 127.800 163.110 128.030 163.210 ;
        RECT 126.160 162.900 128.030 163.110 ;
        RECT 136.440 162.900 136.670 163.210 ;
        RECT 126.160 162.480 128.700 162.900 ;
        RECT 136.070 162.480 136.670 162.900 ;
        RECT 123.930 162.160 124.810 162.310 ;
        RECT 123.940 161.990 124.670 162.160 ;
        RECT 106.460 160.410 118.890 160.430 ;
        RECT 106.730 160.400 112.170 160.410 ;
        RECT 113.170 160.400 118.890 160.410 ;
        RECT 105.930 160.250 106.270 160.360 ;
        RECT 100.370 158.260 101.160 158.290 ;
        RECT 100.370 156.160 101.200 158.260 ;
        RECT 106.870 157.870 108.120 158.310 ;
        RECT 117.950 158.290 118.890 160.400 ;
        RECT 104.810 157.860 110.050 157.870 ;
        RECT 101.860 157.760 117.160 157.860 ;
        RECT 101.860 157.750 117.195 157.760 ;
        RECT 101.820 157.630 117.195 157.750 ;
        RECT 101.820 157.520 105.820 157.630 ;
        RECT 106.870 157.550 108.610 157.630 ;
        RECT 109.190 157.550 117.195 157.630 ;
        RECT 106.870 157.470 108.120 157.550 ;
        RECT 109.195 157.530 117.195 157.550 ;
        RECT 101.430 157.220 101.660 157.470 ;
        RECT 105.980 157.330 106.210 157.470 ;
        RECT 108.760 157.330 108.990 157.480 ;
        RECT 105.980 157.220 108.990 157.330 ;
        RECT 117.400 157.220 117.630 157.480 ;
        RECT 101.430 156.780 117.630 157.220 ;
        RECT 101.430 156.510 101.660 156.780 ;
        RECT 105.980 156.750 117.630 156.780 ;
        RECT 105.980 156.660 108.990 156.750 ;
        RECT 105.980 156.510 106.210 156.660 ;
        RECT 108.760 156.520 108.990 156.660 ;
        RECT 117.400 156.520 117.630 156.750 ;
        RECT 117.950 156.660 118.920 158.290 ;
        RECT 101.820 156.230 105.820 156.460 ;
        RECT 109.195 156.250 117.195 156.470 ;
        RECT 117.960 156.250 118.920 156.660 ;
        RECT 109.195 156.240 118.920 156.250 ;
        RECT 101.820 156.160 105.810 156.230 ;
        RECT 100.370 156.050 105.810 156.160 ;
        RECT 109.250 156.080 118.920 156.240 ;
        RECT 100.370 155.960 103.500 156.050 ;
        RECT 116.990 156.030 118.920 156.080 ;
        RECT 100.370 152.690 101.200 155.960 ;
        RECT 104.850 155.500 110.100 155.510 ;
        RECT 104.850 155.390 117.160 155.500 ;
        RECT 101.880 155.330 117.160 155.390 ;
        RECT 101.880 155.320 117.195 155.330 ;
        RECT 101.820 155.190 117.195 155.320 ;
        RECT 101.820 155.180 106.980 155.190 ;
        RECT 101.820 155.090 105.820 155.180 ;
        RECT 109.195 155.100 117.195 155.190 ;
        RECT 109.280 155.090 117.170 155.100 ;
        RECT 101.430 154.730 101.660 155.040 ;
        RECT 101.880 154.730 105.780 155.090 ;
        RECT 105.980 154.730 106.210 155.040 ;
        RECT 101.430 153.390 106.210 154.730 ;
        RECT 101.430 153.080 101.660 153.390 ;
        RECT 105.980 153.080 106.210 153.390 ;
        RECT 108.760 154.510 108.990 155.050 ;
        RECT 109.800 154.510 110.810 154.540 ;
        RECT 117.400 154.510 117.630 155.050 ;
        RECT 108.760 153.610 117.630 154.510 ;
        RECT 108.760 153.090 108.990 153.610 ;
        RECT 109.800 153.540 110.810 153.610 ;
        RECT 117.400 153.090 117.630 153.610 ;
        RECT 101.820 152.800 105.820 153.030 ;
        RECT 109.195 152.810 117.195 153.040 ;
        RECT 100.370 152.650 101.500 152.690 ;
        RECT 100.370 152.570 101.740 152.650 ;
        RECT 102.110 152.580 105.770 152.800 ;
        RECT 102.110 152.570 103.550 152.580 ;
        RECT 100.370 152.530 103.550 152.570 ;
        RECT 100.370 152.440 103.060 152.530 ;
        RECT 109.260 152.520 117.150 152.810 ;
        RECT 100.370 152.380 102.390 152.440 ;
        RECT 100.370 152.330 102.140 152.380 ;
        RECT 100.370 148.990 101.200 152.330 ;
        RECT 109.250 152.030 117.170 152.040 ;
        RECT 105.480 152.020 117.170 152.030 ;
        RECT 101.860 151.900 117.170 152.020 ;
        RECT 101.860 151.890 117.195 151.900 ;
        RECT 101.820 151.770 117.195 151.890 ;
        RECT 101.820 151.660 105.820 151.770 ;
        RECT 101.430 151.320 101.660 151.610 ;
        RECT 101.880 151.320 105.770 151.660 ;
        RECT 105.980 151.320 106.210 151.610 ;
        RECT 101.430 149.950 106.210 151.320 ;
        RECT 101.430 149.650 101.660 149.950 ;
        RECT 105.980 149.650 106.210 149.950 ;
        RECT 101.820 149.370 105.820 149.600 ;
        RECT 102.070 149.140 105.640 149.370 ;
        RECT 102.070 148.990 105.760 149.140 ;
        RECT 100.370 148.710 105.760 148.990 ;
        RECT 107.010 148.820 107.630 151.770 ;
        RECT 109.195 151.670 117.195 151.770 ;
        RECT 109.250 151.660 117.170 151.670 ;
        RECT 108.760 150.960 108.990 151.620 ;
        RECT 109.770 150.960 110.770 151.050 ;
        RECT 117.400 150.960 117.630 151.620 ;
        RECT 108.760 150.140 117.630 150.960 ;
        RECT 108.760 149.660 108.990 150.140 ;
        RECT 109.770 150.050 110.770 150.140 ;
        RECT 117.400 149.660 117.630 150.140 ;
        RECT 109.195 149.380 117.195 149.610 ;
        RECT 100.370 148.250 105.770 148.710 ;
        RECT 100.370 146.910 102.370 148.250 ;
        RECT 104.120 148.240 105.770 148.250 ;
        RECT 102.810 146.970 103.810 147.690 ;
        RECT 104.120 147.430 104.430 148.240 ;
        RECT 104.890 147.960 105.770 148.240 ;
        RECT 106.010 148.420 107.630 148.820 ;
        RECT 109.280 148.470 117.150 149.380 ;
        RECT 104.830 147.730 105.830 147.960 ;
        RECT 106.010 147.770 106.360 148.420 ;
        RECT 107.010 148.410 107.630 148.420 ;
        RECT 109.195 148.240 117.195 148.470 ;
        RECT 109.280 148.230 117.150 148.240 ;
        RECT 104.890 147.520 105.770 147.540 ;
        RECT 104.160 147.140 104.430 147.430 ;
        RECT 104.830 147.290 105.830 147.520 ;
        RECT 105.990 147.480 106.360 147.770 ;
        RECT 106.020 147.420 106.360 147.480 ;
        RECT 107.120 148.090 107.880 148.140 ;
        RECT 108.760 148.090 108.990 148.190 ;
        RECT 107.120 147.880 108.990 148.090 ;
        RECT 117.400 147.880 117.630 148.190 ;
        RECT 107.120 147.460 109.660 147.880 ;
        RECT 117.030 147.460 117.630 147.880 ;
        RECT 104.890 147.140 105.770 147.290 ;
        RECT 104.900 146.970 105.630 147.140 ;
        RECT 100.380 146.900 102.370 146.910 ;
        RECT 100.380 143.310 101.160 146.900 ;
        RECT 102.780 145.850 105.630 146.970 ;
        RECT 106.020 146.670 106.370 147.420 ;
        RECT 107.120 147.300 108.990 147.460 ;
        RECT 107.120 147.250 107.880 147.300 ;
        RECT 108.760 147.230 108.990 147.300 ;
        RECT 117.400 147.230 117.630 147.460 ;
        RECT 109.195 146.950 117.195 147.180 ;
        RECT 106.020 146.610 106.310 146.670 ;
        RECT 105.930 146.490 106.310 146.610 ;
        RECT 109.290 146.550 117.150 146.950 ;
        RECT 117.960 146.740 118.920 156.030 ;
        RECT 117.910 146.550 118.920 146.740 ;
        RECT 102.720 145.620 105.720 145.850 ;
        RECT 105.930 145.660 106.270 146.490 ;
        RECT 108.280 146.480 118.920 146.550 ;
        RECT 102.770 145.590 105.630 145.620 ;
        RECT 102.770 145.570 103.940 145.590 ;
        RECT 104.900 145.580 105.630 145.590 ;
        RECT 102.720 145.180 105.720 145.410 ;
        RECT 105.925 145.370 106.270 145.660 ;
        RECT 106.460 145.440 118.920 146.480 ;
        RECT 119.380 158.260 120.140 161.920 ;
        RECT 121.820 160.870 124.670 161.990 ;
        RECT 125.060 161.690 125.410 162.440 ;
        RECT 126.160 162.320 128.030 162.480 ;
        RECT 126.160 162.270 126.920 162.320 ;
        RECT 127.800 162.250 128.030 162.320 ;
        RECT 136.440 162.250 136.670 162.480 ;
        RECT 128.235 161.970 136.235 162.200 ;
        RECT 125.060 161.630 125.350 161.690 ;
        RECT 124.970 161.510 125.350 161.630 ;
        RECT 128.330 161.570 136.190 161.970 ;
        RECT 137.000 161.570 137.960 171.050 ;
        RECT 138.360 171.220 139.190 173.320 ;
        RECT 144.860 172.930 146.110 173.370 ;
        RECT 142.800 172.920 148.040 172.930 ;
        RECT 139.850 172.820 155.150 172.920 ;
        RECT 139.850 172.810 155.185 172.820 ;
        RECT 139.810 172.690 155.185 172.810 ;
        RECT 139.810 172.580 143.810 172.690 ;
        RECT 144.860 172.610 146.600 172.690 ;
        RECT 147.180 172.610 155.185 172.690 ;
        RECT 144.860 172.530 146.110 172.610 ;
        RECT 147.185 172.590 155.185 172.610 ;
        RECT 139.420 172.280 139.650 172.530 ;
        RECT 143.970 172.390 144.200 172.530 ;
        RECT 146.750 172.390 146.980 172.540 ;
        RECT 143.970 172.280 146.980 172.390 ;
        RECT 155.390 172.280 155.620 172.540 ;
        RECT 139.420 171.840 155.620 172.280 ;
        RECT 139.420 171.570 139.650 171.840 ;
        RECT 143.970 171.810 155.620 171.840 ;
        RECT 143.970 171.720 146.980 171.810 ;
        RECT 143.970 171.570 144.200 171.720 ;
        RECT 146.750 171.580 146.980 171.720 ;
        RECT 155.390 171.580 155.620 171.810 ;
        RECT 139.810 171.290 143.810 171.520 ;
        RECT 147.185 171.310 155.185 171.530 ;
        RECT 155.950 171.310 156.910 173.350 ;
        RECT 147.185 171.300 156.910 171.310 ;
        RECT 139.810 171.220 143.800 171.290 ;
        RECT 138.360 171.110 143.800 171.220 ;
        RECT 147.240 171.140 156.910 171.300 ;
        RECT 138.360 171.020 141.490 171.110 ;
        RECT 154.980 171.090 156.910 171.140 ;
        RECT 138.360 167.750 139.190 171.020 ;
        RECT 142.840 170.560 148.090 170.570 ;
        RECT 142.840 170.450 155.150 170.560 ;
        RECT 139.870 170.390 155.150 170.450 ;
        RECT 139.870 170.380 155.185 170.390 ;
        RECT 139.810 170.250 155.185 170.380 ;
        RECT 139.810 170.240 144.970 170.250 ;
        RECT 139.810 170.150 143.810 170.240 ;
        RECT 147.185 170.160 155.185 170.250 ;
        RECT 147.270 170.150 155.160 170.160 ;
        RECT 139.420 169.790 139.650 170.100 ;
        RECT 139.870 169.790 143.770 170.150 ;
        RECT 143.970 169.790 144.200 170.100 ;
        RECT 139.420 168.450 144.200 169.790 ;
        RECT 139.420 168.140 139.650 168.450 ;
        RECT 143.970 168.140 144.200 168.450 ;
        RECT 146.750 169.570 146.980 170.110 ;
        RECT 147.790 169.570 148.800 169.600 ;
        RECT 155.390 169.570 155.620 170.110 ;
        RECT 146.750 168.670 155.620 169.570 ;
        RECT 146.750 168.150 146.980 168.670 ;
        RECT 147.790 168.600 148.800 168.670 ;
        RECT 155.390 168.150 155.620 168.670 ;
        RECT 139.810 167.860 143.810 168.090 ;
        RECT 147.185 167.870 155.185 168.100 ;
        RECT 138.360 167.710 139.490 167.750 ;
        RECT 138.360 167.630 139.730 167.710 ;
        RECT 140.100 167.640 143.760 167.860 ;
        RECT 140.100 167.630 141.540 167.640 ;
        RECT 138.360 167.590 141.540 167.630 ;
        RECT 138.360 167.500 141.050 167.590 ;
        RECT 147.250 167.580 155.140 167.870 ;
        RECT 138.360 167.440 140.380 167.500 ;
        RECT 138.360 167.390 140.130 167.440 ;
        RECT 138.360 164.050 139.190 167.390 ;
        RECT 147.240 167.090 155.160 167.100 ;
        RECT 143.470 167.080 155.160 167.090 ;
        RECT 139.850 166.960 155.160 167.080 ;
        RECT 139.850 166.950 155.185 166.960 ;
        RECT 139.810 166.830 155.185 166.950 ;
        RECT 139.810 166.720 143.810 166.830 ;
        RECT 139.420 166.380 139.650 166.670 ;
        RECT 139.870 166.380 143.760 166.720 ;
        RECT 143.970 166.380 144.200 166.670 ;
        RECT 139.420 165.010 144.200 166.380 ;
        RECT 139.420 164.710 139.650 165.010 ;
        RECT 143.970 164.710 144.200 165.010 ;
        RECT 139.810 164.430 143.810 164.660 ;
        RECT 140.060 164.200 143.630 164.430 ;
        RECT 140.060 164.050 143.750 164.200 ;
        RECT 138.360 163.770 143.750 164.050 ;
        RECT 145.000 163.880 145.620 166.830 ;
        RECT 147.185 166.730 155.185 166.830 ;
        RECT 147.240 166.720 155.160 166.730 ;
        RECT 146.750 166.020 146.980 166.680 ;
        RECT 147.760 166.020 148.760 166.110 ;
        RECT 155.390 166.020 155.620 166.680 ;
        RECT 146.750 165.200 155.620 166.020 ;
        RECT 146.750 164.720 146.980 165.200 ;
        RECT 147.760 165.110 148.760 165.200 ;
        RECT 155.390 164.720 155.620 165.200 ;
        RECT 147.185 164.440 155.185 164.670 ;
        RECT 138.360 163.310 143.760 163.770 ;
        RECT 138.360 161.970 140.360 163.310 ;
        RECT 142.110 163.300 143.760 163.310 ;
        RECT 140.800 162.030 141.800 162.750 ;
        RECT 142.110 162.490 142.420 163.300 ;
        RECT 142.880 163.020 143.760 163.300 ;
        RECT 144.000 163.480 145.620 163.880 ;
        RECT 147.270 163.530 155.140 164.440 ;
        RECT 142.820 162.790 143.820 163.020 ;
        RECT 144.000 162.830 144.350 163.480 ;
        RECT 145.000 163.470 145.620 163.480 ;
        RECT 147.185 163.300 155.185 163.530 ;
        RECT 147.270 163.290 155.140 163.300 ;
        RECT 142.880 162.580 143.760 162.600 ;
        RECT 142.150 162.200 142.420 162.490 ;
        RECT 142.820 162.350 143.820 162.580 ;
        RECT 143.980 162.540 144.350 162.830 ;
        RECT 144.010 162.480 144.350 162.540 ;
        RECT 145.110 163.150 145.870 163.200 ;
        RECT 146.750 163.150 146.980 163.250 ;
        RECT 145.110 162.940 146.980 163.150 ;
        RECT 155.390 162.940 155.620 163.250 ;
        RECT 145.110 162.520 147.650 162.940 ;
        RECT 155.020 162.520 155.620 162.940 ;
        RECT 142.880 162.200 143.760 162.350 ;
        RECT 142.890 162.030 143.620 162.200 ;
        RECT 121.760 160.640 124.760 160.870 ;
        RECT 124.970 160.680 125.310 161.510 ;
        RECT 127.320 161.500 137.960 161.570 ;
        RECT 121.810 160.610 124.670 160.640 ;
        RECT 121.810 160.590 122.980 160.610 ;
        RECT 123.940 160.600 124.670 160.610 ;
        RECT 121.760 160.200 124.760 160.430 ;
        RECT 124.965 160.390 125.310 160.680 ;
        RECT 125.500 160.440 137.960 161.500 ;
        RECT 125.770 160.430 131.210 160.440 ;
        RECT 132.210 160.430 137.960 160.440 ;
        RECT 124.970 160.280 125.310 160.390 ;
        RECT 119.380 156.160 120.240 158.260 ;
        RECT 125.910 157.870 127.160 158.310 ;
        RECT 137.020 158.290 137.960 160.430 ;
        RECT 138.440 161.960 140.360 161.970 ;
        RECT 138.440 158.290 139.160 161.960 ;
        RECT 140.770 160.910 143.620 162.030 ;
        RECT 144.010 161.730 144.360 162.480 ;
        RECT 145.110 162.360 146.980 162.520 ;
        RECT 145.110 162.310 145.870 162.360 ;
        RECT 146.750 162.290 146.980 162.360 ;
        RECT 155.390 162.290 155.620 162.520 ;
        RECT 147.185 162.010 155.185 162.240 ;
        RECT 144.010 161.670 144.300 161.730 ;
        RECT 143.920 161.550 144.300 161.670 ;
        RECT 147.280 161.610 155.140 162.010 ;
        RECT 155.950 161.610 156.910 171.090 ;
        RECT 140.710 160.680 143.710 160.910 ;
        RECT 143.920 160.720 144.260 161.550 ;
        RECT 146.270 161.540 156.910 161.610 ;
        RECT 140.760 160.650 143.620 160.680 ;
        RECT 140.760 160.630 141.930 160.650 ;
        RECT 142.890 160.640 143.620 160.650 ;
        RECT 140.710 160.240 143.710 160.470 ;
        RECT 143.915 160.430 144.260 160.720 ;
        RECT 144.450 161.460 156.910 161.540 ;
        RECT 144.450 160.480 156.940 161.460 ;
        RECT 144.720 160.470 150.160 160.480 ;
        RECT 151.160 160.470 156.940 160.480 ;
        RECT 143.920 160.320 144.260 160.430 ;
        RECT 123.850 157.860 129.090 157.870 ;
        RECT 120.900 157.760 136.200 157.860 ;
        RECT 120.900 157.750 136.235 157.760 ;
        RECT 120.860 157.630 136.235 157.750 ;
        RECT 120.860 157.520 124.860 157.630 ;
        RECT 125.910 157.550 127.650 157.630 ;
        RECT 128.230 157.550 136.235 157.630 ;
        RECT 125.910 157.470 127.160 157.550 ;
        RECT 128.235 157.530 136.235 157.550 ;
        RECT 120.470 157.220 120.700 157.470 ;
        RECT 125.020 157.330 125.250 157.470 ;
        RECT 127.800 157.330 128.030 157.480 ;
        RECT 125.020 157.220 128.030 157.330 ;
        RECT 136.440 157.220 136.670 157.480 ;
        RECT 120.470 156.780 136.670 157.220 ;
        RECT 120.470 156.510 120.700 156.780 ;
        RECT 125.020 156.750 136.670 156.780 ;
        RECT 125.020 156.660 128.030 156.750 ;
        RECT 125.020 156.510 125.250 156.660 ;
        RECT 127.800 156.520 128.030 156.660 ;
        RECT 136.440 156.520 136.670 156.750 ;
        RECT 120.860 156.230 124.860 156.460 ;
        RECT 128.235 156.250 136.235 156.470 ;
        RECT 137.000 156.250 137.960 158.290 ;
        RECT 128.235 156.240 137.960 156.250 ;
        RECT 120.860 156.160 124.850 156.230 ;
        RECT 119.380 156.050 124.850 156.160 ;
        RECT 128.290 156.080 137.960 156.240 ;
        RECT 119.380 155.960 122.540 156.050 ;
        RECT 136.030 156.030 137.960 156.080 ;
        RECT 119.380 152.690 120.240 155.960 ;
        RECT 123.890 155.500 129.140 155.510 ;
        RECT 123.890 155.390 136.200 155.500 ;
        RECT 120.920 155.330 136.200 155.390 ;
        RECT 120.920 155.320 136.235 155.330 ;
        RECT 120.860 155.190 136.235 155.320 ;
        RECT 120.860 155.180 126.020 155.190 ;
        RECT 120.860 155.090 124.860 155.180 ;
        RECT 128.235 155.100 136.235 155.190 ;
        RECT 128.320 155.090 136.210 155.100 ;
        RECT 120.470 154.730 120.700 155.040 ;
        RECT 120.920 154.730 124.820 155.090 ;
        RECT 125.020 154.730 125.250 155.040 ;
        RECT 120.470 153.390 125.250 154.730 ;
        RECT 120.470 153.080 120.700 153.390 ;
        RECT 125.020 153.080 125.250 153.390 ;
        RECT 127.800 154.510 128.030 155.050 ;
        RECT 128.840 154.510 129.850 154.540 ;
        RECT 136.440 154.510 136.670 155.050 ;
        RECT 127.800 153.610 136.670 154.510 ;
        RECT 127.800 153.090 128.030 153.610 ;
        RECT 128.840 153.540 129.850 153.610 ;
        RECT 136.440 153.090 136.670 153.610 ;
        RECT 120.860 152.800 124.860 153.030 ;
        RECT 128.235 152.810 136.235 153.040 ;
        RECT 119.380 152.650 120.540 152.690 ;
        RECT 119.380 152.570 120.780 152.650 ;
        RECT 121.150 152.580 124.810 152.800 ;
        RECT 121.150 152.570 122.590 152.580 ;
        RECT 119.380 152.530 122.590 152.570 ;
        RECT 119.380 152.440 122.100 152.530 ;
        RECT 128.300 152.520 136.190 152.810 ;
        RECT 119.380 152.380 121.430 152.440 ;
        RECT 119.380 152.330 121.180 152.380 ;
        RECT 119.380 148.990 120.240 152.330 ;
        RECT 128.290 152.030 136.210 152.040 ;
        RECT 124.520 152.020 136.210 152.030 ;
        RECT 120.900 151.900 136.210 152.020 ;
        RECT 120.900 151.890 136.235 151.900 ;
        RECT 120.860 151.770 136.235 151.890 ;
        RECT 120.860 151.660 124.860 151.770 ;
        RECT 120.470 151.320 120.700 151.610 ;
        RECT 120.920 151.320 124.810 151.660 ;
        RECT 125.020 151.320 125.250 151.610 ;
        RECT 120.470 149.950 125.250 151.320 ;
        RECT 120.470 149.650 120.700 149.950 ;
        RECT 125.020 149.650 125.250 149.950 ;
        RECT 120.860 149.370 124.860 149.600 ;
        RECT 121.110 149.140 124.680 149.370 ;
        RECT 121.110 148.990 124.800 149.140 ;
        RECT 119.380 148.710 124.800 148.990 ;
        RECT 126.050 148.820 126.670 151.770 ;
        RECT 128.235 151.670 136.235 151.770 ;
        RECT 128.290 151.660 136.210 151.670 ;
        RECT 127.800 150.960 128.030 151.620 ;
        RECT 128.810 150.960 129.810 151.050 ;
        RECT 136.440 150.960 136.670 151.620 ;
        RECT 127.800 150.140 136.670 150.960 ;
        RECT 127.800 149.660 128.030 150.140 ;
        RECT 128.810 150.050 129.810 150.140 ;
        RECT 136.440 149.660 136.670 150.140 ;
        RECT 128.235 149.380 136.235 149.610 ;
        RECT 119.380 148.250 124.810 148.710 ;
        RECT 119.380 146.900 121.410 148.250 ;
        RECT 123.160 148.240 124.810 148.250 ;
        RECT 121.850 146.970 122.850 147.690 ;
        RECT 123.160 147.430 123.470 148.240 ;
        RECT 123.930 147.960 124.810 148.240 ;
        RECT 125.050 148.420 126.670 148.820 ;
        RECT 128.320 148.470 136.190 149.380 ;
        RECT 123.870 147.730 124.870 147.960 ;
        RECT 125.050 147.770 125.400 148.420 ;
        RECT 126.050 148.410 126.670 148.420 ;
        RECT 128.235 148.240 136.235 148.470 ;
        RECT 128.320 148.230 136.190 148.240 ;
        RECT 123.930 147.520 124.810 147.540 ;
        RECT 123.200 147.140 123.470 147.430 ;
        RECT 123.870 147.290 124.870 147.520 ;
        RECT 125.030 147.480 125.400 147.770 ;
        RECT 125.060 147.420 125.400 147.480 ;
        RECT 126.160 148.090 126.920 148.140 ;
        RECT 127.800 148.090 128.030 148.190 ;
        RECT 126.160 147.880 128.030 148.090 ;
        RECT 136.440 147.880 136.670 148.190 ;
        RECT 126.160 147.460 128.700 147.880 ;
        RECT 136.070 147.460 136.670 147.880 ;
        RECT 123.930 147.140 124.810 147.290 ;
        RECT 123.940 146.970 124.670 147.140 ;
        RECT 106.460 145.420 118.850 145.440 ;
        RECT 106.730 145.410 112.170 145.420 ;
        RECT 113.170 145.410 118.850 145.420 ;
        RECT 105.930 145.260 106.270 145.370 ;
        RECT 100.370 143.280 101.160 143.310 ;
        RECT 100.370 141.180 101.200 143.280 ;
        RECT 106.870 142.890 108.120 143.330 ;
        RECT 117.910 143.310 118.850 145.410 ;
        RECT 104.810 142.880 110.050 142.890 ;
        RECT 101.860 142.780 117.160 142.880 ;
        RECT 101.860 142.770 117.195 142.780 ;
        RECT 101.820 142.650 117.195 142.770 ;
        RECT 101.820 142.540 105.820 142.650 ;
        RECT 106.870 142.570 108.610 142.650 ;
        RECT 109.190 142.570 117.195 142.650 ;
        RECT 106.870 142.490 108.120 142.570 ;
        RECT 109.195 142.550 117.195 142.570 ;
        RECT 101.430 142.240 101.660 142.490 ;
        RECT 105.980 142.350 106.210 142.490 ;
        RECT 108.760 142.350 108.990 142.500 ;
        RECT 105.980 142.240 108.990 142.350 ;
        RECT 117.400 142.240 117.630 142.500 ;
        RECT 101.430 141.800 117.630 142.240 ;
        RECT 101.430 141.530 101.660 141.800 ;
        RECT 105.980 141.770 117.630 141.800 ;
        RECT 105.980 141.680 108.990 141.770 ;
        RECT 105.980 141.530 106.210 141.680 ;
        RECT 108.760 141.540 108.990 141.680 ;
        RECT 117.400 141.540 117.630 141.770 ;
        RECT 117.910 141.760 118.920 143.310 ;
        RECT 119.380 143.270 120.140 146.900 ;
        RECT 121.820 145.850 124.670 146.970 ;
        RECT 125.060 146.670 125.410 147.420 ;
        RECT 126.160 147.300 128.030 147.460 ;
        RECT 126.160 147.250 126.920 147.300 ;
        RECT 127.800 147.230 128.030 147.300 ;
        RECT 136.440 147.230 136.670 147.460 ;
        RECT 128.235 146.950 136.235 147.180 ;
        RECT 125.060 146.610 125.350 146.670 ;
        RECT 124.970 146.490 125.350 146.610 ;
        RECT 128.330 146.550 136.190 146.950 ;
        RECT 137.000 146.550 137.960 156.030 ;
        RECT 138.410 158.260 139.160 158.290 ;
        RECT 138.410 156.160 139.240 158.260 ;
        RECT 144.910 157.870 146.160 158.310 ;
        RECT 156.000 158.290 156.940 160.470 ;
        RECT 142.850 157.860 148.090 157.870 ;
        RECT 139.900 157.760 155.200 157.860 ;
        RECT 139.900 157.750 155.235 157.760 ;
        RECT 139.860 157.630 155.235 157.750 ;
        RECT 139.860 157.520 143.860 157.630 ;
        RECT 144.910 157.550 146.650 157.630 ;
        RECT 147.230 157.550 155.235 157.630 ;
        RECT 144.910 157.470 146.160 157.550 ;
        RECT 147.235 157.530 155.235 157.550 ;
        RECT 139.470 157.220 139.700 157.470 ;
        RECT 144.020 157.330 144.250 157.470 ;
        RECT 146.800 157.330 147.030 157.480 ;
        RECT 144.020 157.220 147.030 157.330 ;
        RECT 155.440 157.220 155.670 157.480 ;
        RECT 139.470 156.780 155.670 157.220 ;
        RECT 139.470 156.510 139.700 156.780 ;
        RECT 144.020 156.750 155.670 156.780 ;
        RECT 144.020 156.660 147.030 156.750 ;
        RECT 144.020 156.510 144.250 156.660 ;
        RECT 146.800 156.520 147.030 156.660 ;
        RECT 155.440 156.520 155.670 156.750 ;
        RECT 139.860 156.230 143.860 156.460 ;
        RECT 147.235 156.250 155.235 156.470 ;
        RECT 156.000 156.250 156.960 158.290 ;
        RECT 147.235 156.240 156.960 156.250 ;
        RECT 139.860 156.160 143.850 156.230 ;
        RECT 138.410 156.050 143.850 156.160 ;
        RECT 147.290 156.080 156.960 156.240 ;
        RECT 138.410 155.960 141.540 156.050 ;
        RECT 155.030 156.030 156.960 156.080 ;
        RECT 138.410 152.690 139.240 155.960 ;
        RECT 142.890 155.500 148.140 155.510 ;
        RECT 142.890 155.390 155.200 155.500 ;
        RECT 139.920 155.330 155.200 155.390 ;
        RECT 139.920 155.320 155.235 155.330 ;
        RECT 139.860 155.190 155.235 155.320 ;
        RECT 139.860 155.180 145.020 155.190 ;
        RECT 139.860 155.090 143.860 155.180 ;
        RECT 147.235 155.100 155.235 155.190 ;
        RECT 147.320 155.090 155.210 155.100 ;
        RECT 139.470 154.730 139.700 155.040 ;
        RECT 139.920 154.730 143.820 155.090 ;
        RECT 144.020 154.730 144.250 155.040 ;
        RECT 139.470 153.390 144.250 154.730 ;
        RECT 139.470 153.080 139.700 153.390 ;
        RECT 144.020 153.080 144.250 153.390 ;
        RECT 146.800 154.510 147.030 155.050 ;
        RECT 147.840 154.510 148.850 154.540 ;
        RECT 155.440 154.510 155.670 155.050 ;
        RECT 146.800 153.610 155.670 154.510 ;
        RECT 146.800 153.090 147.030 153.610 ;
        RECT 147.840 153.540 148.850 153.610 ;
        RECT 155.440 153.090 155.670 153.610 ;
        RECT 139.860 152.800 143.860 153.030 ;
        RECT 147.235 152.810 155.235 153.040 ;
        RECT 138.410 152.650 139.540 152.690 ;
        RECT 138.410 152.570 139.780 152.650 ;
        RECT 140.150 152.580 143.810 152.800 ;
        RECT 140.150 152.570 141.590 152.580 ;
        RECT 138.410 152.530 141.590 152.570 ;
        RECT 138.410 152.440 141.100 152.530 ;
        RECT 147.300 152.520 155.190 152.810 ;
        RECT 138.410 152.380 140.430 152.440 ;
        RECT 138.410 152.330 140.180 152.380 ;
        RECT 138.410 148.990 139.240 152.330 ;
        RECT 147.290 152.030 155.210 152.040 ;
        RECT 143.520 152.020 155.210 152.030 ;
        RECT 139.900 151.900 155.210 152.020 ;
        RECT 139.900 151.890 155.235 151.900 ;
        RECT 139.860 151.770 155.235 151.890 ;
        RECT 139.860 151.660 143.860 151.770 ;
        RECT 139.470 151.320 139.700 151.610 ;
        RECT 139.920 151.320 143.810 151.660 ;
        RECT 144.020 151.320 144.250 151.610 ;
        RECT 139.470 149.950 144.250 151.320 ;
        RECT 139.470 149.650 139.700 149.950 ;
        RECT 144.020 149.650 144.250 149.950 ;
        RECT 139.860 149.370 143.860 149.600 ;
        RECT 140.110 149.140 143.680 149.370 ;
        RECT 140.110 148.990 143.800 149.140 ;
        RECT 138.410 148.710 143.800 148.990 ;
        RECT 145.050 148.820 145.670 151.770 ;
        RECT 147.235 151.670 155.235 151.770 ;
        RECT 147.290 151.660 155.210 151.670 ;
        RECT 146.800 150.960 147.030 151.620 ;
        RECT 147.810 150.960 148.810 151.050 ;
        RECT 155.440 150.960 155.670 151.620 ;
        RECT 146.800 150.140 155.670 150.960 ;
        RECT 146.800 149.660 147.030 150.140 ;
        RECT 147.810 150.050 148.810 150.140 ;
        RECT 155.440 149.660 155.670 150.140 ;
        RECT 147.235 149.380 155.235 149.610 ;
        RECT 138.410 148.250 143.810 148.710 ;
        RECT 138.410 146.910 140.410 148.250 ;
        RECT 142.160 148.240 143.810 148.250 ;
        RECT 140.850 146.970 141.850 147.690 ;
        RECT 142.160 147.430 142.470 148.240 ;
        RECT 142.930 147.960 143.810 148.240 ;
        RECT 144.050 148.420 145.670 148.820 ;
        RECT 147.320 148.470 155.190 149.380 ;
        RECT 142.870 147.730 143.870 147.960 ;
        RECT 144.050 147.770 144.400 148.420 ;
        RECT 145.050 148.410 145.670 148.420 ;
        RECT 147.235 148.240 155.235 148.470 ;
        RECT 147.320 148.230 155.190 148.240 ;
        RECT 142.930 147.520 143.810 147.540 ;
        RECT 142.200 147.140 142.470 147.430 ;
        RECT 142.870 147.290 143.870 147.520 ;
        RECT 144.030 147.480 144.400 147.770 ;
        RECT 144.060 147.420 144.400 147.480 ;
        RECT 145.160 148.090 145.920 148.140 ;
        RECT 146.800 148.090 147.030 148.190 ;
        RECT 145.160 147.880 147.030 148.090 ;
        RECT 155.440 147.880 155.670 148.190 ;
        RECT 145.160 147.460 147.700 147.880 ;
        RECT 155.070 147.460 155.670 147.880 ;
        RECT 142.930 147.140 143.810 147.290 ;
        RECT 142.940 146.970 143.670 147.140 ;
        RECT 121.760 145.620 124.760 145.850 ;
        RECT 124.970 145.660 125.310 146.490 ;
        RECT 127.320 146.480 137.960 146.550 ;
        RECT 121.810 145.590 124.670 145.620 ;
        RECT 121.810 145.570 122.980 145.590 ;
        RECT 123.940 145.580 124.670 145.590 ;
        RECT 121.760 145.180 124.760 145.410 ;
        RECT 124.965 145.370 125.310 145.660 ;
        RECT 125.500 145.440 137.960 146.480 ;
        RECT 138.430 146.900 140.410 146.910 ;
        RECT 125.500 145.420 137.900 145.440 ;
        RECT 125.770 145.410 131.210 145.420 ;
        RECT 132.210 145.410 137.900 145.420 ;
        RECT 124.970 145.260 125.310 145.370 ;
        RECT 101.820 141.250 105.820 141.480 ;
        RECT 109.195 141.270 117.195 141.490 ;
        RECT 117.960 141.270 118.920 141.760 ;
        RECT 109.195 141.260 118.920 141.270 ;
        RECT 101.820 141.180 105.810 141.250 ;
        RECT 100.370 141.070 105.810 141.180 ;
        RECT 109.250 141.100 118.920 141.260 ;
        RECT 100.370 140.980 103.500 141.070 ;
        RECT 116.990 141.050 118.920 141.100 ;
        RECT 100.370 137.710 101.200 140.980 ;
        RECT 104.850 140.520 110.100 140.530 ;
        RECT 104.850 140.410 117.160 140.520 ;
        RECT 101.880 140.350 117.160 140.410 ;
        RECT 101.880 140.340 117.195 140.350 ;
        RECT 101.820 140.210 117.195 140.340 ;
        RECT 101.820 140.200 106.980 140.210 ;
        RECT 101.820 140.110 105.820 140.200 ;
        RECT 109.195 140.120 117.195 140.210 ;
        RECT 109.280 140.110 117.170 140.120 ;
        RECT 101.430 139.750 101.660 140.060 ;
        RECT 101.880 139.750 105.780 140.110 ;
        RECT 105.980 139.750 106.210 140.060 ;
        RECT 101.430 138.410 106.210 139.750 ;
        RECT 101.430 138.100 101.660 138.410 ;
        RECT 105.980 138.100 106.210 138.410 ;
        RECT 108.760 139.530 108.990 140.070 ;
        RECT 109.800 139.530 110.810 139.560 ;
        RECT 117.400 139.530 117.630 140.070 ;
        RECT 108.760 138.630 117.630 139.530 ;
        RECT 108.760 138.110 108.990 138.630 ;
        RECT 109.800 138.560 110.810 138.630 ;
        RECT 117.400 138.110 117.630 138.630 ;
        RECT 101.820 137.820 105.820 138.050 ;
        RECT 109.195 137.830 117.195 138.060 ;
        RECT 100.370 137.670 101.500 137.710 ;
        RECT 100.370 137.590 101.740 137.670 ;
        RECT 102.110 137.600 105.770 137.820 ;
        RECT 102.110 137.590 103.550 137.600 ;
        RECT 100.370 137.550 103.550 137.590 ;
        RECT 100.370 137.460 103.060 137.550 ;
        RECT 109.260 137.540 117.150 137.830 ;
        RECT 100.370 137.400 102.390 137.460 ;
        RECT 100.370 137.350 102.140 137.400 ;
        RECT 100.370 134.010 101.200 137.350 ;
        RECT 109.250 137.050 117.170 137.060 ;
        RECT 105.480 137.040 117.170 137.050 ;
        RECT 101.860 136.920 117.170 137.040 ;
        RECT 101.860 136.910 117.195 136.920 ;
        RECT 101.820 136.790 117.195 136.910 ;
        RECT 101.820 136.680 105.820 136.790 ;
        RECT 101.430 136.340 101.660 136.630 ;
        RECT 101.880 136.340 105.770 136.680 ;
        RECT 105.980 136.340 106.210 136.630 ;
        RECT 101.430 134.970 106.210 136.340 ;
        RECT 101.430 134.670 101.660 134.970 ;
        RECT 105.980 134.670 106.210 134.970 ;
        RECT 101.820 134.390 105.820 134.620 ;
        RECT 102.070 134.160 105.640 134.390 ;
        RECT 102.070 134.010 105.760 134.160 ;
        RECT 100.370 133.730 105.760 134.010 ;
        RECT 107.010 133.840 107.630 136.790 ;
        RECT 109.195 136.690 117.195 136.790 ;
        RECT 109.250 136.680 117.170 136.690 ;
        RECT 108.760 135.980 108.990 136.640 ;
        RECT 109.770 135.980 110.770 136.070 ;
        RECT 117.400 135.980 117.630 136.640 ;
        RECT 108.760 135.160 117.630 135.980 ;
        RECT 108.760 134.680 108.990 135.160 ;
        RECT 109.770 135.070 110.770 135.160 ;
        RECT 117.400 134.680 117.630 135.160 ;
        RECT 109.195 134.400 117.195 134.630 ;
        RECT 100.370 133.270 105.770 133.730 ;
        RECT 100.370 131.930 102.370 133.270 ;
        RECT 104.120 133.260 105.770 133.270 ;
        RECT 102.810 131.990 103.810 132.710 ;
        RECT 104.120 132.450 104.430 133.260 ;
        RECT 104.890 132.980 105.770 133.260 ;
        RECT 106.010 133.440 107.630 133.840 ;
        RECT 109.280 133.490 117.150 134.400 ;
        RECT 104.830 132.750 105.830 132.980 ;
        RECT 106.010 132.790 106.360 133.440 ;
        RECT 107.010 133.430 107.630 133.440 ;
        RECT 109.195 133.260 117.195 133.490 ;
        RECT 109.280 133.250 117.150 133.260 ;
        RECT 104.890 132.540 105.770 132.560 ;
        RECT 104.160 132.160 104.430 132.450 ;
        RECT 104.830 132.310 105.830 132.540 ;
        RECT 105.990 132.500 106.360 132.790 ;
        RECT 106.020 132.440 106.360 132.500 ;
        RECT 107.120 133.110 107.880 133.160 ;
        RECT 108.760 133.110 108.990 133.210 ;
        RECT 107.120 132.900 108.990 133.110 ;
        RECT 117.400 132.900 117.630 133.210 ;
        RECT 107.120 132.480 109.660 132.900 ;
        RECT 117.030 132.480 117.630 132.900 ;
        RECT 104.890 132.160 105.770 132.310 ;
        RECT 104.900 131.990 105.630 132.160 ;
        RECT 100.380 131.920 102.370 131.930 ;
        RECT 100.380 128.280 101.160 131.920 ;
        RECT 102.780 130.870 105.630 131.990 ;
        RECT 106.020 131.690 106.370 132.440 ;
        RECT 107.120 132.320 108.990 132.480 ;
        RECT 107.120 132.270 107.880 132.320 ;
        RECT 108.760 132.250 108.990 132.320 ;
        RECT 117.400 132.250 117.630 132.480 ;
        RECT 109.195 131.970 117.195 132.200 ;
        RECT 106.020 131.630 106.310 131.690 ;
        RECT 105.930 131.510 106.310 131.630 ;
        RECT 109.290 131.570 117.150 131.970 ;
        RECT 117.960 131.750 118.920 141.050 ;
        RECT 119.360 143.240 120.140 143.270 ;
        RECT 119.360 141.140 120.190 143.240 ;
        RECT 125.860 142.850 127.110 143.290 ;
        RECT 136.960 143.270 137.900 145.410 ;
        RECT 138.430 143.270 139.130 146.900 ;
        RECT 140.820 145.850 143.670 146.970 ;
        RECT 144.060 146.670 144.410 147.420 ;
        RECT 145.160 147.300 147.030 147.460 ;
        RECT 145.160 147.250 145.920 147.300 ;
        RECT 146.800 147.230 147.030 147.300 ;
        RECT 155.440 147.230 155.670 147.460 ;
        RECT 147.235 146.950 155.235 147.180 ;
        RECT 144.060 146.610 144.350 146.670 ;
        RECT 143.970 146.490 144.350 146.610 ;
        RECT 147.330 146.550 155.190 146.950 ;
        RECT 156.000 146.550 156.960 156.030 ;
        RECT 140.760 145.620 143.760 145.850 ;
        RECT 143.970 145.660 144.310 146.490 ;
        RECT 146.320 146.480 156.960 146.550 ;
        RECT 140.810 145.590 143.670 145.620 ;
        RECT 140.810 145.570 141.980 145.590 ;
        RECT 142.940 145.580 143.670 145.590 ;
        RECT 140.760 145.180 143.760 145.410 ;
        RECT 143.965 145.370 144.310 145.660 ;
        RECT 144.500 145.440 156.960 146.480 ;
        RECT 144.500 145.420 156.880 145.440 ;
        RECT 144.770 145.410 150.210 145.420 ;
        RECT 151.210 145.410 156.880 145.420 ;
        RECT 143.970 145.260 144.310 145.370 ;
        RECT 123.800 142.840 129.040 142.850 ;
        RECT 120.850 142.740 136.150 142.840 ;
        RECT 120.850 142.730 136.185 142.740 ;
        RECT 120.810 142.610 136.185 142.730 ;
        RECT 120.810 142.500 124.810 142.610 ;
        RECT 125.860 142.530 127.600 142.610 ;
        RECT 128.180 142.530 136.185 142.610 ;
        RECT 125.860 142.450 127.110 142.530 ;
        RECT 128.185 142.510 136.185 142.530 ;
        RECT 120.420 142.200 120.650 142.450 ;
        RECT 124.970 142.310 125.200 142.450 ;
        RECT 127.750 142.310 127.980 142.460 ;
        RECT 124.970 142.200 127.980 142.310 ;
        RECT 136.390 142.200 136.620 142.460 ;
        RECT 120.420 141.760 136.620 142.200 ;
        RECT 120.420 141.490 120.650 141.760 ;
        RECT 124.970 141.730 136.620 141.760 ;
        RECT 124.970 141.640 127.980 141.730 ;
        RECT 124.970 141.490 125.200 141.640 ;
        RECT 127.750 141.500 127.980 141.640 ;
        RECT 136.390 141.500 136.620 141.730 ;
        RECT 120.810 141.210 124.810 141.440 ;
        RECT 128.185 141.230 136.185 141.450 ;
        RECT 136.950 141.230 137.910 143.270 ;
        RECT 128.185 141.220 137.910 141.230 ;
        RECT 120.810 141.140 124.800 141.210 ;
        RECT 119.360 141.030 124.800 141.140 ;
        RECT 128.240 141.060 137.910 141.220 ;
        RECT 119.360 140.940 122.490 141.030 ;
        RECT 135.980 141.010 137.910 141.060 ;
        RECT 119.360 137.670 120.190 140.940 ;
        RECT 123.840 140.480 129.090 140.490 ;
        RECT 123.840 140.370 136.150 140.480 ;
        RECT 120.870 140.310 136.150 140.370 ;
        RECT 120.870 140.300 136.185 140.310 ;
        RECT 120.810 140.170 136.185 140.300 ;
        RECT 120.810 140.160 125.970 140.170 ;
        RECT 120.810 140.070 124.810 140.160 ;
        RECT 128.185 140.080 136.185 140.170 ;
        RECT 128.270 140.070 136.160 140.080 ;
        RECT 120.420 139.710 120.650 140.020 ;
        RECT 120.870 139.710 124.770 140.070 ;
        RECT 124.970 139.710 125.200 140.020 ;
        RECT 120.420 138.370 125.200 139.710 ;
        RECT 120.420 138.060 120.650 138.370 ;
        RECT 124.970 138.060 125.200 138.370 ;
        RECT 127.750 139.490 127.980 140.030 ;
        RECT 128.790 139.490 129.800 139.520 ;
        RECT 136.390 139.490 136.620 140.030 ;
        RECT 127.750 138.590 136.620 139.490 ;
        RECT 127.750 138.070 127.980 138.590 ;
        RECT 128.790 138.520 129.800 138.590 ;
        RECT 136.390 138.070 136.620 138.590 ;
        RECT 120.810 137.780 124.810 138.010 ;
        RECT 128.185 137.790 136.185 138.020 ;
        RECT 119.360 137.630 120.490 137.670 ;
        RECT 119.360 137.550 120.730 137.630 ;
        RECT 121.100 137.560 124.760 137.780 ;
        RECT 121.100 137.550 122.540 137.560 ;
        RECT 119.360 137.510 122.540 137.550 ;
        RECT 119.360 137.420 122.050 137.510 ;
        RECT 128.250 137.500 136.140 137.790 ;
        RECT 119.360 137.360 121.380 137.420 ;
        RECT 119.360 137.310 121.130 137.360 ;
        RECT 119.360 133.970 120.190 137.310 ;
        RECT 128.240 137.010 136.160 137.020 ;
        RECT 124.470 137.000 136.160 137.010 ;
        RECT 120.850 136.880 136.160 137.000 ;
        RECT 120.850 136.870 136.185 136.880 ;
        RECT 120.810 136.750 136.185 136.870 ;
        RECT 120.810 136.640 124.810 136.750 ;
        RECT 120.420 136.300 120.650 136.590 ;
        RECT 120.870 136.300 124.760 136.640 ;
        RECT 124.970 136.300 125.200 136.590 ;
        RECT 120.420 134.930 125.200 136.300 ;
        RECT 120.420 134.630 120.650 134.930 ;
        RECT 124.970 134.630 125.200 134.930 ;
        RECT 120.810 134.350 124.810 134.580 ;
        RECT 121.060 134.120 124.630 134.350 ;
        RECT 121.060 133.970 124.750 134.120 ;
        RECT 119.360 133.690 124.750 133.970 ;
        RECT 126.000 133.800 126.620 136.750 ;
        RECT 128.185 136.650 136.185 136.750 ;
        RECT 128.240 136.640 136.160 136.650 ;
        RECT 127.750 135.940 127.980 136.600 ;
        RECT 128.760 135.940 129.760 136.030 ;
        RECT 136.390 135.940 136.620 136.600 ;
        RECT 127.750 135.120 136.620 135.940 ;
        RECT 127.750 134.640 127.980 135.120 ;
        RECT 128.760 135.030 129.760 135.120 ;
        RECT 136.390 134.640 136.620 135.120 ;
        RECT 128.185 134.360 136.185 134.590 ;
        RECT 119.360 133.230 124.760 133.690 ;
        RECT 119.360 131.890 121.360 133.230 ;
        RECT 123.110 133.220 124.760 133.230 ;
        RECT 121.800 131.950 122.800 132.670 ;
        RECT 123.110 132.410 123.420 133.220 ;
        RECT 123.880 132.940 124.760 133.220 ;
        RECT 125.000 133.400 126.620 133.800 ;
        RECT 128.270 133.450 136.140 134.360 ;
        RECT 123.820 132.710 124.820 132.940 ;
        RECT 125.000 132.750 125.350 133.400 ;
        RECT 126.000 133.390 126.620 133.400 ;
        RECT 128.185 133.220 136.185 133.450 ;
        RECT 128.270 133.210 136.140 133.220 ;
        RECT 123.880 132.500 124.760 132.520 ;
        RECT 123.150 132.120 123.420 132.410 ;
        RECT 123.820 132.270 124.820 132.500 ;
        RECT 124.980 132.460 125.350 132.750 ;
        RECT 125.010 132.400 125.350 132.460 ;
        RECT 126.110 133.070 126.870 133.120 ;
        RECT 127.750 133.070 127.980 133.170 ;
        RECT 126.110 132.860 127.980 133.070 ;
        RECT 136.390 132.860 136.620 133.170 ;
        RECT 126.110 132.440 128.650 132.860 ;
        RECT 136.020 132.440 136.620 132.860 ;
        RECT 123.880 132.120 124.760 132.270 ;
        RECT 123.890 131.950 124.620 132.120 ;
        RECT 117.950 131.570 118.920 131.750 ;
        RECT 102.720 130.640 105.720 130.870 ;
        RECT 105.930 130.680 106.270 131.510 ;
        RECT 108.280 131.500 118.920 131.570 ;
        RECT 102.770 130.610 105.630 130.640 ;
        RECT 102.770 130.590 103.940 130.610 ;
        RECT 104.900 130.600 105.630 130.610 ;
        RECT 102.720 130.200 105.720 130.430 ;
        RECT 105.925 130.390 106.270 130.680 ;
        RECT 106.460 130.460 118.920 131.500 ;
        RECT 119.380 131.880 121.360 131.890 ;
        RECT 106.460 130.440 118.890 130.460 ;
        RECT 106.730 130.430 112.170 130.440 ;
        RECT 113.170 130.430 118.890 130.440 ;
        RECT 105.930 130.280 106.270 130.390 ;
        RECT 100.370 128.250 101.160 128.280 ;
        RECT 100.370 126.150 101.200 128.250 ;
        RECT 106.870 127.860 108.120 128.300 ;
        RECT 117.950 128.280 118.890 130.430 ;
        RECT 104.810 127.850 110.050 127.860 ;
        RECT 101.860 127.750 117.160 127.850 ;
        RECT 101.860 127.740 117.195 127.750 ;
        RECT 101.820 127.620 117.195 127.740 ;
        RECT 101.820 127.510 105.820 127.620 ;
        RECT 106.870 127.540 108.610 127.620 ;
        RECT 109.190 127.540 117.195 127.620 ;
        RECT 106.870 127.460 108.120 127.540 ;
        RECT 109.195 127.520 117.195 127.540 ;
        RECT 101.430 127.210 101.660 127.460 ;
        RECT 105.980 127.320 106.210 127.460 ;
        RECT 108.760 127.320 108.990 127.470 ;
        RECT 105.980 127.210 108.990 127.320 ;
        RECT 117.400 127.210 117.630 127.470 ;
        RECT 101.430 126.770 117.630 127.210 ;
        RECT 117.950 126.770 118.920 128.280 ;
        RECT 119.380 128.250 120.140 131.880 ;
        RECT 121.770 130.830 124.620 131.950 ;
        RECT 125.010 131.650 125.360 132.400 ;
        RECT 126.110 132.280 127.980 132.440 ;
        RECT 126.110 132.230 126.870 132.280 ;
        RECT 127.750 132.210 127.980 132.280 ;
        RECT 136.390 132.210 136.620 132.440 ;
        RECT 128.185 131.930 136.185 132.160 ;
        RECT 125.010 131.590 125.300 131.650 ;
        RECT 124.920 131.470 125.300 131.590 ;
        RECT 128.280 131.530 136.140 131.930 ;
        RECT 136.950 131.530 137.910 141.010 ;
        RECT 138.360 143.240 139.130 143.270 ;
        RECT 138.360 141.140 139.190 143.240 ;
        RECT 144.860 142.850 146.110 143.290 ;
        RECT 155.940 143.270 156.880 145.410 ;
        RECT 142.800 142.840 148.040 142.850 ;
        RECT 139.850 142.740 155.150 142.840 ;
        RECT 139.850 142.730 155.185 142.740 ;
        RECT 139.810 142.610 155.185 142.730 ;
        RECT 139.810 142.500 143.810 142.610 ;
        RECT 144.860 142.530 146.600 142.610 ;
        RECT 147.180 142.530 155.185 142.610 ;
        RECT 144.860 142.450 146.110 142.530 ;
        RECT 147.185 142.510 155.185 142.530 ;
        RECT 139.420 142.200 139.650 142.450 ;
        RECT 143.970 142.310 144.200 142.450 ;
        RECT 146.750 142.310 146.980 142.460 ;
        RECT 143.970 142.200 146.980 142.310 ;
        RECT 155.390 142.200 155.620 142.460 ;
        RECT 139.420 141.760 155.620 142.200 ;
        RECT 139.420 141.490 139.650 141.760 ;
        RECT 143.970 141.730 155.620 141.760 ;
        RECT 143.970 141.640 146.980 141.730 ;
        RECT 143.970 141.490 144.200 141.640 ;
        RECT 146.750 141.500 146.980 141.640 ;
        RECT 155.390 141.500 155.620 141.730 ;
        RECT 155.940 141.500 156.910 143.270 ;
        RECT 139.810 141.210 143.810 141.440 ;
        RECT 147.185 141.230 155.185 141.450 ;
        RECT 155.950 141.230 156.910 141.500 ;
        RECT 147.185 141.220 156.910 141.230 ;
        RECT 139.810 141.140 143.800 141.210 ;
        RECT 138.360 141.030 143.800 141.140 ;
        RECT 147.240 141.060 156.910 141.220 ;
        RECT 138.360 140.940 141.490 141.030 ;
        RECT 154.980 141.010 156.910 141.060 ;
        RECT 138.360 137.670 139.190 140.940 ;
        RECT 142.840 140.480 148.090 140.490 ;
        RECT 142.840 140.370 155.150 140.480 ;
        RECT 139.870 140.310 155.150 140.370 ;
        RECT 139.870 140.300 155.185 140.310 ;
        RECT 139.810 140.170 155.185 140.300 ;
        RECT 139.810 140.160 144.970 140.170 ;
        RECT 139.810 140.070 143.810 140.160 ;
        RECT 147.185 140.080 155.185 140.170 ;
        RECT 147.270 140.070 155.160 140.080 ;
        RECT 139.420 139.710 139.650 140.020 ;
        RECT 139.870 139.710 143.770 140.070 ;
        RECT 143.970 139.710 144.200 140.020 ;
        RECT 139.420 138.370 144.200 139.710 ;
        RECT 139.420 138.060 139.650 138.370 ;
        RECT 143.970 138.060 144.200 138.370 ;
        RECT 146.750 139.490 146.980 140.030 ;
        RECT 147.790 139.490 148.800 139.520 ;
        RECT 155.390 139.490 155.620 140.030 ;
        RECT 146.750 138.590 155.620 139.490 ;
        RECT 146.750 138.070 146.980 138.590 ;
        RECT 147.790 138.520 148.800 138.590 ;
        RECT 155.390 138.070 155.620 138.590 ;
        RECT 139.810 137.780 143.810 138.010 ;
        RECT 147.185 137.790 155.185 138.020 ;
        RECT 138.360 137.630 139.490 137.670 ;
        RECT 138.360 137.550 139.730 137.630 ;
        RECT 140.100 137.560 143.760 137.780 ;
        RECT 140.100 137.550 141.540 137.560 ;
        RECT 138.360 137.510 141.540 137.550 ;
        RECT 138.360 137.420 141.050 137.510 ;
        RECT 147.250 137.500 155.140 137.790 ;
        RECT 138.360 137.360 140.380 137.420 ;
        RECT 138.360 137.310 140.130 137.360 ;
        RECT 138.360 133.970 139.190 137.310 ;
        RECT 147.240 137.010 155.160 137.020 ;
        RECT 143.470 137.000 155.160 137.010 ;
        RECT 139.850 136.880 155.160 137.000 ;
        RECT 139.850 136.870 155.185 136.880 ;
        RECT 139.810 136.750 155.185 136.870 ;
        RECT 139.810 136.640 143.810 136.750 ;
        RECT 139.420 136.300 139.650 136.590 ;
        RECT 139.870 136.300 143.760 136.640 ;
        RECT 143.970 136.300 144.200 136.590 ;
        RECT 139.420 134.930 144.200 136.300 ;
        RECT 139.420 134.630 139.650 134.930 ;
        RECT 143.970 134.630 144.200 134.930 ;
        RECT 139.810 134.350 143.810 134.580 ;
        RECT 140.060 134.120 143.630 134.350 ;
        RECT 140.060 133.970 143.750 134.120 ;
        RECT 138.360 133.690 143.750 133.970 ;
        RECT 145.000 133.800 145.620 136.750 ;
        RECT 147.185 136.650 155.185 136.750 ;
        RECT 147.240 136.640 155.160 136.650 ;
        RECT 146.750 135.940 146.980 136.600 ;
        RECT 147.760 135.940 148.760 136.030 ;
        RECT 155.390 135.940 155.620 136.600 ;
        RECT 146.750 135.120 155.620 135.940 ;
        RECT 146.750 134.640 146.980 135.120 ;
        RECT 147.760 135.030 148.760 135.120 ;
        RECT 155.390 134.640 155.620 135.120 ;
        RECT 147.185 134.360 155.185 134.590 ;
        RECT 138.360 133.230 143.760 133.690 ;
        RECT 138.360 131.890 140.360 133.230 ;
        RECT 142.110 133.220 143.760 133.230 ;
        RECT 140.800 131.950 141.800 132.670 ;
        RECT 142.110 132.410 142.420 133.220 ;
        RECT 142.880 132.940 143.760 133.220 ;
        RECT 144.000 133.400 145.620 133.800 ;
        RECT 147.270 133.450 155.140 134.360 ;
        RECT 142.820 132.710 143.820 132.940 ;
        RECT 144.000 132.750 144.350 133.400 ;
        RECT 145.000 133.390 145.620 133.400 ;
        RECT 147.185 133.220 155.185 133.450 ;
        RECT 147.270 133.210 155.140 133.220 ;
        RECT 142.880 132.500 143.760 132.520 ;
        RECT 142.150 132.120 142.420 132.410 ;
        RECT 142.820 132.270 143.820 132.500 ;
        RECT 143.980 132.460 144.350 132.750 ;
        RECT 144.010 132.400 144.350 132.460 ;
        RECT 145.110 133.070 145.870 133.120 ;
        RECT 146.750 133.070 146.980 133.170 ;
        RECT 145.110 132.860 146.980 133.070 ;
        RECT 155.390 132.860 155.620 133.170 ;
        RECT 145.110 132.440 147.650 132.860 ;
        RECT 155.020 132.440 155.620 132.860 ;
        RECT 142.880 132.120 143.760 132.270 ;
        RECT 142.890 131.950 143.620 132.120 ;
        RECT 121.710 130.600 124.710 130.830 ;
        RECT 124.920 130.640 125.260 131.470 ;
        RECT 127.270 131.460 137.910 131.530 ;
        RECT 121.760 130.570 124.620 130.600 ;
        RECT 121.760 130.550 122.930 130.570 ;
        RECT 123.890 130.560 124.620 130.570 ;
        RECT 121.710 130.160 124.710 130.390 ;
        RECT 124.915 130.350 125.260 130.640 ;
        RECT 125.450 130.420 137.910 131.460 ;
        RECT 138.430 131.880 140.360 131.890 ;
        RECT 125.450 130.400 137.900 130.420 ;
        RECT 125.720 130.390 131.160 130.400 ;
        RECT 132.160 130.390 137.900 130.400 ;
        RECT 124.920 130.240 125.260 130.350 ;
        RECT 101.430 126.500 101.660 126.770 ;
        RECT 105.980 126.740 117.630 126.770 ;
        RECT 105.980 126.650 108.990 126.740 ;
        RECT 105.980 126.500 106.210 126.650 ;
        RECT 108.760 126.510 108.990 126.650 ;
        RECT 117.400 126.510 117.630 126.740 ;
        RECT 101.820 126.220 105.820 126.450 ;
        RECT 109.195 126.240 117.195 126.460 ;
        RECT 117.960 126.240 118.920 126.770 ;
        RECT 109.195 126.230 118.920 126.240 ;
        RECT 101.820 126.150 105.810 126.220 ;
        RECT 100.370 126.040 105.810 126.150 ;
        RECT 109.250 126.070 118.920 126.230 ;
        RECT 100.370 125.950 103.500 126.040 ;
        RECT 116.990 126.020 118.920 126.070 ;
        RECT 100.370 122.680 101.200 125.950 ;
        RECT 104.850 125.490 110.100 125.500 ;
        RECT 104.850 125.380 117.160 125.490 ;
        RECT 101.880 125.320 117.160 125.380 ;
        RECT 101.880 125.310 117.195 125.320 ;
        RECT 101.820 125.180 117.195 125.310 ;
        RECT 101.820 125.170 106.980 125.180 ;
        RECT 101.820 125.080 105.820 125.170 ;
        RECT 109.195 125.090 117.195 125.180 ;
        RECT 109.280 125.080 117.170 125.090 ;
        RECT 101.430 124.720 101.660 125.030 ;
        RECT 101.880 124.720 105.780 125.080 ;
        RECT 105.980 124.720 106.210 125.030 ;
        RECT 101.430 123.380 106.210 124.720 ;
        RECT 101.430 123.070 101.660 123.380 ;
        RECT 105.980 123.070 106.210 123.380 ;
        RECT 108.760 124.500 108.990 125.040 ;
        RECT 109.800 124.500 110.810 124.530 ;
        RECT 117.400 124.500 117.630 125.040 ;
        RECT 108.760 123.600 117.630 124.500 ;
        RECT 108.760 123.080 108.990 123.600 ;
        RECT 109.800 123.530 110.810 123.600 ;
        RECT 117.400 123.080 117.630 123.600 ;
        RECT 101.820 122.790 105.820 123.020 ;
        RECT 109.195 122.800 117.195 123.030 ;
        RECT 100.370 122.640 101.500 122.680 ;
        RECT 100.370 122.560 101.740 122.640 ;
        RECT 102.110 122.570 105.770 122.790 ;
        RECT 102.110 122.560 103.550 122.570 ;
        RECT 100.370 122.520 103.550 122.560 ;
        RECT 100.370 122.430 103.060 122.520 ;
        RECT 109.260 122.510 117.150 122.800 ;
        RECT 100.370 122.370 102.390 122.430 ;
        RECT 100.370 122.320 102.140 122.370 ;
        RECT 100.370 118.980 101.200 122.320 ;
        RECT 109.250 122.020 117.170 122.030 ;
        RECT 105.480 122.010 117.170 122.020 ;
        RECT 101.860 121.890 117.170 122.010 ;
        RECT 101.860 121.880 117.195 121.890 ;
        RECT 101.820 121.760 117.195 121.880 ;
        RECT 101.820 121.650 105.820 121.760 ;
        RECT 101.430 121.310 101.660 121.600 ;
        RECT 101.880 121.310 105.770 121.650 ;
        RECT 105.980 121.310 106.210 121.600 ;
        RECT 101.430 119.940 106.210 121.310 ;
        RECT 101.430 119.640 101.660 119.940 ;
        RECT 105.980 119.640 106.210 119.940 ;
        RECT 101.820 119.360 105.820 119.590 ;
        RECT 102.070 119.130 105.640 119.360 ;
        RECT 102.070 118.980 105.760 119.130 ;
        RECT 100.370 118.700 105.760 118.980 ;
        RECT 107.010 118.810 107.630 121.760 ;
        RECT 109.195 121.660 117.195 121.760 ;
        RECT 109.250 121.650 117.170 121.660 ;
        RECT 108.760 120.950 108.990 121.610 ;
        RECT 109.770 120.950 110.770 121.040 ;
        RECT 117.400 120.950 117.630 121.610 ;
        RECT 108.760 120.130 117.630 120.950 ;
        RECT 108.760 119.650 108.990 120.130 ;
        RECT 109.770 120.040 110.770 120.130 ;
        RECT 117.400 119.650 117.630 120.130 ;
        RECT 109.195 119.370 117.195 119.600 ;
        RECT 100.370 118.240 105.770 118.700 ;
        RECT 100.370 116.900 102.370 118.240 ;
        RECT 104.120 118.230 105.770 118.240 ;
        RECT 102.810 116.960 103.810 117.680 ;
        RECT 104.120 117.420 104.430 118.230 ;
        RECT 104.890 117.950 105.770 118.230 ;
        RECT 106.010 118.410 107.630 118.810 ;
        RECT 109.280 118.460 117.150 119.370 ;
        RECT 104.830 117.720 105.830 117.950 ;
        RECT 106.010 117.760 106.360 118.410 ;
        RECT 107.010 118.400 107.630 118.410 ;
        RECT 109.195 118.230 117.195 118.460 ;
        RECT 109.280 118.220 117.150 118.230 ;
        RECT 104.890 117.510 105.770 117.530 ;
        RECT 104.160 117.130 104.430 117.420 ;
        RECT 104.830 117.280 105.830 117.510 ;
        RECT 105.990 117.470 106.360 117.760 ;
        RECT 106.020 117.410 106.360 117.470 ;
        RECT 107.120 118.080 107.880 118.130 ;
        RECT 108.760 118.080 108.990 118.180 ;
        RECT 107.120 117.870 108.990 118.080 ;
        RECT 117.400 117.870 117.630 118.180 ;
        RECT 107.120 117.450 109.660 117.870 ;
        RECT 117.030 117.450 117.630 117.870 ;
        RECT 104.890 117.130 105.770 117.280 ;
        RECT 104.900 116.960 105.630 117.130 ;
        RECT 100.380 116.890 102.370 116.900 ;
        RECT 100.380 113.290 101.160 116.890 ;
        RECT 102.780 115.840 105.630 116.960 ;
        RECT 106.020 116.660 106.370 117.410 ;
        RECT 107.120 117.290 108.990 117.450 ;
        RECT 107.120 117.240 107.880 117.290 ;
        RECT 108.760 117.220 108.990 117.290 ;
        RECT 117.400 117.220 117.630 117.450 ;
        RECT 109.195 116.940 117.195 117.170 ;
        RECT 106.020 116.600 106.310 116.660 ;
        RECT 105.930 116.480 106.310 116.600 ;
        RECT 109.290 116.540 117.150 116.940 ;
        RECT 117.960 116.760 118.920 126.020 ;
        RECT 119.360 128.220 120.140 128.250 ;
        RECT 119.360 126.120 120.190 128.220 ;
        RECT 125.860 127.830 127.110 128.270 ;
        RECT 136.960 128.250 137.900 130.390 ;
        RECT 138.430 128.250 139.130 131.880 ;
        RECT 140.770 130.830 143.620 131.950 ;
        RECT 144.010 131.650 144.360 132.400 ;
        RECT 145.110 132.280 146.980 132.440 ;
        RECT 145.110 132.230 145.870 132.280 ;
        RECT 146.750 132.210 146.980 132.280 ;
        RECT 155.390 132.210 155.620 132.440 ;
        RECT 147.185 131.930 155.185 132.160 ;
        RECT 144.010 131.590 144.300 131.650 ;
        RECT 143.920 131.470 144.300 131.590 ;
        RECT 147.280 131.530 155.140 131.930 ;
        RECT 155.950 131.530 156.910 141.010 ;
        RECT 140.710 130.600 143.710 130.830 ;
        RECT 143.920 130.640 144.260 131.470 ;
        RECT 146.270 131.460 156.910 131.530 ;
        RECT 140.760 130.570 143.620 130.600 ;
        RECT 140.760 130.550 141.930 130.570 ;
        RECT 142.890 130.560 143.620 130.570 ;
        RECT 140.710 130.160 143.710 130.390 ;
        RECT 143.915 130.350 144.260 130.640 ;
        RECT 144.450 130.420 156.910 131.460 ;
        RECT 144.450 130.400 156.900 130.420 ;
        RECT 144.720 130.390 150.160 130.400 ;
        RECT 151.160 130.390 156.900 130.400 ;
        RECT 143.920 130.240 144.260 130.350 ;
        RECT 123.800 127.820 129.040 127.830 ;
        RECT 120.850 127.720 136.150 127.820 ;
        RECT 120.850 127.710 136.185 127.720 ;
        RECT 120.810 127.590 136.185 127.710 ;
        RECT 120.810 127.480 124.810 127.590 ;
        RECT 125.860 127.510 127.600 127.590 ;
        RECT 128.180 127.510 136.185 127.590 ;
        RECT 125.860 127.430 127.110 127.510 ;
        RECT 128.185 127.490 136.185 127.510 ;
        RECT 120.420 127.180 120.650 127.430 ;
        RECT 124.970 127.290 125.200 127.430 ;
        RECT 127.750 127.290 127.980 127.440 ;
        RECT 124.970 127.180 127.980 127.290 ;
        RECT 136.390 127.180 136.620 127.440 ;
        RECT 120.420 126.740 136.620 127.180 ;
        RECT 120.420 126.470 120.650 126.740 ;
        RECT 124.970 126.710 136.620 126.740 ;
        RECT 124.970 126.620 127.980 126.710 ;
        RECT 124.970 126.470 125.200 126.620 ;
        RECT 127.750 126.480 127.980 126.620 ;
        RECT 136.390 126.480 136.620 126.710 ;
        RECT 120.810 126.190 124.810 126.420 ;
        RECT 128.185 126.210 136.185 126.430 ;
        RECT 136.950 126.210 137.910 128.250 ;
        RECT 128.185 126.200 137.910 126.210 ;
        RECT 120.810 126.120 124.800 126.190 ;
        RECT 119.360 126.010 124.800 126.120 ;
        RECT 128.240 126.040 137.910 126.200 ;
        RECT 119.360 125.920 122.490 126.010 ;
        RECT 135.980 125.990 137.910 126.040 ;
        RECT 119.360 122.650 120.190 125.920 ;
        RECT 123.840 125.460 129.090 125.470 ;
        RECT 123.840 125.350 136.150 125.460 ;
        RECT 120.870 125.290 136.150 125.350 ;
        RECT 120.870 125.280 136.185 125.290 ;
        RECT 120.810 125.150 136.185 125.280 ;
        RECT 120.810 125.140 125.970 125.150 ;
        RECT 120.810 125.050 124.810 125.140 ;
        RECT 128.185 125.060 136.185 125.150 ;
        RECT 128.270 125.050 136.160 125.060 ;
        RECT 120.420 124.690 120.650 125.000 ;
        RECT 120.870 124.690 124.770 125.050 ;
        RECT 124.970 124.690 125.200 125.000 ;
        RECT 120.420 123.350 125.200 124.690 ;
        RECT 120.420 123.040 120.650 123.350 ;
        RECT 124.970 123.040 125.200 123.350 ;
        RECT 127.750 124.470 127.980 125.010 ;
        RECT 128.790 124.470 129.800 124.500 ;
        RECT 136.390 124.470 136.620 125.010 ;
        RECT 127.750 123.570 136.620 124.470 ;
        RECT 127.750 123.050 127.980 123.570 ;
        RECT 128.790 123.500 129.800 123.570 ;
        RECT 136.390 123.050 136.620 123.570 ;
        RECT 120.810 122.760 124.810 122.990 ;
        RECT 128.185 122.770 136.185 123.000 ;
        RECT 119.360 122.610 120.490 122.650 ;
        RECT 119.360 122.530 120.730 122.610 ;
        RECT 121.100 122.540 124.760 122.760 ;
        RECT 121.100 122.530 122.540 122.540 ;
        RECT 119.360 122.490 122.540 122.530 ;
        RECT 119.360 122.400 122.050 122.490 ;
        RECT 128.250 122.480 136.140 122.770 ;
        RECT 119.360 122.340 121.380 122.400 ;
        RECT 119.360 122.290 121.130 122.340 ;
        RECT 119.360 118.950 120.190 122.290 ;
        RECT 128.240 121.990 136.160 122.000 ;
        RECT 124.470 121.980 136.160 121.990 ;
        RECT 120.850 121.860 136.160 121.980 ;
        RECT 120.850 121.850 136.185 121.860 ;
        RECT 120.810 121.730 136.185 121.850 ;
        RECT 120.810 121.620 124.810 121.730 ;
        RECT 120.420 121.280 120.650 121.570 ;
        RECT 120.870 121.280 124.760 121.620 ;
        RECT 124.970 121.280 125.200 121.570 ;
        RECT 120.420 119.910 125.200 121.280 ;
        RECT 120.420 119.610 120.650 119.910 ;
        RECT 124.970 119.610 125.200 119.910 ;
        RECT 120.810 119.330 124.810 119.560 ;
        RECT 121.060 119.100 124.630 119.330 ;
        RECT 121.060 118.950 124.750 119.100 ;
        RECT 119.360 118.670 124.750 118.950 ;
        RECT 126.000 118.780 126.620 121.730 ;
        RECT 128.185 121.630 136.185 121.730 ;
        RECT 128.240 121.620 136.160 121.630 ;
        RECT 127.750 120.920 127.980 121.580 ;
        RECT 128.760 120.920 129.760 121.010 ;
        RECT 136.390 120.920 136.620 121.580 ;
        RECT 127.750 120.100 136.620 120.920 ;
        RECT 127.750 119.620 127.980 120.100 ;
        RECT 128.760 120.010 129.760 120.100 ;
        RECT 136.390 119.620 136.620 120.100 ;
        RECT 128.185 119.340 136.185 119.570 ;
        RECT 119.360 118.210 124.760 118.670 ;
        RECT 119.360 116.870 121.360 118.210 ;
        RECT 123.110 118.200 124.760 118.210 ;
        RECT 121.800 116.930 122.800 117.650 ;
        RECT 123.110 117.390 123.420 118.200 ;
        RECT 123.880 117.920 124.760 118.200 ;
        RECT 125.000 118.380 126.620 118.780 ;
        RECT 128.270 118.430 136.140 119.340 ;
        RECT 123.820 117.690 124.820 117.920 ;
        RECT 125.000 117.730 125.350 118.380 ;
        RECT 126.000 118.370 126.620 118.380 ;
        RECT 128.185 118.200 136.185 118.430 ;
        RECT 128.270 118.190 136.140 118.200 ;
        RECT 123.880 117.480 124.760 117.500 ;
        RECT 123.150 117.100 123.420 117.390 ;
        RECT 123.820 117.250 124.820 117.480 ;
        RECT 124.980 117.440 125.350 117.730 ;
        RECT 125.010 117.380 125.350 117.440 ;
        RECT 126.110 118.050 126.870 118.100 ;
        RECT 127.750 118.050 127.980 118.150 ;
        RECT 126.110 117.840 127.980 118.050 ;
        RECT 136.390 117.840 136.620 118.150 ;
        RECT 126.110 117.420 128.650 117.840 ;
        RECT 136.020 117.420 136.620 117.840 ;
        RECT 123.880 117.100 124.760 117.250 ;
        RECT 123.890 116.930 124.620 117.100 ;
        RECT 117.940 116.540 118.920 116.760 ;
        RECT 102.720 115.610 105.720 115.840 ;
        RECT 105.930 115.650 106.270 116.480 ;
        RECT 108.280 116.470 118.920 116.540 ;
        RECT 102.770 115.580 105.630 115.610 ;
        RECT 102.770 115.560 103.940 115.580 ;
        RECT 104.900 115.570 105.630 115.580 ;
        RECT 102.720 115.170 105.720 115.400 ;
        RECT 105.925 115.360 106.270 115.650 ;
        RECT 106.460 115.430 118.920 116.470 ;
        RECT 119.380 116.860 121.360 116.870 ;
        RECT 106.460 115.410 118.880 115.430 ;
        RECT 106.730 115.400 112.170 115.410 ;
        RECT 113.170 115.400 118.880 115.410 ;
        RECT 105.930 115.250 106.270 115.360 ;
        RECT 100.370 113.260 101.160 113.290 ;
        RECT 100.370 111.160 101.200 113.260 ;
        RECT 106.870 112.870 108.120 113.310 ;
        RECT 117.940 113.290 118.880 115.400 ;
        RECT 104.810 112.860 110.050 112.870 ;
        RECT 101.860 112.760 117.160 112.860 ;
        RECT 101.860 112.750 117.195 112.760 ;
        RECT 101.820 112.630 117.195 112.750 ;
        RECT 101.820 112.520 105.820 112.630 ;
        RECT 106.870 112.550 108.610 112.630 ;
        RECT 109.190 112.550 117.195 112.630 ;
        RECT 106.870 112.470 108.120 112.550 ;
        RECT 109.195 112.530 117.195 112.550 ;
        RECT 101.430 112.220 101.660 112.470 ;
        RECT 105.980 112.330 106.210 112.470 ;
        RECT 108.760 112.330 108.990 112.480 ;
        RECT 105.980 112.220 108.990 112.330 ;
        RECT 117.400 112.220 117.630 112.480 ;
        RECT 101.430 111.780 117.630 112.220 ;
        RECT 117.940 111.780 118.920 113.290 ;
        RECT 119.380 113.270 120.140 116.860 ;
        RECT 121.770 115.810 124.620 116.930 ;
        RECT 125.010 116.630 125.360 117.380 ;
        RECT 126.110 117.260 127.980 117.420 ;
        RECT 126.110 117.210 126.870 117.260 ;
        RECT 127.750 117.190 127.980 117.260 ;
        RECT 136.390 117.190 136.620 117.420 ;
        RECT 128.185 116.910 136.185 117.140 ;
        RECT 125.010 116.570 125.300 116.630 ;
        RECT 124.920 116.450 125.300 116.570 ;
        RECT 128.280 116.510 136.140 116.910 ;
        RECT 136.950 116.510 137.910 125.990 ;
        RECT 138.360 128.220 139.130 128.250 ;
        RECT 138.360 126.120 139.190 128.220 ;
        RECT 144.860 127.830 146.110 128.270 ;
        RECT 155.960 128.250 156.900 130.390 ;
        RECT 142.800 127.820 148.040 127.830 ;
        RECT 139.850 127.720 155.150 127.820 ;
        RECT 139.850 127.710 155.185 127.720 ;
        RECT 139.810 127.590 155.185 127.710 ;
        RECT 139.810 127.480 143.810 127.590 ;
        RECT 144.860 127.510 146.600 127.590 ;
        RECT 147.180 127.510 155.185 127.590 ;
        RECT 144.860 127.430 146.110 127.510 ;
        RECT 147.185 127.490 155.185 127.510 ;
        RECT 139.420 127.180 139.650 127.430 ;
        RECT 143.970 127.290 144.200 127.430 ;
        RECT 146.750 127.290 146.980 127.440 ;
        RECT 143.970 127.180 146.980 127.290 ;
        RECT 155.390 127.180 155.620 127.440 ;
        RECT 139.420 126.740 155.620 127.180 ;
        RECT 139.420 126.470 139.650 126.740 ;
        RECT 143.970 126.710 155.620 126.740 ;
        RECT 143.970 126.620 146.980 126.710 ;
        RECT 143.970 126.470 144.200 126.620 ;
        RECT 146.750 126.480 146.980 126.620 ;
        RECT 155.390 126.480 155.620 126.710 ;
        RECT 139.810 126.190 143.810 126.420 ;
        RECT 147.185 126.210 155.185 126.430 ;
        RECT 155.950 126.210 156.910 128.250 ;
        RECT 147.185 126.200 156.910 126.210 ;
        RECT 139.810 126.120 143.800 126.190 ;
        RECT 138.360 126.010 143.800 126.120 ;
        RECT 147.240 126.040 156.910 126.200 ;
        RECT 138.360 125.920 141.490 126.010 ;
        RECT 154.980 125.990 156.910 126.040 ;
        RECT 138.360 122.650 139.190 125.920 ;
        RECT 142.840 125.460 148.090 125.470 ;
        RECT 142.840 125.350 155.150 125.460 ;
        RECT 139.870 125.290 155.150 125.350 ;
        RECT 139.870 125.280 155.185 125.290 ;
        RECT 139.810 125.150 155.185 125.280 ;
        RECT 139.810 125.140 144.970 125.150 ;
        RECT 139.810 125.050 143.810 125.140 ;
        RECT 147.185 125.060 155.185 125.150 ;
        RECT 147.270 125.050 155.160 125.060 ;
        RECT 139.420 124.690 139.650 125.000 ;
        RECT 139.870 124.690 143.770 125.050 ;
        RECT 143.970 124.690 144.200 125.000 ;
        RECT 139.420 123.350 144.200 124.690 ;
        RECT 139.420 123.040 139.650 123.350 ;
        RECT 143.970 123.040 144.200 123.350 ;
        RECT 146.750 124.470 146.980 125.010 ;
        RECT 147.790 124.470 148.800 124.500 ;
        RECT 155.390 124.470 155.620 125.010 ;
        RECT 146.750 123.570 155.620 124.470 ;
        RECT 146.750 123.050 146.980 123.570 ;
        RECT 147.790 123.500 148.800 123.570 ;
        RECT 155.390 123.050 155.620 123.570 ;
        RECT 139.810 122.760 143.810 122.990 ;
        RECT 147.185 122.770 155.185 123.000 ;
        RECT 138.360 122.610 139.490 122.650 ;
        RECT 138.360 122.530 139.730 122.610 ;
        RECT 140.100 122.540 143.760 122.760 ;
        RECT 140.100 122.530 141.540 122.540 ;
        RECT 138.360 122.490 141.540 122.530 ;
        RECT 138.360 122.400 141.050 122.490 ;
        RECT 147.250 122.480 155.140 122.770 ;
        RECT 138.360 122.340 140.380 122.400 ;
        RECT 138.360 122.290 140.130 122.340 ;
        RECT 138.360 118.950 139.190 122.290 ;
        RECT 147.240 121.990 155.160 122.000 ;
        RECT 143.470 121.980 155.160 121.990 ;
        RECT 139.850 121.860 155.160 121.980 ;
        RECT 139.850 121.850 155.185 121.860 ;
        RECT 139.810 121.730 155.185 121.850 ;
        RECT 139.810 121.620 143.810 121.730 ;
        RECT 139.420 121.280 139.650 121.570 ;
        RECT 139.870 121.280 143.760 121.620 ;
        RECT 143.970 121.280 144.200 121.570 ;
        RECT 139.420 119.910 144.200 121.280 ;
        RECT 139.420 119.610 139.650 119.910 ;
        RECT 143.970 119.610 144.200 119.910 ;
        RECT 139.810 119.330 143.810 119.560 ;
        RECT 140.060 119.100 143.630 119.330 ;
        RECT 140.060 118.950 143.750 119.100 ;
        RECT 138.360 118.670 143.750 118.950 ;
        RECT 145.000 118.780 145.620 121.730 ;
        RECT 147.185 121.630 155.185 121.730 ;
        RECT 147.240 121.620 155.160 121.630 ;
        RECT 146.750 120.920 146.980 121.580 ;
        RECT 147.760 120.920 148.760 121.010 ;
        RECT 155.390 120.920 155.620 121.580 ;
        RECT 146.750 120.100 155.620 120.920 ;
        RECT 146.750 119.620 146.980 120.100 ;
        RECT 147.760 120.010 148.760 120.100 ;
        RECT 155.390 119.620 155.620 120.100 ;
        RECT 147.185 119.340 155.185 119.570 ;
        RECT 138.360 118.210 143.760 118.670 ;
        RECT 138.360 116.870 140.360 118.210 ;
        RECT 142.110 118.200 143.760 118.210 ;
        RECT 140.800 116.930 141.800 117.650 ;
        RECT 142.110 117.390 142.420 118.200 ;
        RECT 142.880 117.920 143.760 118.200 ;
        RECT 144.000 118.380 145.620 118.780 ;
        RECT 147.270 118.430 155.140 119.340 ;
        RECT 142.820 117.690 143.820 117.920 ;
        RECT 144.000 117.730 144.350 118.380 ;
        RECT 145.000 118.370 145.620 118.380 ;
        RECT 147.185 118.200 155.185 118.430 ;
        RECT 147.270 118.190 155.140 118.200 ;
        RECT 142.880 117.480 143.760 117.500 ;
        RECT 142.150 117.100 142.420 117.390 ;
        RECT 142.820 117.250 143.820 117.480 ;
        RECT 143.980 117.440 144.350 117.730 ;
        RECT 144.010 117.380 144.350 117.440 ;
        RECT 145.110 118.050 145.870 118.100 ;
        RECT 146.750 118.050 146.980 118.150 ;
        RECT 145.110 117.840 146.980 118.050 ;
        RECT 155.390 117.840 155.620 118.150 ;
        RECT 145.110 117.420 147.650 117.840 ;
        RECT 155.020 117.420 155.620 117.840 ;
        RECT 142.880 117.100 143.760 117.250 ;
        RECT 142.890 116.930 143.620 117.100 ;
        RECT 121.710 115.580 124.710 115.810 ;
        RECT 124.920 115.620 125.260 116.450 ;
        RECT 127.270 116.440 137.910 116.510 ;
        RECT 121.760 115.550 124.620 115.580 ;
        RECT 121.760 115.530 122.930 115.550 ;
        RECT 123.890 115.540 124.620 115.550 ;
        RECT 121.710 115.140 124.710 115.370 ;
        RECT 124.915 115.330 125.260 115.620 ;
        RECT 125.450 115.400 137.910 116.440 ;
        RECT 138.430 116.860 140.360 116.870 ;
        RECT 125.450 115.380 137.850 115.400 ;
        RECT 125.720 115.370 131.160 115.380 ;
        RECT 132.160 115.370 137.850 115.380 ;
        RECT 124.920 115.220 125.260 115.330 ;
        RECT 101.430 111.510 101.660 111.780 ;
        RECT 105.980 111.750 117.630 111.780 ;
        RECT 105.980 111.660 108.990 111.750 ;
        RECT 105.980 111.510 106.210 111.660 ;
        RECT 108.760 111.520 108.990 111.660 ;
        RECT 117.400 111.520 117.630 111.750 ;
        RECT 101.820 111.230 105.820 111.460 ;
        RECT 109.195 111.250 117.195 111.470 ;
        RECT 117.960 111.250 118.920 111.780 ;
        RECT 109.195 111.240 118.920 111.250 ;
        RECT 101.820 111.160 105.810 111.230 ;
        RECT 100.370 111.050 105.810 111.160 ;
        RECT 109.250 111.080 118.920 111.240 ;
        RECT 100.370 110.960 103.500 111.050 ;
        RECT 116.990 111.030 118.920 111.080 ;
        RECT 100.370 107.690 101.200 110.960 ;
        RECT 104.850 110.500 110.100 110.510 ;
        RECT 104.850 110.390 117.160 110.500 ;
        RECT 101.880 110.330 117.160 110.390 ;
        RECT 101.880 110.320 117.195 110.330 ;
        RECT 101.820 110.190 117.195 110.320 ;
        RECT 101.820 110.180 106.980 110.190 ;
        RECT 101.820 110.090 105.820 110.180 ;
        RECT 109.195 110.100 117.195 110.190 ;
        RECT 109.280 110.090 117.170 110.100 ;
        RECT 101.430 109.730 101.660 110.040 ;
        RECT 101.880 109.730 105.780 110.090 ;
        RECT 105.980 109.730 106.210 110.040 ;
        RECT 101.430 108.390 106.210 109.730 ;
        RECT 101.430 108.080 101.660 108.390 ;
        RECT 105.980 108.080 106.210 108.390 ;
        RECT 108.760 109.510 108.990 110.050 ;
        RECT 109.800 109.510 110.810 109.540 ;
        RECT 117.400 109.510 117.630 110.050 ;
        RECT 108.760 108.610 117.630 109.510 ;
        RECT 108.760 108.090 108.990 108.610 ;
        RECT 109.800 108.540 110.810 108.610 ;
        RECT 117.400 108.090 117.630 108.610 ;
        RECT 101.820 107.800 105.820 108.030 ;
        RECT 109.195 107.810 117.195 108.040 ;
        RECT 100.370 107.650 101.500 107.690 ;
        RECT 100.370 107.570 101.740 107.650 ;
        RECT 102.110 107.580 105.770 107.800 ;
        RECT 102.110 107.570 103.550 107.580 ;
        RECT 100.370 107.530 103.550 107.570 ;
        RECT 100.370 107.440 103.060 107.530 ;
        RECT 109.260 107.520 117.150 107.810 ;
        RECT 100.370 107.380 102.390 107.440 ;
        RECT 100.370 107.330 102.140 107.380 ;
        RECT 100.370 103.990 101.200 107.330 ;
        RECT 109.250 107.030 117.170 107.040 ;
        RECT 105.480 107.020 117.170 107.030 ;
        RECT 101.860 106.900 117.170 107.020 ;
        RECT 101.860 106.890 117.195 106.900 ;
        RECT 101.820 106.770 117.195 106.890 ;
        RECT 101.820 106.660 105.820 106.770 ;
        RECT 101.430 106.320 101.660 106.610 ;
        RECT 101.880 106.320 105.770 106.660 ;
        RECT 105.980 106.320 106.210 106.610 ;
        RECT 101.430 104.950 106.210 106.320 ;
        RECT 101.430 104.650 101.660 104.950 ;
        RECT 105.980 104.650 106.210 104.950 ;
        RECT 101.820 104.370 105.820 104.600 ;
        RECT 102.070 104.140 105.640 104.370 ;
        RECT 102.070 103.990 105.760 104.140 ;
        RECT 100.370 103.710 105.760 103.990 ;
        RECT 107.010 103.820 107.630 106.770 ;
        RECT 109.195 106.670 117.195 106.770 ;
        RECT 109.250 106.660 117.170 106.670 ;
        RECT 108.760 105.960 108.990 106.620 ;
        RECT 109.770 105.960 110.770 106.050 ;
        RECT 117.400 105.960 117.630 106.620 ;
        RECT 108.760 105.140 117.630 105.960 ;
        RECT 108.760 104.660 108.990 105.140 ;
        RECT 109.770 105.050 110.770 105.140 ;
        RECT 117.400 104.660 117.630 105.140 ;
        RECT 109.195 104.380 117.195 104.610 ;
        RECT 100.370 103.250 105.770 103.710 ;
        RECT 100.370 101.910 102.370 103.250 ;
        RECT 104.120 103.240 105.770 103.250 ;
        RECT 102.810 102.570 103.810 102.690 ;
        RECT 100.390 101.900 102.370 101.910 ;
        RECT 102.780 101.970 103.810 102.570 ;
        RECT 104.120 102.430 104.430 103.240 ;
        RECT 104.890 102.960 105.770 103.240 ;
        RECT 106.010 103.420 107.630 103.820 ;
        RECT 109.280 103.470 117.150 104.380 ;
        RECT 104.830 102.730 105.830 102.960 ;
        RECT 106.010 102.770 106.360 103.420 ;
        RECT 107.010 103.410 107.630 103.420 ;
        RECT 109.195 103.240 117.195 103.470 ;
        RECT 109.280 103.230 117.150 103.240 ;
        RECT 104.890 102.520 105.770 102.540 ;
        RECT 104.160 102.140 104.430 102.430 ;
        RECT 104.830 102.290 105.830 102.520 ;
        RECT 105.990 102.480 106.360 102.770 ;
        RECT 106.020 102.420 106.360 102.480 ;
        RECT 107.120 103.090 107.880 103.140 ;
        RECT 108.760 103.090 108.990 103.190 ;
        RECT 107.120 102.880 108.990 103.090 ;
        RECT 117.400 102.880 117.630 103.190 ;
        RECT 107.120 102.460 109.660 102.880 ;
        RECT 117.030 102.460 117.630 102.880 ;
        RECT 104.890 102.140 105.770 102.290 ;
        RECT 104.900 101.970 105.630 102.140 ;
        RECT 100.390 98.780 101.440 101.900 ;
        RECT 102.780 100.850 105.630 101.970 ;
        RECT 106.020 101.670 106.370 102.420 ;
        RECT 107.120 102.300 108.990 102.460 ;
        RECT 107.120 102.250 107.880 102.300 ;
        RECT 108.760 102.230 108.990 102.300 ;
        RECT 117.400 102.230 117.630 102.460 ;
        RECT 109.195 101.950 117.195 102.180 ;
        RECT 106.020 101.610 106.310 101.670 ;
        RECT 105.930 101.490 106.310 101.610 ;
        RECT 109.290 101.550 117.150 101.950 ;
        RECT 117.960 101.550 118.920 111.030 ;
        RECT 119.360 113.240 120.140 113.270 ;
        RECT 119.360 111.140 120.190 113.240 ;
        RECT 125.860 112.850 127.110 113.290 ;
        RECT 136.910 113.270 137.850 115.370 ;
        RECT 138.430 113.270 139.130 116.860 ;
        RECT 140.770 115.810 143.620 116.930 ;
        RECT 144.010 116.630 144.360 117.380 ;
        RECT 145.110 117.260 146.980 117.420 ;
        RECT 145.110 117.210 145.870 117.260 ;
        RECT 146.750 117.190 146.980 117.260 ;
        RECT 155.390 117.190 155.620 117.420 ;
        RECT 147.185 116.910 155.185 117.140 ;
        RECT 144.010 116.570 144.300 116.630 ;
        RECT 143.920 116.450 144.300 116.570 ;
        RECT 147.280 116.510 155.140 116.910 ;
        RECT 155.950 116.510 156.910 125.990 ;
        RECT 140.710 115.580 143.710 115.810 ;
        RECT 143.920 115.620 144.260 116.450 ;
        RECT 146.270 116.440 156.910 116.510 ;
        RECT 140.760 115.550 143.620 115.580 ;
        RECT 140.760 115.530 141.930 115.550 ;
        RECT 142.890 115.540 143.620 115.550 ;
        RECT 140.710 115.140 143.710 115.370 ;
        RECT 143.915 115.330 144.260 115.620 ;
        RECT 144.450 116.420 156.910 116.440 ;
        RECT 144.450 115.380 156.940 116.420 ;
        RECT 144.720 115.370 150.160 115.380 ;
        RECT 151.160 115.370 156.940 115.380 ;
        RECT 143.920 115.220 144.260 115.330 ;
        RECT 123.800 112.840 129.040 112.850 ;
        RECT 120.850 112.740 136.150 112.840 ;
        RECT 120.850 112.730 136.185 112.740 ;
        RECT 120.810 112.610 136.185 112.730 ;
        RECT 120.810 112.500 124.810 112.610 ;
        RECT 125.860 112.530 127.600 112.610 ;
        RECT 128.180 112.530 136.185 112.610 ;
        RECT 125.860 112.450 127.110 112.530 ;
        RECT 128.185 112.510 136.185 112.530 ;
        RECT 120.420 112.200 120.650 112.450 ;
        RECT 124.970 112.310 125.200 112.450 ;
        RECT 127.750 112.310 127.980 112.460 ;
        RECT 124.970 112.200 127.980 112.310 ;
        RECT 136.390 112.200 136.620 112.460 ;
        RECT 120.420 111.760 136.620 112.200 ;
        RECT 120.420 111.490 120.650 111.760 ;
        RECT 124.970 111.730 136.620 111.760 ;
        RECT 124.970 111.640 127.980 111.730 ;
        RECT 124.970 111.490 125.200 111.640 ;
        RECT 127.750 111.500 127.980 111.640 ;
        RECT 136.390 111.500 136.620 111.730 ;
        RECT 136.910 111.480 137.910 113.270 ;
        RECT 120.810 111.210 124.810 111.440 ;
        RECT 128.185 111.230 136.185 111.450 ;
        RECT 136.950 111.230 137.910 111.480 ;
        RECT 128.185 111.220 137.910 111.230 ;
        RECT 120.810 111.140 124.800 111.210 ;
        RECT 119.360 111.030 124.800 111.140 ;
        RECT 128.240 111.060 137.910 111.220 ;
        RECT 119.360 110.940 122.490 111.030 ;
        RECT 135.980 111.010 137.910 111.060 ;
        RECT 119.360 107.670 120.190 110.940 ;
        RECT 123.840 110.480 129.090 110.490 ;
        RECT 123.840 110.370 136.150 110.480 ;
        RECT 120.870 110.310 136.150 110.370 ;
        RECT 120.870 110.300 136.185 110.310 ;
        RECT 120.810 110.170 136.185 110.300 ;
        RECT 120.810 110.160 125.970 110.170 ;
        RECT 120.810 110.070 124.810 110.160 ;
        RECT 128.185 110.080 136.185 110.170 ;
        RECT 128.270 110.070 136.160 110.080 ;
        RECT 120.420 109.710 120.650 110.020 ;
        RECT 120.870 109.710 124.770 110.070 ;
        RECT 124.970 109.710 125.200 110.020 ;
        RECT 120.420 108.370 125.200 109.710 ;
        RECT 120.420 108.060 120.650 108.370 ;
        RECT 124.970 108.060 125.200 108.370 ;
        RECT 127.750 109.490 127.980 110.030 ;
        RECT 128.790 109.490 129.800 109.520 ;
        RECT 136.390 109.490 136.620 110.030 ;
        RECT 127.750 108.590 136.620 109.490 ;
        RECT 127.750 108.070 127.980 108.590 ;
        RECT 128.790 108.520 129.800 108.590 ;
        RECT 136.390 108.070 136.620 108.590 ;
        RECT 120.810 107.780 124.810 108.010 ;
        RECT 128.185 107.790 136.185 108.020 ;
        RECT 119.360 107.630 120.490 107.670 ;
        RECT 119.360 107.550 120.730 107.630 ;
        RECT 121.100 107.560 124.760 107.780 ;
        RECT 121.100 107.550 122.540 107.560 ;
        RECT 119.360 107.510 122.540 107.550 ;
        RECT 119.360 107.420 122.050 107.510 ;
        RECT 128.250 107.500 136.140 107.790 ;
        RECT 119.360 107.360 121.380 107.420 ;
        RECT 119.360 107.310 121.130 107.360 ;
        RECT 119.360 103.970 120.190 107.310 ;
        RECT 128.240 107.010 136.160 107.020 ;
        RECT 124.470 107.000 136.160 107.010 ;
        RECT 120.850 106.880 136.160 107.000 ;
        RECT 120.850 106.870 136.185 106.880 ;
        RECT 120.810 106.750 136.185 106.870 ;
        RECT 120.810 106.640 124.810 106.750 ;
        RECT 120.420 106.300 120.650 106.590 ;
        RECT 120.870 106.300 124.760 106.640 ;
        RECT 124.970 106.300 125.200 106.590 ;
        RECT 120.420 104.930 125.200 106.300 ;
        RECT 120.420 104.630 120.650 104.930 ;
        RECT 124.970 104.630 125.200 104.930 ;
        RECT 120.810 104.350 124.810 104.580 ;
        RECT 121.060 104.120 124.630 104.350 ;
        RECT 121.060 103.970 124.750 104.120 ;
        RECT 119.360 103.690 124.750 103.970 ;
        RECT 126.000 103.800 126.620 106.750 ;
        RECT 128.185 106.650 136.185 106.750 ;
        RECT 128.240 106.640 136.160 106.650 ;
        RECT 127.750 105.940 127.980 106.600 ;
        RECT 128.760 105.940 129.760 106.030 ;
        RECT 136.390 105.940 136.620 106.600 ;
        RECT 127.750 105.120 136.620 105.940 ;
        RECT 127.750 104.640 127.980 105.120 ;
        RECT 128.760 105.030 129.760 105.120 ;
        RECT 136.390 104.640 136.620 105.120 ;
        RECT 128.185 104.360 136.185 104.590 ;
        RECT 119.360 103.230 124.760 103.690 ;
        RECT 119.360 101.890 121.360 103.230 ;
        RECT 123.110 103.220 124.760 103.230 ;
        RECT 121.800 101.950 122.800 102.670 ;
        RECT 123.110 102.410 123.420 103.220 ;
        RECT 123.880 102.940 124.760 103.220 ;
        RECT 125.000 103.400 126.620 103.800 ;
        RECT 128.270 103.450 136.140 104.360 ;
        RECT 123.820 102.710 124.820 102.940 ;
        RECT 125.000 102.750 125.350 103.400 ;
        RECT 126.000 103.390 126.620 103.400 ;
        RECT 128.185 103.220 136.185 103.450 ;
        RECT 128.270 103.210 136.140 103.220 ;
        RECT 123.880 102.500 124.760 102.520 ;
        RECT 123.150 102.120 123.420 102.410 ;
        RECT 123.820 102.270 124.820 102.500 ;
        RECT 124.980 102.460 125.350 102.750 ;
        RECT 125.010 102.400 125.350 102.460 ;
        RECT 126.110 103.070 126.870 103.120 ;
        RECT 127.750 103.070 127.980 103.170 ;
        RECT 126.110 102.860 127.980 103.070 ;
        RECT 136.390 102.860 136.620 103.170 ;
        RECT 126.110 102.440 128.650 102.860 ;
        RECT 136.020 102.440 136.620 102.860 ;
        RECT 123.880 102.120 124.760 102.270 ;
        RECT 123.890 101.950 124.620 102.120 ;
        RECT 119.440 101.880 121.360 101.890 ;
        RECT 102.720 100.620 105.720 100.850 ;
        RECT 105.930 100.660 106.270 101.490 ;
        RECT 108.280 101.480 118.920 101.550 ;
        RECT 102.770 100.590 105.630 100.620 ;
        RECT 102.770 100.570 103.940 100.590 ;
        RECT 104.900 100.580 105.630 100.590 ;
        RECT 102.720 100.180 105.720 100.410 ;
        RECT 105.925 100.370 106.270 100.660 ;
        RECT 106.460 100.440 118.920 101.480 ;
        RECT 121.770 100.830 124.620 101.950 ;
        RECT 125.010 101.650 125.360 102.400 ;
        RECT 126.110 102.280 127.980 102.440 ;
        RECT 126.110 102.230 126.870 102.280 ;
        RECT 127.750 102.210 127.980 102.280 ;
        RECT 136.390 102.210 136.620 102.440 ;
        RECT 128.185 101.930 136.185 102.160 ;
        RECT 125.010 101.590 125.300 101.650 ;
        RECT 124.920 101.470 125.300 101.590 ;
        RECT 128.280 101.530 136.140 101.930 ;
        RECT 136.950 101.530 137.910 111.010 ;
        RECT 138.410 113.240 139.130 113.270 ;
        RECT 138.410 111.140 139.240 113.240 ;
        RECT 144.910 112.850 146.160 113.290 ;
        RECT 156.000 113.270 156.940 115.370 ;
        RECT 142.850 112.840 148.090 112.850 ;
        RECT 139.900 112.740 155.200 112.840 ;
        RECT 139.900 112.730 155.235 112.740 ;
        RECT 139.860 112.610 155.235 112.730 ;
        RECT 139.860 112.500 143.860 112.610 ;
        RECT 144.910 112.530 146.650 112.610 ;
        RECT 147.230 112.530 155.235 112.610 ;
        RECT 144.910 112.450 146.160 112.530 ;
        RECT 147.235 112.510 155.235 112.530 ;
        RECT 139.470 112.200 139.700 112.450 ;
        RECT 144.020 112.310 144.250 112.450 ;
        RECT 146.800 112.310 147.030 112.460 ;
        RECT 144.020 112.200 147.030 112.310 ;
        RECT 155.440 112.200 155.670 112.460 ;
        RECT 139.470 111.760 155.670 112.200 ;
        RECT 139.470 111.490 139.700 111.760 ;
        RECT 144.020 111.730 155.670 111.760 ;
        RECT 144.020 111.640 147.030 111.730 ;
        RECT 144.020 111.490 144.250 111.640 ;
        RECT 146.800 111.500 147.030 111.640 ;
        RECT 155.440 111.500 155.670 111.730 ;
        RECT 139.860 111.210 143.860 111.440 ;
        RECT 147.235 111.230 155.235 111.450 ;
        RECT 156.000 111.230 156.960 113.270 ;
        RECT 147.235 111.220 156.960 111.230 ;
        RECT 139.860 111.140 143.850 111.210 ;
        RECT 138.410 111.030 143.850 111.140 ;
        RECT 147.290 111.060 156.960 111.220 ;
        RECT 138.410 110.940 141.540 111.030 ;
        RECT 155.030 111.010 156.960 111.060 ;
        RECT 138.410 107.670 139.240 110.940 ;
        RECT 142.890 110.480 148.140 110.490 ;
        RECT 142.890 110.370 155.200 110.480 ;
        RECT 139.920 110.310 155.200 110.370 ;
        RECT 139.920 110.300 155.235 110.310 ;
        RECT 139.860 110.170 155.235 110.300 ;
        RECT 139.860 110.160 145.020 110.170 ;
        RECT 139.860 110.070 143.860 110.160 ;
        RECT 147.235 110.080 155.235 110.170 ;
        RECT 147.320 110.070 155.210 110.080 ;
        RECT 139.470 109.710 139.700 110.020 ;
        RECT 139.920 109.710 143.820 110.070 ;
        RECT 144.020 109.710 144.250 110.020 ;
        RECT 139.470 108.370 144.250 109.710 ;
        RECT 139.470 108.060 139.700 108.370 ;
        RECT 144.020 108.060 144.250 108.370 ;
        RECT 146.800 109.490 147.030 110.030 ;
        RECT 147.840 109.490 148.850 109.520 ;
        RECT 155.440 109.490 155.670 110.030 ;
        RECT 146.800 108.590 155.670 109.490 ;
        RECT 146.800 108.070 147.030 108.590 ;
        RECT 147.840 108.520 148.850 108.590 ;
        RECT 155.440 108.070 155.670 108.590 ;
        RECT 139.860 107.780 143.860 108.010 ;
        RECT 147.235 107.790 155.235 108.020 ;
        RECT 138.410 107.630 139.540 107.670 ;
        RECT 138.410 107.550 139.780 107.630 ;
        RECT 140.150 107.560 143.810 107.780 ;
        RECT 140.150 107.550 141.590 107.560 ;
        RECT 138.410 107.510 141.590 107.550 ;
        RECT 138.410 107.420 141.100 107.510 ;
        RECT 147.300 107.500 155.190 107.790 ;
        RECT 138.410 107.360 140.430 107.420 ;
        RECT 138.410 107.310 140.180 107.360 ;
        RECT 138.410 103.970 139.240 107.310 ;
        RECT 147.290 107.010 155.210 107.020 ;
        RECT 143.520 107.000 155.210 107.010 ;
        RECT 139.900 106.880 155.210 107.000 ;
        RECT 139.900 106.870 155.235 106.880 ;
        RECT 139.860 106.750 155.235 106.870 ;
        RECT 139.860 106.640 143.860 106.750 ;
        RECT 139.470 106.300 139.700 106.590 ;
        RECT 139.920 106.300 143.810 106.640 ;
        RECT 144.020 106.300 144.250 106.590 ;
        RECT 139.470 104.930 144.250 106.300 ;
        RECT 139.470 104.630 139.700 104.930 ;
        RECT 144.020 104.630 144.250 104.930 ;
        RECT 139.860 104.350 143.860 104.580 ;
        RECT 140.110 104.120 143.680 104.350 ;
        RECT 140.110 103.970 143.800 104.120 ;
        RECT 138.410 103.690 143.800 103.970 ;
        RECT 145.050 103.800 145.670 106.750 ;
        RECT 147.235 106.650 155.235 106.750 ;
        RECT 147.290 106.640 155.210 106.650 ;
        RECT 146.800 105.940 147.030 106.600 ;
        RECT 147.810 105.940 148.810 106.030 ;
        RECT 155.440 105.940 155.670 106.600 ;
        RECT 146.800 105.120 155.670 105.940 ;
        RECT 146.800 104.640 147.030 105.120 ;
        RECT 147.810 105.030 148.810 105.120 ;
        RECT 155.440 104.640 155.670 105.120 ;
        RECT 147.235 104.360 155.235 104.590 ;
        RECT 138.410 103.230 143.810 103.690 ;
        RECT 138.410 101.890 140.410 103.230 ;
        RECT 142.160 103.220 143.810 103.230 ;
        RECT 140.850 101.950 141.850 102.670 ;
        RECT 142.160 102.410 142.470 103.220 ;
        RECT 142.930 102.940 143.810 103.220 ;
        RECT 144.050 103.400 145.670 103.800 ;
        RECT 147.320 103.450 155.190 104.360 ;
        RECT 142.870 102.710 143.870 102.940 ;
        RECT 144.050 102.750 144.400 103.400 ;
        RECT 145.050 103.390 145.670 103.400 ;
        RECT 147.235 103.220 155.235 103.450 ;
        RECT 147.320 103.210 155.190 103.220 ;
        RECT 142.930 102.500 143.810 102.520 ;
        RECT 142.200 102.120 142.470 102.410 ;
        RECT 142.870 102.270 143.870 102.500 ;
        RECT 144.030 102.460 144.400 102.750 ;
        RECT 144.060 102.400 144.400 102.460 ;
        RECT 145.160 103.070 145.920 103.120 ;
        RECT 146.800 103.070 147.030 103.170 ;
        RECT 145.160 102.860 147.030 103.070 ;
        RECT 155.440 102.860 155.670 103.170 ;
        RECT 145.160 102.440 147.700 102.860 ;
        RECT 155.070 102.440 155.670 102.860 ;
        RECT 142.930 102.120 143.810 102.270 ;
        RECT 142.940 101.950 143.670 102.120 ;
        RECT 138.490 101.880 140.410 101.890 ;
        RECT 121.710 100.600 124.710 100.830 ;
        RECT 124.920 100.640 125.260 101.470 ;
        RECT 127.270 101.460 137.910 101.530 ;
        RECT 121.760 100.570 124.620 100.600 ;
        RECT 121.760 100.550 122.930 100.570 ;
        RECT 123.890 100.560 124.620 100.570 ;
        RECT 106.460 100.420 118.790 100.440 ;
        RECT 106.730 100.410 112.170 100.420 ;
        RECT 113.170 100.410 118.790 100.420 ;
        RECT 105.930 100.260 106.270 100.370 ;
        RECT 121.710 100.160 124.710 100.390 ;
        RECT 124.915 100.350 125.260 100.640 ;
        RECT 125.450 100.420 137.910 101.460 ;
        RECT 140.820 100.830 143.670 101.950 ;
        RECT 144.060 101.650 144.410 102.400 ;
        RECT 145.160 102.280 147.030 102.440 ;
        RECT 145.160 102.230 145.920 102.280 ;
        RECT 146.800 102.210 147.030 102.280 ;
        RECT 155.440 102.210 155.670 102.440 ;
        RECT 147.235 101.930 155.235 102.160 ;
        RECT 144.060 101.590 144.350 101.650 ;
        RECT 143.970 101.470 144.350 101.590 ;
        RECT 147.330 101.530 155.190 101.930 ;
        RECT 156.000 101.530 156.960 111.010 ;
        RECT 140.760 100.600 143.760 100.830 ;
        RECT 143.970 100.640 144.310 101.470 ;
        RECT 146.320 101.460 156.960 101.530 ;
        RECT 140.810 100.570 143.670 100.600 ;
        RECT 140.810 100.550 141.980 100.570 ;
        RECT 142.940 100.560 143.670 100.570 ;
        RECT 125.450 100.400 137.780 100.420 ;
        RECT 125.720 100.390 131.160 100.400 ;
        RECT 132.160 100.390 137.780 100.400 ;
        RECT 124.920 100.240 125.260 100.350 ;
        RECT 140.760 100.160 143.760 100.390 ;
        RECT 143.965 100.350 144.310 100.640 ;
        RECT 144.500 100.420 156.960 101.460 ;
        RECT 144.500 100.400 156.920 100.420 ;
        RECT 144.770 100.390 150.210 100.400 ;
        RECT 151.210 100.390 156.920 100.400 ;
        RECT 143.970 100.240 144.310 100.350 ;
        RECT 100.390 96.850 102.840 98.780 ;
        RECT 104.720 98.080 105.420 98.100 ;
        RECT 103.020 98.050 105.420 98.080 ;
        RECT 103.020 97.800 105.455 98.050 ;
        RECT 103.020 97.780 105.420 97.800 ;
        RECT 106.040 97.790 108.410 98.090 ;
        RECT 109.070 98.050 111.440 98.090 ;
        RECT 113.520 98.060 114.220 98.100 ;
        RECT 116.680 98.060 117.380 98.070 ;
        RECT 112.050 98.050 114.420 98.060 ;
        RECT 109.070 97.800 111.445 98.050 ;
        RECT 112.035 97.800 114.420 98.050 ;
        RECT 109.070 97.790 111.440 97.800 ;
        RECT 104.720 97.410 105.420 97.780 ;
        RECT 107.300 97.450 108.000 97.790 ;
        RECT 110.700 97.450 111.400 97.790 ;
        RECT 112.050 97.760 114.420 97.800 ;
        RECT 114.980 98.050 117.380 98.060 ;
        RECT 114.980 97.800 117.435 98.050 ;
        RECT 114.980 97.760 117.380 97.800 ;
        RECT 118.000 97.770 120.370 98.070 ;
        RECT 121.000 98.050 123.370 98.080 ;
        RECT 124.060 98.050 126.430 98.110 ;
        RECT 128.630 98.050 129.330 98.070 ;
        RECT 130.010 98.050 132.380 98.090 ;
        RECT 121.000 97.800 123.425 98.050 ;
        RECT 124.015 97.810 126.430 98.050 ;
        RECT 124.015 97.800 126.120 97.810 ;
        RECT 126.980 97.800 129.415 98.050 ;
        RECT 130.005 97.800 132.380 98.050 ;
        RECT 133.300 98.030 135.405 98.050 ;
        RECT 121.000 97.780 123.370 97.800 ;
        RECT 104.720 97.280 106.410 97.410 ;
        RECT 107.300 97.290 109.590 97.450 ;
        RECT 104.720 97.140 106.750 97.280 ;
        RECT 105.160 97.100 106.750 97.140 ;
        RECT 107.300 97.110 110.010 97.290 ;
        RECT 110.700 97.260 112.620 97.450 ;
        RECT 113.520 97.350 114.220 97.760 ;
        RECT 116.680 97.420 117.380 97.760 ;
        RECT 110.700 97.130 112.730 97.260 ;
        RECT 113.520 97.220 115.470 97.350 ;
        RECT 116.680 97.240 118.630 97.420 ;
        RECT 119.540 97.370 120.240 97.770 ;
        RECT 122.540 97.430 123.240 97.780 ;
        RECT 113.520 97.140 115.840 97.220 ;
        RECT 100.390 96.580 103.830 96.850 ;
        RECT 106.050 96.610 106.750 97.100 ;
        RECT 107.770 97.040 110.010 97.110 ;
        RECT 100.390 96.570 105.430 96.580 ;
        RECT 100.390 96.320 105.455 96.570 ;
        RECT 100.390 96.280 105.430 96.320 ;
        RECT 106.040 96.310 108.410 96.610 ;
        RECT 109.310 96.570 110.010 97.040 ;
        RECT 111.110 97.030 112.730 97.130 ;
        RECT 112.030 96.590 112.730 97.030 ;
        RECT 113.960 96.930 115.840 97.140 ;
        RECT 116.680 97.110 118.790 97.240 ;
        RECT 117.120 97.000 118.790 97.110 ;
        RECT 119.540 97.180 121.450 97.370 ;
        RECT 122.540 97.230 124.540 97.430 ;
        RECT 125.240 97.380 125.940 97.800 ;
        RECT 126.980 97.750 129.350 97.800 ;
        RECT 130.010 97.790 132.380 97.800 ;
        RECT 132.990 97.800 135.405 98.030 ;
        RECT 128.630 97.480 129.330 97.750 ;
        RECT 125.240 97.250 127.770 97.380 ;
        RECT 128.630 97.290 130.640 97.480 ;
        RECT 131.480 97.400 132.180 97.790 ;
        RECT 132.990 97.730 135.360 97.800 ;
        RECT 135.980 97.750 138.420 98.100 ;
        RECT 140.640 98.090 141.340 98.120 ;
        RECT 143.900 98.090 145.220 98.100 ;
        RECT 119.540 97.080 121.870 97.180 ;
        RECT 115.140 96.610 115.840 96.930 ;
        RECT 118.090 96.610 118.790 97.000 ;
        RECT 119.940 96.950 121.870 97.080 ;
        RECT 122.540 97.060 124.720 97.230 ;
        RECT 125.240 97.120 127.980 97.250 ;
        RECT 123.030 97.010 124.720 97.060 ;
        RECT 109.060 96.320 111.445 96.570 ;
        RECT 100.390 96.000 103.830 96.280 ;
        RECT 109.060 96.270 111.430 96.320 ;
        RECT 112.030 96.290 114.400 96.590 ;
        RECT 115.060 96.570 117.430 96.610 ;
        RECT 115.060 96.320 117.435 96.570 ;
        RECT 115.060 96.310 117.430 96.320 ;
        RECT 118.020 96.310 120.390 96.610 ;
        RECT 121.170 96.590 121.870 96.950 ;
        RECT 121.010 96.570 123.380 96.590 ;
        RECT 124.020 96.570 124.720 97.010 ;
        RECT 125.600 96.980 127.980 97.120 ;
        RECT 128.630 97.110 130.720 97.290 ;
        RECT 131.480 97.200 133.490 97.400 ;
        RECT 134.660 97.330 135.300 97.730 ;
        RECT 134.660 97.240 136.250 97.330 ;
        RECT 131.480 97.120 133.720 97.200 ;
        RECT 134.660 97.170 136.780 97.240 ;
        RECT 137.100 97.210 138.420 97.750 ;
        RECT 139.260 97.570 141.400 98.090 ;
        RECT 141.980 97.740 147.410 98.090 ;
        RECT 147.980 98.050 153.380 98.090 ;
        RECT 147.975 97.800 153.380 98.050 ;
        RECT 147.980 97.750 153.380 97.800 ;
        RECT 153.960 97.750 156.920 100.390 ;
        RECT 143.900 97.730 145.220 97.740 ;
        RECT 140.760 97.330 141.360 97.570 ;
        RECT 144.300 97.550 144.810 97.730 ;
        RECT 150.420 97.580 150.930 97.750 ;
        RECT 137.100 97.190 139.380 97.210 ;
        RECT 140.760 97.190 142.370 97.330 ;
        RECT 128.720 97.060 130.720 97.110 ;
        RECT 127.280 96.580 127.980 96.980 ;
        RECT 130.020 96.600 130.720 97.060 ;
        RECT 131.570 96.980 133.720 97.120 ;
        RECT 135.190 97.040 136.780 97.170 ;
        RECT 126.980 96.570 129.350 96.580 ;
        RECT 130.010 96.570 132.380 96.600 ;
        RECT 133.020 96.590 133.720 96.980 ;
        RECT 136.040 96.620 136.780 97.040 ;
        RECT 137.950 97.100 139.380 97.190 ;
        RECT 137.950 96.970 140.130 97.100 ;
        RECT 121.010 96.320 123.425 96.570 ;
        RECT 124.015 96.560 126.120 96.570 ;
        RECT 124.015 96.320 126.390 96.560 ;
        RECT 115.140 96.260 115.840 96.310 ;
        RECT 118.090 96.280 118.790 96.310 ;
        RECT 121.010 96.290 123.380 96.320 ;
        RECT 121.170 96.220 121.870 96.290 ;
        RECT 124.020 96.260 126.390 96.320 ;
        RECT 126.980 96.320 129.415 96.570 ;
        RECT 130.005 96.320 132.380 96.570 ;
        RECT 126.980 96.280 129.350 96.320 ;
        RECT 130.010 96.300 132.380 96.320 ;
        RECT 133.010 96.570 135.380 96.590 ;
        RECT 136.000 96.570 138.440 96.620 ;
        RECT 139.080 96.610 140.130 96.970 ;
        RECT 140.850 97.030 142.370 97.190 ;
        RECT 140.850 96.930 144.100 97.030 ;
        RECT 133.010 96.320 135.405 96.570 ;
        RECT 135.995 96.320 138.440 96.570 ;
        RECT 133.010 96.290 135.380 96.320 ;
        RECT 133.020 96.240 133.720 96.290 ;
        RECT 136.000 96.270 138.440 96.320 ;
        RECT 138.960 96.260 141.400 96.610 ;
        RECT 141.960 96.600 144.100 96.930 ;
        RECT 141.960 96.510 144.420 96.600 ;
        RECT 141.980 96.250 144.420 96.510 ;
        RECT 100.390 95.650 102.840 96.000 ;
        RECT 100.390 95.630 101.440 95.650 ;
      LAYER met2 ;
        RECT 69.275 221.420 69.665 221.500 ;
        RECT 69.275 221.280 73.200 221.420 ;
        RECT 69.275 221.200 69.665 221.280 ;
        RECT 73.060 221.240 73.200 221.280 ;
        RECT 73.060 221.100 125.130 221.240 ;
        RECT 71.965 220.960 72.355 221.040 ;
        RECT 71.965 220.820 124.490 220.960 ;
        RECT 71.965 220.740 72.355 220.820 ;
        RECT 74.755 220.560 75.145 220.620 ;
        RECT 123.555 220.560 123.925 220.610 ;
        RECT 74.755 220.380 123.925 220.560 ;
        RECT 74.755 220.320 75.145 220.380 ;
        RECT 123.555 220.330 123.925 220.380 ;
        RECT 124.350 220.370 124.490 220.820 ;
        RECT 124.990 220.650 125.130 221.100 ;
        RECT 124.990 220.510 138.900 220.650 ;
        RECT 138.760 220.480 138.900 220.510 ;
        RECT 147.650 220.480 147.970 220.540 ;
        RECT 124.350 220.230 138.300 220.370 ;
        RECT 138.760 220.340 147.970 220.480 ;
        RECT 147.650 220.280 147.970 220.340 ;
        RECT 80.265 219.985 80.655 220.040 ;
        RECT 137.155 219.985 137.525 220.030 ;
        RECT 80.265 219.830 137.525 219.985 ;
        RECT 80.265 219.795 82.855 219.830 ;
        RECT 83.525 219.795 137.525 219.830 ;
        RECT 138.160 219.940 138.300 220.230 ;
        RECT 147.210 219.940 147.530 220.000 ;
        RECT 138.160 219.800 147.530 219.940 ;
        RECT 80.265 219.740 80.655 219.795 ;
        RECT 137.155 219.750 137.525 219.795 ;
        RECT 147.210 219.740 147.530 219.800 ;
        RECT 82.995 219.610 83.385 219.690 ;
        RECT 82.995 219.470 115.180 219.610 ;
        RECT 82.995 219.390 83.385 219.470 ;
        RECT 115.040 219.450 115.180 219.470 ;
        RECT 146.870 219.450 147.130 219.540 ;
        RECT 115.040 219.310 147.130 219.450 ;
        RECT 114.035 219.260 114.405 219.270 ;
        RECT 85.765 219.220 86.155 219.255 ;
        RECT 113.890 219.220 114.405 219.260 ;
        RECT 146.870 219.220 147.130 219.310 ;
        RECT 85.765 218.990 114.405 219.220 ;
        RECT 85.765 218.955 86.155 218.990 ;
        RECT 146.280 218.960 146.600 219.020 ;
        RECT 115.000 218.820 146.600 218.960 ;
        RECT 94.095 218.740 94.485 218.820 ;
        RECT 115.000 218.740 115.140 218.820 ;
        RECT 146.280 218.760 146.600 218.820 ;
        RECT 94.095 218.600 115.140 218.740 ;
        RECT 91.365 218.415 91.665 218.530 ;
        RECT 94.095 218.520 94.485 218.600 ;
        RECT 130.350 218.565 130.730 218.670 ;
        RECT 115.680 218.415 130.730 218.565 ;
        RECT 91.365 218.360 93.960 218.415 ;
        RECT 94.620 218.400 130.730 218.415 ;
        RECT 94.620 218.360 115.845 218.400 ;
        RECT 91.365 218.250 115.845 218.360 ;
        RECT 130.350 218.290 130.730 218.400 ;
        RECT 140.540 218.510 140.940 218.620 ;
        RECT 143.865 218.510 144.255 218.585 ;
        RECT 140.540 218.355 144.255 218.510 ;
        RECT 140.540 218.250 140.940 218.355 ;
        RECT 143.865 218.285 144.255 218.355 ;
        RECT 91.365 218.140 91.665 218.250 ;
        RECT 93.840 218.220 94.750 218.250 ;
        RECT 88.505 218.010 88.895 218.090 ;
        RECT 88.505 217.990 91.210 218.010 ;
        RECT 91.820 217.990 110.010 218.010 ;
        RECT 88.505 217.870 110.010 217.990 ;
        RECT 88.505 217.790 88.895 217.870 ;
        RECT 90.980 217.830 91.980 217.870 ;
        RECT 77.530 217.660 77.830 217.785 ;
        RECT 77.530 217.650 88.365 217.660 ;
        RECT 89.035 217.650 109.630 217.660 ;
        RECT 77.530 217.520 109.630 217.650 ;
        RECT 77.530 217.395 77.830 217.520 ;
        RECT 88.280 217.510 89.120 217.520 ;
        RECT 66.425 217.260 66.815 217.340 ;
        RECT 66.425 217.250 77.370 217.260 ;
        RECT 77.980 217.250 109.010 217.260 ;
        RECT 66.425 217.120 109.010 217.250 ;
        RECT 66.425 217.040 66.815 217.120 ;
        RECT 77.250 217.110 78.140 217.120 ;
        RECT 63.785 216.900 64.175 216.980 ;
        RECT 63.785 216.760 108.550 216.900 ;
        RECT 63.785 216.680 64.175 216.760 ;
        RECT 108.410 206.130 108.550 216.760 ;
        RECT 108.320 205.870 108.640 206.130 ;
        RECT 108.870 205.580 109.010 217.120 ;
        RECT 108.780 205.320 109.100 205.580 ;
        RECT 109.490 205.090 109.630 217.520 ;
        RECT 109.260 204.860 109.630 205.090 ;
        RECT 109.260 204.830 109.580 204.860 ;
        RECT 99.600 204.020 103.600 204.090 ;
        RECT 109.870 204.020 110.010 217.870 ;
        RECT 119.330 216.900 119.650 216.960 ;
        RECT 123.555 216.900 123.925 216.970 ;
        RECT 119.330 216.760 123.925 216.900 ;
        RECT 119.330 216.700 119.650 216.760 ;
        RECT 123.555 216.690 123.925 216.760 ;
        RECT 126.130 216.900 126.450 216.960 ;
        RECT 130.355 216.900 130.725 216.970 ;
        RECT 137.155 216.960 137.525 216.970 ;
        RECT 126.130 216.760 130.725 216.900 ;
        RECT 126.130 216.700 126.450 216.760 ;
        RECT 130.355 216.690 130.725 216.760 ;
        RECT 137.010 216.700 137.525 216.960 ;
        RECT 137.155 216.690 137.525 216.700 ;
        RECT 114.570 216.440 114.890 216.500 ;
        RECT 117.970 216.440 118.290 216.500 ;
        RECT 119.670 216.440 119.990 216.500 ;
        RECT 114.570 216.300 119.990 216.440 ;
        RECT 114.570 216.240 114.890 216.300 ;
        RECT 117.970 216.240 118.290 216.300 ;
        RECT 119.670 216.240 119.990 216.300 ;
        RECT 122.730 216.440 123.050 216.500 ;
        RECT 124.770 216.440 125.090 216.500 ;
        RECT 122.730 216.300 125.090 216.440 ;
        RECT 122.730 216.240 123.050 216.300 ;
        RECT 124.770 216.240 125.090 216.300 ;
        RECT 125.450 216.440 125.770 216.500 ;
        RECT 128.170 216.440 128.490 216.500 ;
        RECT 129.870 216.440 130.190 216.500 ;
        RECT 125.450 216.300 130.190 216.440 ;
        RECT 125.450 216.240 125.770 216.300 ;
        RECT 128.170 216.240 128.490 216.300 ;
        RECT 129.870 216.240 130.190 216.300 ;
        RECT 131.230 216.440 131.550 216.500 ;
        RECT 132.590 216.440 132.910 216.500 ;
        RECT 131.230 216.300 132.910 216.440 ;
        RECT 131.230 216.240 131.550 216.300 ;
        RECT 132.590 216.240 132.910 216.300 ;
        RECT 137.010 214.600 137.330 214.660 ;
        RECT 138.370 214.600 138.690 214.660 ;
        RECT 137.010 214.460 138.690 214.600 ;
        RECT 137.010 214.400 137.330 214.460 ;
        RECT 138.370 214.400 138.690 214.460 ;
        RECT 122.050 214.140 122.370 214.200 ;
        RECT 124.430 214.140 124.750 214.200 ;
        RECT 122.050 214.000 124.750 214.140 ;
        RECT 122.050 213.940 122.370 214.000 ;
        RECT 124.430 213.940 124.750 214.000 ;
        RECT 133.610 214.140 133.930 214.200 ;
        RECT 135.650 214.140 135.970 214.200 ;
        RECT 133.610 214.000 135.970 214.140 ;
        RECT 133.610 213.940 133.930 214.000 ;
        RECT 135.650 213.940 135.970 214.000 ;
        RECT 115.250 213.680 115.570 213.740 ;
        RECT 116.610 213.680 116.930 213.740 ;
        RECT 115.250 213.540 116.930 213.680 ;
        RECT 115.250 213.480 115.570 213.540 ;
        RECT 116.610 213.480 116.930 213.540 ;
        RECT 142.450 212.300 142.770 212.360 ;
        RECT 144.150 212.300 144.470 212.360 ;
        RECT 142.450 212.160 144.470 212.300 ;
        RECT 142.450 212.100 142.770 212.160 ;
        RECT 144.150 212.100 144.470 212.160 ;
        RECT 115.250 211.840 115.570 211.900 ;
        RECT 118.990 211.840 119.310 211.900 ;
        RECT 115.250 211.700 119.310 211.840 ;
        RECT 115.250 211.640 115.570 211.700 ;
        RECT 118.990 211.640 119.310 211.700 ;
        RECT 128.850 211.840 129.170 211.900 ;
        RECT 132.590 211.840 132.910 211.900 ;
        RECT 128.850 211.700 132.910 211.840 ;
        RECT 128.850 211.640 129.170 211.700 ;
        RECT 132.590 211.640 132.910 211.700 ;
        RECT 115.250 211.380 115.570 211.440 ;
        RECT 119.330 211.380 119.650 211.440 ;
        RECT 125.110 211.380 125.430 211.440 ;
        RECT 115.250 211.240 125.430 211.380 ;
        RECT 115.250 211.180 115.570 211.240 ;
        RECT 119.330 211.180 119.650 211.240 ;
        RECT 125.110 211.180 125.430 211.240 ;
        RECT 126.130 211.380 126.450 211.440 ;
        RECT 127.150 211.380 127.470 211.440 ;
        RECT 126.130 211.240 127.470 211.380 ;
        RECT 126.130 211.180 126.450 211.240 ;
        RECT 127.150 211.180 127.470 211.240 ;
        RECT 125.110 210.920 125.430 210.980 ;
        RECT 132.930 210.920 133.250 210.980 ;
        RECT 135.990 210.920 136.310 210.980 ;
        RECT 125.110 210.780 136.310 210.920 ;
        RECT 125.110 210.720 125.430 210.780 ;
        RECT 132.930 210.720 133.250 210.780 ;
        RECT 135.990 210.720 136.310 210.780 ;
        RECT 117.290 209.540 117.610 209.600 ;
        RECT 122.390 209.540 122.710 209.600 ;
        RECT 117.290 209.400 122.710 209.540 ;
        RECT 117.290 209.340 117.610 209.400 ;
        RECT 122.390 209.340 122.710 209.400 ;
        RECT 130.890 209.540 131.210 209.600 ;
        RECT 133.270 209.540 133.590 209.600 ;
        RECT 130.890 209.400 133.590 209.540 ;
        RECT 130.890 209.340 131.210 209.400 ;
        RECT 133.270 209.340 133.590 209.400 ;
        RECT 136.330 209.540 136.650 209.600 ;
        RECT 138.030 209.540 138.350 209.600 ;
        RECT 136.330 209.400 138.350 209.540 ;
        RECT 136.330 209.340 136.650 209.400 ;
        RECT 138.030 209.340 138.350 209.400 ;
        RECT 115.250 209.080 115.570 209.140 ;
        RECT 119.670 209.080 119.990 209.140 ;
        RECT 115.250 208.940 119.990 209.080 ;
        RECT 115.250 208.880 115.570 208.940 ;
        RECT 119.670 208.880 119.990 208.940 ;
        RECT 137.010 209.080 137.330 209.140 ;
        RECT 138.030 209.080 138.350 209.140 ;
        RECT 137.010 208.940 138.350 209.080 ;
        RECT 137.010 208.880 137.330 208.940 ;
        RECT 138.030 208.880 138.350 208.940 ;
        RECT 120.010 208.620 120.330 208.680 ;
        RECT 123.410 208.620 123.730 208.680 ;
        RECT 127.830 208.620 128.150 208.680 ;
        RECT 120.010 208.480 128.150 208.620 ;
        RECT 120.010 208.420 120.330 208.480 ;
        RECT 123.410 208.420 123.730 208.480 ;
        RECT 127.830 208.420 128.150 208.480 ;
        RECT 142.450 207.700 142.770 207.760 ;
        RECT 144.150 207.700 144.470 207.760 ;
        RECT 142.450 207.560 144.470 207.700 ;
        RECT 142.450 207.500 142.770 207.560 ;
        RECT 144.150 207.500 144.470 207.560 ;
        RECT 141.915 207.240 142.285 207.310 ;
        RECT 144.150 207.240 144.470 207.300 ;
        RECT 141.915 207.100 144.470 207.240 ;
        RECT 141.915 207.030 142.285 207.100 ;
        RECT 144.150 207.040 144.470 207.100 ;
        RECT 111.510 206.780 111.830 206.840 ;
        RECT 115.250 206.780 115.570 206.840 ;
        RECT 111.510 206.640 115.570 206.780 ;
        RECT 111.510 206.580 111.830 206.640 ;
        RECT 115.250 206.580 115.570 206.640 ;
        RECT 133.270 206.780 133.590 206.840 ;
        RECT 137.010 206.780 137.330 206.840 ;
        RECT 138.710 206.780 139.030 206.840 ;
        RECT 140.750 206.780 141.070 206.840 ;
        RECT 133.270 206.640 141.070 206.780 ;
        RECT 133.270 206.580 133.590 206.640 ;
        RECT 137.010 206.580 137.330 206.640 ;
        RECT 138.710 206.580 139.030 206.640 ;
        RECT 140.750 206.580 141.070 206.640 ;
        RECT 131.230 205.860 131.550 205.920 ;
        RECT 140.555 205.860 140.925 205.930 ;
        RECT 131.230 205.720 140.925 205.860 ;
        RECT 131.230 205.660 131.550 205.720 ;
        RECT 140.555 205.650 140.925 205.720 ;
        RECT 142.110 205.400 142.430 205.460 ;
        RECT 143.470 205.400 143.790 205.460 ;
        RECT 142.110 205.260 143.790 205.400 ;
        RECT 142.110 205.200 142.430 205.260 ;
        RECT 143.470 205.200 143.790 205.260 ;
        RECT 114.230 204.940 114.550 205.000 ;
        RECT 119.670 204.940 119.990 205.000 ;
        RECT 125.790 204.940 126.110 205.000 ;
        RECT 114.230 204.800 126.110 204.940 ;
        RECT 114.230 204.740 114.550 204.800 ;
        RECT 119.670 204.740 119.990 204.800 ;
        RECT 125.790 204.740 126.110 204.800 ;
        RECT 133.610 204.480 133.930 204.540 ;
        RECT 137.010 204.480 137.330 204.540 ;
        RECT 133.610 204.340 137.330 204.480 ;
        RECT 133.610 204.280 133.930 204.340 ;
        RECT 137.010 204.280 137.330 204.340 ;
        RECT 139.730 204.480 140.050 204.540 ;
        RECT 141.770 204.480 142.090 204.540 ;
        RECT 139.730 204.340 142.090 204.480 ;
        RECT 139.730 204.280 140.050 204.340 ;
        RECT 141.770 204.280 142.090 204.340 ;
        RECT 110.830 204.020 111.150 204.080 ;
        RECT 99.600 203.880 111.150 204.020 ;
        RECT 99.600 203.810 103.600 203.880 ;
        RECT 110.830 203.820 111.150 203.880 ;
        RECT 145.170 204.020 145.490 204.080 ;
        RECT 147.650 204.020 147.970 204.110 ;
        RECT 153.365 204.020 157.365 204.090 ;
        RECT 145.170 203.880 157.365 204.020 ;
        RECT 145.170 203.820 145.490 203.880 ;
        RECT 147.650 203.790 147.970 203.880 ;
        RECT 153.365 203.810 157.365 203.880 ;
        RECT 122.050 203.560 122.370 203.620 ;
        RECT 124.770 203.560 125.090 203.620 ;
        RECT 122.050 203.420 125.090 203.560 ;
        RECT 122.050 203.360 122.370 203.420 ;
        RECT 124.770 203.360 125.090 203.420 ;
        RECT 125.790 203.560 126.110 203.620 ;
        RECT 128.850 203.560 129.170 203.620 ;
        RECT 134.290 203.560 134.610 203.620 ;
        RECT 137.010 203.560 137.330 203.620 ;
        RECT 125.790 203.420 137.330 203.560 ;
        RECT 125.790 203.360 126.110 203.420 ;
        RECT 128.850 203.360 129.170 203.420 ;
        RECT 134.290 203.360 134.610 203.420 ;
        RECT 137.010 203.360 137.330 203.420 ;
        RECT 109.260 203.080 109.580 203.140 ;
        RECT 126.130 203.100 126.450 203.160 ;
        RECT 127.830 203.100 128.150 203.160 ;
        RECT 109.260 202.880 109.670 203.080 ;
        RECT 126.130 202.960 128.150 203.100 ;
        RECT 126.130 202.900 126.450 202.960 ;
        RECT 127.830 202.900 128.150 202.960 ;
        RECT 128.850 203.100 129.170 203.160 ;
        RECT 141.915 203.100 142.285 203.170 ;
        RECT 128.850 202.960 142.285 203.100 ;
        RECT 128.850 202.900 129.170 202.960 ;
        RECT 141.915 202.890 142.285 202.960 ;
        RECT 109.490 202.750 109.670 202.880 ;
        RECT 109.490 201.260 109.630 202.750 ;
        RECT 111.510 201.520 111.830 201.780 ;
        RECT 110.830 201.260 111.150 201.320 ;
        RECT 105.310 201.120 111.150 201.260 ;
        RECT 99.600 200.800 103.600 200.870 ;
        RECT 105.310 200.800 105.450 201.120 ;
        RECT 110.830 201.060 111.150 201.120 ;
        RECT 99.600 200.660 105.450 200.800 ;
        RECT 99.600 200.590 103.600 200.660 ;
        RECT 111.600 200.340 111.740 201.520 ;
        RECT 113.015 200.890 113.385 202.430 ;
        RECT 118.455 200.890 118.825 202.430 ;
        RECT 123.895 200.890 124.265 202.430 ;
        RECT 129.335 200.890 129.705 202.430 ;
        RECT 134.775 200.890 135.145 202.430 ;
        RECT 140.215 200.890 140.585 202.430 ;
        RECT 145.655 200.890 146.025 202.430 ;
        RECT 153.365 200.800 157.365 200.870 ;
        RECT 146.790 200.660 157.365 200.800 ;
        RECT 115.250 200.340 115.570 200.400 ;
        RECT 118.990 200.340 119.310 200.400 ;
        RECT 111.600 200.200 114.970 200.340 ;
        RECT 114.830 199.480 114.970 200.200 ;
        RECT 115.250 200.200 119.310 200.340 ;
        RECT 115.250 200.140 115.570 200.200 ;
        RECT 118.990 200.140 119.310 200.200 ;
        RECT 127.830 200.340 128.150 200.400 ;
        RECT 138.030 200.340 138.350 200.400 ;
        RECT 127.830 200.200 138.350 200.340 ;
        RECT 127.830 200.140 128.150 200.200 ;
        RECT 138.030 200.140 138.350 200.200 ;
        RECT 138.710 200.340 139.030 200.400 ;
        RECT 143.470 200.340 143.790 200.400 ;
        RECT 138.710 200.200 143.790 200.340 ;
        RECT 138.710 200.140 139.030 200.200 ;
        RECT 143.470 200.140 143.790 200.200 ;
        RECT 116.950 199.880 117.270 199.940 ;
        RECT 129.870 199.880 130.190 199.940 ;
        RECT 136.330 199.880 136.650 199.940 ;
        RECT 116.950 199.740 136.650 199.880 ;
        RECT 116.950 199.680 117.270 199.740 ;
        RECT 129.870 199.680 130.190 199.740 ;
        RECT 136.330 199.680 136.650 199.740 ;
        RECT 137.010 199.880 137.330 199.940 ;
        RECT 138.710 199.880 139.030 199.940 ;
        RECT 137.010 199.740 139.030 199.880 ;
        RECT 137.010 199.680 137.330 199.740 ;
        RECT 138.710 199.680 139.030 199.740 ;
        RECT 141.090 199.880 141.410 199.940 ;
        RECT 146.280 199.880 146.600 199.970 ;
        RECT 146.790 199.880 146.930 200.660 ;
        RECT 153.365 200.590 157.365 200.660 ;
        RECT 141.090 199.740 146.930 199.880 ;
        RECT 141.090 199.680 141.410 199.740 ;
        RECT 146.280 199.650 146.600 199.740 ;
        RECT 111.170 199.420 111.490 199.480 ;
        RECT 113.550 199.420 113.870 199.480 ;
        RECT 111.170 199.280 113.870 199.420 ;
        RECT 114.830 199.420 115.230 199.480 ;
        RECT 117.970 199.420 118.290 199.480 ;
        RECT 120.010 199.420 120.330 199.480 ;
        RECT 121.710 199.420 122.030 199.480 ;
        RECT 114.830 199.280 122.030 199.420 ;
        RECT 111.170 199.220 111.490 199.280 ;
        RECT 113.550 199.220 113.870 199.280 ;
        RECT 114.910 199.220 115.230 199.280 ;
        RECT 117.970 199.220 118.290 199.280 ;
        RECT 120.010 199.220 120.330 199.280 ;
        RECT 121.710 199.220 122.030 199.280 ;
        RECT 127.830 199.420 128.150 199.480 ;
        RECT 130.550 199.420 130.870 199.480 ;
        RECT 135.310 199.420 135.630 199.480 ;
        RECT 127.830 199.280 130.870 199.420 ;
        RECT 127.830 199.220 128.150 199.280 ;
        RECT 130.550 199.220 130.870 199.280 ;
        RECT 131.150 199.280 135.630 199.420 ;
        RECT 106.300 197.880 108.840 198.875 ;
        RECT 99.600 197.580 103.600 197.650 ;
        RECT 110.295 197.590 110.665 199.130 ;
        RECT 115.735 197.590 116.105 199.130 ;
        RECT 121.175 197.590 121.545 199.130 ;
        RECT 126.615 197.590 126.985 199.130 ;
        RECT 128.510 198.960 128.830 199.020 ;
        RECT 131.150 198.960 131.290 199.280 ;
        RECT 135.310 199.220 135.630 199.280 ;
        RECT 139.730 199.420 140.050 199.480 ;
        RECT 144.830 199.420 145.150 199.480 ;
        RECT 139.730 199.280 145.150 199.420 ;
        RECT 139.730 199.220 140.050 199.280 ;
        RECT 144.830 199.220 145.150 199.280 ;
        RECT 128.510 198.820 131.290 198.960 ;
        RECT 128.510 198.760 128.830 198.820 ;
        RECT 132.055 197.590 132.425 199.130 ;
        RECT 137.495 197.590 137.865 199.130 ;
        RECT 138.710 198.960 139.030 199.020 ;
        RECT 141.430 198.960 141.750 199.020 ;
        RECT 138.710 198.820 141.750 198.960 ;
        RECT 138.710 198.760 139.030 198.820 ;
        RECT 141.430 198.760 141.750 198.820 ;
        RECT 142.935 197.590 143.305 199.130 ;
        RECT 145.170 197.580 145.490 197.640 ;
        RECT 146.870 197.580 147.130 197.670 ;
        RECT 153.365 197.580 157.365 197.650 ;
        RECT 99.600 197.440 105.450 197.580 ;
        RECT 99.600 197.370 103.600 197.440 ;
        RECT 105.310 197.120 105.450 197.440 ;
        RECT 145.170 197.440 157.365 197.580 ;
        RECT 145.170 197.380 145.490 197.440 ;
        RECT 146.870 197.350 147.130 197.440 ;
        RECT 153.365 197.370 157.365 197.440 ;
        RECT 109.690 197.120 110.020 197.210 ;
        RECT 110.830 197.120 111.150 197.180 ;
        RECT 105.310 196.980 111.150 197.120 ;
        RECT 109.690 196.890 110.020 196.980 ;
        RECT 110.830 196.920 111.150 196.980 ;
        RECT 125.110 197.120 125.430 197.180 ;
        RECT 132.590 197.120 132.910 197.180 ;
        RECT 134.290 197.120 134.610 197.180 ;
        RECT 138.710 197.120 139.030 197.180 ;
        RECT 125.110 196.980 134.010 197.120 ;
        RECT 125.110 196.920 125.430 196.980 ;
        RECT 132.590 196.920 132.910 196.980 ;
        RECT 112.530 196.660 112.850 196.720 ;
        RECT 121.710 196.660 122.030 196.720 ;
        RECT 125.110 196.660 125.430 196.720 ;
        RECT 112.530 196.520 125.430 196.660 ;
        RECT 112.530 196.460 112.850 196.520 ;
        RECT 121.710 196.460 122.030 196.520 ;
        RECT 125.110 196.460 125.430 196.520 ;
        RECT 131.570 196.660 131.890 196.720 ;
        RECT 132.930 196.660 133.250 196.720 ;
        RECT 131.570 196.520 133.250 196.660 ;
        RECT 133.870 196.660 134.010 196.980 ;
        RECT 134.290 196.980 139.030 197.120 ;
        RECT 134.290 196.920 134.610 196.980 ;
        RECT 138.710 196.920 139.030 196.980 ;
        RECT 142.450 197.120 142.770 197.180 ;
        RECT 144.150 197.120 144.470 197.180 ;
        RECT 142.450 196.980 144.470 197.120 ;
        RECT 142.450 196.920 142.770 196.980 ;
        RECT 144.150 196.920 144.470 196.980 ;
        RECT 138.710 196.660 139.030 196.720 ;
        RECT 133.870 196.520 139.030 196.660 ;
        RECT 131.570 196.460 131.890 196.520 ;
        RECT 132.930 196.460 133.250 196.520 ;
        RECT 138.710 196.460 139.030 196.520 ;
        RECT 142.110 196.660 142.430 196.720 ;
        RECT 143.470 196.660 143.790 196.720 ;
        RECT 142.110 196.520 143.790 196.660 ;
        RECT 142.110 196.460 142.430 196.520 ;
        RECT 143.470 196.460 143.790 196.520 ;
        RECT 122.730 196.200 123.050 196.260 ;
        RECT 122.730 196.000 123.130 196.200 ;
        RECT 126.130 196.000 126.450 196.260 ;
        RECT 133.270 196.200 133.590 196.260 ;
        RECT 135.990 196.200 136.310 196.260 ;
        RECT 133.270 196.060 136.310 196.200 ;
        RECT 133.270 196.000 133.590 196.060 ;
        RECT 135.990 196.000 136.310 196.060 ;
        RECT 139.050 196.200 139.370 196.260 ;
        RECT 140.750 196.200 141.070 196.260 ;
        RECT 139.050 196.060 141.070 196.200 ;
        RECT 139.050 196.000 139.370 196.060 ;
        RECT 140.750 196.000 141.070 196.060 ;
        RECT 122.990 195.740 123.130 196.000 ;
        RECT 126.220 195.740 126.360 196.000 ;
        RECT 128.170 195.740 128.490 195.800 ;
        RECT 133.950 195.740 134.270 195.800 ;
        RECT 122.990 195.600 134.270 195.740 ;
        RECT 128.170 195.540 128.490 195.600 ;
        RECT 133.950 195.540 134.270 195.600 ;
        RECT 138.710 195.740 139.030 195.800 ;
        RECT 141.770 195.740 142.090 195.800 ;
        RECT 138.710 195.600 142.090 195.740 ;
        RECT 138.710 195.540 139.030 195.600 ;
        RECT 141.770 195.540 142.090 195.600 ;
        RECT 123.070 195.280 123.390 195.340 ;
        RECT 132.930 195.280 133.250 195.340 ;
        RECT 123.070 195.140 133.250 195.280 ;
        RECT 123.070 195.080 123.390 195.140 ;
        RECT 132.930 195.080 133.250 195.140 ;
        RECT 115.250 194.820 115.570 194.880 ;
        RECT 120.350 194.820 120.670 194.880 ;
        RECT 124.770 194.820 125.090 194.880 ;
        RECT 115.250 194.680 125.090 194.820 ;
        RECT 115.250 194.620 115.570 194.680 ;
        RECT 120.350 194.620 120.670 194.680 ;
        RECT 124.770 194.620 125.090 194.680 ;
        RECT 128.510 194.820 128.830 194.880 ;
        RECT 129.870 194.820 130.190 194.880 ;
        RECT 136.670 194.820 136.990 194.880 ;
        RECT 141.430 194.820 141.750 194.880 ;
        RECT 128.510 194.680 141.750 194.820 ;
        RECT 128.510 194.620 128.830 194.680 ;
        RECT 129.870 194.620 130.190 194.680 ;
        RECT 136.670 194.620 136.990 194.680 ;
        RECT 141.430 194.620 141.750 194.680 ;
        RECT 131.570 194.360 131.890 194.420 ;
        RECT 135.650 194.360 135.970 194.420 ;
        RECT 138.370 194.360 138.690 194.420 ;
        RECT 139.730 194.360 140.050 194.420 ;
        RECT 141.770 194.360 142.090 194.420 ;
        RECT 131.570 194.220 138.690 194.360 ;
        RECT 131.570 194.160 131.890 194.220 ;
        RECT 135.650 194.160 135.970 194.220 ;
        RECT 138.370 194.160 138.690 194.220 ;
        RECT 139.310 194.220 142.090 194.360 ;
        RECT 114.230 193.900 114.550 193.960 ;
        RECT 120.010 193.900 120.330 193.960 ;
        RECT 123.410 193.900 123.730 193.960 ;
        RECT 139.310 193.900 139.450 194.220 ;
        RECT 139.730 194.160 140.050 194.220 ;
        RECT 141.770 194.160 142.090 194.220 ;
        RECT 144.150 194.360 144.470 194.420 ;
        RECT 146.295 194.360 146.685 194.440 ;
        RECT 153.365 194.360 157.365 194.430 ;
        RECT 144.150 194.220 157.365 194.360 ;
        RECT 144.150 194.160 144.470 194.220 ;
        RECT 146.295 194.140 146.685 194.220 ;
        RECT 153.365 194.150 157.365 194.220 ;
        RECT 114.230 193.760 139.450 193.900 ;
        RECT 114.230 193.700 114.550 193.760 ;
        RECT 120.010 193.700 120.330 193.760 ;
        RECT 123.410 193.700 123.730 193.760 ;
        RECT 111.510 193.440 111.830 193.500 ;
        RECT 112.190 193.440 112.510 193.500 ;
        RECT 114.230 193.440 114.550 193.500 ;
        RECT 111.510 193.300 114.550 193.440 ;
        RECT 111.510 193.240 111.830 193.300 ;
        RECT 112.190 193.240 112.510 193.300 ;
        RECT 114.230 193.240 114.550 193.300 ;
        RECT 138.710 193.440 139.030 193.500 ;
        RECT 140.750 193.440 141.070 193.500 ;
        RECT 138.710 193.300 141.070 193.440 ;
        RECT 138.710 193.240 139.030 193.300 ;
        RECT 140.750 193.240 141.070 193.300 ;
        RECT 118.990 192.980 119.310 193.040 ;
        RECT 119.670 192.980 119.990 193.040 ;
        RECT 127.150 192.980 127.470 193.040 ;
        RECT 118.990 192.840 127.470 192.980 ;
        RECT 118.990 192.780 119.310 192.840 ;
        RECT 119.670 192.780 119.990 192.840 ;
        RECT 127.150 192.780 127.470 192.840 ;
        RECT 113.355 192.520 113.725 192.590 ;
        RECT 116.950 192.520 117.270 192.580 ;
        RECT 113.355 192.380 117.270 192.520 ;
        RECT 113.355 192.310 113.725 192.380 ;
        RECT 116.950 192.320 117.270 192.380 ;
        RECT 125.450 192.520 125.770 192.580 ;
        RECT 128.850 192.520 129.170 192.580 ;
        RECT 135.310 192.520 135.630 192.580 ;
        RECT 125.450 192.380 135.630 192.520 ;
        RECT 125.450 192.320 125.770 192.380 ;
        RECT 128.850 192.320 129.170 192.380 ;
        RECT 135.310 192.320 135.630 192.380 ;
        RECT 141.770 192.520 142.090 192.580 ;
        RECT 144.830 192.520 145.150 192.580 ;
        RECT 141.770 192.380 145.150 192.520 ;
        RECT 141.770 192.320 142.090 192.380 ;
        RECT 144.830 192.320 145.150 192.380 ;
        RECT 130.890 191.600 131.210 191.660 ;
        RECT 132.590 191.600 132.910 191.660 ;
        RECT 130.890 191.460 132.910 191.600 ;
        RECT 130.890 191.400 131.210 191.460 ;
        RECT 132.590 191.400 132.910 191.460 ;
        RECT 99.600 191.140 103.600 191.210 ;
        RECT 109.640 191.140 109.960 191.200 ;
        RECT 110.830 191.140 111.150 191.200 ;
        RECT 99.600 191.000 111.150 191.140 ;
        RECT 99.600 190.930 103.600 191.000 ;
        RECT 109.640 190.940 109.960 191.000 ;
        RECT 110.830 190.940 111.150 191.000 ;
        RECT 116.950 191.140 117.270 191.200 ;
        RECT 123.555 191.140 123.925 191.210 ;
        RECT 116.950 191.000 123.925 191.140 ;
        RECT 116.950 190.940 117.270 191.000 ;
        RECT 123.555 190.930 123.925 191.000 ;
        RECT 145.170 191.140 145.490 191.200 ;
        RECT 146.770 191.140 147.030 191.230 ;
        RECT 153.365 191.140 157.365 191.210 ;
        RECT 145.170 191.000 157.365 191.140 ;
        RECT 145.170 190.940 145.490 191.000 ;
        RECT 146.770 190.910 147.030 191.000 ;
        RECT 153.365 190.930 157.365 191.000 ;
        RECT 111.510 190.680 111.830 190.740 ;
        RECT 118.990 190.680 119.310 190.740 ;
        RECT 122.390 190.680 122.710 190.740 ;
        RECT 111.510 190.540 122.710 190.680 ;
        RECT 111.510 190.480 111.830 190.540 ;
        RECT 118.990 190.480 119.310 190.540 ;
        RECT 122.390 190.480 122.710 190.540 ;
        RECT 130.890 190.680 131.210 190.740 ;
        RECT 136.330 190.680 136.650 190.740 ;
        RECT 143.470 190.680 143.790 190.740 ;
        RECT 130.890 190.540 143.790 190.680 ;
        RECT 130.890 190.480 131.210 190.540 ;
        RECT 136.330 190.480 136.650 190.540 ;
        RECT 143.470 190.480 143.790 190.540 ;
        RECT 125.450 190.220 125.770 190.280 ;
        RECT 127.150 190.220 127.470 190.280 ;
        RECT 125.450 190.080 127.470 190.220 ;
        RECT 125.450 190.020 125.770 190.080 ;
        RECT 127.150 190.020 127.470 190.080 ;
        RECT 136.670 190.220 136.990 190.280 ;
        RECT 136.670 190.080 142.000 190.220 ;
        RECT 136.670 190.020 136.990 190.080 ;
        RECT 141.860 189.830 142.000 190.080 ;
        RECT 116.755 189.820 117.125 189.830 ;
        RECT 141.860 189.820 142.285 189.830 ;
        RECT 116.755 189.560 117.270 189.820 ;
        RECT 120.690 189.760 121.010 189.820 ;
        RECT 121.710 189.760 122.030 189.820 ;
        RECT 120.690 189.620 122.030 189.760 ;
        RECT 120.690 189.560 121.010 189.620 ;
        RECT 121.710 189.560 122.030 189.620 ;
        RECT 127.830 189.760 128.150 189.820 ;
        RECT 133.270 189.760 133.590 189.820 ;
        RECT 135.650 189.760 135.970 189.820 ;
        RECT 136.670 189.760 136.990 189.820 ;
        RECT 127.830 189.620 128.570 189.760 ;
        RECT 127.830 189.560 128.150 189.620 ;
        RECT 116.755 189.550 117.125 189.560 ;
        RECT 126.955 188.840 127.325 188.910 ;
        RECT 127.830 188.840 128.150 188.900 ;
        RECT 126.955 188.700 128.150 188.840 ;
        RECT 128.430 188.840 128.570 189.620 ;
        RECT 133.270 189.620 136.990 189.760 ;
        RECT 133.270 189.560 133.590 189.620 ;
        RECT 135.650 189.560 135.970 189.620 ;
        RECT 136.670 189.560 136.990 189.620 ;
        RECT 141.770 189.560 142.285 189.820 ;
        RECT 141.915 189.550 142.285 189.560 ;
        RECT 139.730 189.300 140.050 189.360 ;
        RECT 141.090 189.300 141.410 189.360 ;
        RECT 144.150 189.300 144.470 189.360 ;
        RECT 139.730 189.160 144.470 189.300 ;
        RECT 139.730 189.100 140.050 189.160 ;
        RECT 141.090 189.100 141.410 189.160 ;
        RECT 144.150 189.100 144.470 189.160 ;
        RECT 133.950 188.840 134.270 188.900 ;
        RECT 128.430 188.700 134.270 188.840 ;
        RECT 126.955 188.630 127.325 188.700 ;
        RECT 127.830 188.640 128.150 188.700 ;
        RECT 133.950 188.640 134.270 188.700 ;
        RECT 111.850 188.380 112.170 188.440 ;
        RECT 114.230 188.380 114.550 188.440 ;
        RECT 116.270 188.380 116.590 188.440 ;
        RECT 111.850 188.240 116.590 188.380 ;
        RECT 111.850 188.180 112.170 188.240 ;
        RECT 114.230 188.180 114.550 188.240 ;
        RECT 116.270 188.180 116.590 188.240 ;
        RECT 122.730 188.380 123.050 188.440 ;
        RECT 125.790 188.380 126.110 188.440 ;
        RECT 127.490 188.380 127.810 188.440 ;
        RECT 129.870 188.380 130.190 188.440 ;
        RECT 122.730 188.240 130.190 188.380 ;
        RECT 122.730 188.180 123.050 188.240 ;
        RECT 125.790 188.180 126.110 188.240 ;
        RECT 127.490 188.180 127.810 188.240 ;
        RECT 129.870 188.180 130.190 188.240 ;
        RECT 109.955 187.920 110.325 187.990 ;
        RECT 111.510 187.920 111.830 187.980 ;
        RECT 109.955 187.780 111.830 187.920 ;
        RECT 109.955 187.710 110.325 187.780 ;
        RECT 111.510 187.720 111.830 187.780 ;
        RECT 114.570 187.920 114.890 187.980 ;
        RECT 116.270 187.920 116.590 187.980 ;
        RECT 114.570 187.780 116.590 187.920 ;
        RECT 114.570 187.720 114.890 187.780 ;
        RECT 116.270 187.720 116.590 187.780 ;
        RECT 117.970 187.920 118.290 187.980 ;
        RECT 119.670 187.920 119.990 187.980 ;
        RECT 122.390 187.920 122.710 187.980 ;
        RECT 117.970 187.780 122.710 187.920 ;
        RECT 117.970 187.720 118.290 187.780 ;
        RECT 119.670 187.720 119.990 187.780 ;
        RECT 122.390 187.720 122.710 187.780 ;
        RECT 123.410 187.920 123.730 187.980 ;
        RECT 133.610 187.920 133.930 187.980 ;
        RECT 123.410 187.780 133.930 187.920 ;
        RECT 123.410 187.720 123.730 187.780 ;
        RECT 133.610 187.720 133.930 187.780 ;
        RECT 120.155 187.520 120.525 187.530 ;
        RECT 112.190 187.460 112.510 187.520 ;
        RECT 117.630 187.460 117.950 187.520 ;
        RECT 112.190 187.320 117.950 187.460 ;
        RECT 112.190 187.260 112.510 187.320 ;
        RECT 117.630 187.260 117.950 187.320 ;
        RECT 120.010 187.260 120.525 187.520 ;
        RECT 138.710 187.460 139.030 187.520 ;
        RECT 140.750 187.460 141.070 187.520 ;
        RECT 138.710 187.320 141.070 187.460 ;
        RECT 138.710 187.260 139.030 187.320 ;
        RECT 140.750 187.260 141.070 187.320 ;
        RECT 120.155 187.250 120.525 187.260 ;
        RECT 112.530 187.000 112.850 187.060 ;
        RECT 116.950 187.000 117.270 187.060 ;
        RECT 118.990 187.000 119.310 187.060 ;
        RECT 125.450 187.000 125.770 187.060 ;
        RECT 112.530 186.860 125.770 187.000 ;
        RECT 112.530 186.800 112.850 186.860 ;
        RECT 116.950 186.800 117.270 186.860 ;
        RECT 118.990 186.800 119.310 186.860 ;
        RECT 125.450 186.800 125.770 186.860 ;
        RECT 133.270 187.000 133.590 187.060 ;
        RECT 136.330 187.000 136.650 187.060 ;
        RECT 137.010 187.000 137.330 187.060 ;
        RECT 143.470 187.000 143.790 187.060 ;
        RECT 133.270 186.860 143.790 187.000 ;
        RECT 133.270 186.800 133.590 186.860 ;
        RECT 136.330 186.800 136.650 186.860 ;
        RECT 137.010 186.800 137.330 186.860 ;
        RECT 143.470 186.800 143.790 186.860 ;
        RECT 117.970 186.540 118.290 186.600 ;
        RECT 125.450 186.540 125.770 186.600 ;
        RECT 117.970 186.400 125.770 186.540 ;
        RECT 117.970 186.340 118.290 186.400 ;
        RECT 125.450 186.340 125.770 186.400 ;
        RECT 126.130 186.540 126.450 186.600 ;
        RECT 127.830 186.540 128.150 186.600 ;
        RECT 126.130 186.400 128.150 186.540 ;
        RECT 126.130 186.340 126.450 186.400 ;
        RECT 127.830 186.340 128.150 186.400 ;
        RECT 128.510 186.540 128.830 186.600 ;
        RECT 133.270 186.540 133.590 186.600 ;
        RECT 139.730 186.540 140.050 186.600 ;
        RECT 141.770 186.540 142.090 186.600 ;
        RECT 128.510 186.400 139.450 186.540 ;
        RECT 128.510 186.340 128.830 186.400 ;
        RECT 133.270 186.340 133.590 186.400 ;
        RECT 116.950 186.080 117.270 186.140 ;
        RECT 120.010 186.080 120.330 186.140 ;
        RECT 116.950 185.940 120.330 186.080 ;
        RECT 116.950 185.880 117.270 185.940 ;
        RECT 120.010 185.880 120.330 185.940 ;
        RECT 120.690 186.080 121.010 186.140 ;
        RECT 125.110 186.080 125.430 186.140 ;
        RECT 120.690 185.940 125.430 186.080 ;
        RECT 120.690 185.880 121.010 185.940 ;
        RECT 125.110 185.880 125.430 185.940 ;
        RECT 127.830 186.080 128.150 186.140 ;
        RECT 130.890 186.080 131.210 186.140 ;
        RECT 127.830 185.940 131.210 186.080 ;
        RECT 127.830 185.880 128.150 185.940 ;
        RECT 130.890 185.880 131.210 185.940 ;
        RECT 133.755 186.080 134.125 186.150 ;
        RECT 138.710 186.080 139.030 186.140 ;
        RECT 133.755 185.940 139.030 186.080 ;
        RECT 139.310 186.080 139.450 186.400 ;
        RECT 139.730 186.400 142.090 186.540 ;
        RECT 139.730 186.340 140.050 186.400 ;
        RECT 141.770 186.340 142.090 186.400 ;
        RECT 144.150 186.540 144.470 186.600 ;
        RECT 147.355 186.540 147.725 186.610 ;
        RECT 144.150 186.400 147.725 186.540 ;
        RECT 144.150 186.340 144.470 186.400 ;
        RECT 147.355 186.330 147.725 186.400 ;
        RECT 141.090 186.080 141.410 186.140 ;
        RECT 139.310 185.940 141.410 186.080 ;
        RECT 133.755 185.870 134.125 185.940 ;
        RECT 138.710 185.880 139.030 185.940 ;
        RECT 141.090 185.880 141.410 185.940 ;
        RECT 120.350 185.620 120.670 185.680 ;
        RECT 122.390 185.620 122.710 185.680 ;
        RECT 127.490 185.620 127.810 185.680 ;
        RECT 120.350 185.480 127.810 185.620 ;
        RECT 120.350 185.420 120.670 185.480 ;
        RECT 122.390 185.420 122.710 185.480 ;
        RECT 127.490 185.420 127.810 185.480 ;
        RECT 134.290 185.620 134.610 185.680 ;
        RECT 136.330 185.620 136.650 185.680 ;
        RECT 134.290 185.480 136.650 185.620 ;
        RECT 134.290 185.420 134.610 185.480 ;
        RECT 136.330 185.420 136.650 185.480 ;
        RECT 143.955 185.220 144.325 185.230 ;
        RECT 115.250 185.160 115.570 185.220 ;
        RECT 122.390 185.160 122.710 185.220 ;
        RECT 115.250 185.020 122.710 185.160 ;
        RECT 115.250 184.960 115.570 185.020 ;
        RECT 122.390 184.960 122.710 185.020 ;
        RECT 128.850 185.160 129.170 185.220 ;
        RECT 133.270 185.160 133.590 185.220 ;
        RECT 138.030 185.160 138.350 185.220 ;
        RECT 128.850 185.020 133.590 185.160 ;
        RECT 128.850 184.960 129.170 185.020 ;
        RECT 133.270 184.960 133.590 185.020 ;
        RECT 133.870 185.020 138.350 185.160 ;
        RECT 112.530 184.700 112.850 184.760 ;
        RECT 116.950 184.700 117.270 184.760 ;
        RECT 112.530 184.560 117.270 184.700 ;
        RECT 112.530 184.500 112.850 184.560 ;
        RECT 116.950 184.500 117.270 184.560 ;
        RECT 119.670 184.700 119.990 184.760 ;
        RECT 125.450 184.700 125.770 184.760 ;
        RECT 119.670 184.560 125.770 184.700 ;
        RECT 119.670 184.500 119.990 184.560 ;
        RECT 125.450 184.500 125.770 184.560 ;
        RECT 130.890 184.700 131.210 184.760 ;
        RECT 133.270 184.700 133.590 184.760 ;
        RECT 133.870 184.700 134.010 185.020 ;
        RECT 138.030 184.960 138.350 185.020 ;
        RECT 143.955 184.960 144.470 185.220 ;
        RECT 143.955 184.950 144.325 184.960 ;
        RECT 130.890 184.560 134.010 184.700 ;
        RECT 137.010 184.700 137.330 184.760 ;
        RECT 138.030 184.700 138.350 184.760 ;
        RECT 137.010 184.560 138.350 184.700 ;
        RECT 130.890 184.500 131.210 184.560 ;
        RECT 133.270 184.500 133.590 184.560 ;
        RECT 137.010 184.500 137.330 184.560 ;
        RECT 138.030 184.500 138.350 184.560 ;
        RECT 106.555 184.265 106.925 184.310 ;
        RECT 101.185 184.240 107.485 184.265 ;
        RECT 117.290 184.240 117.610 184.300 ;
        RECT 101.185 184.100 117.610 184.240 ;
        RECT 101.185 184.075 107.485 184.100 ;
        RECT 101.185 102.165 101.375 184.075 ;
        RECT 106.555 184.030 106.925 184.075 ;
        RECT 117.290 184.040 117.610 184.100 ;
        RECT 133.950 184.240 134.270 184.300 ;
        RECT 136.330 184.240 136.650 184.300 ;
        RECT 143.470 184.240 143.790 184.300 ;
        RECT 133.950 184.100 143.790 184.240 ;
        RECT 133.950 184.040 134.270 184.100 ;
        RECT 136.330 184.040 136.650 184.100 ;
        RECT 143.470 184.040 143.790 184.100 ;
        RECT 114.230 183.780 114.550 183.840 ;
        RECT 116.950 183.780 117.270 183.840 ;
        RECT 119.330 183.780 119.650 183.840 ;
        RECT 114.230 183.640 119.650 183.780 ;
        RECT 114.230 183.580 114.550 183.640 ;
        RECT 116.950 183.580 117.270 183.640 ;
        RECT 119.330 183.580 119.650 183.640 ;
        RECT 130.355 183.780 130.725 183.850 ;
        RECT 130.890 183.780 131.210 183.840 ;
        RECT 130.355 183.640 131.210 183.780 ;
        RECT 130.355 183.570 130.725 183.640 ;
        RECT 130.890 183.580 131.210 183.640 ;
        RECT 137.155 183.780 137.525 183.850 ;
        RECT 138.710 183.780 139.030 183.840 ;
        RECT 137.155 183.640 139.030 183.780 ;
        RECT 137.155 183.570 137.525 183.640 ;
        RECT 138.710 183.580 139.030 183.640 ;
        RECT 140.555 183.780 140.925 183.850 ;
        RECT 141.770 183.780 142.090 183.840 ;
        RECT 140.555 183.640 142.090 183.780 ;
        RECT 140.555 183.570 140.925 183.640 ;
        RECT 141.770 183.580 142.090 183.640 ;
        RECT 144.150 183.780 144.470 183.840 ;
        RECT 150.755 183.780 151.125 183.850 ;
        RECT 144.150 183.640 151.125 183.780 ;
        RECT 144.150 183.580 144.470 183.640 ;
        RECT 116.750 181.695 117.190 181.830 ;
        RECT 101.635 181.520 117.190 181.695 ;
        RECT 146.340 181.670 146.480 183.640 ;
        RECT 150.755 183.570 151.125 183.640 ;
        RECT 101.635 117.240 101.810 181.520 ;
        RECT 116.750 181.390 117.190 181.520 ;
        RECT 141.150 181.530 146.480 181.670 ;
        RECT 120.120 181.145 120.560 181.300 ;
        RECT 102.045 180.970 120.560 181.145 ;
        RECT 102.045 132.280 102.220 180.970 ;
        RECT 120.120 180.860 120.560 180.970 ;
        RECT 123.510 180.750 123.950 181.190 ;
        RECT 113.350 180.630 113.790 180.730 ;
        RECT 102.550 180.425 113.790 180.630 ;
        RECT 123.660 180.610 123.820 180.750 ;
        RECT 102.550 147.295 102.755 180.425 ;
        RECT 113.350 180.290 113.790 180.425 ;
        RECT 119.440 180.450 123.820 180.610 ;
        RECT 126.900 180.590 127.320 181.050 ;
        RECT 130.330 180.670 130.750 181.130 ;
        RECT 133.740 180.820 134.190 181.260 ;
        RECT 140.530 180.830 140.980 181.270 ;
        RECT 109.955 180.005 110.325 180.050 ;
        RECT 103.055 179.815 110.325 180.005 ;
        RECT 103.055 162.300 103.245 179.815 ;
        RECT 109.955 179.770 110.325 179.815 ;
        RECT 107.160 173.250 107.860 173.260 ;
        RECT 106.820 172.510 108.170 173.250 ;
        RECT 107.160 163.080 107.860 172.510 ;
        RECT 118.090 171.510 118.680 173.070 ;
        RECT 116.840 169.115 117.160 169.160 ;
        RECT 116.840 168.945 119.235 169.115 ;
        RECT 116.840 168.900 117.160 168.945 ;
        RECT 109.210 167.560 117.200 167.950 ;
        RECT 109.170 165.675 109.490 165.730 ;
        RECT 108.370 165.525 109.490 165.675 ;
        RECT 103.020 161.980 103.280 162.300 ;
        RECT 107.070 162.290 107.930 163.080 ;
        RECT 107.160 158.260 107.860 158.270 ;
        RECT 106.820 157.520 108.170 158.260 ;
        RECT 107.160 148.090 107.860 157.520 ;
        RECT 108.370 150.655 108.520 165.525 ;
        RECT 109.170 165.470 109.490 165.525 ;
        RECT 111.750 164.500 114.410 167.560 ;
        RECT 109.250 164.050 117.190 164.500 ;
        RECT 116.820 154.090 117.140 154.150 ;
        RECT 116.820 153.950 118.920 154.090 ;
        RECT 116.820 153.890 117.140 153.950 ;
        RECT 109.210 152.570 117.200 152.960 ;
        RECT 109.240 150.655 109.560 150.710 ;
        RECT 108.370 150.505 109.560 150.655 ;
        RECT 103.120 147.295 103.440 147.320 ;
        RECT 107.070 147.300 107.930 148.090 ;
        RECT 102.550 147.090 103.440 147.295 ;
        RECT 103.120 147.060 103.440 147.090 ;
        RECT 107.160 143.280 107.860 143.290 ;
        RECT 106.820 142.540 108.170 143.280 ;
        RECT 107.160 133.110 107.860 142.540 ;
        RECT 108.370 135.665 108.520 150.505 ;
        RECT 109.240 150.450 109.560 150.505 ;
        RECT 111.750 149.510 114.410 152.570 ;
        RECT 109.250 149.060 117.190 149.510 ;
        RECT 116.895 139.165 117.215 139.195 ;
        RECT 116.895 138.970 118.465 139.165 ;
        RECT 116.895 138.935 117.215 138.970 ;
        RECT 109.210 137.590 117.200 137.980 ;
        RECT 109.270 135.665 109.590 135.720 ;
        RECT 108.370 135.515 109.590 135.665 ;
        RECT 107.070 132.320 107.930 133.110 ;
        RECT 103.170 132.280 103.490 132.320 ;
        RECT 102.045 132.105 103.490 132.280 ;
        RECT 103.170 132.060 103.490 132.105 ;
        RECT 107.160 128.250 107.860 128.260 ;
        RECT 106.820 127.510 108.170 128.250 ;
        RECT 107.160 118.080 107.860 127.510 ;
        RECT 108.370 125.015 108.520 135.515 ;
        RECT 109.270 135.460 109.590 135.515 ;
        RECT 111.750 134.530 114.410 137.590 ;
        RECT 109.250 134.080 117.190 134.530 ;
        RECT 108.370 124.865 110.295 125.015 ;
        RECT 109.030 124.210 109.350 124.240 ;
        RECT 108.310 124.010 109.350 124.210 ;
        RECT 107.070 117.290 107.930 118.080 ;
        RECT 103.090 117.240 103.410 117.280 ;
        RECT 101.635 117.065 103.410 117.240 ;
        RECT 103.090 117.020 103.410 117.065 ;
        RECT 107.160 113.260 107.860 113.270 ;
        RECT 106.820 112.520 108.170 113.260 ;
        RECT 107.160 103.090 107.860 112.520 ;
        RECT 108.310 109.590 108.510 124.010 ;
        RECT 109.030 123.980 109.350 124.010 ;
        RECT 110.145 123.615 110.295 124.865 ;
        RECT 108.805 123.465 110.295 123.615 ;
        RECT 108.805 120.695 108.955 123.465 ;
        RECT 109.210 122.560 117.200 122.950 ;
        RECT 109.200 120.695 109.520 120.750 ;
        RECT 108.805 120.545 109.520 120.695 ;
        RECT 108.830 120.490 109.520 120.545 ;
        RECT 108.830 120.410 109.420 120.490 ;
        RECT 108.830 114.240 109.090 120.410 ;
        RECT 111.750 119.500 114.410 122.560 ;
        RECT 109.250 119.050 117.190 119.500 ;
        RECT 108.855 114.090 109.065 114.240 ;
        RECT 117.310 114.090 117.590 114.125 ;
        RECT 108.855 113.790 117.600 114.090 ;
        RECT 108.855 110.765 109.065 113.790 ;
        RECT 117.310 113.755 117.590 113.790 ;
        RECT 108.855 110.555 110.595 110.765 ;
        RECT 108.310 109.390 110.100 109.590 ;
        RECT 109.330 109.220 109.650 109.245 ;
        RECT 108.095 109.015 109.650 109.220 ;
        RECT 102.810 102.165 103.270 102.600 ;
        RECT 107.070 102.300 107.930 103.090 ;
        RECT 101.185 101.975 103.270 102.165 ;
        RECT 102.810 101.540 103.270 101.975 ;
        RECT 108.095 101.470 108.300 109.015 ;
        RECT 109.330 108.985 109.650 109.015 ;
        RECT 109.900 108.750 110.100 109.390 ;
        RECT 106.220 101.265 108.300 101.470 ;
        RECT 108.490 108.550 110.100 108.750 ;
        RECT 106.220 97.090 106.425 101.265 ;
        RECT 108.490 100.980 108.690 108.550 ;
        RECT 110.385 108.370 110.595 110.555 ;
        RECT 108.920 108.255 110.595 108.370 ;
        RECT 108.920 108.230 110.560 108.255 ;
        RECT 108.920 105.580 109.060 108.230 ;
        RECT 109.210 107.570 117.200 107.960 ;
        RECT 109.310 105.580 109.630 105.640 ;
        RECT 108.920 105.440 109.630 105.580 ;
        RECT 109.310 105.380 109.630 105.440 ;
        RECT 111.750 104.510 114.410 107.570 ;
        RECT 109.250 104.060 117.190 104.510 ;
        RECT 118.270 101.295 118.465 138.970 ;
        RECT 107.600 100.780 108.690 100.980 ;
        RECT 110.905 101.100 118.465 101.295 ;
        RECT 107.600 97.770 107.800 100.780 ;
        RECT 107.480 97.210 107.930 97.770 ;
        RECT 110.905 97.760 111.100 101.100 ;
        RECT 118.780 100.700 118.920 153.950 ;
        RECT 113.790 100.560 118.920 100.700 ;
        RECT 110.780 97.200 111.230 97.760 ;
        RECT 113.790 97.710 113.930 100.560 ;
        RECT 119.065 100.255 119.235 168.945 ;
        RECT 119.440 102.400 119.600 180.450 ;
        RECT 127.065 180.240 127.220 180.590 ;
        RECT 119.865 180.085 127.220 180.240 ;
        RECT 119.865 117.270 120.020 180.085 ;
        RECT 130.435 179.830 130.620 180.670 ;
        RECT 120.210 179.645 130.620 179.830 ;
        RECT 120.210 132.445 120.395 179.645 ;
        RECT 133.865 179.400 134.020 180.820 ;
        RECT 120.635 179.245 134.020 179.400 ;
        RECT 120.635 147.340 120.790 179.245 ;
        RECT 140.650 178.990 140.830 180.830 ;
        RECT 120.970 178.810 140.830 178.990 ;
        RECT 120.970 162.360 121.150 178.810 ;
        RECT 141.150 178.580 141.290 181.530 ;
        RECT 143.920 181.075 144.370 181.200 ;
        RECT 147.310 181.115 147.760 181.260 ;
        RECT 139.040 178.440 141.290 178.580 ;
        RECT 141.505 180.880 144.370 181.075 ;
        RECT 126.200 173.280 126.900 173.290 ;
        RECT 125.860 172.540 127.210 173.280 ;
        RECT 126.200 163.110 126.900 172.540 ;
        RECT 137.110 171.290 137.760 172.900 ;
        RECT 135.805 169.165 136.125 169.195 ;
        RECT 135.805 168.970 138.795 169.165 ;
        RECT 135.805 168.935 136.125 168.970 ;
        RECT 128.250 167.590 136.240 167.980 ;
        RECT 128.220 165.725 128.540 165.780 ;
        RECT 127.280 165.575 128.540 165.725 ;
        RECT 122.150 162.360 122.470 162.400 ;
        RECT 120.970 162.180 122.470 162.360 ;
        RECT 126.110 162.320 126.970 163.110 ;
        RECT 122.150 162.140 122.470 162.180 ;
        RECT 127.280 159.925 127.430 165.575 ;
        RECT 128.220 165.520 128.540 165.575 ;
        RECT 130.790 164.530 133.450 167.590 ;
        RECT 128.290 164.080 136.230 164.530 ;
        RECT 127.280 159.610 127.535 159.925 ;
        RECT 126.200 158.260 126.900 158.270 ;
        RECT 125.860 157.520 127.210 158.260 ;
        RECT 126.200 148.090 126.900 157.520 ;
        RECT 127.385 150.635 127.535 159.610 ;
        RECT 135.980 154.145 136.300 154.200 ;
        RECT 135.980 153.995 138.395 154.145 ;
        RECT 135.980 153.940 136.300 153.995 ;
        RECT 128.250 152.570 136.240 152.960 ;
        RECT 128.210 150.635 128.530 150.690 ;
        RECT 127.385 150.485 128.530 150.635 ;
        RECT 122.100 147.340 122.420 147.390 ;
        RECT 120.635 147.185 122.420 147.340 ;
        RECT 126.110 147.300 126.970 148.090 ;
        RECT 122.100 147.130 122.420 147.185 ;
        RECT 126.150 143.240 126.850 143.250 ;
        RECT 125.810 142.500 127.160 143.240 ;
        RECT 126.150 133.070 126.850 142.500 ;
        RECT 127.385 135.645 127.535 150.485 ;
        RECT 128.210 150.430 128.530 150.485 ;
        RECT 130.790 149.510 133.450 152.570 ;
        RECT 128.290 149.060 136.230 149.510 ;
        RECT 135.860 139.115 136.180 139.170 ;
        RECT 135.860 138.965 138.035 139.115 ;
        RECT 135.860 138.910 136.180 138.965 ;
        RECT 128.200 137.550 136.190 137.940 ;
        RECT 128.140 135.645 128.460 135.700 ;
        RECT 127.385 135.495 128.460 135.645 ;
        RECT 120.210 132.430 122.260 132.445 ;
        RECT 120.210 132.260 122.340 132.430 ;
        RECT 126.060 132.280 126.920 133.070 ;
        RECT 120.230 132.230 122.340 132.260 ;
        RECT 122.020 132.170 122.340 132.230 ;
        RECT 126.150 128.220 126.850 128.230 ;
        RECT 125.810 127.480 127.160 128.220 ;
        RECT 126.150 118.050 126.850 127.480 ;
        RECT 127.385 120.635 127.535 135.495 ;
        RECT 128.140 135.440 128.460 135.495 ;
        RECT 130.740 134.490 133.400 137.550 ;
        RECT 128.240 134.040 136.180 134.490 ;
        RECT 135.745 124.170 136.065 124.205 ;
        RECT 135.745 123.985 137.700 124.170 ;
        RECT 135.745 123.945 136.065 123.985 ;
        RECT 128.200 122.530 136.190 122.920 ;
        RECT 128.230 120.635 128.550 120.690 ;
        RECT 127.385 120.485 128.550 120.635 ;
        RECT 122.010 117.270 122.330 117.320 ;
        RECT 119.865 117.115 122.330 117.270 ;
        RECT 126.060 117.260 126.920 118.050 ;
        RECT 122.010 117.060 122.330 117.115 ;
        RECT 127.385 114.695 127.535 120.485 ;
        RECT 128.230 120.430 128.550 120.485 ;
        RECT 130.740 119.470 133.400 122.530 ;
        RECT 128.240 119.020 136.180 119.470 ;
        RECT 127.080 114.395 127.745 114.695 ;
        RECT 127.110 114.090 127.710 114.395 ;
        RECT 136.030 114.090 136.310 114.125 ;
        RECT 120.045 113.790 136.320 114.090 ;
        RECT 126.150 113.240 126.850 113.250 ;
        RECT 125.810 112.500 127.160 113.240 ;
        RECT 126.150 103.070 126.850 112.500 ;
        RECT 127.385 105.635 127.535 113.790 ;
        RECT 136.030 113.755 136.310 113.790 ;
        RECT 135.945 109.090 136.265 109.135 ;
        RECT 135.945 108.925 137.270 109.090 ;
        RECT 135.945 108.875 136.265 108.925 ;
        RECT 128.200 107.550 136.190 107.940 ;
        RECT 128.190 105.635 128.510 105.690 ;
        RECT 127.385 105.485 128.510 105.635 ;
        RECT 128.190 105.430 128.510 105.485 ;
        RECT 130.740 104.490 133.400 107.550 ;
        RECT 128.240 104.040 136.180 104.490 ;
        RECT 122.100 102.400 122.420 102.450 ;
        RECT 119.440 102.240 122.420 102.400 ;
        RECT 126.060 102.280 126.920 103.070 ;
        RECT 122.100 102.190 122.420 102.240 ;
        RECT 137.105 101.300 137.270 108.925 ;
        RECT 116.935 100.085 119.235 100.255 ;
        RECT 119.820 101.135 137.270 101.300 ;
        RECT 116.935 97.760 117.105 100.085 ;
        RECT 113.610 97.150 114.060 97.710 ;
        RECT 116.800 97.200 117.250 97.760 ;
        RECT 119.820 97.670 119.985 101.135 ;
        RECT 137.515 100.830 137.700 123.985 ;
        RECT 122.660 100.645 137.700 100.830 ;
        RECT 122.660 97.690 122.845 100.645 ;
        RECT 137.885 100.395 138.035 138.965 ;
        RECT 125.535 100.245 138.035 100.395 ;
        RECT 125.535 97.690 125.685 100.245 ;
        RECT 138.245 99.985 138.395 153.995 ;
        RECT 128.955 99.835 138.395 99.985 ;
        RECT 128.955 97.740 129.105 99.835 ;
        RECT 138.600 99.625 138.795 168.970 ;
        RECT 139.040 102.260 139.180 178.440 ;
        RECT 141.505 178.220 141.700 180.880 ;
        RECT 143.920 180.760 144.370 180.880 ;
        RECT 144.755 180.940 147.760 181.115 ;
        RECT 144.755 180.450 144.930 180.940 ;
        RECT 147.310 180.820 147.760 180.940 ;
        RECT 139.340 178.060 141.700 178.220 ;
        RECT 139.340 117.270 139.500 178.060 ;
        RECT 141.505 178.045 141.700 178.060 ;
        RECT 141.945 180.275 144.930 180.450 ;
        RECT 141.945 177.830 142.120 180.275 ;
        RECT 146.305 180.200 146.675 180.480 ;
        RECT 146.390 180.005 146.595 180.200 ;
        RECT 139.740 177.455 140.020 177.825 ;
        RECT 140.245 177.655 142.120 177.830 ;
        RECT 142.370 179.800 146.595 180.005 ;
        RECT 139.790 132.320 139.970 177.455 ;
        RECT 140.245 147.250 140.420 177.655 ;
        RECT 142.370 177.455 142.575 179.800 ;
        RECT 140.570 177.250 142.575 177.455 ;
        RECT 140.570 162.425 140.775 177.250 ;
        RECT 145.150 173.320 145.850 173.330 ;
        RECT 144.810 172.580 146.160 173.320 ;
        RECT 145.150 163.150 145.850 172.580 ;
        RECT 156.130 171.410 156.780 173.020 ;
        RECT 154.830 169.185 155.150 169.220 ;
        RECT 154.830 168.995 156.715 169.185 ;
        RECT 154.830 168.960 155.150 168.995 ;
        RECT 147.200 167.630 155.190 168.020 ;
        RECT 147.180 165.725 147.500 165.780 ;
        RECT 146.290 165.575 147.500 165.725 ;
        RECT 141.030 162.425 141.350 162.450 ;
        RECT 140.570 162.220 141.350 162.425 ;
        RECT 145.060 162.360 145.920 163.150 ;
        RECT 141.030 162.190 141.350 162.220 ;
        RECT 146.290 159.585 146.440 165.575 ;
        RECT 147.180 165.520 147.500 165.575 ;
        RECT 149.740 164.570 152.400 167.630 ;
        RECT 147.240 164.120 155.180 164.570 ;
        RECT 146.290 159.330 146.545 159.585 ;
        RECT 145.200 158.260 145.900 158.270 ;
        RECT 144.860 157.520 146.210 158.260 ;
        RECT 145.200 148.090 145.900 157.520 ;
        RECT 146.395 150.515 146.545 159.330 ;
        RECT 154.865 154.080 155.185 154.105 ;
        RECT 154.865 153.875 156.215 154.080 ;
        RECT 154.865 153.845 155.185 153.875 ;
        RECT 147.250 152.570 155.240 152.960 ;
        RECT 147.210 150.515 147.530 150.570 ;
        RECT 146.395 150.365 147.530 150.515 ;
        RECT 145.110 147.300 145.970 148.090 ;
        RECT 141.160 147.250 141.480 147.290 ;
        RECT 140.245 147.075 141.480 147.250 ;
        RECT 141.160 147.030 141.480 147.075 ;
        RECT 145.150 143.240 145.850 143.250 ;
        RECT 144.810 142.500 146.160 143.240 ;
        RECT 145.150 133.070 145.850 142.500 ;
        RECT 146.395 135.575 146.545 150.365 ;
        RECT 147.210 150.310 147.530 150.365 ;
        RECT 149.790 149.510 152.450 152.570 ;
        RECT 147.290 149.060 155.230 149.510 ;
        RECT 156.010 139.830 156.215 153.875 ;
        RECT 156.525 140.395 156.715 168.995 ;
        RECT 156.525 140.205 157.235 140.395 ;
        RECT 156.010 139.625 156.900 139.830 ;
        RECT 154.860 139.105 155.180 139.160 ;
        RECT 154.860 138.955 156.455 139.105 ;
        RECT 154.860 138.900 155.180 138.955 ;
        RECT 147.200 137.550 155.190 137.940 ;
        RECT 147.180 135.575 147.500 135.630 ;
        RECT 146.395 135.425 147.500 135.575 ;
        RECT 141.150 132.320 141.470 132.360 ;
        RECT 139.790 132.140 141.470 132.320 ;
        RECT 145.060 132.280 145.920 133.070 ;
        RECT 141.150 132.100 141.470 132.140 ;
        RECT 145.150 128.220 145.850 128.230 ;
        RECT 144.810 127.480 146.160 128.220 ;
        RECT 145.150 118.050 145.850 127.480 ;
        RECT 146.395 120.575 146.545 135.425 ;
        RECT 147.180 135.370 147.500 135.425 ;
        RECT 149.740 134.490 152.400 137.550 ;
        RECT 147.240 134.040 155.180 134.490 ;
        RECT 154.875 124.080 155.195 124.105 ;
        RECT 154.875 123.875 156.080 124.080 ;
        RECT 154.875 123.845 155.195 123.875 ;
        RECT 147.200 122.530 155.190 122.920 ;
        RECT 147.140 120.575 147.460 120.630 ;
        RECT 146.395 120.425 147.460 120.575 ;
        RECT 141.140 117.270 141.460 117.320 ;
        RECT 139.340 117.110 141.460 117.270 ;
        RECT 145.060 117.260 145.920 118.050 ;
        RECT 141.140 117.060 141.460 117.110 ;
        RECT 139.485 114.015 139.875 114.090 ;
        RECT 146.395 114.015 146.545 120.425 ;
        RECT 147.140 120.370 147.460 120.425 ;
        RECT 149.740 119.470 152.400 122.530 ;
        RECT 147.240 119.020 155.180 119.470 ;
        RECT 139.485 113.865 146.545 114.015 ;
        RECT 139.485 113.790 139.875 113.865 ;
        RECT 145.200 113.240 145.900 113.250 ;
        RECT 144.860 112.500 146.210 113.240 ;
        RECT 145.200 103.070 145.900 112.500 ;
        RECT 146.395 110.275 146.545 113.865 ;
        RECT 146.395 110.125 147.995 110.275 ;
        RECT 147.310 109.170 147.630 109.230 ;
        RECT 146.280 109.030 147.630 109.170 ;
        RECT 141.180 102.260 141.500 102.320 ;
        RECT 145.110 102.280 145.970 103.070 ;
        RECT 139.040 102.120 141.500 102.260 ;
        RECT 141.180 102.060 141.500 102.120 ;
        RECT 146.280 100.870 146.420 109.030 ;
        RECT 147.310 108.970 147.630 109.030 ;
        RECT 147.845 108.555 147.995 110.125 ;
        RECT 146.735 108.405 147.995 108.555 ;
        RECT 146.735 105.645 146.885 108.405 ;
        RECT 147.250 107.550 155.240 107.940 ;
        RECT 147.230 105.645 147.550 105.700 ;
        RECT 146.735 105.495 147.550 105.645 ;
        RECT 147.230 105.440 147.550 105.495 ;
        RECT 149.790 104.490 152.450 107.550 ;
        RECT 147.290 104.040 155.230 104.490 ;
        RECT 131.725 99.430 138.795 99.625 ;
        RECT 139.220 100.730 146.420 100.870 ;
        RECT 119.650 97.200 120.150 97.670 ;
        RECT 122.660 97.540 123.170 97.690 ;
        RECT 122.670 97.220 123.170 97.540 ;
        RECT 125.360 97.220 125.860 97.690 ;
        RECT 128.800 97.270 129.300 97.740 ;
        RECT 131.725 97.720 131.920 99.430 ;
        RECT 139.220 99.210 139.360 100.730 ;
        RECT 155.875 100.280 156.080 123.875 ;
        RECT 134.910 99.070 139.360 99.210 ;
        RECT 139.695 100.075 156.080 100.280 ;
        RECT 131.610 97.250 132.110 97.720 ;
        RECT 134.910 97.680 135.050 99.070 ;
        RECT 139.695 98.740 139.900 100.075 ;
        RECT 156.305 99.785 156.455 138.955 ;
        RECT 137.480 98.535 139.900 98.740 ;
        RECT 140.965 99.635 156.455 99.785 ;
        RECT 134.720 97.210 135.220 97.680 ;
        RECT 137.480 97.670 137.685 98.535 ;
        RECT 137.340 97.200 137.840 97.670 ;
        RECT 140.965 97.640 141.115 99.635 ;
        RECT 156.695 99.400 156.900 139.625 ;
        RECT 144.295 99.195 156.900 99.400 ;
        RECT 144.295 98.050 144.500 99.195 ;
        RECT 157.045 98.995 157.235 140.205 ;
        RECT 150.545 98.805 157.235 98.995 ;
        RECT 150.545 98.060 150.735 98.805 ;
        RECT 144.295 97.715 144.810 98.050 ;
        RECT 119.820 97.180 119.985 97.200 ;
        RECT 140.820 97.170 141.320 97.640 ;
        RECT 144.310 97.580 144.810 97.715 ;
        RECT 150.430 97.590 150.930 98.060 ;
        RECT 106.100 96.620 106.520 97.090 ;
      LAYER met3 ;
        RECT 63.820 225.030 64.140 225.410 ;
        RECT 63.830 217.005 64.130 225.030 ;
        RECT 66.460 224.940 66.780 225.320 ;
        RECT 69.310 225.110 69.630 225.490 ;
        RECT 66.470 217.365 66.770 224.940 ;
        RECT 69.320 221.525 69.620 225.110 ;
        RECT 72.000 224.870 72.320 225.250 ;
        RECT 74.790 224.920 75.110 225.300 ;
        RECT 69.295 221.175 69.645 221.525 ;
        RECT 72.010 221.065 72.310 224.870 ;
        RECT 71.985 220.715 72.335 221.065 ;
        RECT 74.800 220.645 75.100 224.920 ;
        RECT 77.520 224.730 77.840 225.110 ;
        RECT 80.300 224.900 80.620 225.280 ;
        RECT 74.775 220.295 75.125 220.645 ;
        RECT 77.530 217.765 77.830 224.730 ;
        RECT 80.310 220.065 80.610 224.900 ;
        RECT 83.030 224.730 83.350 225.110 ;
        RECT 85.800 224.890 86.120 225.270 ;
        RECT 88.540 224.890 88.860 225.270 ;
        RECT 80.285 219.715 80.635 220.065 ;
        RECT 83.040 219.715 83.340 224.730 ;
        RECT 83.015 219.365 83.365 219.715 ;
        RECT 85.810 219.280 86.110 224.890 ;
        RECT 85.785 218.930 86.135 219.280 ;
        RECT 88.550 218.115 88.850 224.890 ;
        RECT 91.355 224.810 91.675 225.190 ;
        RECT 91.365 218.510 91.665 224.810 ;
        RECT 94.130 224.790 94.450 225.170 ;
        RECT 143.900 225.090 144.220 225.470 ;
        RECT 94.140 218.845 94.440 224.790 ;
        RECT 113.240 219.510 113.840 223.500 ;
        RECT 113.240 219.500 114.370 219.510 ;
        RECT 123.440 219.500 124.040 223.500 ;
        RECT 130.240 219.500 130.840 223.500 ;
        RECT 137.040 219.500 137.640 223.500 ;
        RECT 140.440 219.500 141.040 223.500 ;
        RECT 113.390 219.295 114.370 219.500 ;
        RECT 113.390 219.210 114.385 219.295 ;
        RECT 114.055 218.965 114.385 219.210 ;
        RECT 91.340 218.160 91.690 218.510 ;
        RECT 94.115 218.495 94.465 218.845 ;
        RECT 88.525 217.765 88.875 218.115 ;
        RECT 77.505 217.415 77.855 217.765 ;
        RECT 66.445 217.015 66.795 217.365 ;
        RECT 63.805 216.655 64.155 217.005 ;
        RECT 123.590 216.995 123.890 219.500 ;
        RECT 130.390 218.670 130.690 219.500 ;
        RECT 130.350 218.290 130.730 218.670 ;
        RECT 130.390 216.995 130.690 218.290 ;
        RECT 137.190 216.995 137.490 219.500 ;
        RECT 140.590 218.595 140.890 219.500 ;
        RECT 143.910 218.610 144.210 225.090 ;
        RECT 140.575 218.265 140.905 218.595 ;
        RECT 123.575 216.665 123.905 216.995 ;
        RECT 130.375 216.665 130.705 216.995 ;
        RECT 137.175 216.665 137.505 216.995 ;
        RECT 140.590 205.955 140.890 218.265 ;
        RECT 143.885 218.260 144.235 218.610 ;
        RECT 141.935 207.005 142.265 207.335 ;
        RECT 140.575 205.625 140.905 205.955 ;
        RECT 141.950 203.195 142.250 207.005 ;
        RECT 141.935 202.865 142.265 203.195 ;
        RECT 8.565 202.460 10.155 202.485 ;
        RECT 1.070 200.860 10.160 202.460 ;
        RECT 108.510 202.165 109.525 202.170 ;
        RECT 108.485 201.160 109.550 202.165 ;
        RECT 8.565 200.835 10.155 200.860 ;
        RECT 106.280 197.810 107.410 198.930 ;
        RECT 106.575 184.005 106.905 184.335 ;
        RECT 106.590 180.455 106.890 184.005 ;
        RECT 106.440 176.455 107.040 180.455 ;
        RECT 108.510 173.010 109.525 201.160 ;
        RECT 113.035 200.870 113.365 202.450 ;
        RECT 118.475 200.870 118.805 202.450 ;
        RECT 123.915 200.870 124.245 202.450 ;
        RECT 129.355 200.870 129.685 202.450 ;
        RECT 134.795 200.870 135.125 202.450 ;
        RECT 140.235 200.870 140.565 202.450 ;
        RECT 110.315 197.570 110.645 199.150 ;
        RECT 115.755 197.570 116.085 199.150 ;
        RECT 121.195 197.570 121.525 199.150 ;
        RECT 126.635 197.570 126.965 199.150 ;
        RECT 132.075 197.570 132.405 199.150 ;
        RECT 137.515 197.570 137.845 199.150 ;
        RECT 113.375 192.285 113.705 192.615 ;
        RECT 109.975 187.685 110.305 188.015 ;
        RECT 109.990 180.455 110.290 187.685 ;
        RECT 113.390 180.730 113.690 192.285 ;
        RECT 123.575 190.905 123.905 191.235 ;
        RECT 116.775 189.525 117.105 189.855 ;
        RECT 116.790 181.830 117.090 189.525 ;
        RECT 120.175 187.225 120.505 187.555 ;
        RECT 116.750 181.390 117.190 181.830 ;
        RECT 113.350 180.455 113.790 180.730 ;
        RECT 116.790 180.455 117.090 181.390 ;
        RECT 120.190 181.300 120.490 187.225 ;
        RECT 120.120 180.860 120.560 181.300 ;
        RECT 123.590 181.190 123.890 190.905 ;
        RECT 141.950 189.855 142.250 202.865 ;
        RECT 145.675 200.870 146.005 202.450 ;
        RECT 142.955 197.570 143.285 199.150 ;
        RECT 146.315 194.115 146.665 194.465 ;
        RECT 141.935 189.525 142.265 189.855 ;
        RECT 126.975 188.605 127.305 188.935 ;
        RECT 120.190 180.455 120.490 180.860 ;
        RECT 123.510 180.850 123.950 181.190 ;
        RECT 126.990 181.050 127.290 188.605 ;
        RECT 133.775 185.845 134.105 186.175 ;
        RECT 130.375 183.545 130.705 183.875 ;
        RECT 130.390 181.130 130.690 183.545 ;
        RECT 133.790 181.260 134.090 185.845 ;
        RECT 143.975 184.925 144.305 185.255 ;
        RECT 137.175 183.545 137.505 183.875 ;
        RECT 140.575 183.545 140.905 183.875 ;
        RECT 123.440 180.455 124.000 180.850 ;
        RECT 126.900 180.710 127.320 181.050 ;
        RECT 130.330 180.810 130.780 181.130 ;
        RECT 133.740 180.820 134.190 181.260 ;
        RECT 126.850 180.455 127.390 180.710 ;
        RECT 130.280 180.455 130.840 180.810 ;
        RECT 133.790 180.455 134.090 180.820 ;
        RECT 137.190 180.455 137.490 183.545 ;
        RECT 140.590 181.270 140.890 183.545 ;
        RECT 140.530 180.830 140.980 181.270 ;
        RECT 143.990 181.200 144.290 184.925 ;
        RECT 140.590 180.455 140.890 180.830 ;
        RECT 143.920 180.760 144.370 181.200 ;
        RECT 143.990 180.455 144.290 180.760 ;
        RECT 146.340 180.505 146.640 194.115 ;
        RECT 147.375 186.305 147.705 186.635 ;
        RECT 147.390 181.260 147.690 186.305 ;
        RECT 150.775 183.545 151.105 183.875 ;
        RECT 147.310 180.820 147.760 181.260 ;
        RECT 109.840 176.455 110.440 180.455 ;
        RECT 113.240 176.455 113.840 180.455 ;
        RECT 116.640 176.455 117.240 180.455 ;
        RECT 120.040 176.455 120.640 180.455 ;
        RECT 123.440 176.455 124.040 180.455 ;
        RECT 126.840 176.455 127.440 180.455 ;
        RECT 130.240 176.455 130.840 180.455 ;
        RECT 133.640 176.455 134.240 180.455 ;
        RECT 137.040 177.790 137.640 180.455 ;
        RECT 139.715 177.790 140.045 177.805 ;
        RECT 137.040 177.490 140.045 177.790 ;
        RECT 137.040 176.455 137.640 177.490 ;
        RECT 139.715 177.475 140.045 177.490 ;
        RECT 140.440 176.455 141.040 180.455 ;
        RECT 143.840 176.455 144.440 180.455 ;
        RECT 146.325 180.175 146.655 180.505 ;
        RECT 147.390 180.455 147.690 180.820 ;
        RECT 150.790 180.455 151.090 183.545 ;
        RECT 147.240 176.455 147.840 180.455 ;
        RECT 150.640 176.455 151.240 180.455 ;
        RECT 118.090 173.010 118.680 173.070 ;
        RECT 156.130 173.010 156.780 173.020 ;
        RECT 108.440 171.855 156.795 173.010 ;
        RECT 118.090 171.510 118.680 171.855 ;
        RECT 137.110 171.290 137.760 171.855 ;
        RECT 156.130 171.410 156.780 171.855 ;
        RECT 117.285 114.090 117.615 114.105 ;
        RECT 120.065 114.090 120.415 114.115 ;
        RECT 117.285 113.790 120.415 114.090 ;
        RECT 117.285 113.775 117.615 113.790 ;
        RECT 120.065 113.765 120.415 113.790 ;
        RECT 127.100 113.755 127.725 114.720 ;
        RECT 136.005 114.090 136.335 114.105 ;
        RECT 139.505 114.090 139.855 114.115 ;
        RECT 136.005 113.790 139.855 114.090 ;
        RECT 136.005 113.775 136.335 113.790 ;
        RECT 139.505 113.765 139.855 113.790 ;
        RECT 127.105 113.730 127.720 113.755 ;
      LAYER met4 ;
        RECT 64.090 225.055 64.145 225.385 ;
        RECT 66.455 224.965 66.550 225.295 ;
        RECT 69.305 225.135 69.310 225.465 ;
        RECT 69.610 225.135 69.635 225.465 ;
        RECT 71.995 224.895 72.070 225.225 ;
        RECT 74.785 224.945 74.830 225.275 ;
        RECT 77.515 224.760 77.590 225.085 ;
        RECT 80.295 224.925 80.350 225.255 ;
        RECT 83.025 224.760 83.110 225.085 ;
        RECT 85.795 224.915 85.870 225.245 ;
        RECT 88.535 224.915 88.630 225.245 ;
        RECT 91.350 224.835 91.390 225.165 ;
        RECT 94.125 224.815 94.150 225.145 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 144.130 225.115 144.225 225.445 ;
        RECT 77.515 224.755 77.845 224.760 ;
        RECT 83.025 224.755 83.355 224.760 ;
        RECT 8.560 200.860 146.080 202.460 ;
        RECT 6.000 197.560 146.080 199.160 ;
        RECT 118.090 171.510 118.680 173.070 ;
        RECT 127.100 113.755 152.575 114.380 ;
        RECT 151.950 1.000 152.575 113.755 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

